

module b15_C_gen_AntiSAT_k_256_7 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, 
        keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, 
        keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, 
        keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, 
        keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, 
        keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, 
        keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, 
        keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101, 
        keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105, 
        keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109, 
        keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113, 
        keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117, 
        keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121, 
        keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125, 
        keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67, 
        keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72, 
        keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77, 
        keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82, 
        keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87, 
        keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92, 
        keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97, 
        keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, U3445, U3446, U3447, U3448, U3213, U3212, 
        U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, 
        U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, 
        U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, 
        U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, 
        U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, 
        U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, 
        U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, 
        U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, 
        U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, 
        U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, 
        U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, 
        U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, 
        U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, 
        U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, 
        U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, 
        U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, 
        U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, 
        U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, 
        U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, 
        U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, 
        U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, 
        U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, 
        U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, 
        U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, 
        U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, 
        U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, 
        U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, 
        U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, 
        U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, 
        U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, 
        U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, 
        U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, 
        U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, 
        U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, 
        U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, 
        U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, 
        U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, 
        U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, 
        U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, 
        U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, 
        U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, 
        U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, 
        U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, 
        U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, 
        U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1,
         keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6,
         keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11,
         keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16,
         keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21,
         keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26,
         keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31,
         keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36,
         keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41,
         keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46,
         keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51,
         keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56,
         keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61,
         keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66,
         keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71,
         keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76,
         keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81,
         keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86,
         keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91,
         keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96,
         keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100,
         keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104,
         keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108,
         keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112,
         keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116,
         keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120,
         keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124,
         keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1,
         keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6,
         keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11,
         keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16,
         keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21,
         keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26,
         keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31,
         keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36,
         keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41,
         keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46,
         keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51,
         keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56,
         keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61,
         keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66,
         keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71,
         keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76,
         keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81,
         keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86,
         keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91,
         keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96,
         keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100,
         keyinput_g101, keyinput_g102, keyinput_g103, keyinput_g104,
         keyinput_g105, keyinput_g106, keyinput_g107, keyinput_g108,
         keyinput_g109, keyinput_g110, keyinput_g111, keyinput_g112,
         keyinput_g113, keyinput_g114, keyinput_g115, keyinput_g116,
         keyinput_g117, keyinput_g118, keyinput_g119, keyinput_g120,
         keyinput_g121, keyinput_g122, keyinput_g123, keyinput_g124,
         keyinput_g125, keyinput_g126, keyinput_g127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223;

  OR2_X1 U3597 ( .A1(n5207), .A2(n3179), .ZN(n4798) );
  NAND2_X1 U3598 ( .A1(n5805), .A2(n4693), .ZN(n5630) );
  NAND2_X1 U3599 ( .A1(n4627), .A2(n4628), .ZN(n5817) );
  AOI21_X1 U3600 ( .B1(n4034), .B2(n4648), .A(n4025), .ZN(n4026) );
  INV_X1 U3601 ( .A(n3644), .ZN(n5178) );
  OR2_X1 U3602 ( .A1(n3809), .A2(n3191), .ZN(n3765) );
  CLKBUF_X1 U3603 ( .A(n3571), .Z(n3691) );
  CLKBUF_X2 U3605 ( .A(n5087), .Z(n4882) );
  CLKBUF_X2 U3606 ( .A(n3539), .Z(n5081) );
  AND2_X1 U3607 ( .A1(n3452), .A2(n3629), .ZN(n3510) );
  BUF_X2 U3608 ( .A(n3771), .Z(n5069) );
  BUF_X1 U3609 ( .A(n3437), .Z(n3469) );
  NAND4_X1 U3610 ( .A1(n3382), .A2(n3381), .A3(n3380), .A4(n3379), .ZN(n3460)
         );
  AND2_X1 U3611 ( .A1(n3212), .A2(n3211), .ZN(n3187) );
  AND2_X2 U3612 ( .A1(n3218), .A2(n3920), .ZN(n5068) );
  NOR2_X1 U3613 ( .A1(n3501), .A2(n3500), .ZN(n3575) );
  AND4_X1 U3614 ( .A1(n3274), .A2(n3273), .A3(n3272), .A4(n3271), .ZN(n3292)
         );
  AND4_X1 U3615 ( .A1(n3394), .A2(n3393), .A3(n3392), .A4(n3391), .ZN(n3401)
         );
  AND4_X1 U3616 ( .A1(n3203), .A2(n3202), .A3(n3201), .A4(n3200), .ZN(n3212)
         );
  NAND2_X1 U3617 ( .A1(n3629), .A2(n4086), .ZN(n3644) );
  NAND2_X1 U3618 ( .A1(n3994), .A2(n3833), .ZN(n3868) );
  CLKBUF_X3 U3619 ( .A(n3501), .Z(n4086) );
  AND2_X1 U3620 ( .A1(n3640), .A2(n5178), .ZN(n3846) );
  CLKBUF_X2 U3622 ( .A(n3629), .Z(n4385) );
  INV_X1 U3623 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6828) );
  INV_X1 U3624 ( .A(n5996), .ZN(n5988) );
  AOI211_X1 U3625 ( .C1(INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n5527), .A(n5526), .B(n5525), .ZN(n5532) );
  INV_X1 U3626 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3668) );
  NAND2_X1 U3627 ( .A1(n4175), .A2(n4176), .ZN(n4281) );
  NOR2_X1 U3628 ( .A1(n3252), .A2(n3251), .ZN(n3270) );
  NOR2_X1 U3629 ( .A1(n4795), .A2(n5421), .ZN(n5413) );
  NAND2_X2 U3630 ( .A1(n3808), .A2(n3768), .ZN(n3906) );
  AND2_X1 U3633 ( .A1(n3219), .A2(n3217), .ZN(n3149) );
  OR2_X1 U3634 ( .A1(n3150), .A2(n5652), .ZN(n4781) );
  NAND2_X1 U3635 ( .A1(n3840), .A2(n3841), .ZN(n3984) );
  XNOR2_X1 U3636 ( .A(n3790), .B(n3789), .ZN(n3806) );
  XNOR2_X1 U3637 ( .A(n3922), .B(n6536), .ZN(n3891) );
  OAI211_X1 U3638 ( .C1(n3760), .C2(n3188), .A(n3585), .B(n3584), .ZN(n3758)
         );
  AOI21_X1 U3639 ( .B1(n3614), .B2(n3613), .A(n4282), .ZN(n3793) );
  INV_X1 U3640 ( .A(n3472), .ZN(n5167) );
  INV_X1 U3641 ( .A(n3475), .ZN(n3174) );
  AOI21_X1 U3642 ( .B1(n3598), .B2(INSTQUEUE_REG_13__2__SCAN_IN), .A(n3390), 
        .ZN(n3402) );
  CLKBUF_X2 U3644 ( .A(n3600), .Z(n5070) );
  XNOR2_X1 U3646 ( .A(n4798), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5194)
         );
  OAI21_X1 U3647 ( .B1(n5448), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n5437), 
        .ZN(n5438) );
  AND2_X1 U3648 ( .A1(n5413), .A2(n3158), .ZN(n5207) );
  OR2_X1 U3649 ( .A1(n5465), .A2(n5464), .ZN(n5435) );
  NAND2_X1 U3650 ( .A1(n5323), .A2(n5324), .ZN(n5260) );
  CLKBUF_X1 U3651 ( .A(n5323), .Z(n5417) );
  NOR2_X1 U3652 ( .A1(n5332), .A2(n5334), .ZN(n5333) );
  NAND2_X1 U3654 ( .A1(n5187), .A2(n5186), .ZN(n5257) );
  INV_X2 U3655 ( .A(n5489), .ZN(n3150) );
  OAI21_X2 U3656 ( .B1(n4244), .B2(n4283), .A(n4243), .ZN(n4293) );
  AOI21_X1 U3657 ( .B1(n4297), .B2(n4648), .A(n4268), .ZN(n4274) );
  XNOR2_X1 U3658 ( .A(n4281), .B(n4264), .ZN(n4297) );
  NAND2_X1 U3659 ( .A1(n4015), .A2(n4014), .ZN(n4178) );
  NAND2_X1 U3660 ( .A1(n3804), .A2(n3803), .ZN(n3840) );
  OAI21_X1 U3661 ( .B1(n6806), .B2(n4599), .A(n3839), .ZN(n3841) );
  OR2_X1 U3662 ( .A1(n3802), .A2(n3798), .ZN(n3856) );
  AND2_X1 U3663 ( .A1(n3626), .A2(n3627), .ZN(n3798) );
  NAND2_X2 U3664 ( .A1(n6022), .A2(n4155), .ZN(n6012) );
  NAND2_X1 U3665 ( .A1(n3891), .A2(n6828), .ZN(n3831) );
  BUF_X1 U3666 ( .A(n3792), .Z(n3620) );
  NAND2_X1 U3667 ( .A1(n3977), .A2(n3976), .ZN(n4031) );
  AND2_X1 U3668 ( .A1(n3765), .A2(n3764), .ZN(n3766) );
  NAND2_X1 U3669 ( .A1(n3815), .A2(n3814), .ZN(n6536) );
  OAI21_X1 U3670 ( .B1(n3611), .B2(n3613), .A(n3566), .ZN(n6811) );
  NAND2_X1 U3671 ( .A1(n3498), .A2(n3705), .ZN(n3515) );
  NAND2_X1 U3672 ( .A1(n3564), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3611) );
  AOI22_X1 U3673 ( .A1(n3997), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3788), 
        .B2(n3787), .ZN(n3789) );
  AND2_X1 U3675 ( .A1(n3638), .A2(n3637), .ZN(n3701) );
  INV_X2 U3676 ( .A(n5178), .ZN(n5168) );
  OR2_X1 U3677 ( .A1(n4156), .A2(n3745), .ZN(n3477) );
  AOI21_X1 U3678 ( .B1(n3459), .B2(n4081), .A(n5220), .ZN(n3434) );
  OR2_X1 U3679 ( .A1(n3561), .A2(n3560), .ZN(n3742) );
  AND3_X1 U3680 ( .A1(n3573), .A2(n3572), .A3(n3571), .ZN(n3631) );
  INV_X1 U3681 ( .A(n3475), .ZN(n3842) );
  NAND2_X1 U3682 ( .A1(n3510), .A2(n3572), .ZN(n5157) );
  AND2_X1 U3683 ( .A1(n3469), .A2(n4155), .ZN(n4772) );
  CLKBUF_X1 U3684 ( .A(n3575), .Z(n3576) );
  INV_X1 U3686 ( .A(n3361), .ZN(n3457) );
  INV_X1 U3687 ( .A(n4081), .ZN(n3572) );
  AND4_X2 U3688 ( .A1(n3177), .A2(n3402), .A3(n3401), .A4(n3400), .ZN(n3571)
         );
  AND4_X1 U3689 ( .A1(n3258), .A2(n3257), .A3(n3256), .A4(n3255), .ZN(n3269)
         );
  AND4_X1 U3690 ( .A1(n3399), .A2(n3398), .A3(n3397), .A4(n3396), .ZN(n3400)
         );
  AND4_X1 U3691 ( .A1(n3366), .A2(n3365), .A3(n3364), .A4(n3363), .ZN(n3382)
         );
  AND4_X1 U3692 ( .A1(n3210), .A2(n3209), .A3(n3208), .A4(n3207), .ZN(n3211)
         );
  NAND4_X1 U3693 ( .A1(n3360), .A2(n3359), .A3(n3358), .A4(n3357), .ZN(n3437)
         );
  NAND2_X2 U3694 ( .A1(STATE_REG_2__SCAN_IN), .A2(n7221), .ZN(n6787) );
  AND4_X1 U3695 ( .A1(n3282), .A2(n3281), .A3(n3280), .A4(n3279), .ZN(n3290)
         );
  AND4_X1 U3696 ( .A1(n3262), .A2(n3261), .A3(n3260), .A4(n3259), .ZN(n3268)
         );
  AND4_X1 U3697 ( .A1(n3244), .A2(n3243), .A3(n3242), .A4(n3241), .ZN(n3245)
         );
  AND4_X1 U3698 ( .A1(n3344), .A2(n3343), .A3(n3342), .A4(n3341), .ZN(n3360)
         );
  AND4_X1 U3699 ( .A1(n3348), .A2(n3347), .A3(n3346), .A4(n3345), .ZN(n3359)
         );
  AND4_X1 U3700 ( .A1(n3352), .A2(n3351), .A3(n3350), .A4(n3349), .ZN(n3358)
         );
  AND4_X1 U3701 ( .A1(n3356), .A2(n3355), .A3(n3354), .A4(n3353), .ZN(n3357)
         );
  AND4_X1 U3702 ( .A1(n3411), .A2(n3410), .A3(n3409), .A4(n3408), .ZN(n3426)
         );
  AND4_X1 U3703 ( .A1(n3417), .A2(n3416), .A3(n3415), .A4(n3414), .ZN(n3425)
         );
  AND4_X1 U3704 ( .A1(n3370), .A2(n3369), .A3(n3368), .A4(n3367), .ZN(n3381)
         );
  AND4_X1 U3705 ( .A1(n3406), .A2(n3405), .A3(n3404), .A4(n3403), .ZN(n3427)
         );
  INV_X2 U3706 ( .A(n5074), .ZN(n5018) );
  AND4_X1 U3707 ( .A1(n3423), .A2(n3422), .A3(n3421), .A4(n3420), .ZN(n3424)
         );
  AND4_X1 U3708 ( .A1(n3374), .A2(n3373), .A3(n3372), .A4(n3371), .ZN(n3380)
         );
  AND4_X1 U3709 ( .A1(n3266), .A2(n3265), .A3(n3264), .A4(n3263), .ZN(n3267)
         );
  AND4_X1 U3710 ( .A1(n3224), .A2(n3223), .A3(n3222), .A4(n3221), .ZN(n3225)
         );
  AND4_X1 U3711 ( .A1(n3378), .A2(n3377), .A3(n3376), .A4(n3375), .ZN(n3379)
         );
  CLKBUF_X2 U3712 ( .A(n3598), .Z(n5080) );
  BUF_X2 U3713 ( .A(n3555), .Z(n5075) );
  AND2_X1 U3714 ( .A1(n5051), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3252) );
  OR2_X2 U3715 ( .A1(n6745), .A2(n6802), .ZN(n5512) );
  INV_X2 U3716 ( .A(n7220), .ZN(n7221) );
  AND2_X2 U3717 ( .A1(n3218), .A2(n3220), .ZN(n3597) );
  AND2_X2 U3718 ( .A1(n3218), .A2(n5669), .ZN(n3770) );
  AND2_X1 U3719 ( .A1(n3196), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3220)
         );
  CLKBUF_X1 U3720 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n5197) );
  INV_X1 U3721 ( .A(n3151), .ZN(n3663) );
  NAND2_X1 U3724 ( .A1(n5109), .A2(n5112), .ZN(n5111) );
  OR2_X2 U3725 ( .A1(n4549), .A2(n4548), .ZN(n4564) );
  OAI21_X2 U3726 ( .B1(n5227), .B2(EBX_REG_1__SCAN_IN), .A(n3636), .ZN(n3844)
         );
  NAND2_X1 U3727 ( .A1(n5111), .A2(n3156), .ZN(n3153) );
  AND2_X2 U3728 ( .A1(n3153), .A2(n3154), .ZN(n5496) );
  OR2_X1 U3729 ( .A1(n3155), .A2(n4781), .ZN(n3154) );
  INV_X1 U3730 ( .A(n4782), .ZN(n3155) );
  AND2_X1 U3731 ( .A1(n4780), .A2(n4782), .ZN(n3156) );
  NAND2_X1 U3732 ( .A1(n3508), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3157) );
  AND2_X1 U3733 ( .A1(n5530), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3158)
         );
  NAND4_X1 U3734 ( .A1(n3270), .A2(n3269), .A3(n3268), .A4(n3267), .ZN(n3159)
         );
  NAND2_X1 U3735 ( .A1(n3508), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3760) );
  NAND4_X1 U3736 ( .A1(n3270), .A2(n3269), .A3(n3268), .A4(n3267), .ZN(n3431)
         );
  CLKBUF_X1 U3737 ( .A(n4292), .Z(n3160) );
  CLKBUF_X1 U3738 ( .A(n4238), .Z(n3161) );
  OAI21_X1 U3740 ( .B1(n3868), .B2(n4283), .A(n3867), .ZN(n3163) );
  OAI21_X1 U3741 ( .B1(n3868), .B2(n4283), .A(n3867), .ZN(n3970) );
  OAI21_X2 U3742 ( .B1(n3939), .B2(STATE2_REG_0__SCAN_IN), .A(n3608), .ZN(
        n3168) );
  NOR2_X4 U3743 ( .A1(n4564), .A2(n4565), .ZN(n4627) );
  NOR2_X2 U3744 ( .A1(n4031), .A2(n4032), .ZN(n4277) );
  NAND2_X1 U3745 ( .A1(n3972), .A2(n3971), .ZN(n4043) );
  INV_X1 U3746 ( .A(n5364), .ZN(n3164) );
  NOR2_X2 U3747 ( .A1(n4767), .A2(n3165), .ZN(n5308) );
  NAND2_X1 U3748 ( .A1(n4768), .A2(n3164), .ZN(n3165) );
  AND2_X1 U3749 ( .A1(n4605), .A2(n3167), .ZN(n3166) );
  INV_X1 U3750 ( .A(n4655), .ZN(n3167) );
  NOR2_X1 U3751 ( .A1(n5260), .A2(n5262), .ZN(n3169) );
  NAND2_X1 U3752 ( .A1(n4967), .A2(n4966), .ZN(n3170) );
  NOR2_X2 U3753 ( .A1(n3170), .A2(n3171), .ZN(n5323) );
  OR2_X1 U3754 ( .A1(n3172), .A2(n5334), .ZN(n3171) );
  INV_X1 U3755 ( .A(n5415), .ZN(n3172) );
  XNOR2_X1 U3756 ( .A(n3620), .B(n3791), .ZN(n3173) );
  XNOR2_X1 U3757 ( .A(n3620), .B(n3791), .ZN(n3934) );
  AND2_X1 U3758 ( .A1(n5260), .A2(n5325), .ZN(n5685) );
  NOR2_X1 U3759 ( .A1(n3612), .A2(n6828), .ZN(n4282) );
  NOR2_X1 U3760 ( .A1(n4695), .A2(n6828), .ZN(n5096) );
  NOR2_X1 U3761 ( .A1(n3469), .A2(n6637), .ZN(n4648) );
  INV_X1 U3762 ( .A(n5008), .ZN(n5211) );
  NOR2_X2 U3763 ( .A1(n5260), .A2(n5262), .ZN(n5261) );
  CLKBUF_X1 U3764 ( .A(n3204), .Z(n3188) );
  NAND2_X1 U3765 ( .A1(n3194), .A2(n3193), .ZN(n3303) );
  AND2_X1 U3766 ( .A1(n3303), .A2(n3195), .ZN(n3299) );
  NOR2_X1 U3767 ( .A1(n3299), .A2(n3298), .ZN(n3297) );
  INV_X1 U3768 ( .A(n3787), .ZN(n3870) );
  AOI21_X1 U3769 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n6810), .A(n3297), 
        .ZN(n3294) );
  NOR2_X1 U3770 ( .A1(n4513), .A2(n4512), .ZN(n4514) );
  OR2_X1 U3771 ( .A1(n4511), .A2(n4510), .ZN(n4512) );
  NAND2_X1 U3772 ( .A1(n6637), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4710) );
  NAND2_X1 U3773 ( .A1(n4281), .A2(n4285), .ZN(n4664) );
  OR3_X1 U3774 ( .A1(n3662), .A2(n3661), .A3(n4150), .ZN(n3925) );
  AND2_X1 U3775 ( .A1(n3293), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4261) );
  CLKBUF_X1 U3776 ( .A(n3570), .Z(n3305) );
  OR2_X1 U3777 ( .A1(n4152), .A2(n3577), .ZN(n6062) );
  NOR2_X1 U3778 ( .A1(n5036), .A2(n5408), .ZN(n5040) );
  OAI21_X1 U3779 ( .B1(n5101), .B2(n5397), .A(n5065), .ZN(n5262) );
  AOI21_X1 U3780 ( .B1(n5039), .B2(n5038), .A(n5037), .ZN(n5324) );
  AND2_X1 U3781 ( .A1(n4694), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4761)
         );
  NOR2_X1 U3782 ( .A1(n3150), .A2(n4678), .ZN(n4778) );
  AOI21_X1 U3783 ( .B1(n3985), .B2(n4648), .A(n3991), .ZN(n4122) );
  OR2_X1 U3784 ( .A1(n3150), .A2(n4665), .ZN(n4675) );
  NAND2_X1 U3785 ( .A1(n3696), .A2(n6738), .ZN(n3722) );
  CLKBUF_X1 U3786 ( .A(n3173), .Z(n3935) );
  NOR2_X1 U3787 ( .A1(n6427), .A2(n6811), .ZN(n6395) );
  OR2_X1 U3788 ( .A1(n3809), .A2(n3903), .ZN(n3815) );
  INV_X1 U3789 ( .A(n5934), .ZN(n5977) );
  AND2_X1 U3790 ( .A1(n5931), .A2(n4377), .ZN(n5996) );
  NAND2_X1 U3791 ( .A1(n5786), .A2(n6116), .ZN(n6111) );
  AND2_X1 U3792 ( .A1(n6714), .A2(n6738), .ZN(n6115) );
  INV_X1 U3793 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6819) );
  AND2_X1 U3794 ( .A1(n3305), .A2(n3306), .ZN(n3318) );
  NAND2_X2 U3795 ( .A1(n3894), .A2(n5669), .ZN(n4947) );
  AOI21_X1 U3796 ( .B1(n3573), .B2(n3503), .A(n3502), .ZN(n3504) );
  NAND2_X1 U3797 ( .A1(n3438), .A2(n3460), .ZN(n3496) );
  NAND2_X1 U3798 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6819), .ZN(n3313) );
  AND2_X1 U3799 ( .A1(n3309), .A2(n3190), .ZN(n3302) );
  NAND2_X1 U3800 ( .A1(n4281), .A2(n4179), .ZN(n4244) );
  NAND2_X1 U3801 ( .A1(n4178), .A2(n4177), .ZN(n4179) );
  OR2_X1 U3802 ( .A1(n4011), .A2(n4010), .ZN(n4038) );
  OR2_X1 U3803 ( .A1(n3963), .A2(n3962), .ZN(n4035) );
  NAND2_X1 U3804 ( .A1(n3717), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3786) );
  AND2_X2 U3805 ( .A1(n3197), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3217)
         );
  NAND2_X1 U3806 ( .A1(n3457), .A2(n3432), .ZN(n3430) );
  NAND2_X1 U3807 ( .A1(n3591), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3208)
         );
  NAND2_X1 U3808 ( .A1(n3206), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3210)
         );
  NAND2_X1 U3809 ( .A1(n3771), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3213) );
  NAND2_X1 U3810 ( .A1(n5087), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3221) );
  OR2_X1 U3811 ( .A1(n3528), .A2(n3283), .ZN(n3288) );
  INV_X1 U3812 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3283) );
  OR2_X1 U3813 ( .A1(n3528), .A2(n3253), .ZN(n3258) );
  INV_X1 U3814 ( .A(n4263), .ZN(n3997) );
  AOI211_X1 U3815 ( .C1(n3299), .C2(n3298), .A(n3297), .B(n3296), .ZN(n3445)
         );
  AND2_X1 U3816 ( .A1(n3295), .A2(n5831), .ZN(n3296) );
  NAND2_X1 U3817 ( .A1(n3583), .A2(n3181), .ZN(n3586) );
  BUF_X1 U3818 ( .A(n3429), .Z(n3573) );
  INV_X1 U3819 ( .A(n5342), .ZN(n4966) );
  INV_X1 U3820 ( .A(n4771), .ZN(n4768) );
  INV_X1 U3821 ( .A(n4648), .ZN(n4599) );
  AOI21_X1 U3822 ( .B1(n5443), .B2(n4793), .A(n3185), .ZN(n5402) );
  OR2_X1 U3823 ( .A1(n3150), .A2(n5497), .ZN(n4783) );
  AND2_X1 U3824 ( .A1(n3150), .A2(n5497), .ZN(n4784) );
  NAND2_X1 U3825 ( .A1(n5178), .A2(n3842), .ZN(n5170) );
  INV_X1 U3826 ( .A(n5227), .ZN(n5171) );
  NAND2_X1 U3827 ( .A1(n3796), .A2(n3795), .ZN(n3805) );
  AND2_X1 U3828 ( .A1(n3517), .A2(n3516), .ZN(n3518) );
  AND2_X2 U3829 ( .A1(n3917), .A2(n5669), .ZN(n3591) );
  AND2_X1 U3830 ( .A1(n3811), .A2(n6634), .ZN(n6397) );
  OAI21_X1 U3831 ( .B1(n6747), .B2(n3890), .A(n6733), .ZN(n4079) );
  INV_X1 U3832 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6704) );
  INV_X1 U3833 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3903) );
  AND2_X1 U3834 ( .A1(n3710), .A2(n3683), .ZN(n3893) );
  AND2_X1 U3835 ( .A1(n4916), .A2(n4915), .ZN(n5280) );
  CLKBUF_X1 U3836 ( .A(n3510), .Z(n5239) );
  AOI21_X1 U3837 ( .B1(n5104), .B2(n5103), .A(n5102), .ZN(n5209) );
  AND2_X1 U3838 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n4368), .ZN(n5012)
         );
  NOR2_X1 U3839 ( .A1(n4935), .A2(n4367), .ZN(n4962) );
  CLKBUF_X1 U3840 ( .A(n5339), .Z(n5340) );
  NOR2_X1 U3841 ( .A1(n4879), .A2(n5459), .ZN(n4913) );
  CLKBUF_X1 U3842 ( .A(n5278), .Z(n5279) );
  AND2_X1 U3843 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n4366), .ZN(n4857)
         );
  NAND2_X1 U3844 ( .A1(n4857), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4879)
         );
  CLKBUF_X1 U3845 ( .A(n5292), .Z(n5293) );
  AND2_X1 U3846 ( .A1(n4839), .A2(n4838), .ZN(n5310) );
  NOR2_X1 U3847 ( .A1(n4760), .A2(n4365), .ZN(n4799) );
  CLKBUF_X1 U3848 ( .A(n5308), .Z(n5309) );
  CLKBUF_X1 U3849 ( .A(n4767), .Z(n4766) );
  NOR2_X1 U3850 ( .A1(n4635), .A2(n4364), .ZN(n4694) );
  CLKBUF_X1 U3851 ( .A(n4741), .Z(n4716) );
  CLKBUF_X1 U3852 ( .A(n4715), .Z(n4657) );
  NOR2_X1 U3853 ( .A1(n4516), .A2(n4363), .ZN(n4582) );
  INV_X1 U3854 ( .A(n4555), .ZN(n4578) );
  NOR2_X1 U3855 ( .A1(n4504), .A2(n4362), .ZN(n4470) );
  AND2_X1 U3856 ( .A1(n4457), .A2(n4508), .ZN(n4558) );
  NAND2_X1 U3857 ( .A1(n4361), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4394)
         );
  INV_X1 U3858 ( .A(n4360), .ZN(n4361) );
  NOR2_X1 U3859 ( .A1(n4415), .A2(n4510), .ZN(n4457) );
  NAND2_X1 U3860 ( .A1(n4265), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4360)
         );
  CLKBUF_X1 U3861 ( .A(n4469), .Z(n4272) );
  AND2_X1 U3862 ( .A1(n4182), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4265)
         );
  INV_X1 U3863 ( .A(n4122), .ZN(n3992) );
  INV_X1 U3864 ( .A(n3834), .ZN(n3835) );
  NAND2_X1 U3865 ( .A1(n3835), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3988)
         );
  OAI211_X1 U3866 ( .C1(n3801), .C2(n3191), .A(n3800), .B(n3799), .ZN(n3857)
         );
  NAND2_X1 U3867 ( .A1(n5367), .A2(n5152), .ZN(n5299) );
  NAND2_X1 U3868 ( .A1(n5149), .A2(n5148), .ZN(n5151) );
  AND2_X1 U3869 ( .A1(n5629), .A2(n5368), .ZN(n5367) );
  CLKBUF_X1 U3870 ( .A(n5443), .Z(n5444) );
  NOR2_X2 U3871 ( .A1(n5630), .A2(n5631), .ZN(n5629) );
  CLKBUF_X1 U3872 ( .A(n5477), .Z(n5478) );
  AND2_X1 U3873 ( .A1(n3150), .A2(n4538), .ZN(n4661) );
  OR2_X1 U3874 ( .A1(n3150), .A2(n4538), .ZN(n4660) );
  NAND2_X1 U3875 ( .A1(n4315), .A2(n4314), .ZN(n4549) );
  NOR2_X1 U3876 ( .A1(n5677), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3813) );
  OR2_X1 U3877 ( .A1(n3722), .A2(n3711), .ZN(n5649) );
  OR2_X1 U3878 ( .A1(n3722), .A2(n5666), .ZN(n4048) );
  NAND2_X1 U3879 ( .A1(n5167), .A2(n3842), .ZN(n5234) );
  CLKBUF_X1 U3880 ( .A(n3906), .Z(n3907) );
  AND2_X1 U3881 ( .A1(n6217), .A2(n6812), .ZN(n6219) );
  CLKBUF_X1 U3882 ( .A(n3891), .Z(n6319) );
  INV_X1 U3883 ( .A(n3571), .ZN(n4108) );
  AND2_X1 U3884 ( .A1(n3933), .A2(n6188), .ZN(n6640) );
  NAND2_X1 U3885 ( .A1(n3338), .A2(n3337), .ZN(n3735) );
  INV_X1 U3886 ( .A(n5101), .ZN(n5060) );
  INV_X1 U3887 ( .A(n5997), .ZN(n5872) );
  INV_X1 U3888 ( .A(n5992), .ZN(n5965) );
  OR3_X1 U3889 ( .A1(n6830), .A2(n4387), .A3(n4386), .ZN(n5934) );
  CLKBUF_X1 U3890 ( .A(n3939), .Z(n3940) );
  AND2_X1 U3891 ( .A1(n5931), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5997) );
  AND2_X1 U3892 ( .A1(n4372), .A2(n5937), .ZN(n5994) );
  INV_X1 U3893 ( .A(n6033), .ZN(n6026) );
  AND2_X1 U3894 ( .A1(n6032), .A2(n4772), .ZN(n6029) );
  AND2_X1 U3895 ( .A1(n5219), .A2(n4157), .ZN(n6030) );
  INV_X1 U3896 ( .A(n6030), .ZN(n5391) );
  NOR2_X1 U3897 ( .A1(n6037), .A2(n4063), .ZN(n6047) );
  CLKBUF_X1 U3899 ( .A(n6093), .Z(n6097) );
  OR2_X1 U3900 ( .A1(n5100), .A2(n5252), .ZN(n4370) );
  AOI21_X1 U3901 ( .B1(n5262), .B2(n5260), .A(n3169), .ZN(n5399) );
  CLKBUF_X1 U3902 ( .A(n5496), .Z(n5499) );
  CLKBUF_X1 U3903 ( .A(n4779), .Z(n4677) );
  INV_X1 U3904 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4127) );
  INV_X1 U3905 ( .A(n6111), .ZN(n5781) );
  INV_X2 U3906 ( .A(n5512), .ZN(n6113) );
  AND2_X1 U3907 ( .A1(n5580), .A2(n5582), .ZN(n5575) );
  OR2_X1 U3908 ( .A1(n6138), .A2(n5595), .ZN(n5634) );
  INV_X1 U3909 ( .A(n6163), .ZN(n6172) );
  CLKBUF_X1 U3910 ( .A(n3932), .Z(n3933) );
  INV_X1 U3911 ( .A(n6812), .ZN(n6802) );
  INV_X1 U3912 ( .A(n6808), .ZN(n6818) );
  BUF_X1 U3913 ( .A(n3657), .Z(n5825) );
  OR2_X1 U3914 ( .A1(n6406), .A2(n6405), .ZN(n6424) );
  OR2_X1 U3915 ( .A1(n6540), .A2(n6539), .ZN(n6558) );
  NAND2_X1 U3916 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n3735), .ZN(n6733) );
  CLKBUF_X1 U3917 ( .A(n6789), .Z(n6788) );
  AOI21_X1 U3918 ( .B1(n5377), .B2(n6113), .A(n5107), .ZN(n5108) );
  INV_X1 U3919 ( .A(n3437), .ZN(n3432) );
  AND2_X2 U3920 ( .A1(n3920), .A2(n3217), .ZN(n3555) );
  OR2_X1 U3921 ( .A1(n3150), .A2(n6146), .ZN(n3175) );
  INV_X1 U3922 ( .A(n3431), .ZN(n3429) );
  INV_X1 U3923 ( .A(n6025), .ZN(n6032) );
  OAI211_X1 U3924 ( .C1(n3663), .C2(n4154), .A(n4153), .B(n6102), .ZN(n5219)
         );
  NAND2_X1 U3925 ( .A1(n4190), .A2(n4189), .ZN(n4192) );
  INV_X1 U3926 ( .A(n4664), .ZN(n5489) );
  BUF_X1 U3927 ( .A(n4664), .Z(n5432) );
  INV_X1 U3928 ( .A(n3458), .ZN(n3512) );
  CLKBUF_X1 U3929 ( .A(n3157), .Z(n3809) );
  XNOR2_X1 U3930 ( .A(n5261), .B(n5105), .ZN(n5377) );
  NAND2_X1 U3931 ( .A1(n4578), .A2(n4577), .ZN(n4579) );
  OR2_X1 U3932 ( .A1(n5514), .A2(n4797), .ZN(n3176) );
  AND4_X1 U3933 ( .A1(n3386), .A2(n3385), .A3(n3384), .A4(n3383), .ZN(n3177)
         );
  AND4_X1 U3934 ( .A1(n3216), .A2(n3215), .A3(n3214), .A4(n3213), .ZN(n3178)
         );
  AND2_X1 U3935 ( .A1(n5401), .A2(n4796), .ZN(n3179) );
  AND3_X1 U3936 ( .A1(n3150), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3180) );
  OR2_X1 U3937 ( .A1(n3582), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3181)
         );
  AND2_X1 U3938 ( .A1(n5366), .A2(n3174), .ZN(n3182) );
  NOR2_X1 U3939 ( .A1(n5417), .A2(n5416), .ZN(n3183) );
  AND2_X1 U3940 ( .A1(n5432), .A2(n5431), .ZN(n3184) );
  AND2_X1 U3941 ( .A1(n3619), .A2(n3618), .ZN(n3791) );
  AND2_X1 U3942 ( .A1(n5489), .A2(n4792), .ZN(n3185) );
  AND2_X1 U3943 ( .A1(n5489), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3186)
         );
  INV_X1 U3944 ( .A(n3496), .ZN(n3470) );
  INV_X1 U3945 ( .A(n6404), .ZN(n6256) );
  INV_X1 U3946 ( .A(n3318), .ZN(n3327) );
  INV_X1 U3947 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3199) );
  OR2_X1 U3948 ( .A1(n3606), .A2(n3605), .ZN(n3743) );
  OR2_X1 U3949 ( .A1(n3785), .A2(n3784), .ZN(n3787) );
  NAND2_X1 U3950 ( .A1(n3429), .A2(n3437), .ZN(n3455) );
  INV_X1 U3951 ( .A(n3302), .ZN(n3194) );
  AND2_X1 U3952 ( .A1(n4013), .A2(n4012), .ZN(n4016) );
  OR2_X1 U3953 ( .A1(n4947), .A2(n3340), .ZN(n3341) );
  INV_X1 U3954 ( .A(n4176), .ZN(n4177) );
  INV_X1 U3955 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3197) );
  AND4_X1 U3956 ( .A1(n3533), .A2(n3532), .A3(n3531), .A4(n3530), .ZN(n3537)
         );
  OR2_X1 U3957 ( .A1(n3307), .A2(n3313), .ZN(n3309) );
  NAND2_X1 U3958 ( .A1(n5087), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3392) );
  NAND2_X1 U3959 ( .A1(n3254), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3257) );
  INV_X1 U3960 ( .A(n4274), .ZN(n4270) );
  INV_X1 U3961 ( .A(n5295), .ZN(n4860) );
  INV_X1 U3962 ( .A(n5779), .ZN(n4764) );
  OR2_X1 U3963 ( .A1(n4947), .A2(n3413), .ZN(n3414) );
  OR2_X1 U3964 ( .A1(n3829), .A2(n3828), .ZN(n3866) );
  AND4_X1 U3965 ( .A1(n3288), .A2(n3287), .A3(n3286), .A4(n3285), .ZN(n3289)
         );
  AND4_X1 U3966 ( .A1(n3278), .A2(n3277), .A3(n3276), .A4(n3275), .ZN(n3291)
         );
  NAND2_X1 U3967 ( .A1(n3723), .A2(n3452), .ZN(n3570) );
  AND2_X1 U3968 ( .A1(n5014), .A2(n5013), .ZN(n5415) );
  INV_X1 U3969 ( .A(n4837), .ZN(n4366) );
  INV_X1 U3970 ( .A(n5096), .ZN(n5063) );
  OR2_X1 U3971 ( .A1(n4155), .A2(n6478), .ZN(n5008) );
  INV_X1 U3972 ( .A(n4949), .ZN(n5082) );
  INV_X1 U3973 ( .A(n3634), .ZN(n3475) );
  NAND2_X1 U3974 ( .A1(n4385), .A2(n4091), .ZN(n3293) );
  NAND2_X1 U3975 ( .A1(n4081), .A2(n3501), .ZN(n3634) );
  NOR2_X1 U3976 ( .A1(n5151), .A2(n3182), .ZN(n5152) );
  NAND2_X1 U3977 ( .A1(n4913), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4935)
         );
  NAND2_X1 U3978 ( .A1(n4438), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4504)
         );
  NAND2_X1 U3979 ( .A1(n5345), .A2(n5335), .ZN(n5543) );
  INV_X1 U3980 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5433) );
  INV_X1 U3981 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3881) );
  CLKBUF_X1 U3982 ( .A(n3920), .Z(n5670) );
  OR2_X1 U3983 ( .A1(n3293), .A2(n6828), .ZN(n4263) );
  AND2_X1 U3984 ( .A1(n4080), .A2(n4079), .ZN(n4114) );
  NAND2_X1 U3985 ( .A1(n5012), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5036)
         );
  NOR2_X1 U3986 ( .A1(n6983), .A2(n5860), .ZN(n5747) );
  AND2_X1 U3987 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n4019), .ZN(n4182)
         );
  NOR2_X1 U3988 ( .A1(n3988), .A2(n4127), .ZN(n4019) );
  OR2_X1 U3989 ( .A1(n4547), .A2(n4546), .ZN(n4548) );
  INV_X1 U3990 ( .A(n5209), .ZN(n5105) );
  NOR2_X1 U3991 ( .A1(n4394), .A2(n4422), .ZN(n4438) );
  INV_X1 U3992 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4797) );
  NAND2_X1 U3993 ( .A1(n3882), .A2(n3881), .ZN(n6104) );
  OR2_X1 U3994 ( .A1(n3722), .A2(n3702), .ZN(n5645) );
  OR2_X1 U3995 ( .A1(n4208), .A2(n6811), .ZN(n6251) );
  OR2_X1 U3996 ( .A1(n6279), .A2(n6589), .ZN(n6326) );
  INV_X1 U3997 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6400) );
  OR2_X1 U3998 ( .A1(n6806), .A2(n3933), .ZN(n6427) );
  INV_X1 U3999 ( .A(n6319), .ZN(n6804) );
  NAND2_X1 U4000 ( .A1(n6828), .A2(n4079), .ZN(n6404) );
  NOR2_X1 U4001 ( .A1(n6783), .A2(n5314), .ZN(n5297) );
  NAND2_X1 U4002 ( .A1(n4761), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4760)
         );
  NAND2_X1 U4003 ( .A1(n6830), .A2(n4359), .ZN(n5931) );
  INV_X1 U4004 ( .A(n5937), .ZN(n5951) );
  INV_X1 U4005 ( .A(n6000), .ZN(n5980) );
  AND2_X1 U4006 ( .A1(n6062), .A2(n3494), .ZN(n6830) );
  NOR2_X2 U4007 ( .A1(n5350), .A2(n5349), .ZN(n5351) );
  INV_X1 U4008 ( .A(n6011), .ZN(n6018) );
  BUF_X1 U4009 ( .A(n3460), .Z(n4155) );
  INV_X1 U4010 ( .A(n5219), .ZN(n6025) );
  AND2_X1 U4011 ( .A1(n3440), .A2(n4380), .ZN(n6037) );
  NAND2_X1 U4012 ( .A1(n3735), .A2(n6738), .ZN(n4152) );
  NAND2_X1 U4013 ( .A1(n4962), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4989)
         );
  NAND2_X1 U4014 ( .A1(n4799), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4837)
         );
  AND2_X1 U4015 ( .A1(n4558), .A2(n4557), .ZN(n4560) );
  NAND2_X1 U4016 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3834) );
  INV_X1 U4017 ( .A(n5786), .ZN(n6117) );
  OAI211_X1 U4018 ( .C1(n5191), .C2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n3176), .B(n5190), .ZN(n5192) );
  AND2_X1 U4019 ( .A1(n5575), .A2(n5133), .ZN(n5792) );
  NAND2_X1 U4020 ( .A1(n5435), .A2(n5434), .ZN(n5457) );
  INV_X1 U4021 ( .A(n6125), .ZN(n6175) );
  INV_X1 U4022 ( .A(n5197), .ZN(n3191) );
  INV_X1 U4023 ( .A(n6251), .ZN(n6274) );
  INV_X1 U4024 ( .A(n4236), .ZN(n4118) );
  OR2_X1 U4025 ( .A1(n6351), .A2(n3935), .ZN(n6279) );
  INV_X1 U4026 ( .A(n6326), .ZN(n6343) );
  INV_X1 U4027 ( .A(n6401), .ZN(n6423) );
  INV_X1 U4028 ( .A(n3935), .ZN(n6394) );
  INV_X1 U4029 ( .A(n6593), .ZN(n6628) );
  AND2_X1 U4030 ( .A1(n6640), .A2(n6811), .ZN(n6690) );
  INV_X1 U4031 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6728) );
  INV_X1 U4032 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6912) );
  OR3_X1 U4033 ( .A1(n6830), .A2(n5168), .A3(n4375), .ZN(n5992) );
  NAND2_X1 U4034 ( .A1(n5931), .A2(n4371), .ZN(n5937) );
  OR2_X1 U4035 ( .A1(n6830), .A2(n4383), .ZN(n6000) );
  OR2_X1 U4036 ( .A1(n4558), .A2(n4458), .ZN(n5910) );
  NAND2_X1 U4037 ( .A1(n6032), .A2(n4158), .ZN(n4659) );
  INV_X1 U4038 ( .A(n6037), .ZN(n6061) );
  OR2_X1 U4039 ( .A1(n6115), .A2(n3736), .ZN(n5786) );
  OR2_X1 U4040 ( .A1(n4560), .A2(n4559), .ZN(n4672) );
  INV_X1 U4041 ( .A(n6115), .ZN(n5835) );
  NOR2_X1 U4042 ( .A1(n5651), .A2(n6121), .ZN(n6138) );
  OR2_X1 U4043 ( .A1(n3722), .A2(n3721), .ZN(n6125) );
  OR2_X1 U4044 ( .A1(n3722), .A2(n3699), .ZN(n6163) );
  INV_X1 U4045 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6810) );
  OR2_X1 U4046 ( .A1(n6216), .A2(n6811), .ZN(n6243) );
  OR2_X1 U4047 ( .A1(n6216), .A2(n6589), .ZN(n6278) );
  OR2_X1 U4048 ( .A1(n4208), .A2(n6589), .ZN(n4236) );
  OR2_X1 U4049 ( .A1(n6279), .A2(n6811), .ZN(n6316) );
  OR3_X1 U4050 ( .A1(n6351), .A2(n6394), .A3(n6811), .ZN(n6386) );
  NAND2_X1 U4051 ( .A1(n6395), .A2(n6394), .ZN(n6464) );
  NAND2_X1 U4052 ( .A1(n6434), .A2(n6428), .ZN(n6516) );
  NAND2_X1 U4053 ( .A1(n6395), .A2(n3935), .ZN(n6530) );
  OR2_X1 U4054 ( .A1(n6568), .A2(n6811), .ZN(n6588) );
  NAND2_X1 U4055 ( .A1(n6640), .A2(n6589), .ZN(n6695) );
  INV_X1 U4056 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6798) );
  NAND2_X1 U4057 ( .A1(n6400), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3190) );
  INV_X2 U4058 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3204) );
  NAND2_X1 U4059 ( .A1(n3188), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3189) );
  NAND2_X1 U4060 ( .A1(n3190), .A2(n3189), .ZN(n3307) );
  NAND2_X1 U4061 ( .A1(n6704), .A2(n5197), .ZN(n3195) );
  NAND2_X1 U4062 ( .A1(n3191), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3192) );
  NAND2_X1 U4063 ( .A1(n3195), .A2(n3192), .ZN(n3301) );
  INV_X1 U4064 ( .A(n3301), .ZN(n3193) );
  XNOR2_X1 U4065 ( .A(n3903), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3298)
         );
  INV_X1 U4066 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5831) );
  AOI222_X1 U4067 ( .A1(n3294), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B1(
        n3294), .B2(n5831), .C1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n5831), 
        .ZN(n3443) );
  AND2_X4 U4068 ( .A1(n3204), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3219)
         );
  NAND2_X2 U4069 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3205) );
  INV_X2 U4070 ( .A(n3205), .ZN(n3917) );
  AND2_X4 U4071 ( .A1(n3219), .A2(n3917), .ZN(n3598) );
  NAND2_X1 U4072 ( .A1(n3598), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3203)
         );
  AND2_X4 U4073 ( .A1(n3198), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3218)
         );
  INV_X1 U4074 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3196) );
  NAND2_X1 U4075 ( .A1(n3597), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3202)
         );
  NOR2_X4 U4076 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3920) );
  NAND2_X1 U4077 ( .A1(n3555), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3201) );
  INV_X2 U4078 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3198) );
  AND2_X4 U4079 ( .A1(n3199), .A2(n3198), .ZN(n3894) );
  AND2_X2 U4080 ( .A1(n3894), .A2(n3920), .ZN(n3407) );
  NAND2_X1 U4081 ( .A1(n3407), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3200) );
  NOR2_X2 U4082 ( .A1(n3205), .A2(n3204), .ZN(n3899) );
  NAND2_X2 U4083 ( .A1(n3899), .A2(n3668), .ZN(n3528) );
  INV_X1 U4084 ( .A(n3528), .ZN(n3206) );
  NAND2_X1 U4086 ( .A1(n3770), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3209)
         );
  AND2_X2 U4087 ( .A1(n3917), .A2(n3920), .ZN(n3419) );
  NAND2_X1 U4088 ( .A1(n3419), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3207)
         );
  NAND2_X1 U4090 ( .A1(n3149), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3216) );
  NAND2_X1 U4091 ( .A1(n5068), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3215) );
  AND2_X2 U4092 ( .A1(n3217), .A2(n5669), .ZN(n3600) );
  NAND2_X1 U4093 ( .A1(n3600), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3214) );
  AND2_X2 U4094 ( .A1(n3217), .A2(n3220), .ZN(n3539) );
  NAND2_X1 U4095 ( .A1(n3539), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3224) );
  AND2_X4 U4096 ( .A1(n3219), .A2(n3218), .ZN(n5051) );
  NAND2_X1 U4097 ( .A1(n5051), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3223) );
  AND2_X4 U4098 ( .A1(n3894), .A2(n3219), .ZN(n3412) );
  NAND2_X1 U4099 ( .A1(n3412), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3222) );
  NAND3_X2 U4101 ( .A1(n3187), .A2(n3178), .A3(n3225), .ZN(n3629) );
  INV_X1 U4102 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3226) );
  OR2_X1 U4103 ( .A1(n3528), .A2(n3226), .ZN(n3230) );
  NAND2_X1 U4104 ( .A1(n3597), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3229)
         );
  NAND2_X1 U4105 ( .A1(n3539), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3228) );
  NAND2_X1 U4106 ( .A1(n3407), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3227) );
  NAND2_X1 U4108 ( .A1(n3600), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3234) );
  NAND2_X1 U4109 ( .A1(n3598), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3233)
         );
  NAND2_X1 U4110 ( .A1(n3412), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3232) );
  NAND2_X1 U4111 ( .A1(n3419), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3231)
         );
  AND2_X2 U4113 ( .A1(n3236), .A2(n3235), .ZN(n3247) );
  NAND2_X1 U4114 ( .A1(n3776), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3240) );
  NAND2_X1 U4115 ( .A1(n5068), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3239) );
  NAND2_X1 U4116 ( .A1(n3770), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3238)
         );
  INV_X2 U4117 ( .A(n4947), .ZN(n3771) );
  NAND2_X1 U4118 ( .A1(n3771), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3237) );
  AND4_X2 U4119 ( .A1(n3240), .A2(n3239), .A3(n3238), .A4(n3237), .ZN(n3246)
         );
  NAND2_X1 U4120 ( .A1(n5051), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3244) );
  NAND2_X1 U4121 ( .A1(n3555), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3243) );
  NAND2_X1 U4122 ( .A1(n5087), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3242) );
  NAND2_X1 U4123 ( .A1(n3591), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3241)
         );
  AND3_X4 U4124 ( .A1(n3247), .A2(n3246), .A3(n3245), .ZN(n3361) );
  NAND2_X1 U4125 ( .A1(n3407), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3250) );
  NAND2_X1 U4126 ( .A1(n5068), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3249) );
  NAND2_X1 U4127 ( .A1(n3597), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3248)
         );
  NAND3_X1 U4128 ( .A1(n3250), .A2(n3249), .A3(n3248), .ZN(n3251) );
  INV_X1 U4129 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3253) );
  INV_X1 U4130 ( .A(n4947), .ZN(n3254) );
  NAND2_X1 U4131 ( .A1(n3600), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3256) );
  NAND2_X1 U4132 ( .A1(n5087), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3255) );
  NAND2_X1 U4133 ( .A1(n3776), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3262) );
  NAND2_X1 U4134 ( .A1(n3555), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3261) );
  NAND2_X1 U4135 ( .A1(n3770), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3260)
         );
  NAND2_X1 U4136 ( .A1(n3419), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3259)
         );
  NAND2_X1 U4137 ( .A1(n3598), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3266)
         );
  NAND2_X1 U4138 ( .A1(n3539), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3265) );
  NAND2_X1 U4139 ( .A1(n3412), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3264) );
  NAND2_X1 U4140 ( .A1(n3591), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3263)
         );
  NAND2_X1 U4141 ( .A1(n3600), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3274) );
  NAND2_X1 U4142 ( .A1(n3598), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3273)
         );
  NAND2_X1 U4143 ( .A1(n3412), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3272) );
  NAND2_X1 U4144 ( .A1(n3419), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3271)
         );
  NAND2_X1 U4145 ( .A1(n5051), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3278) );
  NAND2_X1 U4146 ( .A1(n3776), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3277) );
  NAND2_X1 U4147 ( .A1(n3555), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3276) );
  NAND2_X1 U4148 ( .A1(n5087), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3275) );
  NAND2_X1 U4149 ( .A1(n3597), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3282)
         );
  NAND2_X1 U4150 ( .A1(n3539), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3281) );
  NAND2_X1 U4151 ( .A1(n3407), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3280) );
  NAND2_X1 U4152 ( .A1(n3591), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3279)
         );
  NAND2_X1 U4153 ( .A1(n5068), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3287) );
  NAND2_X1 U4154 ( .A1(n3770), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3286)
         );
  INV_X1 U4155 ( .A(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3284) );
  OR2_X2 U4156 ( .A1(n4947), .A2(n3284), .ZN(n3285) );
  NAND4_X4 U4157 ( .A1(n3292), .A2(n3291), .A3(n3290), .A4(n3289), .ZN(n3501)
         );
  NAND2_X1 U4158 ( .A1(n4773), .A2(n4086), .ZN(n4283) );
  NOR2_X1 U4159 ( .A1(n4263), .A2(n4283), .ZN(n3311) );
  NAND2_X1 U4160 ( .A1(n3443), .A2(n3311), .ZN(n3338) );
  AND2_X1 U4161 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n3294), .ZN(n3295)
         );
  INV_X1 U4162 ( .A(n3445), .ZN(n3300) );
  AOI22_X1 U4163 ( .A1(n3311), .A2(n3300), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6828), .ZN(n3334) );
  NAND2_X1 U4164 ( .A1(n3302), .A2(n3301), .ZN(n3304) );
  NAND2_X1 U4165 ( .A1(n3304), .A2(n3303), .ZN(n3441) );
  INV_X2 U4166 ( .A(n3629), .ZN(n3723) );
  INV_X2 U4167 ( .A(n3501), .ZN(n3452) );
  NAND2_X1 U4168 ( .A1(n3452), .A2(n4773), .ZN(n3306) );
  AOI21_X1 U4169 ( .B1(n3997), .B2(n3441), .A(n3327), .ZN(n3331) );
  AOI21_X1 U4170 ( .B1(n4261), .B2(n4086), .A(n3573), .ZN(n3312) );
  NAND2_X1 U4171 ( .A1(n3307), .A2(n3313), .ZN(n3308) );
  NAND2_X1 U4172 ( .A1(n3309), .A2(n3308), .ZN(n3442) );
  NOR3_X1 U4173 ( .A1(n3312), .A2(n3442), .A3(n6828), .ZN(n3310) );
  NOR2_X1 U4174 ( .A1(n3311), .A2(n3310), .ZN(n3325) );
  INV_X1 U4175 ( .A(n3442), .ZN(n3320) );
  INV_X1 U4176 ( .A(n3312), .ZN(n3322) );
  INV_X1 U4177 ( .A(n4261), .ZN(n3314) );
  OAI21_X1 U4178 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6819), .A(n3313), 
        .ZN(n3315) );
  NOR2_X1 U4179 ( .A1(n3314), .A2(n3315), .ZN(n3319) );
  NAND2_X1 U4180 ( .A1(n3361), .A2(n4773), .ZN(n3497) );
  INV_X1 U4181 ( .A(n3497), .ZN(n3316) );
  OAI21_X1 U4182 ( .B1(n3316), .B2(n3315), .A(n4385), .ZN(n3317) );
  NAND2_X1 U4183 ( .A1(n3318), .A2(n3317), .ZN(n3321) );
  OAI211_X1 U4184 ( .C1(n3320), .C2(n3322), .A(n3319), .B(n3321), .ZN(n3324)
         );
  NOR3_X1 U4185 ( .A1(n3322), .A2(n3321), .A3(n3442), .ZN(n3323) );
  AOI21_X1 U4186 ( .B1(n3325), .B2(n3324), .A(n3323), .ZN(n3328) );
  INV_X1 U4187 ( .A(n3328), .ZN(n3330) );
  INV_X1 U4188 ( .A(n3441), .ZN(n3326) );
  OAI211_X1 U4189 ( .C1(n3328), .C2(n3327), .A(n4261), .B(n3326), .ZN(n3329)
         );
  OAI21_X1 U4190 ( .B1(n3331), .B2(n3330), .A(n3329), .ZN(n3332) );
  OAI21_X1 U4191 ( .B1(n3997), .B2(n3445), .A(n3332), .ZN(n3333) );
  NAND2_X1 U4192 ( .A1(n3334), .A2(n3333), .ZN(n3335) );
  AOI21_X1 U4193 ( .B1(n4261), .B2(n3443), .A(n3335), .ZN(n3336) );
  INV_X1 U4194 ( .A(n3336), .ZN(n3337) );
  NAND2_X1 U4195 ( .A1(n6728), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3812) );
  OR2_X1 U4196 ( .A1(n3812), .A2(n6828), .ZN(n6736) );
  INV_X1 U4197 ( .A(n6736), .ZN(n6738) );
  INV_X1 U4198 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3339) );
  OR2_X1 U4199 ( .A1(n3528), .A2(n3339), .ZN(n3344) );
  NAND2_X1 U4200 ( .A1(n5068), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3343) );
  NAND2_X1 U4201 ( .A1(n3770), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3342)
         );
  INV_X1 U4202 ( .A(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3340) );
  NAND2_X1 U4203 ( .A1(n5051), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3348) );
  NAND2_X1 U4204 ( .A1(n3149), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3347) );
  NAND2_X1 U4205 ( .A1(n3555), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3346) );
  NAND2_X1 U4206 ( .A1(n5087), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3345) );
  NAND2_X1 U4207 ( .A1(n3598), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3352)
         );
  NAND2_X1 U4208 ( .A1(n3600), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3351) );
  NAND2_X1 U4209 ( .A1(n3412), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3350) );
  NAND2_X1 U4210 ( .A1(n3419), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3349)
         );
  NAND2_X1 U4211 ( .A1(n3591), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3356)
         );
  NAND2_X1 U4212 ( .A1(n3539), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3355) );
  NAND2_X1 U4213 ( .A1(n3407), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3354) );
  NAND2_X1 U4214 ( .A1(n3597), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3353)
         );
  INV_X1 U4216 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3362) );
  OR2_X1 U4217 ( .A1(n3528), .A2(n3362), .ZN(n3366) );
  NAND2_X1 U4218 ( .A1(n5068), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3365) );
  NAND2_X1 U4219 ( .A1(n3770), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3364)
         );
  NAND2_X1 U4220 ( .A1(n3771), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3363) );
  NAND2_X1 U4221 ( .A1(n5051), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3370) );
  NAND2_X1 U4222 ( .A1(n3776), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3369) );
  NAND2_X1 U4223 ( .A1(n3555), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3368) );
  NAND2_X1 U4224 ( .A1(n5087), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3367) );
  NAND2_X1 U4225 ( .A1(n3600), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3374) );
  NAND2_X1 U4226 ( .A1(n3598), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3373)
         );
  NAND2_X1 U4227 ( .A1(n3412), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3372) );
  NAND2_X1 U4228 ( .A1(n3419), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3371)
         );
  NAND2_X1 U4229 ( .A1(n3597), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3378)
         );
  NAND2_X1 U4230 ( .A1(n3539), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3377) );
  NAND2_X1 U4231 ( .A1(n3407), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3376) );
  NAND2_X1 U4232 ( .A1(n3591), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3375)
         );
  NAND2_X1 U4233 ( .A1(n3412), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3386) );
  NAND2_X1 U4234 ( .A1(n5051), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3385) );
  NAND2_X1 U4235 ( .A1(n5068), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3384) );
  NAND2_X1 U4236 ( .A1(n3407), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3383) );
  NAND2_X1 U4237 ( .A1(n3539), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3389) );
  NAND2_X1 U4238 ( .A1(n3591), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3388)
         );
  NAND2_X1 U4239 ( .A1(n3597), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3387)
         );
  NAND3_X1 U4240 ( .A1(n3389), .A2(n3388), .A3(n3387), .ZN(n3390) );
  NAND2_X1 U4241 ( .A1(n3776), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3394) );
  NAND2_X1 U4242 ( .A1(n3600), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3393) );
  NAND2_X1 U4243 ( .A1(n3419), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3391)
         );
  INV_X1 U4244 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3395) );
  OR2_X1 U4245 ( .A1(n3528), .A2(n3395), .ZN(n3399) );
  NAND2_X1 U4246 ( .A1(n3555), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3398) );
  NAND2_X1 U4247 ( .A1(n3770), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3397)
         );
  NAND2_X1 U4248 ( .A1(n3771), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3396) );
  NAND2_X1 U4249 ( .A1(n3539), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3406) );
  NAND2_X1 U4250 ( .A1(n3776), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3405) );
  NAND2_X1 U4251 ( .A1(n3600), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3404) );
  NAND2_X1 U4252 ( .A1(n3591), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3403)
         );
  NAND2_X1 U4253 ( .A1(n3598), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3411)
         );
  NAND2_X1 U4254 ( .A1(n5051), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3410) );
  NAND2_X1 U4255 ( .A1(n3555), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3409) );
  NAND2_X1 U4256 ( .A1(n3407), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3408) );
  NAND2_X1 U4257 ( .A1(n5068), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3417) );
  NAND2_X1 U4258 ( .A1(n3597), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3416)
         );
  NAND2_X1 U4259 ( .A1(n3412), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3415) );
  INV_X1 U4260 ( .A(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3413) );
  INV_X1 U4261 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3418) );
  OR2_X1 U4262 ( .A1(n3528), .A2(n3418), .ZN(n3423) );
  NAND2_X1 U4263 ( .A1(n3770), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3422)
         );
  NAND2_X1 U4264 ( .A1(n5087), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3421) );
  NAND2_X1 U4265 ( .A1(n3419), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3420)
         );
  NAND4_X4 U4266 ( .A1(n3427), .A2(n3426), .A3(n3425), .A4(n3424), .ZN(n4081)
         );
  NAND2_X2 U4267 ( .A1(n3571), .A2(n4081), .ZN(n3502) );
  NOR2_X2 U4268 ( .A1(n3502), .A2(n4773), .ZN(n3643) );
  NAND2_X2 U4270 ( .A1(n3470), .A2(n3428), .ZN(n3577) );
  OR2_X1 U4271 ( .A1(n6062), .A2(n4086), .ZN(n6064) );
  NAND2_X1 U4272 ( .A1(n3430), .A2(n4773), .ZN(n3435) );
  BUF_X1 U4273 ( .A(n3431), .Z(n3433) );
  NAND2_X2 U4274 ( .A1(n3433), .A2(n3432), .ZN(n3459) );
  OAI21_X1 U4276 ( .B1(n3435), .B2(n4108), .A(n3434), .ZN(n3436) );
  INV_X1 U4277 ( .A(n3436), .ZN(n3568) );
  NAND2_X1 U4278 ( .A1(n3438), .A2(n3469), .ZN(n3465) );
  NOR2_X1 U4279 ( .A1(n3465), .A2(n4385), .ZN(n3569) );
  AND2_X1 U4280 ( .A1(n3568), .A2(n3569), .ZN(n3651) );
  NAND2_X1 U4281 ( .A1(n3651), .A2(n4086), .ZN(n5666) );
  OR2_X1 U4282 ( .A1(n4152), .A2(n5666), .ZN(n3439) );
  NAND2_X1 U4283 ( .A1(n6064), .A2(n3439), .ZN(n3440) );
  NAND2_X1 U4284 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6749) );
  OAI21_X1 U4285 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .A(
        n6749), .ZN(n3499) );
  OR2_X1 U4286 ( .A1(n3499), .A2(STATE_REG_0__SCAN_IN), .ZN(n6755) );
  INV_X1 U4287 ( .A(n6755), .ZN(n4380) );
  NOR2_X1 U4288 ( .A1(n6728), .A2(n6637), .ZN(n3890) );
  INV_X1 U4289 ( .A(n3890), .ZN(n6723) );
  OR2_X1 U4290 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6723), .ZN(n6832) );
  INV_X1 U4291 ( .A(n6832), .ZN(n4063) );
  AND2_X1 U4292 ( .A1(n6058), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  OR2_X1 U4293 ( .A1(n3735), .A2(n3574), .ZN(n3448) );
  NOR2_X1 U4294 ( .A1(n3442), .A2(n3441), .ZN(n3444) );
  AOI21_X1 U4295 ( .B1(n3445), .B2(n3444), .A(n3443), .ZN(n3658) );
  AND2_X1 U4296 ( .A1(n3658), .A2(n3651), .ZN(n3486) );
  INV_X1 U4297 ( .A(n3486), .ZN(n3446) );
  NAND2_X1 U4298 ( .A1(n3446), .A2(n3577), .ZN(n3447) );
  AND2_X1 U4299 ( .A1(n3448), .A2(n3447), .ZN(n3454) );
  AND2_X1 U4300 ( .A1(n3454), .A2(n6738), .ZN(n3451) );
  INV_X1 U4301 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n3450) );
  NOR2_X2 U4302 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6812) );
  AND2_X1 U4303 ( .A1(n6812), .A2(n6728), .ZN(n3487) );
  NAND2_X1 U4304 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n3487), .ZN(n3449) );
  OAI21_X1 U4305 ( .B1(n3451), .B2(n3450), .A(n3449), .ZN(U2790) );
  AND2_X1 U4306 ( .A1(n3723), .A2(n4086), .ZN(n4373) );
  OR2_X1 U4307 ( .A1(n5239), .A2(n4373), .ZN(n3495) );
  NAND2_X1 U4308 ( .A1(n3495), .A2(n6755), .ZN(n6826) );
  INV_X1 U4309 ( .A(READY_N), .ZN(n7199) );
  NAND2_X1 U4310 ( .A1(n6826), .A2(n7199), .ZN(n3453) );
  AND2_X1 U4311 ( .A1(n3454), .A2(n3453), .ZN(n6716) );
  NOR2_X1 U4312 ( .A1(n6716), .A2(n6736), .ZN(n5836) );
  INV_X1 U4313 ( .A(MORE_REG_SCAN_IN), .ZN(n7029) );
  INV_X1 U4314 ( .A(n3651), .ZN(n3484) );
  AND2_X1 U4315 ( .A1(n3455), .A2(n3460), .ZN(n3456) );
  OAI21_X1 U4316 ( .B1(n3459), .B2(n3457), .A(n3456), .ZN(n3458) );
  BUF_X2 U4317 ( .A(n3459), .Z(n4156) );
  NAND2_X1 U4318 ( .A1(n4091), .A2(n4155), .ZN(n3461) );
  OR2_X1 U4319 ( .A1(n4156), .A2(n3461), .ZN(n4695) );
  AOI21_X1 U4320 ( .B1(n4695), .B2(n3723), .A(n3502), .ZN(n3462) );
  NAND2_X1 U4321 ( .A1(n3512), .A2(n3462), .ZN(n3650) );
  NOR2_X1 U4322 ( .A1(n3650), .A2(n3305), .ZN(n3892) );
  NOR2_X1 U4323 ( .A1(n3650), .A2(n3497), .ZN(n3734) );
  OR2_X1 U4324 ( .A1(n3892), .A2(n3734), .ZN(n3719) );
  INV_X1 U4325 ( .A(n3577), .ZN(n3463) );
  NOR2_X1 U4326 ( .A1(n3719), .A2(n3463), .ZN(n3464) );
  OR2_X1 U4327 ( .A1(n3735), .A2(n3464), .ZN(n3483) );
  AOI21_X1 U4328 ( .B1(n3465), .B2(n4108), .A(n4086), .ZN(n3466) );
  NAND2_X1 U4329 ( .A1(n3568), .A2(n3466), .ZN(n3467) );
  NAND2_X1 U4330 ( .A1(n3467), .A2(n3723), .ZN(n3506) );
  NOR2_X1 U4331 ( .A1(n4283), .A2(n4091), .ZN(n3468) );
  OR2_X1 U4332 ( .A1(n3506), .A2(n3468), .ZN(n3519) );
  INV_X1 U4333 ( .A(n4156), .ZN(n3471) );
  OR3_X1 U4334 ( .A1(n3470), .A2(n3723), .A3(n3471), .ZN(n3474) );
  AND2_X1 U4335 ( .A1(n4373), .A2(n3691), .ZN(n3654) );
  NAND2_X1 U4336 ( .A1(n3572), .A2(n4385), .ZN(n4249) );
  INV_X1 U4337 ( .A(n4249), .ZN(n3472) );
  OAI21_X1 U4338 ( .B1(n3654), .B2(n5234), .A(n3502), .ZN(n3473) );
  OAI211_X1 U4339 ( .C1(n3691), .C2(n4772), .A(n3474), .B(n3473), .ZN(n3648)
         );
  INV_X1 U4340 ( .A(n3510), .ZN(n3745) );
  NAND2_X1 U4341 ( .A1(n4385), .A2(n4108), .ZN(n3476) );
  NAND2_X1 U4342 ( .A1(n3477), .A2(n3476), .ZN(n3649) );
  INV_X1 U4343 ( .A(n3649), .ZN(n3478) );
  OAI21_X1 U4344 ( .B1(n3512), .B2(n3174), .A(n3478), .ZN(n3480) );
  NOR2_X1 U4345 ( .A1(n3648), .A2(n3480), .ZN(n3481) );
  AND2_X1 U4346 ( .A1(n3519), .A2(n3481), .ZN(n3710) );
  NOR2_X1 U4347 ( .A1(n4695), .A2(n3452), .ZN(n3683) );
  NAND2_X1 U4348 ( .A1(n3735), .A2(n3893), .ZN(n3482) );
  OAI211_X1 U4349 ( .C1(n3658), .C2(n3484), .A(n3483), .B(n3482), .ZN(n6713)
         );
  NAND2_X1 U4350 ( .A1(n5836), .A2(n6713), .ZN(n3485) );
  OAI21_X1 U4351 ( .B1(n5836), .B2(n7029), .A(n3485), .ZN(U3471) );
  NAND2_X1 U4352 ( .A1(n3486), .A2(n6738), .ZN(n3494) );
  INV_X1 U4353 ( .A(n3494), .ZN(n3490) );
  INV_X1 U4354 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n7062) );
  INV_X1 U4355 ( .A(n3487), .ZN(n3488) );
  NAND2_X1 U4356 ( .A1(n6062), .A2(n3488), .ZN(n3491) );
  INV_X1 U4357 ( .A(n3491), .ZN(n3489) );
  OAI21_X1 U4358 ( .B1(n3490), .B2(n7062), .A(n3489), .ZN(U2788) );
  INV_X1 U4359 ( .A(n3495), .ZN(n3492) );
  OAI22_X1 U4360 ( .A1(n6830), .A2(n3492), .B1(n3491), .B2(
        READREQUEST_REG_SCAN_IN), .ZN(n3493) );
  OAI21_X1 U4361 ( .B1(n3495), .B2(n3494), .A(n3493), .ZN(U3474) );
  NAND2_X1 U4362 ( .A1(n3496), .A2(n3510), .ZN(n3498) );
  OR2_X2 U4363 ( .A1(n3497), .A2(n3634), .ZN(n3705) );
  INV_X1 U4364 ( .A(n3499), .ZN(n3500) );
  INV_X1 U4365 ( .A(n3575), .ZN(n3503) );
  NAND2_X1 U4366 ( .A1(n4156), .A2(n4091), .ZN(n3513) );
  NAND3_X1 U4367 ( .A1(n3512), .A2(n3504), .A3(n3513), .ZN(n3505) );
  NOR2_X1 U4368 ( .A1(n3515), .A2(n3505), .ZN(n3507) );
  NAND2_X1 U4369 ( .A1(n3507), .A2(n3506), .ZN(n3508) );
  NAND2_X1 U4370 ( .A1(n6798), .A2(n6728), .ZN(n5677) );
  MUX2_X1 U4371 ( .A(n3812), .B(n3813), .S(n6819), .Z(n3609) );
  INV_X1 U4372 ( .A(n3609), .ZN(n3509) );
  OAI21_X2 U4373 ( .B1(n3157), .B2(n3668), .A(n3509), .ZN(n3521) );
  NAND3_X1 U4374 ( .A1(n3572), .A2(n3691), .A3(n3723), .ZN(n3703) );
  NOR2_X1 U4375 ( .A1(n5677), .A2(n6828), .ZN(n6739) );
  OAI211_X1 U4376 ( .C1(n3703), .C2(n3469), .A(n6739), .B(n5157), .ZN(n3511)
         );
  NOR2_X1 U4377 ( .A1(n3511), .A2(n3649), .ZN(n3520) );
  NAND2_X1 U4378 ( .A1(n3513), .A2(n4081), .ZN(n3514) );
  OAI21_X1 U4379 ( .B1(n3458), .B2(n3514), .A(n4086), .ZN(n3517) );
  INV_X1 U4380 ( .A(n3515), .ZN(n3516) );
  NAND3_X1 U4381 ( .A1(n3520), .A2(n3519), .A3(n3518), .ZN(n3522) );
  NAND2_X1 U4382 ( .A1(n3521), .A2(n3522), .ZN(n3756) );
  OAI21_X1 U4383 ( .B1(n3521), .B2(n3522), .A(n3756), .ZN(n6430) );
  OR2_X1 U4384 ( .A1(n6430), .A2(n4599), .ZN(n3527) );
  AND2_X1 U4385 ( .A1(n4772), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3986) );
  INV_X1 U4386 ( .A(EAX_REG_0__SCAN_IN), .ZN(n3524) );
  INV_X1 U4387 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n3523) );
  OAI22_X1 U4388 ( .A1(n5008), .A2(n3524), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3523), .ZN(n3525) );
  AOI21_X1 U4389 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n3986), .A(n3525), 
        .ZN(n3526) );
  NAND2_X1 U4390 ( .A1(n3527), .A2(n3526), .ZN(n3860) );
  NAND2_X1 U4391 ( .A1(n6637), .A2(n6912), .ZN(n5101) );
  INV_X1 U4392 ( .A(n3528), .ZN(n5074) );
  INV_X1 U4393 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3529) );
  OR2_X1 U4394 ( .A1(n5018), .A2(n3529), .ZN(n3533) );
  NAND2_X1 U4395 ( .A1(n5050), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3532) );
  NAND2_X1 U4396 ( .A1(n3770), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3531)
         );
  NAND2_X1 U4397 ( .A1(n5069), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3530) );
  AOI22_X1 U4398 ( .A1(n5051), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3555), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3536) );
  AOI22_X1 U4399 ( .A1(n3776), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4882), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3535) );
  NAND3_X1 U4400 ( .A1(n3537), .A2(n3536), .A3(n3535), .ZN(n3546) );
  BUF_X2 U4401 ( .A(n3412), .Z(n5076) );
  AOI22_X1 U4402 ( .A1(n5076), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3544) );
  INV_X1 U4403 ( .A(n3419), .ZN(n4949) );
  INV_X1 U4404 ( .A(n4949), .ZN(n3547) );
  AOI22_X1 U4405 ( .A1(n3600), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3543) );
  AOI22_X1 U4408 ( .A1(n3538), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3599), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3542) );
  INV_X1 U4409 ( .A(n3591), .ZN(n3540) );
  AOI22_X1 U4410 ( .A1(n5081), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3541) );
  NAND4_X1 U4411 ( .A1(n3544), .A2(n3543), .A3(n3542), .A4(n3541), .ZN(n3545)
         );
  OR2_X2 U4412 ( .A1(n3546), .A2(n3545), .ZN(n4298) );
  NAND2_X1 U4413 ( .A1(n3717), .A2(n4298), .ZN(n3612) );
  INV_X1 U4414 ( .A(n3612), .ZN(n3563) );
  NOR2_X1 U4415 ( .A1(n4298), .A2(n4091), .ZN(n3562) );
  AOI22_X1 U4416 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n3149), .B1(n3538), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3554) );
  AOI22_X1 U4417 ( .A1(n5051), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3553) );
  NAND2_X1 U4418 ( .A1(n4882), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3550) );
  NAND2_X1 U4419 ( .A1(n3547), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3549)
         );
  NAND2_X1 U4420 ( .A1(n5069), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3548) );
  AND3_X1 U4421 ( .A1(n3550), .A2(n3549), .A3(n3548), .ZN(n3552) );
  INV_X1 U4422 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4897) );
  OR2_X1 U4423 ( .A1(n5018), .A2(n4897), .ZN(n3551) );
  NAND4_X1 U4424 ( .A1(n3554), .A2(n3553), .A3(n3552), .A4(n3551), .ZN(n3561)
         );
  AOI22_X1 U4425 ( .A1(n5081), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3559) );
  AOI22_X1 U4426 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n5050), .B1(n3555), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3558) );
  AOI22_X1 U4427 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n3600), .B1(n5083), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3557) );
  AOI22_X1 U4428 ( .A1(n3599), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3556) );
  NAND4_X1 U4429 ( .A1(n3559), .A2(n3558), .A3(n3557), .A4(n3556), .ZN(n3560)
         );
  MUX2_X1 U4430 ( .A(n3563), .B(n3562), .S(n3742), .Z(n3564) );
  INV_X1 U4431 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4896) );
  AOI21_X1 U4432 ( .B1(n3723), .B2(n3742), .A(n6828), .ZN(n3565) );
  OAI211_X1 U4433 ( .C1(n4263), .C2(n4896), .A(n3565), .B(n3612), .ZN(n3613)
         );
  OAI211_X1 U4434 ( .C1(n3609), .C2(STATE2_REG_0__SCAN_IN), .A(n3611), .B(
        n3613), .ZN(n3566) );
  OR2_X1 U4435 ( .A1(n6811), .A2(n3469), .ZN(n3567) );
  AND2_X1 U4436 ( .A1(n3567), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3861) );
  NAND2_X1 U4437 ( .A1(n3860), .A2(n3861), .ZN(n3864) );
  OAI21_X1 U4438 ( .B1(n3860), .B2(n5101), .A(n3864), .ZN(n3627) );
  NAND3_X1 U4439 ( .A1(n3569), .A2(n3568), .A3(n3452), .ZN(n3657) );
  INV_X1 U4440 ( .A(n3570), .ZN(n3574) );
  NAND2_X1 U4442 ( .A1(n3657), .A2(n3716), .ZN(n3579) );
  NOR2_X2 U4443 ( .A1(n3577), .A2(n3576), .ZN(n3578) );
  OAI21_X2 U4444 ( .B1(n3579), .B2(n3578), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n3585) );
  INV_X1 U4445 ( .A(n3585), .ZN(n3583) );
  NAND2_X1 U4446 ( .A1(n6819), .A2(n6400), .ZN(n3580) );
  NAND2_X1 U4447 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3762) );
  AND2_X1 U4448 ( .A1(n3580), .A2(n3762), .ZN(n6480) );
  AND2_X1 U4449 ( .A1(n3812), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3581)
         );
  AOI21_X1 U4450 ( .B1(n3813), .B2(n6480), .A(n3581), .ZN(n3584) );
  INV_X1 U4451 ( .A(n3584), .ZN(n3582) );
  NAND2_X1 U4452 ( .A1(n3586), .A2(n3758), .ZN(n3755) );
  XNOR2_X1 U4453 ( .A(n3755), .B(n3756), .ZN(n3939) );
  INV_X1 U4454 ( .A(n3786), .ZN(n3607) );
  NAND2_X1 U4455 ( .A1(n3534), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3589) );
  NAND2_X1 U4456 ( .A1(n5076), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3588) );
  NAND2_X1 U4457 ( .A1(n5083), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3587)
         );
  AND3_X1 U4458 ( .A1(n3589), .A2(n3588), .A3(n3587), .ZN(n3596) );
  INV_X1 U4459 ( .A(n5068), .ZN(n3590) );
  INV_X2 U4460 ( .A(n3590), .ZN(n5050) );
  AOI22_X1 U4461 ( .A1(n5050), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4882), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3595) );
  AOI22_X1 U4462 ( .A1(n5075), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3594) );
  INV_X1 U4463 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3592) );
  OR2_X1 U4464 ( .A1(n5018), .A2(n3592), .ZN(n3593) );
  NAND4_X1 U4465 ( .A1(n3596), .A2(n3595), .A3(n3594), .A4(n3593), .ZN(n3606)
         );
  BUF_X1 U4466 ( .A(n3597), .Z(n5026) );
  AOI22_X1 U4467 ( .A1(n5026), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3604) );
  AOI22_X1 U4469 ( .A1(n5051), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5069), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3603) );
  AOI22_X1 U4470 ( .A1(n5081), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3599), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3602) );
  AOI22_X1 U4471 ( .A1(n5070), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3601) );
  NAND4_X1 U4472 ( .A1(n3604), .A2(n3603), .A3(n3602), .A4(n3601), .ZN(n3605)
         );
  NAND2_X1 U4473 ( .A1(n3607), .A2(n3743), .ZN(n3608) );
  OR2_X1 U4474 ( .A1(n3609), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3610) );
  NAND2_X1 U4475 ( .A1(n3611), .A2(n3610), .ZN(n3614) );
  XNOR2_X1 U4476 ( .A(n3168), .B(n3793), .ZN(n3792) );
  NAND2_X1 U4477 ( .A1(n3997), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3619) );
  INV_X1 U4478 ( .A(n3743), .ZN(n3616) );
  NOR2_X1 U4479 ( .A1(n4385), .A2(n6828), .ZN(n3788) );
  INV_X1 U4480 ( .A(n3788), .ZN(n3615) );
  OAI22_X1 U4481 ( .A1(n3616), .A2(n3615), .B1(n3786), .B2(n4298), .ZN(n3617)
         );
  INV_X1 U4482 ( .A(n3617), .ZN(n3618) );
  NAND2_X1 U4483 ( .A1(n3934), .A2(n4648), .ZN(n3624) );
  INV_X1 U4484 ( .A(EAX_REG_1__SCAN_IN), .ZN(n3621) );
  INV_X1 U4485 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3740) );
  OAI22_X1 U4486 ( .A1(n5008), .A2(n3621), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3740), .ZN(n3622) );
  AOI21_X1 U4487 ( .B1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n3986), .A(n3622), 
        .ZN(n3623) );
  NAND2_X1 U4488 ( .A1(n3624), .A2(n3623), .ZN(n3626) );
  INV_X1 U4489 ( .A(n3798), .ZN(n3625) );
  OAI21_X1 U4490 ( .B1(n3627), .B2(n3626), .A(n3625), .ZN(n4393) );
  NAND2_X1 U4491 ( .A1(n3893), .A2(n6738), .ZN(n3628) );
  OR2_X1 U4492 ( .A1(n3628), .A2(n3735), .ZN(n3633) );
  NAND4_X1 U4493 ( .A1(n3717), .A2(n5220), .A3(n6738), .A4(n3469), .ZN(n4154)
         );
  INV_X1 U4494 ( .A(n4154), .ZN(n3630) );
  NAND3_X1 U4495 ( .A1(n3631), .A2(n3630), .A3(n5178), .ZN(n3632) );
  NAND2_X2 U4496 ( .A1(n3633), .A2(n3632), .ZN(n6022) );
  NAND2_X1 U4497 ( .A1(n6022), .A2(n5220), .ZN(n6011) );
  OR2_X2 U4498 ( .A1(n3634), .A2(n3644), .ZN(n5227) );
  INV_X1 U4499 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3876) );
  NAND2_X1 U4500 ( .A1(n4249), .A2(n3876), .ZN(n3635) );
  OAI211_X1 U4501 ( .C1(n3644), .C2(EBX_REG_1__SCAN_IN), .A(n3635), .B(n3634), 
        .ZN(n3636) );
  NAND2_X1 U4502 ( .A1(n4249), .A2(EBX_REG_0__SCAN_IN), .ZN(n3638) );
  INV_X1 U4503 ( .A(EBX_REG_0__SCAN_IN), .ZN(n6001) );
  NAND2_X1 U4504 ( .A1(n3634), .A2(n6001), .ZN(n3637) );
  INV_X1 U4505 ( .A(n3701), .ZN(n3639) );
  XNOR2_X1 U4506 ( .A(n3844), .B(n3639), .ZN(n3640) );
  NOR2_X1 U4507 ( .A1(n3640), .A2(n5178), .ZN(n3641) );
  OR2_X1 U4508 ( .A1(n3846), .A2(n3641), .ZN(n6173) );
  INV_X1 U4509 ( .A(n6022), .ZN(n5371) );
  AOI22_X1 U4510 ( .A1(n6018), .A2(n6173), .B1(n5371), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n3642) );
  OAI21_X1 U4511 ( .B1(n4393), .B2(n6012), .A(n3642), .ZN(U2858) );
  NAND2_X1 U4512 ( .A1(n6828), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6796) );
  INV_X1 U4513 ( .A(n6796), .ZN(n4080) );
  INV_X1 U4514 ( .A(n3893), .ZN(n3702) );
  NOR2_X1 U4515 ( .A1(n3702), .A2(n3735), .ZN(n3662) );
  NAND2_X1 U4516 ( .A1(n3470), .A2(n3643), .ZN(n3697) );
  INV_X1 U4517 ( .A(n3697), .ZN(n3647) );
  INV_X1 U4518 ( .A(n5666), .ZN(n3646) );
  OR2_X1 U4519 ( .A1(n3697), .A2(n5168), .ZN(n4151) );
  AOI21_X1 U4520 ( .B1(n4151), .B2(n6755), .A(READY_N), .ZN(n3645) );
  OAI211_X1 U4521 ( .C1(n3647), .C2(n3646), .A(n3735), .B(n3645), .ZN(n3656)
         );
  INV_X1 U4522 ( .A(n3648), .ZN(n3653) );
  NOR2_X1 U4523 ( .A1(n3650), .A2(n3649), .ZN(n3652) );
  AOI21_X1 U4524 ( .B1(n3653), .B2(n3652), .A(n3651), .ZN(n3682) );
  NOR2_X1 U4525 ( .A1(n3682), .A2(n3654), .ZN(n3655) );
  NAND2_X1 U4526 ( .A1(n3656), .A2(n3655), .ZN(n3661) );
  NAND2_X1 U4527 ( .A1(n3735), .A2(n3892), .ZN(n3660) );
  NAND2_X1 U4528 ( .A1(n3658), .A2(n7199), .ZN(n3685) );
  OR2_X1 U4529 ( .A1(n5825), .A2(n3685), .ZN(n3659) );
  NAND2_X1 U4530 ( .A1(n3660), .A2(n3659), .ZN(n4150) );
  INV_X1 U4531 ( .A(n3925), .ZN(n6700) );
  INV_X1 U4532 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6712) );
  NOR2_X1 U4533 ( .A1(n6828), .A2(n6723), .ZN(n3930) );
  INV_X1 U4534 ( .A(n3930), .ZN(n6795) );
  OAI22_X1 U4535 ( .A1(n6700), .A2(n6736), .B1(n6712), .B2(n6795), .ZN(n5826)
         );
  NOR2_X1 U4536 ( .A1(n4080), .A2(n5826), .ZN(n5679) );
  INV_X1 U4537 ( .A(n5679), .ZN(n5832) );
  AND4_X1 U4538 ( .A1(n5825), .A2(n3705), .A3(n3697), .A4(n3663), .ZN(n3664)
         );
  AND2_X1 U4539 ( .A1(n3710), .A2(n3664), .ZN(n3914) );
  OAI22_X1 U4540 ( .A1(n6430), .A2(n3914), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n4695), .ZN(n6698) );
  AOI21_X1 U4541 ( .B1(n6698), .B2(n6798), .A(STATE2_REG_1__SCAN_IN), .ZN(
        n3665) );
  NAND2_X1 U4542 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5196) );
  INV_X1 U4543 ( .A(n5196), .ZN(n5672) );
  OAI22_X1 U4544 ( .A1(n3665), .A2(n5672), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6733), .ZN(n3666) );
  INV_X1 U4545 ( .A(n5677), .ZN(n5827) );
  NOR2_X1 U4546 ( .A1(n5666), .A2(n3668), .ZN(n6697) );
  AOI22_X1 U4547 ( .A1(n5832), .A2(n3666), .B1(n5827), .B2(n6697), .ZN(n3667)
         );
  OAI21_X1 U4548 ( .B1(n3668), .B2(n5832), .A(n3667), .ZN(U3461) );
  INV_X1 U4549 ( .A(EAX_REG_30__SCAN_IN), .ZN(n3670) );
  NAND2_X1 U4550 ( .A1(n6037), .A2(n4385), .ZN(n4072) );
  AOI22_X1 U4551 ( .A1(n4063), .A2(UWORD_REG_14__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n3669) );
  OAI21_X1 U4552 ( .B1(n3670), .B2(n4072), .A(n3669), .ZN(U2893) );
  INV_X1 U4553 ( .A(EAX_REG_28__SCAN_IN), .ZN(n3672) );
  AOI22_X1 U4554 ( .A1(n4063), .A2(UWORD_REG_12__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n3671) );
  OAI21_X1 U4555 ( .B1(n3672), .B2(n4072), .A(n3671), .ZN(U2895) );
  INV_X1 U4556 ( .A(EAX_REG_29__SCAN_IN), .ZN(n3674) );
  AOI22_X1 U4557 ( .A1(n4063), .A2(UWORD_REG_13__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n3673) );
  OAI21_X1 U4558 ( .B1(n3674), .B2(n4072), .A(n3673), .ZN(U2894) );
  AOI22_X1 U4559 ( .A1(n4063), .A2(UWORD_REG_10__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n3675) );
  OAI21_X1 U4560 ( .B1(n4985), .B2(n4072), .A(n3675), .ZN(U2897) );
  INV_X1 U4561 ( .A(EAX_REG_24__SCAN_IN), .ZN(n3677) );
  AOI22_X1 U4562 ( .A1(n4063), .A2(UWORD_REG_8__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n3676) );
  OAI21_X1 U4563 ( .B1(n3677), .B2(n4072), .A(n3676), .ZN(U2899) );
  INV_X1 U4564 ( .A(EAX_REG_25__SCAN_IN), .ZN(n3679) );
  AOI22_X1 U4565 ( .A1(n4063), .A2(UWORD_REG_9__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n3678) );
  OAI21_X1 U4566 ( .B1(n3679), .B2(n4072), .A(n3678), .ZN(U2898) );
  INV_X1 U4567 ( .A(EAX_REG_27__SCAN_IN), .ZN(n3681) );
  AOI22_X1 U4568 ( .A1(n4063), .A2(UWORD_REG_11__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n3680) );
  OAI21_X1 U4569 ( .B1(n3681), .B2(n4072), .A(n3680), .ZN(U2896) );
  INV_X1 U4570 ( .A(n3735), .ZN(n3684) );
  AOI21_X1 U4571 ( .B1(n3684), .B2(n3683), .A(n3682), .ZN(n3695) );
  NAND2_X1 U4572 ( .A1(n4086), .A2(n6755), .ZN(n3687) );
  INV_X1 U4573 ( .A(n3685), .ZN(n3686) );
  NAND2_X1 U4574 ( .A1(n3687), .A2(n3686), .ZN(n3693) );
  NOR2_X1 U4575 ( .A1(n4086), .A2(n4380), .ZN(n4387) );
  OR3_X1 U4576 ( .A1(n3697), .A2(n4387), .A3(READY_N), .ZN(n3689) );
  NOR2_X1 U4577 ( .A1(n4772), .A2(n3723), .ZN(n3688) );
  NAND2_X1 U4578 ( .A1(n3689), .A2(n3688), .ZN(n3690) );
  NAND2_X1 U4579 ( .A1(n3735), .A2(n3690), .ZN(n3692) );
  MUX2_X1 U4580 ( .A(n3693), .B(n3692), .S(n3691), .Z(n3694) );
  NAND2_X1 U4581 ( .A1(n3695), .A2(n3694), .ZN(n3696) );
  OR2_X1 U4582 ( .A1(n3697), .A2(n3745), .ZN(n6726) );
  OAI21_X1 U4583 ( .B1(n3716), .B2(n4091), .A(n6726), .ZN(n3698) );
  INV_X1 U4584 ( .A(n3698), .ZN(n3699) );
  NOR2_X1 U4585 ( .A1(n5234), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3700)
         );
  OR2_X1 U4586 ( .A1(n3701), .A2(n3700), .ZN(n5991) );
  INV_X1 U4587 ( .A(n4695), .ZN(n5664) );
  INV_X1 U4588 ( .A(n3703), .ZN(n3704) );
  NAND2_X1 U4589 ( .A1(n5664), .A2(n3704), .ZN(n3908) );
  INV_X1 U4590 ( .A(n3705), .ZN(n3706) );
  NAND2_X1 U4591 ( .A1(n3706), .A2(n3723), .ZN(n3707) );
  OAI211_X1 U4592 ( .C1(n3663), .C2(n3469), .A(n3908), .B(n3707), .ZN(n3708)
         );
  INV_X1 U4593 ( .A(n3708), .ZN(n3709) );
  AND2_X1 U4594 ( .A1(n3710), .A2(n3709), .ZN(n3711) );
  AND2_X1 U4595 ( .A1(n5645), .A2(n5649), .ZN(n5639) );
  INV_X1 U4596 ( .A(n5639), .ZN(n3715) );
  INV_X1 U4597 ( .A(n4048), .ZN(n5648) );
  INV_X1 U4598 ( .A(n5645), .ZN(n6161) );
  INV_X1 U4599 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3885) );
  OR2_X1 U4600 ( .A1(n5649), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3713)
         );
  AND2_X1 U4601 ( .A1(n3813), .A2(n6478), .ZN(n6176) );
  INV_X1 U4602 ( .A(n6176), .ZN(n5819) );
  NAND2_X1 U4603 ( .A1(n3722), .A2(n5819), .ZN(n3712) );
  NAND2_X1 U4604 ( .A1(n3713), .A2(n3712), .ZN(n5641) );
  AOI21_X1 U4605 ( .B1(n6161), .B2(n3885), .A(n5641), .ZN(n6178) );
  INV_X1 U4606 ( .A(n6178), .ZN(n3714) );
  OAI22_X1 U4607 ( .A1(n3715), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .B1(n5648), 
        .B2(n3714), .ZN(n3733) );
  OAI21_X1 U4608 ( .B1(n3717), .B2(n3716), .A(n4151), .ZN(n3718) );
  NOR2_X1 U4609 ( .A1(n3719), .A2(n3718), .ZN(n3720) );
  AND2_X1 U4610 ( .A1(n3720), .A2(n5825), .ZN(n3721) );
  INV_X1 U4611 ( .A(n4283), .ZN(n4296) );
  NAND2_X1 U4612 ( .A1(n6811), .A2(n4296), .ZN(n3727) );
  AND2_X1 U4613 ( .A1(n3723), .A2(n4081), .ZN(n3872) );
  INV_X1 U4614 ( .A(n3872), .ZN(n3724) );
  OAI21_X1 U4615 ( .B1(n3745), .B2(n3742), .A(n3724), .ZN(n3725) );
  INV_X1 U4616 ( .A(n3725), .ZN(n3726) );
  NAND2_X1 U4617 ( .A1(n3727), .A2(n3726), .ZN(n3728) );
  INV_X1 U4618 ( .A(n3728), .ZN(n3730) );
  NAND2_X1 U4619 ( .A1(n3728), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3877)
         );
  INV_X1 U4620 ( .A(n3877), .ZN(n3729) );
  AOI21_X1 U4621 ( .B1(n3730), .B2(n3885), .A(n3729), .ZN(n6114) );
  NAND2_X1 U4622 ( .A1(n6176), .A2(REIP_REG_0__SCAN_IN), .ZN(n6119) );
  INV_X1 U4623 ( .A(n6119), .ZN(n3731) );
  AOI21_X1 U4624 ( .B1(n6175), .B2(n6114), .A(n3731), .ZN(n3732) );
  OAI211_X1 U4625 ( .C1(n6163), .C2(n5991), .A(n3733), .B(n3732), .ZN(U3018)
         );
  AND2_X1 U4626 ( .A1(n6828), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4358) );
  NAND2_X1 U4627 ( .A1(n4358), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6745) );
  AND2_X1 U4628 ( .A1(n3735), .A2(n3734), .ZN(n6714) );
  NOR2_X1 U4629 ( .A1(n3813), .A2(n6812), .ZN(n6831) );
  NOR2_X1 U4630 ( .A1(n6831), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3736) );
  NAND2_X1 U4631 ( .A1(n6828), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3738) );
  NAND2_X1 U4632 ( .A1(n6912), .A2(STATE2_REG_1__SCAN_IN), .ZN(n3737) );
  NAND2_X1 U4633 ( .A1(n3738), .A2(n3737), .ZN(n6116) );
  INV_X1 U4634 ( .A(REIP_REG_1__SCAN_IN), .ZN(n3739) );
  OAI22_X1 U4635 ( .A1(n5786), .A2(n3740), .B1(n5819), .B2(n3739), .ZN(n3741)
         );
  AOI21_X1 U4636 ( .B1(n5781), .B2(n3740), .A(n3741), .ZN(n3754) );
  NAND2_X1 U4637 ( .A1(n3173), .A2(n4296), .ZN(n3749) );
  NAND2_X1 U4638 ( .A1(n3742), .A2(n3743), .ZN(n3871) );
  OAI21_X1 U4639 ( .B1(n3743), .B2(n3742), .A(n3871), .ZN(n3746) );
  INV_X1 U4640 ( .A(n3502), .ZN(n3744) );
  OAI211_X1 U4641 ( .C1(n3746), .C2(n3745), .A(n3744), .B(n4773), .ZN(n3747)
         );
  INV_X1 U4642 ( .A(n3747), .ZN(n3748) );
  NAND2_X1 U4643 ( .A1(n3749), .A2(n3748), .ZN(n3751) );
  XNOR2_X1 U4644 ( .A(n3877), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3750)
         );
  NAND2_X1 U4645 ( .A1(n3751), .A2(n3750), .ZN(n3879) );
  OR2_X1 U4646 ( .A1(n3751), .A2(n3750), .ZN(n3752) );
  AND2_X1 U4647 ( .A1(n3879), .A2(n3752), .ZN(n6174) );
  NAND2_X1 U4648 ( .A1(n6174), .A2(n6115), .ZN(n3753) );
  OAI211_X1 U4649 ( .C1(n4393), .C2(n5512), .A(n3754), .B(n3753), .ZN(U2985)
         );
  INV_X1 U4650 ( .A(n3755), .ZN(n3757) );
  NAND2_X1 U4651 ( .A1(n3757), .A2(n3756), .ZN(n3759) );
  NAND2_X1 U4652 ( .A1(n3759), .A2(n3758), .ZN(n3767) );
  INV_X1 U4653 ( .A(n3762), .ZN(n3761) );
  NAND2_X1 U4654 ( .A1(n3761), .A2(n6704), .ZN(n4200) );
  NAND2_X1 U4655 ( .A1(n3762), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3763) );
  NAND2_X1 U4656 ( .A1(n4200), .A2(n3763), .ZN(n4078) );
  AOI22_X1 U4657 ( .A1(n3813), .A2(n4078), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3812), .ZN(n3764) );
  OR2_X2 U4658 ( .A1(n3767), .A2(n3766), .ZN(n3808) );
  NAND2_X1 U4659 ( .A1(n3767), .A2(n3766), .ZN(n3768) );
  INV_X1 U4660 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3769) );
  OR2_X1 U4661 ( .A1(n5018), .A2(n3769), .ZN(n3775) );
  NAND2_X1 U4662 ( .A1(n5050), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3774) );
  INV_X1 U4663 ( .A(n3770), .ZN(n5044) );
  INV_X2 U4664 ( .A(n5044), .ZN(n5083) );
  NAND2_X1 U4665 ( .A1(n5083), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3773)
         );
  NAND2_X1 U4666 ( .A1(n5069), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3772) );
  AND4_X1 U4667 ( .A1(n3775), .A2(n3774), .A3(n3773), .A4(n3772), .ZN(n3779)
         );
  AOI22_X1 U4668 ( .A1(n5085), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4669 ( .A1(n3534), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4882), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3777) );
  NAND3_X1 U4670 ( .A1(n3779), .A2(n3778), .A3(n3777), .ZN(n3785) );
  AOI22_X1 U4671 ( .A1(n5076), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3783) );
  AOI22_X1 U4672 ( .A1(n5070), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n5082), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3782) );
  AOI22_X1 U4673 ( .A1(n5026), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3599), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3781) );
  AOI22_X1 U4674 ( .A1(n5081), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3780) );
  NAND4_X1 U4675 ( .A1(n3783), .A2(n3782), .A3(n3781), .A4(n3780), .ZN(n3784)
         );
  OAI22_X2 U4676 ( .A1(n3906), .A2(STATE2_REG_0__SCAN_IN), .B1(n3870), .B2(
        n3786), .ZN(n3790) );
  NAND2_X1 U4677 ( .A1(n3792), .A2(n3791), .ZN(n3796) );
  INV_X1 U4678 ( .A(n3168), .ZN(n3794) );
  NAND2_X1 U4679 ( .A1(n3794), .A2(n3793), .ZN(n3795) );
  XNOR2_X1 U4680 ( .A(n3806), .B(n3805), .ZN(n3932) );
  NAND2_X1 U4681 ( .A1(n3932), .A2(n4648), .ZN(n3797) );
  NAND2_X1 U4682 ( .A1(n3797), .A2(n4710), .ZN(n3802) );
  INV_X1 U4683 ( .A(n3986), .ZN(n3801) );
  OAI21_X1 U4684 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3834), .ZN(n6110) );
  INV_X1 U4685 ( .A(n4710), .ZN(n5210) );
  AOI22_X1 U4686 ( .A1(n5060), .A2(n6110), .B1(n5210), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3800) );
  NAND2_X1 U4687 ( .A1(n5211), .A2(EAX_REG_2__SCAN_IN), .ZN(n3799) );
  NAND2_X1 U4688 ( .A1(n3856), .A2(n3857), .ZN(n3804) );
  NAND2_X1 U4689 ( .A1(n3802), .A2(n3798), .ZN(n3803) );
  INV_X1 U4690 ( .A(n3805), .ZN(n3807) );
  AND2_X2 U4691 ( .A1(n3807), .A2(n3806), .ZN(n3832) );
  BUF_X2 U4692 ( .A(n3808), .Z(n3922) );
  NOR3_X1 U4693 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6704), .A3(n6400), 
        .ZN(n6357) );
  NAND2_X1 U4694 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6357), .ZN(n6387) );
  NAND2_X1 U4695 ( .A1(n6810), .A2(n6387), .ZN(n3811) );
  NAND3_X1 U4696 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n6641) );
  INV_X1 U4697 ( .A(n6641), .ZN(n3810) );
  NAND2_X1 U4698 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3810), .ZN(n6634) );
  AOI22_X1 U4699 ( .A1(n3813), .A2(n6397), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3812), .ZN(n3814) );
  INV_X1 U4700 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3816) );
  OR2_X1 U4701 ( .A1(n5018), .A2(n3816), .ZN(n3820) );
  NAND2_X1 U4702 ( .A1(n5050), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3819) );
  NAND2_X1 U4703 ( .A1(n5083), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3818)
         );
  NAND2_X1 U4704 ( .A1(n5069), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3817) );
  AND4_X1 U4705 ( .A1(n3820), .A2(n3819), .A3(n3818), .A4(n3817), .ZN(n3823)
         );
  AOI22_X1 U4706 ( .A1(n5085), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4707 ( .A1(n3534), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4882), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3821) );
  NAND3_X1 U4708 ( .A1(n3823), .A2(n3822), .A3(n3821), .ZN(n3829) );
  AOI22_X1 U4709 ( .A1(n5076), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4710 ( .A1(n5070), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n5082), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4711 ( .A1(n5026), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3599), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4712 ( .A1(n5081), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3824) );
  NAND4_X1 U4713 ( .A1(n3827), .A2(n3826), .A3(n3825), .A4(n3824), .ZN(n3828)
         );
  AOI22_X1 U4714 ( .A1(n3997), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4261), 
        .B2(n3866), .ZN(n3830) );
  NAND2_X2 U4715 ( .A1(n3831), .A2(n3830), .ZN(n6187) );
  NAND2_X2 U4716 ( .A1(n3832), .A2(n6187), .ZN(n3994) );
  OR2_X2 U4717 ( .A1(n3832), .A2(n6187), .ZN(n3833) );
  INV_X1 U4718 ( .A(EAX_REG_3__SCAN_IN), .ZN(n3837) );
  OAI21_X1 U4719 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3835), .A(n3988), 
        .ZN(n4461) );
  AOI22_X1 U4720 ( .A1(n5060), .A2(n4461), .B1(n5210), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3836) );
  OAI21_X1 U4721 ( .B1(n5008), .B2(n3837), .A(n3836), .ZN(n3838) );
  AOI21_X1 U4722 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n3986), .A(n3838), 
        .ZN(n3839) );
  OAI21_X1 U4723 ( .B1(n3840), .B2(n3841), .A(n3984), .ZN(n4468) );
  MUX2_X1 U4724 ( .A(n5170), .B(n3842), .S(EBX_REG_3__SCAN_IN), .Z(n3843) );
  OAI21_X1 U4725 ( .B1(n5234), .B2(INSTADDRPOINTER_REG_3__SCAN_IN), .A(n3843), 
        .ZN(n3850) );
  INV_X1 U4726 ( .A(n3844), .ZN(n3845) );
  NOR2_X2 U4727 ( .A1(n3846), .A2(n3845), .ZN(n3853) );
  INV_X1 U4728 ( .A(EBX_REG_2__SCAN_IN), .ZN(n3859) );
  NAND2_X1 U4729 ( .A1(n5171), .A2(n3859), .ZN(n3849) );
  OR2_X1 U4730 ( .A1(n5167), .A2(n3859), .ZN(n3848) );
  NAND2_X1 U4731 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n5168), .ZN(n3847)
         );
  NAND4_X1 U4732 ( .A1(n3849), .A2(n5157), .A3(n3848), .A4(n3847), .ZN(n3852)
         );
  NAND2_X1 U4733 ( .A1(n3853), .A2(n3852), .ZN(n3854) );
  NOR2_X2 U4734 ( .A1(n3854), .A2(n3850), .ZN(n3977) );
  AOI21_X1 U4735 ( .B1(n3850), .B2(n3854), .A(n3977), .ZN(n4459) );
  AOI22_X1 U4736 ( .A1(n6018), .A2(n4459), .B1(n5371), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n3851) );
  OAI21_X1 U4737 ( .B1(n4468), .B2(n6012), .A(n3851), .ZN(U2856) );
  OR2_X1 U4738 ( .A1(n3853), .A2(n3852), .ZN(n3855) );
  NAND2_X1 U4739 ( .A1(n3855), .A2(n3854), .ZN(n6164) );
  NOR2_X1 U4740 ( .A1(n3856), .A2(n3857), .ZN(n3858) );
  NOR2_X1 U4741 ( .A1(n3840), .A2(n3858), .ZN(n6107) );
  INV_X1 U4742 ( .A(n6107), .ZN(n4159) );
  OAI222_X1 U4743 ( .A1(n6164), .A2(n6011), .B1(n3859), .B2(n6022), .C1(n4159), 
        .C2(n6012), .ZN(U2857) );
  INV_X1 U4744 ( .A(n3860), .ZN(n3863) );
  INV_X1 U4745 ( .A(n3861), .ZN(n3862) );
  NAND2_X1 U4746 ( .A1(n3863), .A2(n3862), .ZN(n3865) );
  AND2_X1 U4747 ( .A1(n3865), .A2(n3864), .ZN(n6112) );
  INV_X1 U4748 ( .A(n6112), .ZN(n5993) );
  OAI222_X1 U4749 ( .A1(n5991), .A2(n6011), .B1(n6022), .B2(n6001), .C1(n6012), 
        .C2(n5993), .ZN(U2859) );
  NAND2_X1 U4750 ( .A1(n3871), .A2(n3870), .ZN(n3869) );
  NAND2_X1 U4751 ( .A1(n3869), .A2(n3866), .ZN(n4037) );
  OAI211_X1 U4752 ( .C1(n3866), .C2(n3869), .A(n4037), .B(n5239), .ZN(n3867)
         );
  INV_X1 U4753 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3886) );
  XNOR2_X1 U4754 ( .A(n3970), .B(n3886), .ZN(n3969) );
  NAND2_X1 U4755 ( .A1(n3932), .A2(n4296), .ZN(n3875) );
  OAI21_X1 U4756 ( .B1(n3871), .B2(n3870), .A(n3869), .ZN(n3873) );
  AOI21_X1 U4757 ( .B1(n3873), .B2(n5239), .A(n3872), .ZN(n3874) );
  NAND2_X1 U4758 ( .A1(n3875), .A2(n3874), .ZN(n3880) );
  NAND2_X1 U4759 ( .A1(n3880), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6103)
         );
  OR2_X1 U4760 ( .A1(n3877), .A2(n3876), .ZN(n3878) );
  AND2_X1 U4761 ( .A1(n3879), .A2(n3878), .ZN(n6106) );
  NAND2_X1 U4762 ( .A1(n6103), .A2(n6106), .ZN(n3883) );
  INV_X1 U4763 ( .A(n3880), .ZN(n3882) );
  AND2_X1 U4764 ( .A1(n3883), .A2(n6104), .ZN(n3968) );
  XNOR2_X1 U4765 ( .A(n3969), .B(n3968), .ZN(n3949) );
  NAND2_X1 U4766 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6159) );
  NAND2_X1 U4767 ( .A1(n3881), .A2(n6159), .ZN(n6158) );
  NAND2_X1 U4768 ( .A1(n4048), .A2(n5649), .ZN(n5643) );
  NAND2_X1 U4769 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3884) );
  AOI21_X1 U4770 ( .B1(n5643), .B2(n3884), .A(n5641), .ZN(n6168) );
  OAI21_X1 U4771 ( .B1(n5645), .B2(n6158), .A(n6168), .ZN(n3982) );
  NAND2_X1 U4772 ( .A1(n4048), .A2(n3885), .ZN(n6171) );
  NAND2_X1 U4773 ( .A1(n5643), .A2(n6171), .ZN(n5134) );
  INV_X1 U4774 ( .A(n5134), .ZN(n6157) );
  NAND3_X1 U4775 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n6157), .ZN(n4053) );
  NAND2_X1 U4776 ( .A1(n5645), .A2(n4053), .ZN(n4317) );
  NAND2_X1 U4777 ( .A1(n6158), .A2(n4317), .ZN(n4254) );
  INV_X1 U4778 ( .A(n4254), .ZN(n3887) );
  AOI22_X1 U4779 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n3982), .B1(n3887), 
        .B2(n3886), .ZN(n3889) );
  AND2_X1 U4780 ( .A1(n5969), .A2(REIP_REG_3__SCAN_IN), .ZN(n3944) );
  AOI21_X1 U4781 ( .B1(n6172), .B2(n4459), .A(n3944), .ZN(n3888) );
  OAI211_X1 U4782 ( .C1(n3949), .C2(n6125), .A(n3889), .B(n3888), .ZN(U3015)
         );
  NAND2_X1 U4783 ( .A1(n6728), .A2(n6478), .ZN(n6827) );
  INV_X1 U4784 ( .A(n6827), .ZN(n6747) );
  INV_X1 U4785 ( .A(n3914), .ZN(n5668) );
  OAI21_X1 U4786 ( .B1(n5070), .B2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n3540), 
        .ZN(n5676) );
  OR2_X1 U4787 ( .A1(n3893), .A2(n3892), .ZN(n3912) );
  MUX2_X1 U4788 ( .A(n3894), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n5669), 
        .Z(n3895) );
  NOR2_X1 U4789 ( .A1(n3895), .A2(n3917), .ZN(n3896) );
  NAND2_X1 U4790 ( .A1(n3912), .A2(n3896), .ZN(n3901) );
  AND2_X1 U4791 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n5197), .ZN(n3897)
         );
  NOR2_X1 U4792 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n3897), .ZN(n3898)
         );
  OR3_X1 U4793 ( .A1(n5666), .A2(n3899), .A3(n3898), .ZN(n3900) );
  OAI211_X1 U4794 ( .C1(n3908), .C2(n5676), .A(n3901), .B(n3900), .ZN(n3902)
         );
  AOI21_X1 U4795 ( .B1(n6319), .B2(n5668), .A(n3902), .ZN(n5678) );
  NAND2_X1 U4796 ( .A1(n5678), .A2(n3925), .ZN(n3905) );
  NAND2_X1 U4797 ( .A1(n6700), .A2(n3903), .ZN(n3904) );
  NAND2_X1 U4798 ( .A1(n3905), .A2(n3904), .ZN(n6711) );
  XNOR2_X1 U4799 ( .A(n5669), .B(n5197), .ZN(n3911) );
  XNOR2_X1 U4800 ( .A(n5197), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3909)
         );
  OAI22_X1 U4801 ( .A1(n5666), .A2(n3909), .B1(n3908), .B2(n3911), .ZN(n3910)
         );
  AOI21_X1 U4802 ( .B1(n3912), .B2(n3911), .A(n3910), .ZN(n3913) );
  OAI21_X1 U4803 ( .B1(n3907), .B2(n3914), .A(n3913), .ZN(n5200) );
  NOR2_X1 U4804 ( .A1(n3925), .A2(n3191), .ZN(n3915) );
  AOI21_X1 U4805 ( .B1(n5200), .B2(n3925), .A(n3915), .ZN(n6707) );
  OR3_X1 U4806 ( .A1(n6711), .A2(STATE2_REG_1__SCAN_IN), .A3(n6707), .ZN(n3919) );
  NOR2_X1 U4807 ( .A1(FLUSH_REG_SCAN_IN), .A2(n6728), .ZN(n3916) );
  NAND2_X1 U4808 ( .A1(n3917), .A2(n3916), .ZN(n3918) );
  NAND2_X1 U4809 ( .A1(n3919), .A2(n3918), .ZN(n6720) );
  INV_X1 U4810 ( .A(n5670), .ZN(n5663) );
  NAND2_X1 U4811 ( .A1(n6720), .A2(n5663), .ZN(n3929) );
  INV_X1 U4812 ( .A(n6536), .ZN(n3921) );
  NOR2_X1 U4813 ( .A1(n3922), .A2(n3921), .ZN(n3923) );
  XNOR2_X1 U4814 ( .A(n3923), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5966)
         );
  OR2_X1 U4815 ( .A1(n5825), .A2(STATE2_REG_1__SCAN_IN), .ZN(n3924) );
  OR2_X1 U4816 ( .A1(n5966), .A2(n3924), .ZN(n3928) );
  MUX2_X1 U4817 ( .A(n3925), .B(FLUSH_REG_SCAN_IN), .S(STATE2_REG_1__SCAN_IN), 
        .Z(n3926) );
  OR2_X1 U4818 ( .A1(n3926), .A2(n5831), .ZN(n3927) );
  AND2_X1 U4819 ( .A1(n3928), .A2(n3927), .ZN(n6718) );
  NAND2_X1 U4820 ( .A1(n3929), .A2(n6718), .ZN(n6724) );
  OAI21_X1 U4821 ( .B1(n6724), .B2(FLUSH_REG_SCAN_IN), .A(n3930), .ZN(n3931)
         );
  NAND2_X1 U4822 ( .A1(n6404), .A2(n3931), .ZN(n6808) );
  NAND2_X1 U4823 ( .A1(n3935), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6347) );
  XNOR2_X1 U4824 ( .A(n3933), .B(n6347), .ZN(n3936) );
  INV_X1 U4825 ( .A(n3907), .ZN(n6182) );
  NOR2_X1 U4826 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6728), .ZN(n6803) );
  INV_X1 U4827 ( .A(n6803), .ZN(n6813) );
  AOI22_X1 U4828 ( .A1(n3936), .A2(n6812), .B1(n6182), .B2(n6813), .ZN(n3938)
         );
  NAND2_X1 U4829 ( .A1(n6818), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3937) );
  OAI21_X1 U4830 ( .B1(n6818), .B2(n3938), .A(n3937), .ZN(U3463) );
  AOI21_X1 U4831 ( .B1(n6394), .B2(n6912), .A(n6802), .ZN(n3941) );
  INV_X1 U4832 ( .A(n3940), .ZN(n6181) );
  AOI22_X1 U4833 ( .A1(n3941), .A2(n6347), .B1(n6181), .B2(n6813), .ZN(n3943)
         );
  NAND2_X1 U4834 ( .A1(n6818), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3942) );
  OAI21_X1 U4835 ( .B1(n6818), .B2(n3943), .A(n3942), .ZN(U3464) );
  INV_X1 U4836 ( .A(n4468), .ZN(n3947) );
  AOI21_X1 U4837 ( .B1(n6117), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n3944), 
        .ZN(n3945) );
  OAI21_X1 U4838 ( .B1(n4461), .B2(n6111), .A(n3945), .ZN(n3946) );
  AOI21_X1 U4839 ( .B1(n3947), .B2(n6113), .A(n3946), .ZN(n3948) );
  OAI21_X1 U4840 ( .B1(n3949), .B2(n5835), .A(n3948), .ZN(U2983) );
  INV_X1 U4841 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4474) );
  INV_X1 U4842 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3950) );
  OR2_X1 U4843 ( .A1(n5018), .A2(n3950), .ZN(n3954) );
  NAND2_X1 U4844 ( .A1(n5050), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3953) );
  NAND2_X1 U4845 ( .A1(n5083), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3952)
         );
  NAND2_X1 U4846 ( .A1(n5069), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3951) );
  AND4_X1 U4847 ( .A1(n3954), .A2(n3953), .A3(n3952), .A4(n3951), .ZN(n3957)
         );
  AOI22_X1 U4848 ( .A1(n5085), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3956) );
  AOI22_X1 U4849 ( .A1(n3534), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4882), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3955) );
  NAND3_X1 U4850 ( .A1(n3957), .A2(n3956), .A3(n3955), .ZN(n3963) );
  AOI22_X1 U4851 ( .A1(n5076), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3961) );
  AOI22_X1 U4852 ( .A1(n5070), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n5082), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3960) );
  AOI22_X1 U4853 ( .A1(n5026), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3599), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3959) );
  INV_X2 U4854 ( .A(n3540), .ZN(n5086) );
  AOI22_X1 U4855 ( .A1(n5081), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3958) );
  NAND4_X1 U4856 ( .A1(n3961), .A2(n3960), .A3(n3959), .A4(n3958), .ZN(n3962)
         );
  NAND2_X1 U4857 ( .A1(n4261), .A2(n4035), .ZN(n3964) );
  OAI21_X1 U4858 ( .B1(n4263), .B2(n4474), .A(n3964), .ZN(n3995) );
  XNOR2_X1 U4859 ( .A(n3994), .B(n3995), .ZN(n3985) );
  NAND2_X1 U4860 ( .A1(n3985), .A2(n4296), .ZN(n3967) );
  XNOR2_X1 U4861 ( .A(n4037), .B(n4035), .ZN(n3965) );
  NAND2_X1 U4862 ( .A1(n3965), .A2(n5239), .ZN(n3966) );
  NAND2_X1 U4863 ( .A1(n3967), .A2(n3966), .ZN(n4044) );
  INV_X1 U4864 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3973) );
  XNOR2_X1 U4865 ( .A(n4044), .B(n3973), .ZN(n4042) );
  NAND2_X1 U4866 ( .A1(n3969), .A2(n3968), .ZN(n3972) );
  NAND2_X1 U4867 ( .A1(n3163), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3971)
         );
  XNOR2_X1 U4868 ( .A(n4042), .B(n4043), .ZN(n4130) );
  NAND2_X1 U4869 ( .A1(n5167), .A2(n3973), .ZN(n3974) );
  OAI211_X1 U4870 ( .C1(n5168), .C2(EBX_REG_4__SCAN_IN), .A(n3974), .B(n3842), 
        .ZN(n3975) );
  OAI21_X1 U4871 ( .B1(n5227), .B2(EBX_REG_4__SCAN_IN), .A(n3975), .ZN(n3976)
         );
  OR2_X1 U4872 ( .A1(n3976), .A2(n3977), .ZN(n3978) );
  NAND2_X1 U4873 ( .A1(n3978), .A2(n4031), .ZN(n4123) );
  NAND2_X1 U4874 ( .A1(n5969), .A2(REIP_REG_4__SCAN_IN), .ZN(n4125) );
  OAI21_X1 U4875 ( .B1(n6163), .B2(n4123), .A(n4125), .ZN(n3981) );
  NAND2_X1 U4876 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4054) );
  OAI21_X1 U4877 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4054), .ZN(n3979) );
  NOR2_X1 U4878 ( .A1(n4254), .A2(n3979), .ZN(n3980) );
  AOI211_X1 U4879 ( .C1(n3982), .C2(INSTADDRPOINTER_REG_4__SCAN_IN), .A(n3981), 
        .B(n3980), .ZN(n3983) );
  OAI21_X1 U4880 ( .B1(n6125), .B2(n4130), .A(n3983), .ZN(U3014) );
  INV_X1 U4881 ( .A(n3984), .ZN(n3993) );
  NAND2_X1 U4882 ( .A1(n3986), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3990) );
  AOI21_X1 U4883 ( .B1(n4127), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3987) );
  AOI21_X1 U4884 ( .B1(n5211), .B2(EAX_REG_4__SCAN_IN), .A(n3987), .ZN(n3989)
         );
  AOI21_X1 U4885 ( .B1(n4127), .B2(n3988), .A(n4019), .ZN(n5970) );
  AOI22_X1 U4886 ( .A1(n3990), .A2(n3989), .B1(n5060), .B2(n5970), .ZN(n3991)
         );
  NAND2_X1 U4887 ( .A1(n3993), .A2(n3992), .ZN(n4027) );
  INV_X1 U4888 ( .A(n3994), .ZN(n3996) );
  NAND2_X1 U4889 ( .A1(n3996), .A2(n3995), .ZN(n4017) );
  INV_X1 U4890 ( .A(n4017), .ZN(n4015) );
  NAND2_X1 U4891 ( .A1(n3997), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4013) );
  INV_X1 U4892 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3998) );
  OR2_X1 U4893 ( .A1(n5018), .A2(n3998), .ZN(n4002) );
  NAND2_X1 U4894 ( .A1(n5050), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4001) );
  NAND2_X1 U4895 ( .A1(n5070), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4000) );
  NAND2_X1 U4896 ( .A1(n5082), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3999)
         );
  AND4_X1 U4897 ( .A1(n4002), .A2(n4001), .A3(n4000), .A4(n3999), .ZN(n4005)
         );
  AOI22_X1 U4898 ( .A1(n5085), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3534), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4004) );
  AOI22_X1 U4899 ( .A1(n5076), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4882), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4003) );
  NAND3_X1 U4900 ( .A1(n4005), .A2(n4004), .A3(n4003), .ZN(n4011) );
  AOI22_X1 U4901 ( .A1(n5026), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4009) );
  AOI22_X1 U4902 ( .A1(n5081), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3599), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U4903 ( .A1(n5083), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5069), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4007) );
  AOI22_X1 U4904 ( .A1(n5075), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4006) );
  NAND4_X1 U4905 ( .A1(n4009), .A2(n4008), .A3(n4007), .A4(n4006), .ZN(n4010)
         );
  NAND2_X1 U4906 ( .A1(n4261), .A2(n4038), .ZN(n4012) );
  INV_X1 U4907 ( .A(n4016), .ZN(n4014) );
  NAND2_X1 U4908 ( .A1(n4017), .A2(n4016), .ZN(n4018) );
  AND2_X2 U4909 ( .A1(n4178), .A2(n4018), .ZN(n4034) );
  INV_X1 U4910 ( .A(EAX_REG_5__SCAN_IN), .ZN(n4024) );
  INV_X1 U4911 ( .A(n4182), .ZN(n4184) );
  INV_X1 U4912 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4021) );
  INV_X1 U4913 ( .A(n4019), .ZN(n4020) );
  NAND2_X1 U4914 ( .A1(n4021), .A2(n4020), .ZN(n4022) );
  NAND2_X1 U4915 ( .A1(n4184), .A2(n4022), .ZN(n5954) );
  AOI22_X1 U4916 ( .A1(n5954), .A2(n5060), .B1(n5210), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4023) );
  OAI21_X1 U4917 ( .B1(n5008), .B2(n4024), .A(n4023), .ZN(n4025) );
  AND2_X1 U4918 ( .A1(n4027), .A2(n4026), .ZN(n4029) );
  NOR2_X2 U4919 ( .A1(n4027), .A2(n4026), .ZN(n4191) );
  CLKBUF_X1 U4920 ( .A(n4191), .Z(n4028) );
  OR2_X1 U4921 ( .A1(n4029), .A2(n4028), .ZN(n5955) );
  MUX2_X1 U4922 ( .A(n5170), .B(n3842), .S(EBX_REG_5__SCAN_IN), .Z(n4030) );
  OAI21_X1 U4923 ( .B1(n5234), .B2(INSTADDRPOINTER_REG_5__SCAN_IN), .A(n4030), 
        .ZN(n4032) );
  AOI21_X1 U4924 ( .B1(n4032), .B2(n4031), .A(n4277), .ZN(n5957) );
  AOI22_X1 U4925 ( .A1(n6018), .A2(n5957), .B1(n5371), .B2(EBX_REG_5__SCAN_IN), 
        .ZN(n4033) );
  OAI21_X1 U4926 ( .B1(n5955), .B2(n6012), .A(n4033), .ZN(U2854) );
  NAND2_X1 U4927 ( .A1(n4034), .A2(n4296), .ZN(n4041) );
  INV_X1 U4928 ( .A(n4035), .ZN(n4036) );
  NOR2_X1 U4929 ( .A1(n4037), .A2(n4036), .ZN(n4039) );
  NAND2_X1 U4930 ( .A1(n4039), .A2(n4038), .ZN(n4288) );
  OAI211_X1 U4931 ( .C1(n4039), .C2(n4038), .A(n4288), .B(n5239), .ZN(n4040)
         );
  NAND2_X1 U4932 ( .A1(n4041), .A2(n4040), .ZN(n4239) );
  INV_X1 U4933 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4051) );
  XNOR2_X1 U4934 ( .A(n4239), .B(n4051), .ZN(n4237) );
  NAND2_X1 U4935 ( .A1(n4043), .A2(n4042), .ZN(n4046) );
  NAND2_X1 U4936 ( .A1(n4044), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4045)
         );
  NAND2_X1 U4937 ( .A1(n4046), .A2(n4045), .ZN(n4238) );
  XNOR2_X1 U4938 ( .A(n4237), .B(n3161), .ZN(n4149) );
  INV_X1 U4939 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6768) );
  NOR2_X1 U4940 ( .A1(n5819), .A2(n6768), .ZN(n4144) );
  INV_X1 U4941 ( .A(n4054), .ZN(n4047) );
  NAND3_X1 U4942 ( .A1(n6161), .A2(n4047), .A3(n6158), .ZN(n4050) );
  NOR2_X1 U4943 ( .A1(n4051), .A2(n4054), .ZN(n4253) );
  NAND2_X1 U4944 ( .A1(n4253), .A2(n6158), .ZN(n4307) );
  NAND2_X1 U4945 ( .A1(n5639), .A2(n4048), .ZN(n6170) );
  INV_X1 U4946 ( .A(n6168), .ZN(n4049) );
  AOI21_X1 U4947 ( .B1(n4307), .B2(n6170), .A(n4049), .ZN(n4255) );
  AOI21_X1 U4948 ( .B1(n4051), .B2(n4050), .A(n4255), .ZN(n4052) );
  AOI211_X1 U4949 ( .C1(n6172), .C2(n5957), .A(n4144), .B(n4052), .ZN(n4056)
         );
  OR3_X1 U4950 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n4054), .A3(n4053), 
        .ZN(n4055) );
  OAI211_X1 U4951 ( .C1(n6125), .C2(n4149), .A(n4056), .B(n4055), .ZN(U3013)
         );
  INV_X1 U4952 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4058) );
  AOI22_X1 U4953 ( .A1(n4063), .A2(UWORD_REG_4__SCAN_IN), .B1(n6058), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4057) );
  OAI21_X1 U4954 ( .B1(n4058), .B2(n4072), .A(n4057), .ZN(U2903) );
  INV_X1 U4955 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4060) );
  AOI22_X1 U4956 ( .A1(n4063), .A2(UWORD_REG_5__SCAN_IN), .B1(n6058), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4059) );
  OAI21_X1 U4957 ( .B1(n4060), .B2(n4072), .A(n4059), .ZN(U2902) );
  INV_X1 U4958 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4062) );
  AOI22_X1 U4959 ( .A1(n4063), .A2(UWORD_REG_7__SCAN_IN), .B1(n6058), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4061) );
  OAI21_X1 U4960 ( .B1(n4062), .B2(n4072), .A(n4061), .ZN(U2900) );
  INV_X1 U4961 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4065) );
  AOI22_X1 U4962 ( .A1(n4063), .A2(UWORD_REG_6__SCAN_IN), .B1(n6058), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4064) );
  OAI21_X1 U4963 ( .B1(n4065), .B2(n4072), .A(n4064), .ZN(U2901) );
  INV_X1 U4964 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4067) );
  INV_X1 U4965 ( .A(n6832), .ZN(n6059) );
  AOI22_X1 U4966 ( .A1(n6059), .A2(UWORD_REG_1__SCAN_IN), .B1(n6058), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4066) );
  OAI21_X1 U4967 ( .B1(n4067), .B2(n4072), .A(n4066), .ZN(U2906) );
  INV_X1 U4968 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4069) );
  AOI22_X1 U4969 ( .A1(n6059), .A2(UWORD_REG_3__SCAN_IN), .B1(n6058), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4068) );
  OAI21_X1 U4970 ( .B1(n4069), .B2(n4072), .A(n4068), .ZN(U2904) );
  AOI22_X1 U4971 ( .A1(n6059), .A2(UWORD_REG_2__SCAN_IN), .B1(n6058), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4070) );
  OAI21_X1 U4972 ( .B1(n4735), .B2(n4072), .A(n4070), .ZN(U2905) );
  INV_X1 U4973 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4073) );
  AOI22_X1 U4974 ( .A1(n6059), .A2(UWORD_REG_0__SCAN_IN), .B1(n6058), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4071) );
  OAI21_X1 U4975 ( .B1(n4073), .B2(n4072), .A(n4071), .ZN(U2907) );
  INV_X1 U4976 ( .A(n6187), .ZN(n4194) );
  NAND2_X1 U4977 ( .A1(n3933), .A2(n4194), .ZN(n6351) );
  INV_X1 U4978 ( .A(DATAI_19_), .ZN(n7047) );
  NOR2_X1 U4979 ( .A1(n5512), .A2(n7047), .ZN(n6664) );
  INV_X1 U4980 ( .A(n6664), .ZN(n6613) );
  OR2_X1 U4981 ( .A1(n6279), .A2(n6912), .ZN(n4074) );
  NAND2_X1 U4982 ( .A1(n4074), .A2(n6812), .ZN(n6288) );
  INV_X1 U4983 ( .A(n3933), .ZN(n6180) );
  NAND3_X1 U4984 ( .A1(n6806), .A2(n6180), .A3(n3935), .ZN(n4208) );
  INV_X1 U4985 ( .A(n6811), .ZN(n6589) );
  AND2_X1 U4986 ( .A1(n6812), .A2(n6912), .ZN(n6252) );
  OR2_X1 U4987 ( .A1(n3907), .A2(n6181), .ZN(n6281) );
  OAI22_X1 U4988 ( .A1(n4236), .A2(n6252), .B1(n6536), .B2(n6281), .ZN(n4076)
         );
  NAND2_X1 U4989 ( .A1(n6400), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6562) );
  OR2_X1 U4990 ( .A1(n6562), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6287)
         );
  OR2_X1 U4991 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6287), .ZN(n4115)
         );
  INV_X1 U4992 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6637) );
  NOR2_X1 U4993 ( .A1(n4078), .A2(n6637), .ZN(n6324) );
  NOR2_X1 U4994 ( .A1(n6480), .A2(n6397), .ZN(n6183) );
  OAI21_X1 U4995 ( .B1(n6183), .B2(n6478), .A(n6256), .ZN(n6185) );
  AOI211_X1 U4996 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4115), .A(n6324), .B(
        n6185), .ZN(n4075) );
  OAI21_X1 U4997 ( .B1(n6288), .B2(n4076), .A(n4075), .ZN(n4112) );
  NAND2_X1 U4998 ( .A1(n4112), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4084) );
  INV_X1 U4999 ( .A(DATAI_27_), .ZN(n4077) );
  NOR2_X1 U5000 ( .A1(n5512), .A2(n4077), .ZN(n6610) );
  INV_X1 U5001 ( .A(DATAI_3_), .ZN(n6934) );
  NOR2_X2 U5002 ( .A1(n6934), .A2(n6404), .ZN(n6663) );
  INV_X1 U5003 ( .A(n6663), .ZN(n6373) );
  NOR2_X1 U5004 ( .A1(n6281), .A2(n6802), .ZN(n6531) );
  AND2_X1 U5005 ( .A1(n4078), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6317) );
  AOI22_X1 U5006 ( .A1(n6531), .A2(n6804), .B1(n6317), .B2(n6183), .ZN(n4116)
         );
  NAND2_X1 U5007 ( .A1(n4114), .A2(n4081), .ZN(n6493) );
  OAI22_X1 U5008 ( .A1(n6373), .A2(n4116), .B1(n6493), .B2(n4115), .ZN(n4082)
         );
  AOI21_X1 U5009 ( .B1(n4118), .B2(n6610), .A(n4082), .ZN(n4083) );
  OAI211_X1 U5010 ( .C1(n6316), .C2(n6613), .A(n4084), .B(n4083), .ZN(U3055)
         );
  INV_X1 U5011 ( .A(DATAI_17_), .ZN(n7198) );
  NOR2_X1 U5012 ( .A1(n5512), .A2(n7198), .ZN(n6652) );
  INV_X1 U5013 ( .A(n6652), .ZN(n6605) );
  NAND2_X1 U5014 ( .A1(n4112), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4089) );
  INV_X1 U5015 ( .A(DATAI_25_), .ZN(n4085) );
  NOR2_X1 U5016 ( .A1(n5512), .A2(n4085), .ZN(n6602) );
  INV_X1 U5017 ( .A(DATAI_1_), .ZN(n7170) );
  NOR2_X2 U5018 ( .A1(n7170), .A2(n6404), .ZN(n6651) );
  INV_X1 U5019 ( .A(n6651), .ZN(n6365) );
  NAND2_X1 U5020 ( .A1(n4114), .A2(n4086), .ZN(n6485) );
  OAI22_X1 U5021 ( .A1(n6365), .A2(n4116), .B1(n6485), .B2(n4115), .ZN(n4087)
         );
  AOI21_X1 U5022 ( .B1(n4118), .B2(n6602), .A(n4087), .ZN(n4088) );
  OAI211_X1 U5023 ( .C1(n6316), .C2(n6605), .A(n4089), .B(n4088), .ZN(U3053)
         );
  INV_X1 U5024 ( .A(DATAI_20_), .ZN(n7059) );
  NOR2_X1 U5025 ( .A1(n5512), .A2(n7059), .ZN(n6670) );
  INV_X1 U5026 ( .A(n6670), .ZN(n6617) );
  NAND2_X1 U5027 ( .A1(n4112), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4094) );
  INV_X1 U5028 ( .A(DATAI_28_), .ZN(n4090) );
  NOR2_X1 U5029 ( .A1(n5512), .A2(n4090), .ZN(n6614) );
  INV_X1 U5030 ( .A(DATAI_4_), .ZN(n6972) );
  NOR2_X2 U5031 ( .A1(n6972), .A2(n6404), .ZN(n6669) );
  INV_X1 U5032 ( .A(n6669), .ZN(n6377) );
  NAND2_X1 U5033 ( .A1(n4114), .A2(n4091), .ZN(n6497) );
  OAI22_X1 U5034 ( .A1(n6377), .A2(n4116), .B1(n6497), .B2(n4115), .ZN(n4092)
         );
  AOI21_X1 U5035 ( .B1(n4118), .B2(n6614), .A(n4092), .ZN(n4093) );
  OAI211_X1 U5036 ( .C1(n6316), .C2(n6617), .A(n4094), .B(n4093), .ZN(U3056)
         );
  INV_X1 U5037 ( .A(DATAI_16_), .ZN(n7044) );
  NOR2_X1 U5038 ( .A1(n5512), .A2(n7044), .ZN(n6646) );
  INV_X1 U5039 ( .A(n6646), .ZN(n6601) );
  NAND2_X1 U5040 ( .A1(n4112), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4098) );
  INV_X1 U5041 ( .A(DATAI_24_), .ZN(n4095) );
  NOR2_X1 U5042 ( .A1(n5512), .A2(n4095), .ZN(n6598) );
  INV_X1 U5043 ( .A(DATAI_0_), .ZN(n6081) );
  NOR2_X2 U5044 ( .A1(n6081), .A2(n6404), .ZN(n6639) );
  INV_X1 U5045 ( .A(n6639), .ZN(n6360) );
  NAND2_X1 U5046 ( .A1(n4114), .A2(n4385), .ZN(n6471) );
  OAI22_X1 U5047 ( .A1(n6360), .A2(n4116), .B1(n6471), .B2(n4115), .ZN(n4096)
         );
  AOI21_X1 U5048 ( .B1(n4118), .B2(n6598), .A(n4096), .ZN(n4097) );
  OAI211_X1 U5049 ( .C1(n6601), .C2(n6316), .A(n4098), .B(n4097), .ZN(U3052)
         );
  INV_X1 U5050 ( .A(DATAI_22_), .ZN(n7153) );
  NOR2_X1 U5051 ( .A1(n5512), .A2(n7153), .ZN(n6682) );
  INV_X1 U5052 ( .A(n6682), .ZN(n6625) );
  NAND2_X1 U5053 ( .A1(n4112), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4102) );
  INV_X1 U5054 ( .A(DATAI_30_), .ZN(n4099) );
  NOR2_X1 U5055 ( .A1(n5512), .A2(n4099), .ZN(n6622) );
  INV_X1 U5056 ( .A(DATAI_6_), .ZN(n6995) );
  NOR2_X2 U5057 ( .A1(n6995), .A2(n6404), .ZN(n6681) );
  INV_X1 U5058 ( .A(n6681), .ZN(n6385) );
  NAND2_X1 U5059 ( .A1(n4114), .A2(n3469), .ZN(n6505) );
  OAI22_X1 U5060 ( .A1(n6385), .A2(n4116), .B1(n6505), .B2(n4115), .ZN(n4100)
         );
  AOI21_X1 U5061 ( .B1(n4118), .B2(n6622), .A(n4100), .ZN(n4101) );
  OAI211_X1 U5062 ( .C1(n6316), .C2(n6625), .A(n4102), .B(n4101), .ZN(U3058)
         );
  INV_X1 U5063 ( .A(DATAI_21_), .ZN(n7151) );
  NOR2_X1 U5064 ( .A1(n5512), .A2(n7151), .ZN(n6676) );
  INV_X1 U5065 ( .A(n6676), .ZN(n6621) );
  NAND2_X1 U5066 ( .A1(n4112), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4106) );
  INV_X1 U5067 ( .A(DATAI_29_), .ZN(n4103) );
  NOR2_X1 U5068 ( .A1(n5512), .A2(n4103), .ZN(n6618) );
  INV_X1 U5069 ( .A(DATAI_5_), .ZN(n7161) );
  NOR2_X2 U5070 ( .A1(n7161), .A2(n6404), .ZN(n6675) );
  INV_X1 U5071 ( .A(n6675), .ZN(n6381) );
  NAND2_X1 U5072 ( .A1(n4114), .A2(n4773), .ZN(n6501) );
  OAI22_X1 U5073 ( .A1(n6381), .A2(n4116), .B1(n6501), .B2(n4115), .ZN(n4104)
         );
  AOI21_X1 U5074 ( .B1(n4118), .B2(n6618), .A(n4104), .ZN(n4105) );
  OAI211_X1 U5075 ( .C1(n6316), .C2(n6621), .A(n4106), .B(n4105), .ZN(U3057)
         );
  INV_X1 U5076 ( .A(DATAI_18_), .ZN(n4107) );
  NOR2_X1 U5077 ( .A1(n5512), .A2(n4107), .ZN(n6658) );
  INV_X1 U5078 ( .A(n6658), .ZN(n6609) );
  NAND2_X1 U5079 ( .A1(n4112), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4111) );
  NOR2_X1 U5080 ( .A1(n5512), .A2(n7037), .ZN(n6606) );
  INV_X1 U5081 ( .A(DATAI_2_), .ZN(n7145) );
  NOR2_X2 U5082 ( .A1(n7145), .A2(n6404), .ZN(n6657) );
  INV_X1 U5083 ( .A(n6657), .ZN(n6369) );
  NAND2_X1 U5084 ( .A1(n4114), .A2(n4108), .ZN(n6489) );
  OAI22_X1 U5085 ( .A1(n6369), .A2(n4116), .B1(n6489), .B2(n4115), .ZN(n4109)
         );
  AOI21_X1 U5086 ( .B1(n4118), .B2(n6606), .A(n4109), .ZN(n4110) );
  OAI211_X1 U5087 ( .C1(n6316), .C2(n6609), .A(n4111), .B(n4110), .ZN(U3054)
         );
  INV_X1 U5088 ( .A(DATAI_23_), .ZN(n7147) );
  NOR2_X1 U5089 ( .A1(n5512), .A2(n7147), .ZN(n6691) );
  INV_X1 U5090 ( .A(n6691), .ZN(n6633) );
  NAND2_X1 U5091 ( .A1(n4112), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4120) );
  INV_X1 U5092 ( .A(DATAI_31_), .ZN(n4113) );
  NOR2_X1 U5093 ( .A1(n5512), .A2(n4113), .ZN(n6629) );
  INV_X1 U5094 ( .A(DATAI_7_), .ZN(n6991) );
  NOR2_X2 U5095 ( .A1(n6991), .A2(n6404), .ZN(n6689) );
  INV_X1 U5096 ( .A(n6689), .ZN(n6392) );
  NAND2_X1 U5097 ( .A1(n4114), .A2(n4155), .ZN(n6510) );
  OAI22_X1 U5098 ( .A1(n6392), .A2(n4116), .B1(n6510), .B2(n4115), .ZN(n4117)
         );
  AOI21_X1 U5099 ( .B1(n4118), .B2(n6629), .A(n4117), .ZN(n4119) );
  OAI211_X1 U5100 ( .C1(n6316), .C2(n6633), .A(n4120), .B(n4119), .ZN(U3059)
         );
  INV_X1 U5101 ( .A(n4027), .ZN(n4121) );
  AOI21_X1 U5102 ( .B1(n4122), .B2(n3984), .A(n4121), .ZN(n5971) );
  INV_X1 U5103 ( .A(n5971), .ZN(n4160) );
  INV_X1 U5104 ( .A(n4123), .ZN(n5964) );
  AOI22_X1 U5105 ( .A1(n6018), .A2(n5964), .B1(n5371), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4124) );
  OAI21_X1 U5106 ( .B1(n4160), .B2(n6012), .A(n4124), .ZN(U2855) );
  NAND2_X1 U5107 ( .A1(n5781), .A2(n5970), .ZN(n4126) );
  OAI211_X1 U5108 ( .C1(n5786), .C2(n4127), .A(n4126), .B(n4125), .ZN(n4128)
         );
  AOI21_X1 U5109 ( .B1(n5971), .B2(n6113), .A(n4128), .ZN(n4129) );
  OAI21_X1 U5110 ( .B1(n5835), .B2(n4130), .A(n4129), .ZN(U2982) );
  INV_X1 U5111 ( .A(n6629), .ZN(n6696) );
  OAI21_X1 U5112 ( .B1(n6427), .B2(n6347), .A(n6812), .ZN(n4137) );
  NAND2_X1 U5113 ( .A1(n3907), .A2(n6181), .ZN(n4199) );
  INV_X1 U5114 ( .A(n4199), .ZN(n4131) );
  NAND2_X1 U5115 ( .A1(n4131), .A2(n6319), .ZN(n6481) );
  OR2_X1 U5116 ( .A1(n6481), .A2(n6430), .ZN(n4133) );
  NOR2_X1 U5117 ( .A1(n4200), .A2(n6810), .ZN(n6525) );
  INV_X1 U5118 ( .A(n6525), .ZN(n4132) );
  AND2_X1 U5119 ( .A1(n4133), .A2(n4132), .ZN(n4136) );
  INV_X1 U5120 ( .A(n4136), .ZN(n4135) );
  NAND3_X1 U5121 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6704), .ZN(n6470) );
  OAI21_X1 U5122 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6798), .A(n6256), 
        .ZN(n6284) );
  AOI21_X1 U5123 ( .B1(n6802), .B2(n6470), .A(n6284), .ZN(n4134) );
  OAI21_X1 U5124 ( .B1(n4137), .B2(n4135), .A(n4134), .ZN(n6527) );
  OAI22_X1 U5125 ( .A1(n4137), .A2(n4136), .B1(n6478), .B2(n6470), .ZN(n6526)
         );
  AOI22_X1 U5126 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6527), .B1(n6689), 
        .B2(n6526), .ZN(n4139) );
  INV_X1 U5127 ( .A(n6510), .ZN(n6686) );
  NAND2_X1 U5128 ( .A1(n3935), .A2(n6811), .ZN(n6350) );
  NOR2_X2 U5129 ( .A1(n6427), .A2(n6350), .ZN(n6557) );
  AOI22_X1 U5130 ( .A1(n6686), .A2(n6525), .B1(n6557), .B2(n6691), .ZN(n4138)
         );
  OAI211_X1 U5131 ( .C1(n6696), .C2(n6530), .A(n4139), .B(n4138), .ZN(U3115)
         );
  INV_X1 U5132 ( .A(n6622), .ZN(n6685) );
  AOI22_X1 U5133 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6527), .B1(n6681), 
        .B2(n6526), .ZN(n4141) );
  INV_X1 U5134 ( .A(n6505), .ZN(n6680) );
  AOI22_X1 U5135 ( .A1(n6680), .A2(n6525), .B1(n6557), .B2(n6682), .ZN(n4140)
         );
  OAI211_X1 U5136 ( .C1(n6685), .C2(n6530), .A(n4141), .B(n4140), .ZN(U3114)
         );
  INV_X1 U5137 ( .A(n6618), .ZN(n6679) );
  AOI22_X1 U5138 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6527), .B1(n6675), 
        .B2(n6526), .ZN(n4143) );
  INV_X1 U5139 ( .A(n6501), .ZN(n6674) );
  AOI22_X1 U5140 ( .A1(n6674), .A2(n6525), .B1(n6557), .B2(n6676), .ZN(n4142)
         );
  OAI211_X1 U5141 ( .C1(n6679), .C2(n6530), .A(n4143), .B(n4142), .ZN(U3113)
         );
  INV_X1 U5142 ( .A(n5955), .ZN(n4147) );
  AOI21_X1 U5143 ( .B1(n6117), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n4144), 
        .ZN(n4145) );
  OAI21_X1 U5144 ( .B1(n5954), .B2(n6111), .A(n4145), .ZN(n4146) );
  AOI21_X1 U5145 ( .B1(n4147), .B2(n6113), .A(n4146), .ZN(n4148) );
  OAI21_X1 U5146 ( .B1(n5835), .B2(n4149), .A(n4148), .ZN(U2981) );
  NAND2_X1 U5147 ( .A1(n4150), .A2(n6738), .ZN(n4153) );
  OR3_X2 U5148 ( .A1(n4152), .A2(n4151), .A3(READY_N), .ZN(n6102) );
  NAND2_X1 U5149 ( .A1(n4156), .A2(n4155), .ZN(n4157) );
  INV_X1 U5150 ( .A(n4157), .ZN(n4158) );
  INV_X1 U5151 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6056) );
  OAI222_X1 U5152 ( .A1(n4159), .A2(n5391), .B1(n4659), .B2(n7145), .C1(n5219), 
        .C2(n6056), .ZN(U2889) );
  OAI222_X1 U5153 ( .A1(n4468), .A2(n5391), .B1(n4659), .B2(n6934), .C1(n6032), 
        .C2(n3837), .ZN(U2888) );
  INV_X1 U5154 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6053) );
  OAI222_X1 U5155 ( .A1(n4160), .A2(n5391), .B1(n4659), .B2(n6972), .C1(n5219), 
        .C2(n6053), .ZN(U2887) );
  OAI222_X1 U5156 ( .A1(n5955), .A2(n5391), .B1(n4659), .B2(n7161), .C1(n5219), 
        .C2(n4024), .ZN(U2886) );
  INV_X1 U5157 ( .A(n4178), .ZN(n4175) );
  INV_X1 U5158 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4591) );
  INV_X1 U5159 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n5043) );
  OR2_X1 U5160 ( .A1(n5018), .A2(n5043), .ZN(n4164) );
  NAND2_X1 U5161 ( .A1(n5050), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4163) );
  NAND2_X1 U5162 ( .A1(n5083), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4162)
         );
  NAND2_X1 U5163 ( .A1(n5069), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4161) );
  AND4_X1 U5164 ( .A1(n4164), .A2(n4163), .A3(n4162), .A4(n4161), .ZN(n4167)
         );
  AOI22_X1 U5165 ( .A1(n5085), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4166) );
  AOI22_X1 U5166 ( .A1(n3534), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4882), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4165) );
  NAND3_X1 U5167 ( .A1(n4167), .A2(n4166), .A3(n4165), .ZN(n4173) );
  AOI22_X1 U5168 ( .A1(n5076), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4171) );
  AOI22_X1 U5169 ( .A1(n5070), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n5082), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4170) );
  AOI22_X1 U5170 ( .A1(n5026), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3599), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4169) );
  AOI22_X1 U5171 ( .A1(n5081), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4168) );
  NAND4_X1 U5172 ( .A1(n4171), .A2(n4170), .A3(n4169), .A4(n4168), .ZN(n4172)
         );
  OR2_X1 U5173 ( .A1(n4173), .A2(n4172), .ZN(n4286) );
  NAND2_X1 U5174 ( .A1(n4261), .A2(n4286), .ZN(n4174) );
  OAI21_X1 U5175 ( .B1(n4263), .B2(n4591), .A(n4174), .ZN(n4176) );
  INV_X1 U5176 ( .A(n4244), .ZN(n4180) );
  NAND2_X1 U5177 ( .A1(n4180), .A2(n4648), .ZN(n4190) );
  INV_X1 U5178 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4181) );
  INV_X1 U5179 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4183) );
  OAI22_X1 U5180 ( .A1(n5008), .A2(n4181), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4183), .ZN(n4188) );
  INV_X1 U5181 ( .A(n4265), .ZN(n4186) );
  NAND2_X1 U5182 ( .A1(n4184), .A2(n4183), .ZN(n4185) );
  NAND2_X1 U5183 ( .A1(n4186), .A2(n4185), .ZN(n5953) );
  AND2_X1 U5184 ( .A1(n5953), .A2(n5060), .ZN(n4187) );
  AOI21_X1 U5185 ( .B1(n4188), .B2(n5101), .A(n4187), .ZN(n4189) );
  NAND2_X1 U5186 ( .A1(n4192), .A2(n4191), .ZN(n4269) );
  CLKBUF_X1 U5187 ( .A(n4269), .Z(n4193) );
  OAI21_X1 U5188 ( .B1(n4028), .B2(n4192), .A(n4193), .ZN(n4245) );
  OAI222_X1 U5189 ( .A1(n4245), .A2(n5391), .B1(n4659), .B2(n6995), .C1(n6032), 
        .C2(n4181), .ZN(U2885) );
  OAI222_X1 U5190 ( .A1(n4393), .A2(n5391), .B1(n4659), .B2(n7170), .C1(n6032), 
        .C2(n3621), .ZN(U2890) );
  OAI222_X1 U5191 ( .A1(n5993), .A2(n5391), .B1(n4659), .B2(n6081), .C1(n5219), 
        .C2(n3524), .ZN(U2891) );
  NOR2_X1 U5192 ( .A1(n3935), .A2(n4194), .ZN(n4195) );
  NAND2_X1 U5193 ( .A1(n3933), .A2(n4195), .ZN(n6568) );
  INV_X1 U5194 ( .A(n6568), .ZN(n4196) );
  NAND2_X1 U5195 ( .A1(n4196), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6564) );
  NAND2_X1 U5196 ( .A1(n6564), .A2(n6427), .ZN(n6800) );
  INV_X1 U5197 ( .A(n6347), .ZN(n4197) );
  NAND2_X1 U5198 ( .A1(n6180), .A2(n4197), .ZN(n4198) );
  OAI21_X1 U5199 ( .B1(n6800), .B2(n4198), .A(n6812), .ZN(n4206) );
  OR2_X1 U5200 ( .A1(n6319), .A2(n4199), .ZN(n6254) );
  INV_X1 U5201 ( .A(n6254), .ZN(n4203) );
  INV_X1 U5202 ( .A(n6430), .ZN(n6814) );
  INV_X1 U5203 ( .A(n4200), .ZN(n4201) );
  NAND2_X1 U5204 ( .A1(n4201), .A2(n6810), .ZN(n4232) );
  INV_X1 U5205 ( .A(n4232), .ZN(n4202) );
  AOI21_X1 U5206 ( .B1(n4203), .B2(n6814), .A(n4202), .ZN(n4207) );
  INV_X1 U5207 ( .A(n4207), .ZN(n4205) );
  NAND3_X1 U5208 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6810), .A3(n6704), .ZN(n6250) );
  AOI21_X1 U5209 ( .B1(n6802), .B2(n6250), .A(n6284), .ZN(n4204) );
  OAI21_X1 U5210 ( .B1(n4206), .B2(n4205), .A(n4204), .ZN(n4231) );
  INV_X1 U5211 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6478) );
  OAI22_X1 U5212 ( .A1(n4207), .A2(n4206), .B1(n6478), .B2(n6250), .ZN(n4230)
         );
  AOI22_X1 U5213 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n4231), .B1(n6669), 
        .B2(n4230), .ZN(n4211) );
  INV_X1 U5214 ( .A(n6614), .ZN(n6673) );
  OAI22_X1 U5215 ( .A1(n6497), .A2(n4232), .B1(n6251), .B2(n6673), .ZN(n4209)
         );
  INV_X1 U5216 ( .A(n4209), .ZN(n4210) );
  OAI211_X1 U5217 ( .C1(n4236), .C2(n6617), .A(n4211), .B(n4210), .ZN(U3048)
         );
  AOI22_X1 U5218 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n4231), .B1(n6675), 
        .B2(n4230), .ZN(n4214) );
  OAI22_X1 U5219 ( .A1(n6501), .A2(n4232), .B1(n6251), .B2(n6679), .ZN(n4212)
         );
  INV_X1 U5220 ( .A(n4212), .ZN(n4213) );
  OAI211_X1 U5221 ( .C1(n4236), .C2(n6621), .A(n4214), .B(n4213), .ZN(U3049)
         );
  AOI22_X1 U5222 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n4231), .B1(n6681), 
        .B2(n4230), .ZN(n4217) );
  OAI22_X1 U5223 ( .A1(n6505), .A2(n4232), .B1(n6251), .B2(n6685), .ZN(n4215)
         );
  INV_X1 U5224 ( .A(n4215), .ZN(n4216) );
  OAI211_X1 U5225 ( .C1(n4236), .C2(n6625), .A(n4217), .B(n4216), .ZN(U3050)
         );
  AOI22_X1 U5226 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n4231), .B1(n6689), 
        .B2(n4230), .ZN(n4220) );
  OAI22_X1 U5227 ( .A1(n6510), .A2(n4232), .B1(n6251), .B2(n6696), .ZN(n4218)
         );
  INV_X1 U5228 ( .A(n4218), .ZN(n4219) );
  OAI211_X1 U5229 ( .C1(n4236), .C2(n6633), .A(n4220), .B(n4219), .ZN(U3051)
         );
  AOI22_X1 U5230 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n4231), .B1(n6639), 
        .B2(n4230), .ZN(n4223) );
  INV_X1 U5231 ( .A(n6598), .ZN(n6649) );
  OAI22_X1 U5232 ( .A1(n6471), .A2(n4232), .B1(n6251), .B2(n6649), .ZN(n4221)
         );
  INV_X1 U5233 ( .A(n4221), .ZN(n4222) );
  OAI211_X1 U5234 ( .C1(n6601), .C2(n4236), .A(n4223), .B(n4222), .ZN(U3044)
         );
  AOI22_X1 U5235 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n4231), .B1(n6651), 
        .B2(n4230), .ZN(n4226) );
  INV_X1 U5236 ( .A(n6602), .ZN(n6655) );
  OAI22_X1 U5237 ( .A1(n6485), .A2(n4232), .B1(n6251), .B2(n6655), .ZN(n4224)
         );
  INV_X1 U5238 ( .A(n4224), .ZN(n4225) );
  OAI211_X1 U5239 ( .C1(n4236), .C2(n6605), .A(n4226), .B(n4225), .ZN(U3045)
         );
  AOI22_X1 U5240 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n4231), .B1(n6657), 
        .B2(n4230), .ZN(n4229) );
  INV_X1 U5241 ( .A(n6606), .ZN(n6661) );
  OAI22_X1 U5242 ( .A1(n6489), .A2(n4232), .B1(n6251), .B2(n6661), .ZN(n4227)
         );
  INV_X1 U5243 ( .A(n4227), .ZN(n4228) );
  OAI211_X1 U5244 ( .C1(n4236), .C2(n6609), .A(n4229), .B(n4228), .ZN(U3046)
         );
  AOI22_X1 U5245 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n4231), .B1(n6663), 
        .B2(n4230), .ZN(n4235) );
  INV_X1 U5246 ( .A(n6610), .ZN(n6667) );
  OAI22_X1 U5247 ( .A1(n6493), .A2(n4232), .B1(n6251), .B2(n6667), .ZN(n4233)
         );
  INV_X1 U5248 ( .A(n4233), .ZN(n4234) );
  OAI211_X1 U5249 ( .C1(n4236), .C2(n6613), .A(n4235), .B(n4234), .ZN(U3047)
         );
  NAND2_X1 U5250 ( .A1(n4238), .A2(n4237), .ZN(n4241) );
  NAND2_X1 U5251 ( .A1(n4239), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4240)
         );
  NAND2_X1 U5252 ( .A1(n4241), .A2(n4240), .ZN(n4292) );
  XNOR2_X1 U5253 ( .A(n4288), .B(n4286), .ZN(n4242) );
  NAND2_X1 U5254 ( .A1(n4242), .A2(n5239), .ZN(n4243) );
  INV_X1 U5255 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4309) );
  XNOR2_X1 U5256 ( .A(n4293), .B(n4309), .ZN(n4291) );
  XNOR2_X1 U5257 ( .A(n3160), .B(n4291), .ZN(n4260) );
  INV_X1 U5258 ( .A(n4245), .ZN(n6020) );
  AOI22_X1 U5259 ( .A1(n6117), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .B1(n5969), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n4246) );
  OAI21_X1 U5260 ( .B1(n5953), .B2(n6111), .A(n4246), .ZN(n4247) );
  AOI21_X1 U5261 ( .B1(n6020), .B2(n6113), .A(n4247), .ZN(n4248) );
  OAI21_X1 U5262 ( .B1(n5835), .B2(n4260), .A(n4248), .ZN(U2980) );
  NAND2_X1 U5263 ( .A1(n5167), .A2(n4309), .ZN(n4250) );
  OAI211_X1 U5264 ( .C1(n5168), .C2(EBX_REG_6__SCAN_IN), .A(n4250), .B(n3174), 
        .ZN(n4251) );
  OAI21_X1 U5265 ( .B1(n5227), .B2(EBX_REG_6__SCAN_IN), .A(n4251), .ZN(n4276)
         );
  INV_X1 U5266 ( .A(n4277), .ZN(n4252) );
  XNOR2_X1 U5267 ( .A(n4276), .B(n4252), .ZN(n6017) );
  INV_X1 U5268 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6770) );
  NOR2_X1 U5269 ( .A1(n5819), .A2(n6770), .ZN(n4258) );
  INV_X1 U5271 ( .A(n4253), .ZN(n4308) );
  OAI33_X1 U5272 ( .A1(1'b0), .A2(n4255), .A3(n4309), .B1(
        INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n4308), .B3(n4254), .ZN(n4257) );
  AOI211_X1 U5273 ( .C1(n6172), .C2(n6017), .A(n4258), .B(n4257), .ZN(n4259)
         );
  OAI21_X1 U5274 ( .B1(n6125), .B2(n4260), .A(n4259), .ZN(U3012) );
  INV_X1 U5275 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4643) );
  NAND2_X1 U5276 ( .A1(n4261), .A2(n4298), .ZN(n4262) );
  OAI21_X1 U5277 ( .B1(n4643), .B2(n4263), .A(n4262), .ZN(n4264) );
  INV_X1 U5278 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4267) );
  OAI21_X1 U5279 ( .B1(n4265), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n4360), 
        .ZN(n5945) );
  AOI22_X1 U5280 ( .A1(n5945), .A2(n5060), .B1(n5210), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4266) );
  OAI21_X1 U5281 ( .B1(n5008), .B2(n4267), .A(n4266), .ZN(n4268) );
  INV_X1 U5282 ( .A(n4269), .ZN(n4271) );
  NAND2_X1 U5283 ( .A1(n4271), .A2(n4270), .ZN(n4469) );
  INV_X1 U5284 ( .A(n4272), .ZN(n4273) );
  AOI21_X1 U5285 ( .B1(n4274), .B2(n4193), .A(n4273), .ZN(n4328) );
  INV_X1 U5286 ( .A(n4328), .ZN(n5938) );
  OAI222_X1 U5287 ( .A1(n5938), .A2(n5391), .B1(n4659), .B2(n6991), .C1(n6032), 
        .C2(n4267), .ZN(U2884) );
  MUX2_X1 U5288 ( .A(n5170), .B(n3174), .S(EBX_REG_7__SCAN_IN), .Z(n4275) );
  OAI21_X1 U5289 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n5234), .A(n4275), 
        .ZN(n4279) );
  NAND2_X1 U5290 ( .A1(n4277), .A2(n4276), .ZN(n4278) );
  NOR2_X2 U5291 ( .A1(n4278), .A2(n4279), .ZN(n4315) );
  AOI21_X1 U5292 ( .B1(n4279), .B2(n4278), .A(n4315), .ZN(n6148) );
  INV_X1 U5293 ( .A(n6148), .ZN(n4280) );
  INV_X1 U5294 ( .A(EBX_REG_7__SCAN_IN), .ZN(n5936) );
  OAI222_X1 U5295 ( .A1(n4280), .A2(n6011), .B1(n5936), .B2(n6022), .C1(n5938), 
        .C2(n6012), .ZN(U2852) );
  INV_X1 U5296 ( .A(n4282), .ZN(n4284) );
  NOR2_X1 U5297 ( .A1(n4284), .A2(n4283), .ZN(n4285) );
  INV_X1 U5298 ( .A(n4286), .ZN(n4287) );
  OR2_X1 U5299 ( .A1(n4288), .A2(n4287), .ZN(n4299) );
  INV_X1 U5300 ( .A(n4299), .ZN(n4289) );
  NAND3_X1 U5301 ( .A1(n4289), .A2(n5239), .A3(n4298), .ZN(n4290) );
  NAND2_X1 U5302 ( .A1(n4664), .A2(n4290), .ZN(n4430) );
  INV_X1 U5303 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4318) );
  XNOR2_X1 U5304 ( .A(n4430), .B(n4318), .ZN(n4428) );
  NAND2_X1 U5305 ( .A1(n4292), .A2(n4291), .ZN(n4295) );
  NAND2_X1 U5306 ( .A1(n4293), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4294)
         );
  NAND2_X1 U5307 ( .A1(n4295), .A2(n4294), .ZN(n4323) );
  NAND2_X1 U5308 ( .A1(n4297), .A2(n4296), .ZN(n4302) );
  XNOR2_X1 U5309 ( .A(n4299), .B(n4298), .ZN(n4300) );
  NAND2_X1 U5310 ( .A1(n4300), .A2(n5239), .ZN(n4301) );
  NAND2_X1 U5311 ( .A1(n4302), .A2(n4301), .ZN(n4303) );
  INV_X1 U5312 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6155) );
  XNOR2_X1 U5313 ( .A(n4303), .B(n6155), .ZN(n4325) );
  NAND2_X1 U5314 ( .A1(n4323), .A2(n4325), .ZN(n4305) );
  NAND2_X1 U5315 ( .A1(n4303), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4304)
         );
  NAND2_X1 U5316 ( .A1(n4305), .A2(n4304), .ZN(n4429) );
  CLKBUF_X1 U5317 ( .A(n4429), .Z(n4306) );
  XNOR2_X1 U5318 ( .A(n4428), .B(n4306), .ZN(n4357) );
  NOR2_X1 U5319 ( .A1(n4309), .A2(n4307), .ZN(n5120) );
  INV_X1 U5320 ( .A(n5643), .ZN(n4310) );
  NOR4_X1 U5321 ( .A1(n3881), .A2(n3876), .A3(n4309), .A4(n4308), .ZN(n5121)
         );
  OAI22_X1 U5322 ( .A1(n5120), .A2(n5645), .B1(n4310), .B2(n5121), .ZN(n4311)
         );
  NOR2_X1 U5323 ( .A1(n5641), .A2(n4311), .ZN(n6156) );
  INV_X1 U5324 ( .A(n6156), .ZN(n4321) );
  NAND2_X1 U5325 ( .A1(n5167), .A2(n4318), .ZN(n4312) );
  OAI211_X1 U5326 ( .C1(n5168), .C2(EBX_REG_8__SCAN_IN), .A(n4312), .B(n3174), 
        .ZN(n4313) );
  OAI21_X1 U5327 ( .B1(n5227), .B2(EBX_REG_8__SCAN_IN), .A(n4313), .ZN(n4314)
         );
  OR2_X1 U5328 ( .A1(n4314), .A2(n4315), .ZN(n4316) );
  NAND2_X1 U5329 ( .A1(n4316), .A2(n4549), .ZN(n4350) );
  INV_X1 U5330 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6773) );
  OAI22_X1 U5331 ( .A1(n6163), .A2(n4350), .B1(n6773), .B2(n5819), .ZN(n4320)
         );
  NAND2_X1 U5332 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5119) );
  INV_X1 U5333 ( .A(n5119), .ZN(n4541) );
  NAND2_X1 U5334 ( .A1(n5120), .A2(n4317), .ZN(n6151) );
  AOI211_X1 U5335 ( .C1(n6155), .C2(n4318), .A(n4541), .B(n6151), .ZN(n4319)
         );
  AOI211_X1 U5336 ( .C1(INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n4321), .A(n4320), 
        .B(n4319), .ZN(n4322) );
  OAI21_X1 U5337 ( .B1(n6125), .B2(n4357), .A(n4322), .ZN(U3010) );
  CLKBUF_X1 U5338 ( .A(n4323), .Z(n4324) );
  XOR2_X1 U5339 ( .A(n4325), .B(n4324), .Z(n6153) );
  INV_X1 U5340 ( .A(n6153), .ZN(n4330) );
  NAND2_X1 U5341 ( .A1(n6176), .A2(REIP_REG_7__SCAN_IN), .ZN(n6149) );
  NAND2_X1 U5342 ( .A1(n6117), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4326)
         );
  OAI211_X1 U5343 ( .C1(n6111), .C2(n5945), .A(n6149), .B(n4326), .ZN(n4327)
         );
  AOI21_X1 U5344 ( .B1(n4328), .B2(n6113), .A(n4327), .ZN(n4329) );
  OAI21_X1 U5345 ( .B1(n4330), .B2(n5835), .A(n4329), .ZN(U2979) );
  AOI22_X1 U5346 ( .A1(n5076), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n5070), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4334) );
  AOI22_X1 U5347 ( .A1(n3538), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4333) );
  AOI22_X1 U5348 ( .A1(n5085), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4332) );
  AOI22_X1 U5349 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n5083), .B1(n3599), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4331) );
  NAND4_X1 U5350 ( .A1(n4334), .A2(n4333), .A3(n4332), .A4(n4331), .ZN(n4343)
         );
  AOI22_X1 U5351 ( .A1(n5081), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4882), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4341) );
  NAND2_X1 U5352 ( .A1(n5050), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4337)
         );
  NAND2_X1 U5353 ( .A1(n5082), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4336)
         );
  NAND2_X1 U5354 ( .A1(n5069), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4335) );
  AND3_X1 U5355 ( .A1(n4337), .A2(n4336), .A3(n4335), .ZN(n4340) );
  AOI22_X1 U5356 ( .A1(n3534), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4339) );
  OR2_X1 U5357 ( .A1(n5018), .A2(n4896), .ZN(n4338) );
  NAND4_X1 U5358 ( .A1(n4341), .A2(n4340), .A3(n4339), .A4(n4338), .ZN(n4342)
         );
  NOR2_X1 U5359 ( .A1(n4343), .A2(n4342), .ZN(n4345) );
  XNOR2_X1 U5360 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n4360), .ZN(n5926) );
  INV_X1 U5361 ( .A(n5926), .ZN(n4354) );
  AOI22_X1 U5362 ( .A1(n5210), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n5060), 
        .B2(n4354), .ZN(n4344) );
  OAI21_X1 U5363 ( .B1(n4599), .B2(n4345), .A(n4344), .ZN(n4348) );
  INV_X1 U5364 ( .A(EAX_REG_8__SCAN_IN), .ZN(n4346) );
  NOR2_X1 U5365 ( .A1(n5008), .A2(n4346), .ZN(n4347) );
  NOR2_X1 U5366 ( .A1(n4348), .A2(n4347), .ZN(n4513) );
  OR2_X1 U5367 ( .A1(n4272), .A2(n4513), .ZN(n4415) );
  NAND2_X1 U5368 ( .A1(n4272), .A2(n4513), .ZN(n4349) );
  AND2_X1 U5369 ( .A1(n4415), .A2(n4349), .ZN(n5927) );
  INV_X1 U5370 ( .A(n5927), .ZN(n4352) );
  INV_X1 U5371 ( .A(n4350), .ZN(n5921) );
  AOI22_X1 U5372 ( .A1(n6018), .A2(n5921), .B1(n5371), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n4351) );
  OAI21_X1 U5373 ( .B1(n4352), .B2(n6012), .A(n4351), .ZN(U2851) );
  INV_X1 U5374 ( .A(DATAI_8_), .ZN(n7196) );
  OAI222_X1 U5375 ( .A1(n4352), .A2(n5391), .B1(n4659), .B2(n7196), .C1(n5219), 
        .C2(n4346), .ZN(U2883) );
  AOI22_X1 U5376 ( .A1(n6117), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n5969), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n4353) );
  OAI21_X1 U5377 ( .B1(n6111), .B2(n4354), .A(n4353), .ZN(n4355) );
  AOI21_X1 U5378 ( .B1(n5927), .B2(n6113), .A(n4355), .ZN(n4356) );
  OAI21_X1 U5379 ( .B1(n4357), .B2(n5835), .A(n4356), .ZN(U2978) );
  OR2_X1 U5380 ( .A1(n6830), .A2(n3305), .ZN(n4372) );
  NAND3_X1 U5381 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), 
        .A3(n6747), .ZN(n6729) );
  NAND2_X1 U5382 ( .A1(n5060), .A2(n4358), .ZN(n6742) );
  AND3_X1 U5383 ( .A1(n5819), .A2(n6729), .A3(n6742), .ZN(n4359) );
  INV_X1 U5384 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4422) );
  INV_X1 U5385 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4362) );
  NAND2_X1 U5386 ( .A1(n4470), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4516)
         );
  INV_X1 U5387 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4363) );
  NAND2_X1 U5388 ( .A1(n4582), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4635)
         );
  INV_X1 U5389 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4364) );
  INV_X1 U5390 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4365) );
  INV_X1 U5391 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5459) );
  INV_X1 U5392 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4367) );
  INV_X1 U5393 ( .A(n4989), .ZN(n4368) );
  INV_X1 U5394 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5408) );
  NAND2_X1 U5395 ( .A1(n5040), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5100)
         );
  INV_X1 U5396 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5252) );
  INV_X1 U5397 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4369) );
  XNOR2_X1 U5398 ( .A(n4370), .B(n4369), .ZN(n5216) );
  NOR2_X1 U5399 ( .A1(n5216), .A2(n6728), .ZN(n4371) );
  INV_X1 U5400 ( .A(n4373), .ZN(n4374) );
  OR2_X1 U5401 ( .A1(n6830), .A2(n4374), .ZN(n5981) );
  OR2_X1 U5402 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4381) );
  NAND2_X1 U5403 ( .A1(EBX_REG_31__SCAN_IN), .A2(n4381), .ZN(n4375) );
  INV_X1 U5404 ( .A(n3640), .ZN(n4376) );
  OAI22_X1 U5405 ( .A1(n3940), .A2(n5981), .B1(n5992), .B2(n4376), .ZN(n4391)
         );
  AND2_X1 U5406 ( .A1(n5216), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4377) );
  INV_X1 U5407 ( .A(n5931), .ZN(n4378) );
  AOI22_X1 U5408 ( .A1(n5997), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n4378), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n4379) );
  OAI21_X1 U5409 ( .B1(n5988), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4379), 
        .ZN(n4390) );
  INV_X1 U5410 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4388) );
  NAND3_X1 U5411 ( .A1(n4380), .A2(n7199), .A3(n6912), .ZN(n6725) );
  INV_X1 U5412 ( .A(n4381), .ZN(n4384) );
  NOR2_X1 U5413 ( .A1(EBX_REG_31__SCAN_IN), .A2(n4384), .ZN(n4382) );
  AOI22_X1 U5414 ( .A1(n5239), .A2(n6725), .B1(n4382), .B2(n4385), .ZN(n4383)
         );
  NAND2_X1 U5415 ( .A1(n4385), .A2(n4384), .ZN(n4386) );
  OAI22_X1 U5416 ( .A1(n4388), .A2(n6000), .B1(n5934), .B2(REIP_REG_1__SCAN_IN), .ZN(n4389) );
  NOR3_X1 U5417 ( .A1(n4391), .A2(n4390), .A3(n4389), .ZN(n4392) );
  OAI21_X1 U5418 ( .B1(n4393), .B2(n5994), .A(n4392), .ZN(U2826) );
  INV_X1 U5419 ( .A(EAX_REG_9__SCAN_IN), .ZN(n4397) );
  INV_X1 U5420 ( .A(n4394), .ZN(n4395) );
  XNOR2_X1 U5421 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n4395), .ZN(n4426) );
  AOI22_X1 U5422 ( .A1(n5060), .A2(n4426), .B1(n5210), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4396) );
  OAI21_X1 U5423 ( .B1(n5008), .B2(n4397), .A(n4396), .ZN(n4414) );
  NAND2_X1 U5424 ( .A1(n5081), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4400) );
  NAND2_X1 U5425 ( .A1(n5075), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4399) );
  NAND2_X1 U5426 ( .A1(n5069), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4398) );
  AND3_X1 U5427 ( .A1(n4400), .A2(n4399), .A3(n4398), .ZN(n4405) );
  AOI22_X1 U5428 ( .A1(n3534), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4404) );
  AOI22_X1 U5429 ( .A1(n5070), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4882), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4403) );
  INV_X1 U5430 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4401) );
  OR2_X1 U5431 ( .A1(n5018), .A2(n4401), .ZN(n4402) );
  NAND4_X1 U5432 ( .A1(n4405), .A2(n4404), .A3(n4403), .A4(n4402), .ZN(n4411)
         );
  AOI22_X1 U5433 ( .A1(n5085), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n5026), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4409) );
  AOI22_X1 U5434 ( .A1(n5076), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n5083), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4408) );
  AOI22_X1 U5435 ( .A1(n5050), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3599), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4407) );
  AOI22_X1 U5436 ( .A1(n5082), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4406) );
  NAND4_X1 U5437 ( .A1(n4409), .A2(n4408), .A3(n4407), .A4(n4406), .ZN(n4410)
         );
  NOR2_X1 U5438 ( .A1(n4411), .A2(n4410), .ZN(n4412) );
  NOR2_X1 U5439 ( .A1(n4599), .A2(n4412), .ZN(n4413) );
  NOR2_X1 U5440 ( .A1(n4414), .A2(n4413), .ZN(n4510) );
  AOI21_X1 U5441 ( .B1(n4510), .B2(n4415), .A(n4457), .ZN(n4416) );
  INV_X1 U5442 ( .A(n4416), .ZN(n4437) );
  MUX2_X1 U5443 ( .A(n5170), .B(n3174), .S(EBX_REG_9__SCAN_IN), .Z(n4417) );
  OAI21_X1 U5444 ( .B1(n5234), .B2(INSTADDRPOINTER_REG_9__SCAN_IN), .A(n4417), 
        .ZN(n4546) );
  NOR2_X1 U5445 ( .A1(n4546), .A2(n4549), .ZN(n4550) );
  AOI21_X1 U5446 ( .B1(n4546), .B2(n4549), .A(n4550), .ZN(n6141) );
  AOI22_X1 U5447 ( .A1(n6018), .A2(n6141), .B1(n5371), .B2(EBX_REG_9__SCAN_IN), 
        .ZN(n4418) );
  OAI21_X1 U5448 ( .B1(n4437), .B2(n6012), .A(n4418), .ZN(U2850) );
  INV_X1 U5449 ( .A(n4426), .ZN(n4424) );
  INV_X1 U5450 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6766) );
  INV_X1 U5451 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6765) );
  NOR3_X1 U5452 ( .A1(n3739), .A2(n6766), .A3(n6765), .ZN(n5972) );
  NAND2_X1 U5453 ( .A1(REIP_REG_4__SCAN_IN), .A2(n5972), .ZN(n5933) );
  NOR2_X1 U5454 ( .A1(n6768), .A2(n5933), .ZN(n5932) );
  NAND3_X1 U5455 ( .A1(n5932), .A2(REIP_REG_7__SCAN_IN), .A3(
        REIP_REG_6__SCAN_IN), .ZN(n5923) );
  NOR2_X1 U5456 ( .A1(n6773), .A2(n5923), .ZN(n4567) );
  INV_X1 U5457 ( .A(n4567), .ZN(n4419) );
  NAND2_X1 U5458 ( .A1(n5977), .A2(n4419), .ZN(n5922) );
  NAND2_X1 U5459 ( .A1(n5922), .A2(n5931), .ZN(n5920) );
  AOI22_X1 U5460 ( .A1(n5965), .A2(n6141), .B1(REIP_REG_9__SCAN_IN), .B2(n5920), .ZN(n4421) );
  INV_X1 U5461 ( .A(n5819), .ZN(n5969) );
  OR2_X1 U5462 ( .A1(n5934), .A2(n4419), .ZN(n5914) );
  NOR2_X1 U5463 ( .A1(REIP_REG_9__SCAN_IN), .A2(n5914), .ZN(n5913) );
  AOI211_X1 U5464 ( .C1(n5980), .C2(EBX_REG_9__SCAN_IN), .A(n5969), .B(n5913), 
        .ZN(n4420) );
  OAI211_X1 U5465 ( .C1(n4422), .C2(n5872), .A(n4421), .B(n4420), .ZN(n4423)
         );
  AOI21_X1 U5466 ( .B1(n5996), .B2(n4424), .A(n4423), .ZN(n4425) );
  OAI21_X1 U5467 ( .B1(n4437), .B2(n5937), .A(n4425), .ZN(U2818) );
  INV_X1 U5468 ( .A(DATAI_9_), .ZN(n6091) );
  OAI222_X1 U5469 ( .A1(n4437), .A2(n5391), .B1(n4659), .B2(n6091), .C1(n5219), 
        .C2(n4397), .ZN(U2882) );
  AND2_X1 U5470 ( .A1(n5969), .A2(REIP_REG_9__SCAN_IN), .ZN(n6140) );
  NOR2_X1 U5471 ( .A1(n6111), .A2(n4426), .ZN(n4427) );
  AOI211_X1 U5472 ( .C1(n6117), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6140), 
        .B(n4427), .ZN(n4436) );
  NAND2_X1 U5473 ( .A1(n4429), .A2(n4428), .ZN(n4432) );
  NAND2_X1 U5474 ( .A1(n4430), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4431)
         );
  NAND2_X1 U5475 ( .A1(n4432), .A2(n4431), .ZN(n4533) );
  CLKBUF_X1 U5476 ( .A(n4533), .Z(n4433) );
  INV_X1 U5477 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6146) );
  XNOR2_X1 U5478 ( .A(n5432), .B(n6146), .ZN(n4434) );
  XNOR2_X1 U5479 ( .A(n4433), .B(n4434), .ZN(n6143) );
  NAND2_X1 U5480 ( .A1(n6143), .A2(n6115), .ZN(n4435) );
  OAI211_X1 U5481 ( .C1(n4437), .C2(n5512), .A(n4436), .B(n4435), .ZN(U2977)
         );
  XOR2_X1 U5482 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n4438), .Z(n5911) );
  AOI22_X1 U5483 ( .A1(n5070), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4442) );
  AOI22_X1 U5484 ( .A1(n3534), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n5081), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4441) );
  AOI22_X1 U5485 ( .A1(n5076), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4440) );
  AOI22_X1 U5486 ( .A1(n5083), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3599), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4439) );
  NAND4_X1 U5487 ( .A1(n4442), .A2(n4441), .A3(n4440), .A4(n4439), .ZN(n4451)
         );
  AOI22_X1 U5488 ( .A1(n5085), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n5050), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4449) );
  NAND2_X1 U5489 ( .A1(n4882), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4445) );
  NAND2_X1 U5490 ( .A1(n5082), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4444)
         );
  NAND2_X1 U5491 ( .A1(n5069), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4443) );
  AND3_X1 U5492 ( .A1(n4445), .A2(n4444), .A3(n4443), .ZN(n4448) );
  AOI22_X1 U5493 ( .A1(n5026), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4447) );
  INV_X1 U5494 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4948) );
  OR2_X1 U5495 ( .A1(n5018), .A2(n4948), .ZN(n4446) );
  NAND4_X1 U5496 ( .A1(n4449), .A2(n4448), .A3(n4447), .A4(n4446), .ZN(n4450)
         );
  NOR2_X1 U5497 ( .A1(n4451), .A2(n4450), .ZN(n4452) );
  INV_X1 U5498 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4630) );
  OAI22_X1 U5499 ( .A1(n4599), .A2(n4452), .B1(n4710), .B2(n4630), .ZN(n4455)
         );
  INV_X1 U5500 ( .A(EAX_REG_10__SCAN_IN), .ZN(n4453) );
  NOR2_X1 U5501 ( .A1(n5008), .A2(n4453), .ZN(n4454) );
  NOR2_X1 U5502 ( .A1(n4455), .A2(n4454), .ZN(n4456) );
  OAI21_X1 U5503 ( .B1(n5911), .B2(n5101), .A(n4456), .ZN(n4508) );
  NOR2_X1 U5504 ( .A1(n4457), .A2(n4508), .ZN(n4458) );
  INV_X1 U5505 ( .A(DATAI_10_), .ZN(n6921) );
  OAI222_X1 U5506 ( .A1(n5910), .A2(n5391), .B1(n4659), .B2(n6921), .C1(n5219), 
        .C2(n4453), .ZN(U2881) );
  INV_X1 U5507 ( .A(n4459), .ZN(n4460) );
  OAI22_X1 U5508 ( .A1(n6804), .A2(n5981), .B1(n5992), .B2(n4460), .ZN(n4464)
         );
  INV_X1 U5509 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4462) );
  OAI22_X1 U5510 ( .A1(n4462), .A2(n5872), .B1(n5988), .B2(n4461), .ZN(n4463)
         );
  AOI211_X1 U5511 ( .C1(n5980), .C2(EBX_REG_3__SCAN_IN), .A(n4464), .B(n4463), 
        .ZN(n4467) );
  NAND2_X1 U5512 ( .A1(n5934), .A2(n5931), .ZN(n5989) );
  INV_X1 U5513 ( .A(n5989), .ZN(n5303) );
  AOI21_X1 U5514 ( .B1(n5931), .B2(REIP_REG_1__SCAN_IN), .A(n5303), .ZN(n4465)
         );
  NOR2_X1 U5515 ( .A1(n4465), .A2(n6765), .ZN(n5979) );
  OAI21_X1 U5516 ( .B1(n5934), .B2(n5972), .A(n5931), .ZN(n5963) );
  OAI21_X1 U5517 ( .B1(n5979), .B2(REIP_REG_3__SCAN_IN), .A(n5963), .ZN(n4466)
         );
  OAI211_X1 U5518 ( .C1(n4468), .C2(n5994), .A(n4467), .B(n4466), .ZN(U2824)
         );
  INV_X1 U5519 ( .A(n4469), .ZN(n4515) );
  XOR2_X1 U5520 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n4470), .Z(n5902) );
  NAND2_X1 U5521 ( .A1(n5050), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4473)
         );
  NAND2_X1 U5522 ( .A1(n5083), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4472)
         );
  NAND2_X1 U5523 ( .A1(n5069), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4471) );
  AND3_X1 U5524 ( .A1(n4473), .A2(n4472), .A3(n4471), .ZN(n4478) );
  AOI22_X1 U5525 ( .A1(n5085), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3534), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4477) );
  AOI22_X1 U5526 ( .A1(n5076), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4476) );
  OR2_X1 U5527 ( .A1(n5018), .A2(n4474), .ZN(n4475) );
  NAND4_X1 U5528 ( .A1(n4478), .A2(n4477), .A3(n4476), .A4(n4475), .ZN(n4484)
         );
  AOI22_X1 U5529 ( .A1(n5026), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4482) );
  AOI22_X1 U5530 ( .A1(n5070), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4882), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4481) );
  AOI22_X1 U5531 ( .A1(n5080), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3599), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4480) );
  AOI22_X1 U5532 ( .A1(n5081), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n5082), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4479) );
  NAND4_X1 U5533 ( .A1(n4482), .A2(n4481), .A3(n4480), .A4(n4479), .ZN(n4483)
         );
  NOR2_X1 U5534 ( .A1(n4484), .A2(n4483), .ZN(n4485) );
  INV_X1 U5535 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4682) );
  OAI22_X1 U5536 ( .A1(n4599), .A2(n4485), .B1(n4710), .B2(n4682), .ZN(n4488)
         );
  INV_X1 U5537 ( .A(EAX_REG_12__SCAN_IN), .ZN(n4486) );
  NOR2_X1 U5538 ( .A1(n5008), .A2(n4486), .ZN(n4487) );
  NOR2_X1 U5539 ( .A1(n4488), .A2(n4487), .ZN(n4489) );
  OAI21_X1 U5540 ( .B1(n5902), .B2(n5101), .A(n4489), .ZN(n4556) );
  NAND2_X1 U5541 ( .A1(n5075), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4492) );
  NAND2_X1 U5542 ( .A1(n5070), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4491) );
  NAND2_X1 U5543 ( .A1(n5069), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4490) );
  AND3_X1 U5544 ( .A1(n4492), .A2(n4491), .A3(n4490), .ZN(n4497) );
  AOI22_X1 U5545 ( .A1(n5026), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4882), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4496) );
  AOI22_X1 U5546 ( .A1(n5050), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3599), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4495) );
  INV_X1 U5547 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4493) );
  OR2_X1 U5548 ( .A1(n5018), .A2(n4493), .ZN(n4494) );
  NAND4_X1 U5549 ( .A1(n4497), .A2(n4496), .A3(n4495), .A4(n4494), .ZN(n4503)
         );
  AOI22_X1 U5550 ( .A1(n5085), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n5081), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4501) );
  AOI22_X1 U5551 ( .A1(n5076), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4500) );
  AOI22_X1 U5552 ( .A1(n3534), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4499) );
  AOI22_X1 U5553 ( .A1(n5083), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n5082), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4498) );
  NAND4_X1 U5554 ( .A1(n4501), .A2(n4500), .A3(n4499), .A4(n4498), .ZN(n4502)
         );
  NOR2_X1 U5555 ( .A1(n4503), .A2(n4502), .ZN(n4507) );
  XNOR2_X1 U5556 ( .A(n4504), .B(n4362), .ZN(n4667) );
  NAND2_X1 U5557 ( .A1(n4667), .A2(n5060), .ZN(n4506) );
  AOI22_X1 U5558 ( .A1(n5211), .A2(EAX_REG_11__SCAN_IN), .B1(n5210), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4505) );
  OAI211_X1 U5559 ( .C1(n4507), .C2(n4599), .A(n4506), .B(n4505), .ZN(n4557)
         );
  AND2_X1 U5560 ( .A1(n4556), .A2(n4557), .ZN(n4509) );
  NAND2_X1 U5561 ( .A1(n4509), .A2(n4508), .ZN(n4511) );
  NAND2_X1 U5562 ( .A1(n4515), .A2(n4514), .ZN(n4555) );
  XNOR2_X1 U5563 ( .A(n4516), .B(n4363), .ZN(n5891) );
  INV_X1 U5564 ( .A(EAX_REG_13__SCAN_IN), .ZN(n4517) );
  OAI22_X1 U5565 ( .A1(n5008), .A2(n4517), .B1(n4710), .B2(n4363), .ZN(n4518)
         );
  AOI21_X1 U5566 ( .B1(n5891), .B2(n5060), .A(n4518), .ZN(n4576) );
  XNOR2_X1 U5567 ( .A(n4555), .B(n4576), .ZN(n4580) );
  AOI22_X1 U5568 ( .A1(n5076), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4522) );
  AOI22_X1 U5569 ( .A1(n5070), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n5082), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4521) );
  AOI22_X1 U5570 ( .A1(n5026), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3599), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4520) );
  AOI22_X1 U5571 ( .A1(n5081), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4519) );
  NAND4_X1 U5572 ( .A1(n4522), .A2(n4521), .A3(n4520), .A4(n4519), .ZN(n4532)
         );
  NAND2_X1 U5573 ( .A1(n5050), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4525)
         );
  NAND2_X1 U5574 ( .A1(n5083), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4524)
         );
  NAND2_X1 U5575 ( .A1(n5069), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4523) );
  AND3_X1 U5576 ( .A1(n4525), .A2(n4524), .A3(n4523), .ZN(n4530) );
  AOI22_X1 U5577 ( .A1(n5085), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4529) );
  AOI22_X1 U5578 ( .A1(n3534), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4882), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4528) );
  INV_X1 U5579 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4526) );
  OR2_X1 U5580 ( .A1(n5018), .A2(n4526), .ZN(n4527) );
  NAND4_X1 U5581 ( .A1(n4530), .A2(n4529), .A3(n4528), .A4(n4527), .ZN(n4531)
         );
  OAI21_X1 U5582 ( .B1(n4532), .B2(n4531), .A(n4648), .ZN(n4581) );
  XNOR2_X1 U5583 ( .A(n4580), .B(n4581), .ZN(n6013) );
  INV_X1 U5584 ( .A(DATAI_13_), .ZN(n6993) );
  OAI222_X1 U5585 ( .A1(n5391), .A2(n6013), .B1(n4659), .B2(n6993), .C1(n5219), 
        .C2(n4517), .ZN(U2878) );
  INV_X1 U5586 ( .A(n4533), .ZN(n4534) );
  NAND2_X1 U5587 ( .A1(n4534), .A2(n3175), .ZN(n4536) );
  NAND2_X1 U5588 ( .A1(n3150), .A2(n6146), .ZN(n4535) );
  NAND2_X1 U5589 ( .A1(n4536), .A2(n4535), .ZN(n4662) );
  CLKBUF_X1 U5590 ( .A(n4662), .Z(n4537) );
  INV_X1 U5591 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4538) );
  INV_X1 U5592 ( .A(n4661), .ZN(n4539) );
  NAND2_X1 U5593 ( .A1(n4539), .A2(n4660), .ZN(n4540) );
  XNOR2_X1 U5594 ( .A(n4537), .B(n4540), .ZN(n4634) );
  NOR2_X1 U5595 ( .A1(n5119), .A2(n6151), .ZN(n6142) );
  NAND2_X1 U5596 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5118) );
  OAI211_X1 U5597 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6142), .B(n5118), .ZN(n4554) );
  INV_X1 U5598 ( .A(n6170), .ZN(n5598) );
  OAI21_X1 U5599 ( .B1(n4541), .B2(n5598), .A(n6156), .ZN(n6139) );
  INV_X1 U5600 ( .A(EBX_REG_10__SCAN_IN), .ZN(n4542) );
  NAND2_X1 U5601 ( .A1(n5171), .A2(n4542), .ZN(n4545) );
  OR2_X1 U5602 ( .A1(n5167), .A2(n4542), .ZN(n4544) );
  NAND2_X1 U5603 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n5168), .ZN(n4543) );
  NAND4_X1 U5604 ( .A1(n4545), .A2(n5157), .A3(n4544), .A4(n4543), .ZN(n4551)
         );
  INV_X1 U5605 ( .A(n4551), .ZN(n4547) );
  OAI21_X1 U5606 ( .B1(n4551), .B2(n4550), .A(n4564), .ZN(n5908) );
  INV_X1 U5607 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6775) );
  OAI22_X1 U5608 ( .A1(n6163), .A2(n5908), .B1(n6775), .B2(n5819), .ZN(n4552)
         );
  AOI21_X1 U5609 ( .B1(n6139), .B2(INSTADDRPOINTER_REG_10__SCAN_IN), .A(n4552), 
        .ZN(n4553) );
  OAI211_X1 U5610 ( .C1(n4634), .C2(n6125), .A(n4554), .B(n4553), .ZN(U3008)
         );
  OAI21_X1 U5611 ( .B1(n4560), .B2(n4556), .A(n4555), .ZN(n5901) );
  INV_X1 U5612 ( .A(DATAI_12_), .ZN(n7186) );
  OAI222_X1 U5613 ( .A1(n5901), .A2(n5391), .B1(n4659), .B2(n7186), .C1(n6032), 
        .C2(n4486), .ZN(U2879) );
  OAI222_X1 U5614 ( .A1(n5908), .A2(n6011), .B1(n6022), .B2(n4542), .C1(n6012), 
        .C2(n5910), .ZN(U2849) );
  NOR2_X1 U5615 ( .A1(n4558), .A2(n4557), .ZN(n4559) );
  INV_X1 U5616 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4665) );
  INV_X1 U5617 ( .A(EBX_REG_11__SCAN_IN), .ZN(n4561) );
  NAND2_X1 U5618 ( .A1(n5178), .A2(n4561), .ZN(n4562) );
  OAI211_X1 U5619 ( .C1(n3475), .C2(n4665), .A(n4562), .B(n5167), .ZN(n4563)
         );
  OAI21_X1 U5620 ( .B1(EBX_REG_11__SCAN_IN), .B2(n5170), .A(n4563), .ZN(n4565)
         );
  AOI21_X1 U5621 ( .B1(n4565), .B2(n4564), .A(n4627), .ZN(n6133) );
  AOI22_X1 U5622 ( .A1(n6018), .A2(n6133), .B1(n5371), .B2(EBX_REG_11__SCAN_IN), .ZN(n4566) );
  OAI21_X1 U5623 ( .B1(n4672), .B2(n6012), .A(n4566), .ZN(U2848) );
  INV_X1 U5624 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6776) );
  NAND3_X1 U5625 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .A3(
        n4567), .ZN(n4572) );
  NOR2_X1 U5626 ( .A1(n6776), .A2(n4572), .ZN(n4607) );
  INV_X1 U5627 ( .A(n4607), .ZN(n4568) );
  NAND2_X1 U5628 ( .A1(n5977), .A2(n4568), .ZN(n4571) );
  NAND2_X1 U5629 ( .A1(n4571), .A2(n5931), .ZN(n5898) );
  INV_X1 U5630 ( .A(n6133), .ZN(n4569) );
  OAI22_X1 U5631 ( .A1(n5988), .A2(n4667), .B1(n5992), .B2(n4569), .ZN(n4574)
         );
  AOI22_X1 U5632 ( .A1(EBX_REG_11__SCAN_IN), .A2(n5980), .B1(
        PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n5997), .ZN(n4570) );
  OAI211_X1 U5633 ( .C1(n4572), .C2(n4571), .A(n4570), .B(n5819), .ZN(n4573)
         );
  AOI211_X1 U5634 ( .C1(REIP_REG_11__SCAN_IN), .C2(n5898), .A(n4574), .B(n4573), .ZN(n4575) );
  OAI21_X1 U5635 ( .B1(n4672), .B2(n5937), .A(n4575), .ZN(U2816) );
  INV_X1 U5636 ( .A(n4576), .ZN(n4577) );
  OAI21_X2 U5637 ( .B1(n4581), .B2(n4580), .A(n4579), .ZN(n4604) );
  XNOR2_X1 U5638 ( .A(n4582), .B(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5507)
         );
  NAND2_X1 U5639 ( .A1(n5507), .A2(n5060), .ZN(n4603) );
  INV_X1 U5640 ( .A(EAX_REG_14__SCAN_IN), .ZN(n4583) );
  INV_X1 U5641 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4619) );
  OAI22_X1 U5642 ( .A1(n5008), .A2(n4583), .B1(n4710), .B2(n4619), .ZN(n4601)
         );
  AOI22_X1 U5643 ( .A1(n5076), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4587) );
  AOI22_X1 U5644 ( .A1(n5085), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4586) );
  AOI22_X1 U5645 ( .A1(n5081), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n5083), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4585) );
  AOI22_X1 U5646 ( .A1(n5069), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4584) );
  NAND4_X1 U5647 ( .A1(n4587), .A2(n4586), .A3(n4585), .A4(n4584), .ZN(n4597)
         );
  NAND2_X1 U5648 ( .A1(n5050), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4590)
         );
  NAND2_X1 U5649 ( .A1(n5070), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4589) );
  NAND2_X1 U5650 ( .A1(n5082), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4588)
         );
  AND3_X1 U5651 ( .A1(n4590), .A2(n4589), .A3(n4588), .ZN(n4595) );
  AOI22_X1 U5652 ( .A1(n3538), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4882), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4594) );
  AOI22_X1 U5653 ( .A1(n3534), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3599), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4593) );
  OR2_X1 U5654 ( .A1(n5018), .A2(n4591), .ZN(n4592) );
  NAND4_X1 U5655 ( .A1(n4595), .A2(n4594), .A3(n4593), .A4(n4592), .ZN(n4596)
         );
  NOR2_X1 U5656 ( .A1(n4597), .A2(n4596), .ZN(n4598) );
  NOR2_X1 U5657 ( .A1(n4599), .A2(n4598), .ZN(n4600) );
  NOR2_X1 U5658 ( .A1(n4601), .A2(n4600), .ZN(n4602) );
  NAND2_X1 U5659 ( .A1(n4603), .A2(n4602), .ZN(n4605) );
  NAND2_X1 U5660 ( .A1(n4604), .A2(n4605), .ZN(n4656) );
  OAI21_X1 U5661 ( .B1(n4604), .B2(n4605), .A(n4656), .ZN(n5511) );
  NAND2_X1 U5662 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .ZN(
        n4606) );
  NAND2_X1 U5663 ( .A1(n5977), .A2(n4607), .ZN(n5893) );
  INV_X1 U5664 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6778) );
  OAI21_X1 U5665 ( .B1(n4606), .B2(n5893), .A(n6778), .ZN(n4625) );
  NAND4_X1 U5666 ( .A1(REIP_REG_14__SCAN_IN), .A2(n4607), .A3(
        REIP_REG_13__SCAN_IN), .A4(REIP_REG_12__SCAN_IN), .ZN(n5868) );
  INV_X1 U5667 ( .A(n5868), .ZN(n4608) );
  OAI21_X1 U5668 ( .B1(n5934), .B2(n4608), .A(n5931), .ZN(n5880) );
  INV_X1 U5669 ( .A(EBX_REG_14__SCAN_IN), .ZN(n4623) );
  INV_X1 U5670 ( .A(n5507), .ZN(n4621) );
  NAND2_X1 U5671 ( .A1(n5171), .A2(n4623), .ZN(n4611) );
  OR2_X1 U5672 ( .A1(n5167), .A2(n4623), .ZN(n4610) );
  NAND2_X1 U5673 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5168), .ZN(n4609) );
  NAND4_X1 U5674 ( .A1(n4611), .A2(n5157), .A3(n4610), .A4(n4609), .ZN(n4618)
         );
  INV_X1 U5675 ( .A(EBX_REG_12__SCAN_IN), .ZN(n4629) );
  NAND2_X1 U5676 ( .A1(n5171), .A2(n4629), .ZN(n4614) );
  OR2_X1 U5677 ( .A1(n5167), .A2(n4629), .ZN(n4613) );
  NAND2_X1 U5678 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n5168), .ZN(n4612) );
  NAND4_X1 U5679 ( .A1(n4614), .A2(n5157), .A3(n4613), .A4(n4612), .ZN(n4628)
         );
  OR2_X1 U5680 ( .A1(n5170), .A2(EBX_REG_13__SCAN_IN), .ZN(n4617) );
  NAND2_X1 U5681 ( .A1(n3174), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4615) );
  OAI211_X1 U5682 ( .C1(n5168), .C2(EBX_REG_13__SCAN_IN), .A(n5167), .B(n4615), 
        .ZN(n4616) );
  NAND2_X1 U5683 ( .A1(n4617), .A2(n4616), .ZN(n5818) );
  NOR2_X4 U5684 ( .A1(n5817), .A2(n5818), .ZN(n5816) );
  NAND2_X2 U5685 ( .A1(n5816), .A2(n4618), .ZN(n5806) );
  OAI21_X1 U5686 ( .B1(n4618), .B2(n5816), .A(n5806), .ZN(n5655) );
  OAI22_X1 U5687 ( .A1(n4619), .A2(n5872), .B1(n5992), .B2(n5655), .ZN(n4620)
         );
  AOI211_X1 U5688 ( .C1(n5996), .C2(n4621), .A(n4620), .B(n5969), .ZN(n4622)
         );
  OAI21_X1 U5689 ( .B1(n6000), .B2(n4623), .A(n4622), .ZN(n4624) );
  AOI21_X1 U5690 ( .B1(n4625), .B2(n5880), .A(n4624), .ZN(n4626) );
  OAI21_X1 U5691 ( .B1(n5511), .B2(n5937), .A(n4626), .ZN(U2813) );
  INV_X1 U5692 ( .A(DATAI_11_), .ZN(n7040) );
  INV_X1 U5693 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6044) );
  OAI222_X1 U5694 ( .A1(n4672), .A2(n5391), .B1(n4659), .B2(n7040), .C1(n6032), 
        .C2(n6044), .ZN(U2880) );
  OAI21_X1 U5695 ( .B1(n4628), .B2(n4627), .A(n5817), .ZN(n6124) );
  OAI222_X1 U5696 ( .A1(n6124), .A2(n6011), .B1(n4629), .B2(n6022), .C1(n6012), 
        .C2(n5901), .ZN(U2847) );
  INV_X1 U5697 ( .A(DATAI_14_), .ZN(n6099) );
  OAI222_X1 U5698 ( .A1(n5511), .A2(n5391), .B1(n4659), .B2(n6099), .C1(n6032), 
        .C2(n4583), .ZN(U2877) );
  OAI222_X1 U5699 ( .A1(n5655), .A2(n6011), .B1(n6022), .B2(n4623), .C1(n6012), 
        .C2(n5511), .ZN(U2845) );
  OAI22_X1 U5700 ( .A1(n5786), .A2(n4630), .B1(n5819), .B2(n6775), .ZN(n4632)
         );
  NOR2_X1 U5701 ( .A1(n5910), .A2(n5512), .ZN(n4631) );
  AOI211_X1 U5702 ( .C1(n5781), .C2(n5911), .A(n4632), .B(n4631), .ZN(n4633)
         );
  OAI21_X1 U5703 ( .B1(n5835), .B2(n4634), .A(n4633), .ZN(U2976) );
  XNOR2_X1 U5704 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n4635), .ZN(n5886)
         );
  INV_X1 U5705 ( .A(n5886), .ZN(n5501) );
  AOI22_X1 U5706 ( .A1(n5081), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4639) );
  AOI22_X1 U5707 ( .A1(n5050), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4638) );
  AOI22_X1 U5708 ( .A1(n5070), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n5083), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4637) );
  AOI22_X1 U5709 ( .A1(n5085), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4882), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4636) );
  NAND4_X1 U5710 ( .A1(n4639), .A2(n4638), .A3(n4637), .A4(n4636), .ZN(n4650)
         );
  AOI22_X1 U5711 ( .A1(n3534), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3538), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4647) );
  AOI22_X1 U5712 ( .A1(n5076), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3599), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4646) );
  NAND2_X1 U5713 ( .A1(n5082), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4642)
         );
  NAND2_X1 U5714 ( .A1(n5069), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4641) );
  NAND2_X1 U5715 ( .A1(n5086), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4640) );
  AND3_X1 U5716 ( .A1(n4642), .A2(n4641), .A3(n4640), .ZN(n4645) );
  OR2_X1 U5717 ( .A1(n5018), .A2(n4643), .ZN(n4644) );
  NAND4_X1 U5718 ( .A1(n4647), .A2(n4646), .A3(n4645), .A4(n4644), .ZN(n4649)
         );
  OAI21_X1 U5719 ( .B1(n4650), .B2(n4649), .A(n4648), .ZN(n4653) );
  NAND2_X1 U5720 ( .A1(n5211), .A2(EAX_REG_15__SCAN_IN), .ZN(n4652) );
  NAND2_X1 U5721 ( .A1(n5210), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4651)
         );
  NAND3_X1 U5722 ( .A1(n4653), .A2(n4652), .A3(n4651), .ZN(n4654) );
  AOI21_X1 U5723 ( .B1(n5501), .B2(n5060), .A(n4654), .ZN(n4655) );
  AND2_X1 U5724 ( .A1(n4656), .A2(n4655), .ZN(n4658) );
  OR2_X1 U5725 ( .A1(n4658), .A2(n4657), .ZN(n6006) );
  INV_X1 U5726 ( .A(DATAI_15_), .ZN(n7028) );
  INV_X1 U5727 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6039) );
  OAI222_X1 U5728 ( .A1(n6006), .A2(n5391), .B1(n4659), .B2(n7028), .C1(n6032), 
        .C2(n6039), .ZN(U2876) );
  OAI21_X2 U5729 ( .B1(n4662), .B2(n4661), .A(n4660), .ZN(n4674) );
  CLKBUF_X1 U5730 ( .A(n4674), .Z(n4663) );
  NAND2_X1 U5731 ( .A1(n5432), .A2(n4665), .ZN(n4673) );
  NAND2_X1 U5732 ( .A1(n4675), .A2(n4673), .ZN(n4666) );
  XNOR2_X1 U5733 ( .A(n4663), .B(n4666), .ZN(n6135) );
  NAND2_X1 U5734 ( .A1(n6135), .A2(n6115), .ZN(n4671) );
  INV_X1 U5735 ( .A(n4667), .ZN(n4669) );
  NAND2_X1 U5736 ( .A1(n6176), .A2(REIP_REG_11__SCAN_IN), .ZN(n6131) );
  OAI21_X1 U5737 ( .B1(n5786), .B2(n4362), .A(n6131), .ZN(n4668) );
  AOI21_X1 U5738 ( .B1(n5781), .B2(n4669), .A(n4668), .ZN(n4670) );
  OAI211_X1 U5739 ( .C1(n5512), .C2(n4672), .A(n4671), .B(n4670), .ZN(U2975)
         );
  NAND2_X1 U5740 ( .A1(n4674), .A2(n4673), .ZN(n4676) );
  NAND2_X1 U5741 ( .A1(n4676), .A2(n4675), .ZN(n4779) );
  INV_X1 U5742 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4678) );
  NAND2_X1 U5743 ( .A1(n5432), .A2(n4678), .ZN(n4777) );
  INV_X1 U5744 ( .A(n4777), .ZN(n4679) );
  NOR2_X1 U5745 ( .A1(n4778), .A2(n4679), .ZN(n4680) );
  XNOR2_X1 U5746 ( .A(n4677), .B(n4680), .ZN(n6126) );
  INV_X1 U5747 ( .A(REIP_REG_12__SCAN_IN), .ZN(n4681) );
  OAI22_X1 U5748 ( .A1(n5786), .A2(n4682), .B1(n5819), .B2(n4681), .ZN(n4684)
         );
  NOR2_X1 U5749 ( .A1(n5901), .A2(n5512), .ZN(n4683) );
  AOI211_X1 U5750 ( .C1(n5781), .C2(n5902), .A(n4684), .B(n4683), .ZN(n4685)
         );
  OAI21_X1 U5751 ( .B1(n6126), .B2(n5835), .A(n4685), .ZN(U2974) );
  INV_X1 U5752 ( .A(EBX_REG_16__SCAN_IN), .ZN(n4686) );
  NAND2_X1 U5753 ( .A1(n5171), .A2(n4686), .ZN(n4689) );
  OR2_X1 U5754 ( .A1(n5167), .A2(n4686), .ZN(n4688) );
  NAND2_X1 U5755 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n5168), .ZN(n4687) );
  NAND4_X1 U5756 ( .A1(n4689), .A2(n5157), .A3(n4688), .A4(n4687), .ZN(n4693)
         );
  OR2_X1 U5757 ( .A1(n5170), .A2(EBX_REG_15__SCAN_IN), .ZN(n4692) );
  NAND2_X1 U5758 ( .A1(n3174), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4690) );
  OAI211_X1 U5759 ( .C1(n5168), .C2(EBX_REG_15__SCAN_IN), .A(n5167), .B(n4690), 
        .ZN(n4691) );
  NAND2_X1 U5760 ( .A1(n4692), .A2(n4691), .ZN(n5807) );
  NOR2_X4 U5761 ( .A1(n5806), .A2(n5807), .ZN(n5805) );
  OAI21_X1 U5762 ( .B1(n4693), .B2(n5805), .A(n5630), .ZN(n5879) );
  XNOR2_X1 U5763 ( .A(n4694), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5875)
         );
  NAND2_X1 U5764 ( .A1(n5875), .A2(n5060), .ZN(n4714) );
  NAND2_X1 U5765 ( .A1(n5075), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4698) );
  NAND2_X1 U5766 ( .A1(n5076), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4697) );
  NAND2_X1 U5767 ( .A1(n5083), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4696)
         );
  AND3_X1 U5768 ( .A1(n4698), .A2(n4697), .A3(n4696), .ZN(n4703) );
  AOI22_X1 U5769 ( .A1(n3534), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3599), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4702) );
  AOI22_X1 U5770 ( .A1(n5070), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4701) );
  INV_X1 U5771 ( .A(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4699) );
  OR2_X1 U5772 ( .A1(n5018), .A2(n4699), .ZN(n4700) );
  NAND4_X1 U5773 ( .A1(n4703), .A2(n4702), .A3(n4701), .A4(n4700), .ZN(n4709)
         );
  AOI22_X1 U5774 ( .A1(n5085), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n5026), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4707) );
  AOI22_X1 U5775 ( .A1(n5081), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n5050), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4706) );
  AOI22_X1 U5776 ( .A1(n4882), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n5082), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4705) );
  AOI22_X1 U5777 ( .A1(n5080), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n5069), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4704) );
  NAND4_X1 U5778 ( .A1(n4707), .A2(n4706), .A3(n4705), .A4(n4704), .ZN(n4708)
         );
  OR2_X1 U5779 ( .A1(n4709), .A2(n4708), .ZN(n4712) );
  INV_X1 U5780 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5871) );
  OAI22_X1 U5781 ( .A1(n5008), .A2(n4073), .B1(n4710), .B2(n5871), .ZN(n4711)
         );
  AOI21_X1 U5782 ( .B1(n5096), .B2(n4712), .A(n4711), .ZN(n4713) );
  NAND2_X1 U5783 ( .A1(n4714), .A2(n4713), .ZN(n4717) );
  NAND2_X1 U5784 ( .A1(n4715), .A2(n4717), .ZN(n4741) );
  OR2_X1 U5785 ( .A1(n4657), .A2(n4717), .ZN(n4718) );
  AND2_X1 U5786 ( .A1(n4716), .A2(n4718), .ZN(n6031) );
  INV_X1 U5787 ( .A(n6031), .ZN(n4719) );
  OAI222_X1 U5788 ( .A1(n5879), .A2(n6011), .B1(n6022), .B2(n4686), .C1(n6012), 
        .C2(n4719), .ZN(U2843) );
  AOI22_X1 U5789 ( .A1(n3534), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n5026), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4727) );
  AOI22_X1 U5790 ( .A1(n5081), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n5070), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4726) );
  NAND2_X1 U5791 ( .A1(n5080), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4722) );
  NAND2_X1 U5792 ( .A1(n3599), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4721) );
  NAND2_X1 U5793 ( .A1(n5069), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4720) );
  AND3_X1 U5794 ( .A1(n4722), .A2(n4721), .A3(n4720), .ZN(n4725) );
  INV_X1 U5795 ( .A(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4723) );
  OR2_X1 U5796 ( .A1(n5018), .A2(n4723), .ZN(n4724) );
  NAND4_X1 U5797 ( .A1(n4727), .A2(n4726), .A3(n4725), .A4(n4724), .ZN(n4733)
         );
  AOI22_X1 U5798 ( .A1(n5076), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n5083), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4731) );
  AOI22_X1 U5799 ( .A1(n5085), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4882), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4730) );
  AOI22_X1 U5800 ( .A1(n5050), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4729) );
  AOI22_X1 U5801 ( .A1(n5075), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n5082), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4728) );
  NAND4_X1 U5802 ( .A1(n4731), .A2(n4730), .A3(n4729), .A4(n4728), .ZN(n4732)
         );
  NOR2_X1 U5803 ( .A1(n4733), .A2(n4732), .ZN(n4738) );
  INV_X1 U5804 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4735) );
  NAND2_X1 U5805 ( .A1(n6478), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4734)
         );
  OAI211_X1 U5806 ( .C1(n5008), .C2(n4735), .A(n5101), .B(n4734), .ZN(n4736)
         );
  INV_X1 U5807 ( .A(n4736), .ZN(n4737) );
  OAI21_X1 U5808 ( .B1(n5063), .B2(n4738), .A(n4737), .ZN(n4740) );
  XNOR2_X1 U5809 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n4760), .ZN(n5857)
         );
  NAND2_X1 U5810 ( .A1(n5857), .A2(n5060), .ZN(n4739) );
  NAND2_X1 U5811 ( .A1(n4740), .A2(n4739), .ZN(n4771) );
  INV_X1 U5812 ( .A(n4741), .ZN(n4765) );
  AOI22_X1 U5813 ( .A1(n5070), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4745) );
  AOI22_X1 U5814 ( .A1(n5085), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3538), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4744) );
  AOI22_X1 U5815 ( .A1(n3534), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4743) );
  AOI22_X1 U5816 ( .A1(n5076), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n5083), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4742) );
  NAND4_X1 U5817 ( .A1(n4745), .A2(n4744), .A3(n4743), .A4(n4742), .ZN(n4755)
         );
  NAND2_X1 U5818 ( .A1(n4882), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4748) );
  NAND2_X1 U5819 ( .A1(n5082), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4747)
         );
  NAND2_X1 U5820 ( .A1(n5069), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4746) );
  AND3_X1 U5821 ( .A1(n4748), .A2(n4747), .A3(n4746), .ZN(n4753) );
  AOI22_X1 U5822 ( .A1(n5050), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3599), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4752) );
  AOI22_X1 U5823 ( .A1(n5081), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4751) );
  INV_X1 U5824 ( .A(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4749) );
  OR2_X1 U5825 ( .A1(n5018), .A2(n4749), .ZN(n4750) );
  NAND4_X1 U5826 ( .A1(n4753), .A2(n4752), .A3(n4751), .A4(n4750), .ZN(n4754)
         );
  NOR2_X1 U5827 ( .A1(n4755), .A2(n4754), .ZN(n4759) );
  NAND2_X1 U5828 ( .A1(n6637), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4756)
         );
  OAI211_X1 U5829 ( .C1(n5008), .C2(n4067), .A(n5101), .B(n4756), .ZN(n4757)
         );
  INV_X1 U5830 ( .A(n4757), .ZN(n4758) );
  OAI21_X1 U5831 ( .B1(n5063), .B2(n4759), .A(n4758), .ZN(n4763) );
  OAI21_X1 U5832 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n4761), .A(n4760), 
        .ZN(n5867) );
  OR2_X1 U5833 ( .A1(n5101), .A2(n5867), .ZN(n4762) );
  NAND2_X1 U5834 ( .A1(n4763), .A2(n4762), .ZN(n5779) );
  NAND2_X1 U5835 ( .A1(n4765), .A2(n4764), .ZN(n4767) );
  INV_X1 U5836 ( .A(n4767), .ZN(n4769) );
  NAND2_X1 U5837 ( .A1(n4769), .A2(n4768), .ZN(n4819) );
  INV_X1 U5838 ( .A(n4819), .ZN(n4770) );
  AOI21_X1 U5839 ( .B1(n4771), .B2(n4766), .A(n4770), .ZN(n5487) );
  INV_X1 U5840 ( .A(n5487), .ZN(n5855) );
  AOI22_X1 U5841 ( .A1(n6029), .A2(DATAI_18_), .B1(n6025), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n4776) );
  NOR2_X1 U5842 ( .A1(n5220), .A2(n4773), .ZN(n4774) );
  NAND2_X1 U5843 ( .A1(n6032), .A2(n4774), .ZN(n6033) );
  NAND2_X1 U5844 ( .A1(n6026), .A2(DATAI_2_), .ZN(n4775) );
  OAI211_X1 U5845 ( .C1(n5855), .C2(n5391), .A(n4776), .B(n4775), .ZN(U2873)
         );
  OAI21_X1 U5846 ( .B1(n4779), .B2(n4778), .A(n4777), .ZN(n5109) );
  XNOR2_X1 U5847 ( .A(n5432), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5112)
         );
  INV_X1 U5848 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5814) );
  NAND2_X1 U5849 ( .A1(n5432), .A2(n5814), .ZN(n4780) );
  NAND2_X1 U5850 ( .A1(n3152), .A2(n4780), .ZN(n5505) );
  INV_X1 U5851 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5652) );
  NAND2_X1 U5852 ( .A1(n5432), .A2(n5652), .ZN(n4782) );
  INV_X1 U5853 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5497) );
  OAI21_X2 U5854 ( .B1(n5496), .B2(n4784), .A(n4783), .ZN(n5477) );
  INV_X1 U5855 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4786) );
  NAND2_X1 U5856 ( .A1(n5432), .A2(n4786), .ZN(n4785) );
  NAND2_X1 U5857 ( .A1(n5477), .A2(n4785), .ZN(n5479) );
  INV_X1 U5858 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5481) );
  INV_X1 U5859 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5482) );
  AND3_X1 U5860 ( .A1(n4786), .A2(n5481), .A3(n5482), .ZN(n4787) );
  NAND2_X1 U5861 ( .A1(n5479), .A2(n4787), .ZN(n4788) );
  NAND2_X1 U5862 ( .A1(n4788), .A2(n5489), .ZN(n4791) );
  INV_X1 U5863 ( .A(n5479), .ZN(n4789) );
  NAND2_X1 U5864 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5603) );
  NAND2_X1 U5865 ( .A1(n4789), .A2(n5611), .ZN(n4790) );
  NAND2_X2 U5866 ( .A1(n4791), .A2(n4790), .ZN(n5443) );
  AND2_X1 U5867 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5582) );
  AND2_X1 U5868 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5604) );
  NAND2_X1 U5869 ( .A1(n5582), .A2(n5604), .ZN(n5445) );
  NAND2_X1 U5870 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5123) );
  OAI21_X1 U5871 ( .B1(n5445), .B2(n5123), .A(n3150), .ZN(n4793) );
  NOR2_X1 U5872 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5605) );
  NOR2_X1 U5873 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5581) );
  INV_X1 U5874 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5574) );
  INV_X1 U5875 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5562) );
  NAND4_X1 U5876 ( .A1(n5605), .A2(n5581), .A3(n5574), .A4(n5562), .ZN(n4792)
         );
  XNOR2_X1 U5877 ( .A(n5432), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5769)
         );
  NAND2_X1 U5878 ( .A1(n5402), .A2(n5769), .ZN(n5203) );
  INV_X1 U5879 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5791) );
  NAND2_X1 U5880 ( .A1(n5432), .A2(n5791), .ZN(n4794) );
  NAND2_X1 U5881 ( .A1(n5203), .A2(n4794), .ZN(n4795) );
  NAND2_X1 U5882 ( .A1(n5432), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5421) );
  AND2_X1 U5883 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5530) );
  NAND2_X1 U5884 ( .A1(n5413), .A2(n5530), .ZN(n5392) );
  INV_X1 U5885 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5529) );
  BUF_X2 U5886 ( .A(n4795), .Z(n5401) );
  OR2_X1 U5887 ( .A1(n3150), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5422)
         );
  INV_X1 U5888 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5550) );
  INV_X1 U5889 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5172) );
  NAND2_X1 U5890 ( .A1(n5550), .A2(n5172), .ZN(n5538) );
  NOR2_X1 U5891 ( .A1(n5422), .A2(n5538), .ZN(n5393) );
  NAND2_X1 U5892 ( .A1(n5393), .A2(n5529), .ZN(n5205) );
  INV_X1 U5893 ( .A(n5205), .ZN(n4796) );
  OR2_X1 U5894 ( .A1(n4799), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4800)
         );
  NAND2_X1 U5895 ( .A1(n4800), .A2(n4837), .ZN(n5778) );
  AOI22_X1 U5896 ( .A1(n5081), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n5026), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4804) );
  AOI22_X1 U5897 ( .A1(n3534), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4803) );
  AOI22_X1 U5898 ( .A1(n5051), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3599), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4802) );
  AOI22_X1 U5899 ( .A1(n5070), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n5082), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4801) );
  NAND4_X1 U5900 ( .A1(n4804), .A2(n4803), .A3(n4802), .A4(n4801), .ZN(n4814)
         );
  INV_X1 U5901 ( .A(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4805) );
  OR2_X1 U5902 ( .A1(n5018), .A2(n4805), .ZN(n4809) );
  NAND2_X1 U5903 ( .A1(n5083), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4808)
         );
  NAND2_X1 U5904 ( .A1(n4882), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4807) );
  NAND2_X1 U5905 ( .A1(n5069), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4806) );
  AND4_X1 U5906 ( .A1(n4809), .A2(n4808), .A3(n4807), .A4(n4806), .ZN(n4812)
         );
  AOI22_X1 U5907 ( .A1(n5076), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4811) );
  AOI22_X1 U5908 ( .A1(n5050), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4810) );
  NAND3_X1 U5909 ( .A1(n4812), .A2(n4811), .A3(n4810), .ZN(n4813) );
  OAI21_X1 U5910 ( .B1(n4814), .B2(n4813), .A(n5096), .ZN(n4817) );
  NAND2_X1 U5911 ( .A1(n5211), .A2(EAX_REG_19__SCAN_IN), .ZN(n4816) );
  NAND2_X1 U5912 ( .A1(n6478), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4815)
         );
  NAND4_X1 U5913 ( .A1(n4817), .A2(n5101), .A3(n4816), .A4(n4815), .ZN(n4818)
         );
  OAI21_X1 U5914 ( .B1(n5778), .B2(n5101), .A(n4818), .ZN(n5364) );
  NAND2_X1 U5915 ( .A1(n5050), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4822)
         );
  NAND2_X1 U5916 ( .A1(n5083), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4821)
         );
  NAND2_X1 U5917 ( .A1(n5069), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4820) );
  AND3_X1 U5918 ( .A1(n4822), .A2(n4821), .A3(n4820), .ZN(n4827) );
  AOI22_X1 U5919 ( .A1(n5051), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4826) );
  AOI22_X1 U5920 ( .A1(n3534), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4882), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4825) );
  INV_X1 U5921 ( .A(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4823) );
  OR2_X1 U5922 ( .A1(n5018), .A2(n4823), .ZN(n4824) );
  NAND4_X1 U5923 ( .A1(n4827), .A2(n4826), .A3(n4825), .A4(n4824), .ZN(n4833)
         );
  AOI22_X1 U5924 ( .A1(n5076), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4831) );
  AOI22_X1 U5925 ( .A1(n5070), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4830) );
  AOI22_X1 U5926 ( .A1(n5026), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3599), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4829) );
  AOI22_X1 U5927 ( .A1(n5081), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4828) );
  NAND4_X1 U5928 ( .A1(n4831), .A2(n4830), .A3(n4829), .A4(n4828), .ZN(n4832)
         );
  NOR2_X1 U5929 ( .A1(n4833), .A2(n4832), .ZN(n4836) );
  NAND2_X1 U5930 ( .A1(n5211), .A2(EAX_REG_20__SCAN_IN), .ZN(n4835) );
  OAI21_X1 U5931 ( .B1(n6912), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n6637), 
        .ZN(n4834) );
  OAI211_X1 U5932 ( .C1(n5063), .C2(n4836), .A(n4835), .B(n4834), .ZN(n4839)
         );
  XNOR2_X1 U5933 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .B(n4837), .ZN(n5472)
         );
  NAND2_X1 U5934 ( .A1(n5472), .A2(n5060), .ZN(n4838) );
  NAND2_X1 U5935 ( .A1(n5308), .A2(n5310), .ZN(n5294) );
  INV_X1 U5936 ( .A(n5294), .ZN(n4861) );
  NAND2_X1 U5937 ( .A1(n5051), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4842)
         );
  NAND2_X1 U5938 ( .A1(n5080), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4841) );
  NAND2_X1 U5939 ( .A1(n5069), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4840) );
  AND3_X1 U5940 ( .A1(n4842), .A2(n4841), .A3(n4840), .ZN(n4847) );
  AOI22_X1 U5941 ( .A1(n3534), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n5081), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4846) );
  AOI22_X1 U5942 ( .A1(n5076), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n5070), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4845) );
  INV_X1 U5943 ( .A(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4843) );
  OR2_X1 U5944 ( .A1(n5018), .A2(n4843), .ZN(n4844) );
  NAND4_X1 U5945 ( .A1(n4847), .A2(n4846), .A3(n4845), .A4(n4844), .ZN(n4853)
         );
  AOI22_X1 U5946 ( .A1(n5050), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4851) );
  AOI22_X1 U5947 ( .A1(n5026), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3599), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4850) );
  AOI22_X1 U5948 ( .A1(n5083), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n5082), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4849) );
  AOI22_X1 U5949 ( .A1(n4882), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4848) );
  NAND4_X1 U5950 ( .A1(n4851), .A2(n4850), .A3(n4849), .A4(n4848), .ZN(n4852)
         );
  NOR2_X1 U5951 ( .A1(n4853), .A2(n4852), .ZN(n4856) );
  INV_X1 U5952 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5301) );
  OAI21_X1 U5953 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5301), .A(n5101), .ZN(
        n4854) );
  AOI21_X1 U5954 ( .B1(n5211), .B2(EAX_REG_21__SCAN_IN), .A(n4854), .ZN(n4855)
         );
  OAI21_X1 U5955 ( .B1(n5063), .B2(n4856), .A(n4855), .ZN(n4859) );
  OAI21_X1 U5956 ( .B1(n4857), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n4879), 
        .ZN(n5467) );
  OR2_X1 U5957 ( .A1(n5467), .A2(n5101), .ZN(n4858) );
  NAND2_X1 U5958 ( .A1(n4859), .A2(n4858), .ZN(n5295) );
  NAND2_X1 U5959 ( .A1(n4861), .A2(n4860), .ZN(n5292) );
  AOI22_X1 U5960 ( .A1(n5085), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4865) );
  AOI22_X1 U5961 ( .A1(n5081), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4864) );
  AOI22_X1 U5962 ( .A1(n5050), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4882), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4863) );
  AOI22_X1 U5963 ( .A1(n5070), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n5082), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4862) );
  NAND4_X1 U5964 ( .A1(n4865), .A2(n4864), .A3(n4863), .A4(n4862), .ZN(n4875)
         );
  NAND2_X1 U5965 ( .A1(n5075), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4868) );
  NAND2_X1 U5966 ( .A1(n5083), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4867)
         );
  NAND2_X1 U5967 ( .A1(n5069), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4866) );
  AND3_X1 U5968 ( .A1(n4868), .A2(n4867), .A3(n4866), .ZN(n4873) );
  AOI22_X1 U5969 ( .A1(n3534), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3599), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4872) );
  AOI22_X1 U5970 ( .A1(n5026), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4871) );
  INV_X1 U5971 ( .A(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4869) );
  OR2_X1 U5972 ( .A1(n5018), .A2(n4869), .ZN(n4870) );
  NAND4_X1 U5973 ( .A1(n4873), .A2(n4872), .A3(n4871), .A4(n4870), .ZN(n4874)
         );
  NOR2_X1 U5974 ( .A1(n4875), .A2(n4874), .ZN(n4878) );
  OAI21_X1 U5975 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5459), .A(n5101), .ZN(
        n4876) );
  AOI21_X1 U5976 ( .B1(n5211), .B2(EAX_REG_22__SCAN_IN), .A(n4876), .ZN(n4877)
         );
  OAI21_X1 U5977 ( .B1(n5063), .B2(n4878), .A(n4877), .ZN(n4881) );
  XNOR2_X1 U5978 ( .A(n4879), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5729)
         );
  NAND2_X1 U5979 ( .A1(n5729), .A2(n5060), .ZN(n4880) );
  NAND2_X1 U5980 ( .A1(n4881), .A2(n4880), .ZN(n5358) );
  NOR2_X2 U5981 ( .A1(n5292), .A2(n5358), .ZN(n5278) );
  AOI22_X1 U5982 ( .A1(n5081), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4884) );
  AOI22_X1 U5983 ( .A1(n3534), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4882), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4883) );
  AND2_X1 U5984 ( .A1(n4884), .A2(n4883), .ZN(n4889) );
  AOI22_X1 U5985 ( .A1(n5069), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n5082), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4888) );
  NAND2_X1 U5986 ( .A1(n5050), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4887)
         );
  INV_X1 U5987 ( .A(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4885) );
  OR2_X1 U5988 ( .A1(n5018), .A2(n4885), .ZN(n4886) );
  NAND4_X1 U5989 ( .A1(n4889), .A2(n4888), .A3(n4887), .A4(n4886), .ZN(n4895)
         );
  AOI22_X1 U5990 ( .A1(n5070), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n5083), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4893) );
  AOI22_X1 U5991 ( .A1(n5076), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4892) );
  AOI22_X1 U5992 ( .A1(n3538), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3599), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4891) );
  AOI22_X1 U5993 ( .A1(n5085), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4890) );
  NAND4_X1 U5994 ( .A1(n4893), .A2(n4892), .A3(n4891), .A4(n4890), .ZN(n4894)
         );
  NOR2_X1 U5995 ( .A1(n4895), .A2(n4894), .ZN(n4917) );
  OAI22_X1 U5996 ( .A1(n5044), .A2(n4897), .B1(n4949), .B2(n4896), .ZN(n4898)
         );
  AOI21_X1 U5997 ( .B1(n5050), .B2(INSTQUEUE_REG_12__0__SCAN_IN), .A(n4898), 
        .ZN(n4902) );
  AOI22_X1 U5998 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n3534), .B1(n5026), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4901) );
  AOI22_X1 U5999 ( .A1(n5076), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4900) );
  NAND2_X1 U6000 ( .A1(n5074), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4899) );
  NAND4_X1 U6001 ( .A1(n4902), .A2(n4901), .A3(n4900), .A4(n4899), .ZN(n4908)
         );
  AOI22_X1 U6002 ( .A1(n5081), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4906) );
  AOI22_X1 U6003 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n5075), .B1(n4882), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4905) );
  AOI22_X1 U6004 ( .A1(n5070), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n5069), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4904) );
  AOI22_X1 U6005 ( .A1(n5085), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3599), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4903) );
  NAND4_X1 U6006 ( .A1(n4906), .A2(n4905), .A3(n4904), .A4(n4903), .ZN(n4907)
         );
  NOR2_X1 U6007 ( .A1(n4908), .A2(n4907), .ZN(n4918) );
  XNOR2_X1 U6008 ( .A(n4917), .B(n4918), .ZN(n4912) );
  NAND2_X1 U6009 ( .A1(n6637), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4909)
         );
  OAI211_X1 U6010 ( .C1(n5008), .C2(n4062), .A(n5101), .B(n4909), .ZN(n4910)
         );
  INV_X1 U6011 ( .A(n4910), .ZN(n4911) );
  OAI21_X1 U6012 ( .B1(n4912), .B2(n5063), .A(n4911), .ZN(n4916) );
  OR2_X1 U6013 ( .A1(n4913), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4914)
         );
  NAND2_X1 U6014 ( .A1(n4935), .A2(n4914), .ZN(n5452) );
  OR2_X1 U6015 ( .A1(n5452), .A2(n5101), .ZN(n4915) );
  AND2_X2 U6016 ( .A1(n5278), .A2(n5280), .ZN(n5277) );
  NOR2_X1 U6017 ( .A1(n4918), .A2(n4917), .ZN(n4942) );
  INV_X1 U6018 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4919) );
  OR2_X1 U6019 ( .A1(n5018), .A2(n4919), .ZN(n4923) );
  NAND2_X1 U6020 ( .A1(n5050), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4922)
         );
  NAND2_X1 U6021 ( .A1(n5083), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4921)
         );
  NAND2_X1 U6022 ( .A1(n5069), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4920) );
  AND4_X1 U6023 ( .A1(n4923), .A2(n4922), .A3(n4921), .A4(n4920), .ZN(n4926)
         );
  AOI22_X1 U6024 ( .A1(n5085), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4925) );
  AOI22_X1 U6025 ( .A1(n3534), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4882), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4924) );
  NAND3_X1 U6026 ( .A1(n4926), .A2(n4925), .A3(n4924), .ZN(n4932) );
  AOI22_X1 U6027 ( .A1(n5076), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4930) );
  AOI22_X1 U6028 ( .A1(n5070), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4929) );
  AOI22_X1 U6029 ( .A1(n3538), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3599), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4928) );
  AOI22_X1 U6030 ( .A1(n5081), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4927) );
  NAND4_X1 U6031 ( .A1(n4930), .A2(n4929), .A3(n4928), .A4(n4927), .ZN(n4931)
         );
  OR2_X1 U6032 ( .A1(n4932), .A2(n4931), .ZN(n4941) );
  INV_X1 U6033 ( .A(n4941), .ZN(n4933) );
  XNOR2_X1 U6034 ( .A(n4942), .B(n4933), .ZN(n4934) );
  NAND2_X1 U6035 ( .A1(n4934), .A2(n5096), .ZN(n4940) );
  NAND2_X1 U6036 ( .A1(n5210), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4937)
         );
  XNOR2_X1 U6037 ( .A(n4935), .B(n4367), .ZN(n5717) );
  NAND2_X1 U6038 ( .A1(n5717), .A2(n5060), .ZN(n4936) );
  OAI211_X1 U6039 ( .C1(n5008), .C2(n3677), .A(n4937), .B(n4936), .ZN(n4938)
         );
  INV_X1 U6040 ( .A(n4938), .ZN(n4939) );
  NAND2_X1 U6041 ( .A1(n4940), .A2(n4939), .ZN(n5348) );
  NAND2_X1 U6042 ( .A1(n5277), .A2(n5348), .ZN(n5339) );
  INV_X1 U6043 ( .A(n5339), .ZN(n4967) );
  NAND2_X1 U6044 ( .A1(n4942), .A2(n4941), .ZN(n4968) );
  AOI22_X1 U6045 ( .A1(n5076), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n5083), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4946) );
  AOI22_X1 U6046 ( .A1(n5026), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4945) );
  AOI22_X1 U6047 ( .A1(n3534), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4944) );
  AOI22_X1 U6048 ( .A1(n5051), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4882), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4943) );
  NAND4_X1 U6049 ( .A1(n4946), .A2(n4945), .A3(n4944), .A4(n4943), .ZN(n4957)
         );
  INV_X1 U6050 ( .A(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4950) );
  OAI22_X1 U6051 ( .A1(n4947), .A2(n4950), .B1(n4949), .B2(n4948), .ZN(n4951)
         );
  AOI21_X1 U6052 ( .B1(n5086), .B2(INSTQUEUE_REG_3__2__SCAN_IN), .A(n4951), 
        .ZN(n4955) );
  AOI22_X1 U6053 ( .A1(n5081), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5050), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4954) );
  AOI22_X1 U6054 ( .A1(n5070), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3599), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4953) );
  NAND2_X1 U6055 ( .A1(n5074), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4952) );
  NAND4_X1 U6056 ( .A1(n4955), .A2(n4954), .A3(n4953), .A4(n4952), .ZN(n4956)
         );
  NOR2_X1 U6057 ( .A1(n4957), .A2(n4956), .ZN(n4969) );
  XNOR2_X1 U6058 ( .A(n4968), .B(n4969), .ZN(n4961) );
  NAND2_X1 U6059 ( .A1(n6637), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4958)
         );
  OAI211_X1 U6060 ( .C1(n5008), .C2(n3679), .A(n5101), .B(n4958), .ZN(n4959)
         );
  INV_X1 U6061 ( .A(n4959), .ZN(n4960) );
  OAI21_X1 U6062 ( .B1(n4961), .B2(n5063), .A(n4960), .ZN(n4965) );
  OR2_X1 U6063 ( .A1(n4962), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4963)
         );
  NAND2_X1 U6064 ( .A1(n4963), .A2(n4989), .ZN(n5773) );
  OR2_X1 U6065 ( .A1(n5773), .A2(n5101), .ZN(n4964) );
  NAND2_X1 U6066 ( .A1(n4965), .A2(n4964), .ZN(n5342) );
  NAND2_X1 U6067 ( .A1(n4967), .A2(n4966), .ZN(n5332) );
  NOR2_X1 U6068 ( .A1(n4969), .A2(n4968), .ZN(n5006) );
  INV_X1 U6069 ( .A(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4970) );
  OR2_X1 U6070 ( .A1(n5018), .A2(n4970), .ZN(n4974) );
  NAND2_X1 U6071 ( .A1(n5050), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4973)
         );
  NAND2_X1 U6072 ( .A1(n5083), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4972)
         );
  NAND2_X1 U6073 ( .A1(n5069), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4971) );
  AND4_X1 U6074 ( .A1(n4974), .A2(n4973), .A3(n4972), .A4(n4971), .ZN(n4977)
         );
  AOI22_X1 U6075 ( .A1(n5085), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4976) );
  AOI22_X1 U6076 ( .A1(n3534), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4882), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4975) );
  NAND3_X1 U6077 ( .A1(n4977), .A2(n4976), .A3(n4975), .ZN(n4983) );
  AOI22_X1 U6078 ( .A1(n5076), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4981) );
  AOI22_X1 U6079 ( .A1(n5070), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4980) );
  AOI22_X1 U6080 ( .A1(n5026), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3599), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4979) );
  AOI22_X1 U6081 ( .A1(n5081), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4978) );
  NAND4_X1 U6082 ( .A1(n4981), .A2(n4980), .A3(n4979), .A4(n4978), .ZN(n4982)
         );
  OR2_X1 U6083 ( .A1(n4983), .A2(n4982), .ZN(n5005) );
  XNOR2_X1 U6084 ( .A(n5006), .B(n5005), .ZN(n4988) );
  INV_X1 U6085 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4985) );
  NAND2_X1 U6086 ( .A1(n6637), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4984)
         );
  OAI211_X1 U6087 ( .C1(n5008), .C2(n4985), .A(n5101), .B(n4984), .ZN(n4986)
         );
  INV_X1 U6088 ( .A(n4986), .ZN(n4987) );
  OAI21_X1 U6089 ( .B1(n4988), .B2(n5063), .A(n4987), .ZN(n4991) );
  XNOR2_X1 U6090 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .B(n4989), .ZN(n5698)
         );
  NAND2_X1 U6091 ( .A1(n5698), .A2(n5060), .ZN(n4990) );
  NAND2_X1 U6092 ( .A1(n4991), .A2(n4990), .ZN(n5334) );
  INV_X1 U6093 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4994) );
  AOI22_X1 U6094 ( .A1(n5083), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n5082), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4993) );
  NAND2_X1 U6095 ( .A1(n4882), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4992) );
  OAI211_X1 U6096 ( .C1(n4994), .C2(n5018), .A(n4993), .B(n4992), .ZN(n4995)
         );
  INV_X1 U6097 ( .A(n4995), .ZN(n4998) );
  AOI22_X1 U6098 ( .A1(n5076), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4997) );
  AOI22_X1 U6099 ( .A1(n5075), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3599), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4996) );
  NAND3_X1 U6100 ( .A1(n4998), .A2(n4997), .A3(n4996), .ZN(n5004) );
  AOI22_X1 U6101 ( .A1(n5026), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n5002) );
  AOI22_X1 U6102 ( .A1(n5051), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n5081), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5001) );
  AOI22_X1 U6103 ( .A1(n3534), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n5050), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5000) );
  AOI22_X1 U6104 ( .A1(n5070), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n5069), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4999) );
  NAND4_X1 U6105 ( .A1(n5002), .A2(n5001), .A3(n5000), .A4(n4999), .ZN(n5003)
         );
  NOR2_X1 U6106 ( .A1(n5004), .A2(n5003), .ZN(n5016) );
  NAND2_X1 U6107 ( .A1(n5006), .A2(n5005), .ZN(n5015) );
  XNOR2_X1 U6108 ( .A(n5016), .B(n5015), .ZN(n5011) );
  NAND2_X1 U6109 ( .A1(n6637), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5007)
         );
  OAI211_X1 U6110 ( .C1(n5008), .C2(n3681), .A(n5101), .B(n5007), .ZN(n5009)
         );
  INV_X1 U6111 ( .A(n5009), .ZN(n5010) );
  OAI21_X1 U6112 ( .B1(n5011), .B2(n5063), .A(n5010), .ZN(n5014) );
  OAI21_X1 U6113 ( .B1(n5012), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5036), 
        .ZN(n5690) );
  OR2_X1 U6114 ( .A1(n5690), .A2(n5101), .ZN(n5013) );
  NOR2_X1 U6115 ( .A1(n5016), .A2(n5015), .ZN(n5059) );
  INV_X1 U6116 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5017) );
  OR2_X1 U6117 ( .A1(n5018), .A2(n5017), .ZN(n5022) );
  NAND2_X1 U6118 ( .A1(n5050), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5021)
         );
  NAND2_X1 U6119 ( .A1(n5083), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n5020)
         );
  NAND2_X1 U6120 ( .A1(n5069), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n5019) );
  AND4_X1 U6121 ( .A1(n5022), .A2(n5021), .A3(n5020), .A4(n5019), .ZN(n5025)
         );
  AOI22_X1 U6122 ( .A1(n5085), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5024) );
  AOI22_X1 U6123 ( .A1(n3534), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4882), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n5023) );
  NAND3_X1 U6124 ( .A1(n5025), .A2(n5024), .A3(n5023), .ZN(n5032) );
  AOI22_X1 U6125 ( .A1(n5076), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n5030) );
  AOI22_X1 U6126 ( .A1(n5070), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n5082), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5029) );
  AOI22_X1 U6127 ( .A1(n5026), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3599), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5028) );
  AOI22_X1 U6128 ( .A1(n5081), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n5027) );
  NAND4_X1 U6129 ( .A1(n5030), .A2(n5029), .A3(n5028), .A4(n5027), .ZN(n5031)
         );
  OR2_X1 U6130 ( .A1(n5032), .A2(n5031), .ZN(n5058) );
  INV_X1 U6131 ( .A(n5058), .ZN(n5033) );
  XNOR2_X1 U6132 ( .A(n5059), .B(n5033), .ZN(n5034) );
  NAND2_X1 U6133 ( .A1(n5034), .A2(n5096), .ZN(n5039) );
  OAI21_X1 U6134 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5408), .A(n5101), .ZN(
        n5035) );
  AOI21_X1 U6135 ( .B1(n5211), .B2(EAX_REG_28__SCAN_IN), .A(n5035), .ZN(n5038)
         );
  XNOR2_X1 U6136 ( .A(n5036), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5682)
         );
  AND2_X1 U6137 ( .A1(n5682), .A2(n5060), .ZN(n5037) );
  OR2_X1 U6138 ( .A1(n5040), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5041)
         );
  NAND2_X1 U6139 ( .A1(n5100), .A2(n5041), .ZN(n5397) );
  INV_X1 U6140 ( .A(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n5042) );
  OAI22_X1 U6141 ( .A1(n5044), .A2(n5043), .B1(n4947), .B2(n5042), .ZN(n5045)
         );
  AOI21_X1 U6142 ( .B1(n5081), .B2(INSTQUEUE_REG_10__6__SCAN_IN), .A(n5045), 
        .ZN(n5049) );
  AOI22_X1 U6143 ( .A1(n3534), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n5048) );
  AOI22_X1 U6144 ( .A1(n5076), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5047) );
  NAND2_X1 U6145 ( .A1(n5074), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5046) );
  NAND4_X1 U6146 ( .A1(n5049), .A2(n5048), .A3(n5047), .A4(n5046), .ZN(n5057)
         );
  AOI22_X1 U6147 ( .A1(n3538), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n5070), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n5055) );
  AOI22_X1 U6148 ( .A1(n5050), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5054) );
  AOI22_X1 U6149 ( .A1(n5051), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3599), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5053) );
  AOI22_X1 U6150 ( .A1(n4882), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n5052) );
  NAND4_X1 U6151 ( .A1(n5055), .A2(n5054), .A3(n5053), .A4(n5052), .ZN(n5056)
         );
  NOR2_X1 U6152 ( .A1(n5057), .A2(n5056), .ZN(n5067) );
  NAND2_X1 U6153 ( .A1(n5059), .A2(n5058), .ZN(n5066) );
  XNOR2_X1 U6154 ( .A(n5067), .B(n5066), .ZN(n5064) );
  AOI21_X1 U6155 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6637), .A(n5060), 
        .ZN(n5062) );
  NAND2_X1 U6156 ( .A1(n5211), .A2(EAX_REG_29__SCAN_IN), .ZN(n5061) );
  OAI211_X1 U6157 ( .C1(n5064), .C2(n5063), .A(n5062), .B(n5061), .ZN(n5065)
         );
  NOR2_X1 U6158 ( .A1(n5067), .A2(n5066), .ZN(n5095) );
  INV_X1 U6159 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5072) );
  AOI22_X1 U6160 ( .A1(n5070), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5069), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n5071) );
  OAI21_X1 U6161 ( .B1(n3590), .B2(n5072), .A(n5071), .ZN(n5073) );
  AOI21_X1 U6162 ( .B1(n5074), .B2(INSTQUEUE_REG_2__7__SCAN_IN), .A(n5073), 
        .ZN(n5079) );
  AOI22_X1 U6163 ( .A1(n5076), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5078) );
  AOI22_X1 U6164 ( .A1(n3534), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n5026), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5077) );
  NAND3_X1 U6165 ( .A1(n5079), .A2(n5078), .A3(n5077), .ZN(n5093) );
  AOI22_X1 U6166 ( .A1(n5081), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n5091) );
  AOI22_X1 U6167 ( .A1(n5083), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n5082), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5090) );
  AOI22_X1 U6168 ( .A1(n5085), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3599), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5089) );
  AOI22_X1 U6169 ( .A1(n5087), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5088) );
  NAND4_X1 U6170 ( .A1(n5091), .A2(n5090), .A3(n5089), .A4(n5088), .ZN(n5092)
         );
  NOR2_X1 U6171 ( .A1(n5093), .A2(n5092), .ZN(n5094) );
  XNOR2_X1 U6172 ( .A(n5095), .B(n5094), .ZN(n5097) );
  NAND2_X1 U6173 ( .A1(n5097), .A2(n5096), .ZN(n5104) );
  OAI21_X1 U6174 ( .B1(n6912), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n6637), 
        .ZN(n5098) );
  OAI21_X1 U6175 ( .B1(n5008), .B2(n3670), .A(n5098), .ZN(n5099) );
  INV_X1 U6176 ( .A(n5099), .ZN(n5103) );
  XNOR2_X1 U6177 ( .A(n5100), .B(n5252), .ZN(n5251) );
  NOR2_X1 U6178 ( .A1(n5251), .A2(n5101), .ZN(n5102) );
  NAND2_X1 U6179 ( .A1(n6176), .A2(REIP_REG_30__SCAN_IN), .ZN(n5188) );
  NAND2_X1 U6180 ( .A1(n6117), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5106)
         );
  OAI211_X1 U6181 ( .C1(n6111), .C2(n5251), .A(n5188), .B(n5106), .ZN(n5107)
         );
  OAI21_X1 U6182 ( .B1(n5194), .B2(n5835), .A(n5108), .ZN(U2956) );
  CLKBUF_X1 U6183 ( .A(n5109), .Z(n5110) );
  OAI21_X1 U6184 ( .B1(n5110), .B2(n5112), .A(n3152), .ZN(n5822) );
  NAND2_X1 U6185 ( .A1(n5822), .A2(n6115), .ZN(n5117) );
  INV_X1 U6186 ( .A(n5891), .ZN(n5115) );
  INV_X1 U6187 ( .A(REIP_REG_13__SCAN_IN), .ZN(n5113) );
  OAI22_X1 U6188 ( .A1(n5786), .A2(n4363), .B1(n5819), .B2(n5113), .ZN(n5114)
         );
  AOI21_X1 U6189 ( .B1(n5781), .B2(n5115), .A(n5114), .ZN(n5116) );
  OAI211_X1 U6190 ( .C1(n6013), .C2(n5512), .A(n5117), .B(n5116), .ZN(U2973)
         );
  NOR2_X1 U6191 ( .A1(n5119), .A2(n5118), .ZN(n5122) );
  NAND2_X1 U6192 ( .A1(n5120), .A2(n5122), .ZN(n5640) );
  NOR2_X1 U6193 ( .A1(n5645), .A2(n5640), .ZN(n5651) );
  NAND2_X1 U6194 ( .A1(n5122), .A2(n5121), .ZN(n5642) );
  NOR2_X1 U6195 ( .A1(n5134), .A2(n5642), .ZN(n6121) );
  NAND2_X1 U6196 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6122) );
  INV_X1 U6197 ( .A(n6122), .ZN(n5813) );
  NAND2_X1 U6198 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5813), .ZN(n5654) );
  NOR2_X1 U6199 ( .A1(n5652), .A2(n5654), .ZN(n5797) );
  NAND3_X1 U6200 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5797), .ZN(n5595) );
  INV_X1 U6201 ( .A(n5603), .ZN(n5611) );
  NAND2_X1 U6202 ( .A1(n5611), .A2(n5604), .ZN(n5127) );
  NOR2_X1 U6203 ( .A1(n5634), .A2(n5127), .ZN(n5580) );
  INV_X1 U6204 ( .A(n5123), .ZN(n5133) );
  AND2_X1 U6205 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5554) );
  NAND2_X1 U6206 ( .A1(n5792), .A2(n5554), .ZN(n5528) );
  INV_X1 U6207 ( .A(n5530), .ZN(n5537) );
  NOR3_X1 U6208 ( .A1(n5528), .A2(n5537), .A3(n5529), .ZN(n5519) );
  INV_X1 U6209 ( .A(n5519), .ZN(n5191) );
  NOR2_X1 U6210 ( .A1(n5640), .A2(n5595), .ZN(n5597) );
  INV_X1 U6211 ( .A(n5127), .ZN(n5124) );
  AND2_X1 U6212 ( .A1(n5597), .A2(n5124), .ZN(n5125) );
  NOR2_X1 U6213 ( .A1(n5645), .A2(n5125), .ZN(n5126) );
  NOR2_X1 U6214 ( .A1(n5641), .A2(n5126), .ZN(n5130) );
  OR3_X1 U6215 ( .A1(n5642), .A2(n5595), .A3(n5127), .ZN(n5128) );
  NAND2_X1 U6216 ( .A1(n5643), .A2(n5128), .ZN(n5129) );
  AND2_X1 U6217 ( .A1(n5130), .A2(n5129), .ZN(n5578) );
  INV_X1 U6218 ( .A(n5582), .ZN(n5131) );
  NAND2_X1 U6219 ( .A1(n6170), .A2(n5131), .ZN(n5132) );
  NAND2_X1 U6220 ( .A1(n5578), .A2(n5132), .ZN(n5569) );
  AOI21_X1 U6221 ( .B1(n5134), .B2(n5645), .A(n5133), .ZN(n5135) );
  OR2_X1 U6222 ( .A1(n5569), .A2(n5135), .ZN(n5790) );
  INV_X1 U6223 ( .A(n5554), .ZN(n5136) );
  AND2_X1 U6224 ( .A1(n6170), .A2(n5136), .ZN(n5137) );
  NOR2_X1 U6225 ( .A1(n5790), .A2(n5137), .ZN(n5548) );
  NAND2_X1 U6226 ( .A1(n6170), .A2(n5537), .ZN(n5138) );
  NAND2_X1 U6227 ( .A1(n5548), .A2(n5138), .ZN(n5527) );
  AOI21_X1 U6228 ( .B1(n5529), .B2(n6170), .A(n5527), .ZN(n5514) );
  OR2_X1 U6229 ( .A1(n5170), .A2(EBX_REG_17__SCAN_IN), .ZN(n5141) );
  NAND2_X1 U6230 ( .A1(n3174), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5139) );
  OAI211_X1 U6231 ( .C1(n5168), .C2(EBX_REG_17__SCAN_IN), .A(n5167), .B(n5139), 
        .ZN(n5140) );
  NAND2_X1 U6232 ( .A1(n5141), .A2(n5140), .ZN(n5631) );
  INV_X1 U6233 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5609) );
  NAND2_X1 U6234 ( .A1(n5167), .A2(n5609), .ZN(n5143) );
  INV_X1 U6235 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5744) );
  NAND2_X1 U6236 ( .A1(n5178), .A2(n5744), .ZN(n5142) );
  NAND3_X1 U6237 ( .A1(n5143), .A2(n3174), .A3(n5142), .ZN(n5144) );
  OAI21_X1 U6238 ( .B1(n5227), .B2(EBX_REG_19__SCAN_IN), .A(n5144), .ZN(n5368)
         );
  OR2_X1 U6239 ( .A1(n5234), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5145)
         );
  INV_X1 U6240 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5851) );
  NAND2_X1 U6241 ( .A1(n5178), .A2(n5851), .ZN(n5365) );
  AND2_X1 U6242 ( .A1(n5145), .A2(n5365), .ZN(n5150) );
  OR2_X1 U6243 ( .A1(n5234), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5147)
         );
  INV_X1 U6244 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5362) );
  NAND2_X1 U6245 ( .A1(n5178), .A2(n5362), .ZN(n5146) );
  NAND2_X1 U6246 ( .A1(n5147), .A2(n5146), .ZN(n5311) );
  NAND2_X1 U6247 ( .A1(n5150), .A2(n5311), .ZN(n5149) );
  NAND2_X1 U6248 ( .A1(n3475), .A2(EBX_REG_20__SCAN_IN), .ZN(n5148) );
  INV_X1 U6249 ( .A(n5150), .ZN(n5366) );
  MUX2_X1 U6250 ( .A(n5170), .B(n3842), .S(EBX_REG_21__SCAN_IN), .Z(n5153) );
  OAI21_X1 U6251 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n5234), .A(n5153), 
        .ZN(n5298) );
  NOR2_X2 U6252 ( .A1(n5299), .A2(n5298), .ZN(n5356) );
  AOI22_X1 U6253 ( .A1(n3472), .A2(EBX_REG_22__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5168), .ZN(n5154) );
  OAI211_X1 U6254 ( .C1(EBX_REG_22__SCAN_IN), .C2(n5227), .A(n5154), .B(n5157), 
        .ZN(n5355) );
  NAND2_X1 U6255 ( .A1(n5356), .A2(n5355), .ZN(n5283) );
  NAND2_X1 U6256 ( .A1(n3842), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5155) );
  OAI211_X1 U6257 ( .C1(n5168), .C2(EBX_REG_23__SCAN_IN), .A(n5167), .B(n5155), 
        .ZN(n5156) );
  OAI21_X1 U6258 ( .B1(n5170), .B2(EBX_REG_23__SCAN_IN), .A(n5156), .ZN(n5284)
         );
  OR2_X2 U6259 ( .A1(n5283), .A2(n5284), .ZN(n5350) );
  INV_X1 U6260 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5721) );
  OAI21_X1 U6261 ( .B1(n5721), .B2(n5167), .A(n5157), .ZN(n5160) );
  NAND2_X1 U6262 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n5168), .ZN(n5158) );
  OAI21_X1 U6263 ( .B1(n5227), .B2(EBX_REG_24__SCAN_IN), .A(n5158), .ZN(n5159)
         );
  NOR2_X1 U6264 ( .A1(n5160), .A2(n5159), .ZN(n5349) );
  MUX2_X1 U6265 ( .A(n5170), .B(n3842), .S(EBX_REG_25__SCAN_IN), .Z(n5162) );
  OR2_X1 U6266 ( .A1(n5234), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5161)
         );
  AND2_X1 U6267 ( .A1(n5162), .A2(n5161), .ZN(n5343) );
  AND2_X2 U6268 ( .A1(n5351), .A2(n5343), .ZN(n5345) );
  INV_X1 U6269 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5555) );
  NAND2_X1 U6270 ( .A1(n5167), .A2(n5555), .ZN(n5164) );
  INV_X1 U6271 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5707) );
  NAND2_X1 U6272 ( .A1(n5178), .A2(n5707), .ZN(n5163) );
  NAND3_X1 U6273 ( .A1(n5164), .A2(n3842), .A3(n5163), .ZN(n5165) );
  OAI21_X1 U6274 ( .B1(n5227), .B2(EBX_REG_26__SCAN_IN), .A(n5165), .ZN(n5335)
         );
  NAND2_X1 U6275 ( .A1(n3842), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5166) );
  OAI211_X1 U6276 ( .C1(n5168), .C2(EBX_REG_27__SCAN_IN), .A(n5167), .B(n5166), 
        .ZN(n5169) );
  OAI21_X1 U6277 ( .B1(n5170), .B2(EBX_REG_27__SCAN_IN), .A(n5169), .ZN(n5542)
         );
  OR2_X2 U6278 ( .A1(n5543), .A2(n5542), .ZN(n5545) );
  INV_X1 U6279 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5329) );
  NAND2_X1 U6280 ( .A1(n5171), .A2(n5329), .ZN(n5176) );
  NAND2_X1 U6281 ( .A1(n5167), .A2(n5172), .ZN(n5174) );
  NAND2_X1 U6282 ( .A1(n5178), .A2(n5329), .ZN(n5173) );
  NAND3_X1 U6283 ( .A1(n5174), .A2(n3174), .A3(n5173), .ZN(n5175) );
  AND2_X1 U6284 ( .A1(n5176), .A2(n5175), .ZN(n5326) );
  OR2_X2 U6285 ( .A1(n5545), .A2(n5326), .ZN(n5328) );
  OR2_X1 U6286 ( .A1(n5234), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5180)
         );
  INV_X1 U6287 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5177) );
  NAND2_X1 U6288 ( .A1(n5178), .A2(n5177), .ZN(n5179) );
  NAND2_X1 U6289 ( .A1(n5180), .A2(n5179), .ZN(n5263) );
  NOR2_X2 U6290 ( .A1(n5328), .A2(n5263), .ZN(n5226) );
  INV_X1 U6291 ( .A(n5226), .ZN(n5185) );
  NAND2_X1 U6292 ( .A1(n5185), .A2(n3174), .ZN(n5232) );
  NAND2_X1 U6293 ( .A1(n5234), .A2(EBX_REG_30__SCAN_IN), .ZN(n5182) );
  NAND2_X1 U6294 ( .A1(n5168), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5181) );
  AND2_X1 U6295 ( .A1(n5182), .A2(n5181), .ZN(n5231) );
  INV_X1 U6296 ( .A(n5231), .ZN(n5184) );
  OR2_X1 U6297 ( .A1(n5226), .A2(n5328), .ZN(n5183) );
  NAND3_X1 U6298 ( .A1(n5232), .A2(n5184), .A3(n5183), .ZN(n5187) );
  INV_X1 U6299 ( .A(n5328), .ZN(n5228) );
  OAI211_X1 U6300 ( .C1(n5228), .C2(n3174), .A(n5185), .B(n5231), .ZN(n5186)
         );
  OAI21_X1 U6301 ( .B1(n5257), .B2(n6163), .A(n5188), .ZN(n5189) );
  INV_X1 U6302 ( .A(n5189), .ZN(n5190) );
  INV_X1 U6303 ( .A(n5192), .ZN(n5193) );
  OAI21_X1 U6304 ( .B1(n5194), .B2(n6125), .A(n5193), .ZN(U2988) );
  INV_X1 U6305 ( .A(n5669), .ZN(n5662) );
  INV_X1 U6306 ( .A(n6733), .ZN(n5195) );
  AOI21_X1 U6307 ( .B1(n5662), .B2(n5195), .A(n5679), .ZN(n5202) );
  INV_X1 U6308 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5518) );
  AOI22_X1 U6309 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5518), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n3876), .ZN(n5673) );
  NOR2_X1 U6310 ( .A1(n5673), .A2(n5196), .ZN(n5199) );
  NOR3_X1 U6311 ( .A1(n5662), .A2(n5197), .A3(n6733), .ZN(n5198) );
  AOI211_X1 U6312 ( .C1(n5200), .C2(n5827), .A(n5199), .B(n5198), .ZN(n5201)
         );
  OAI22_X1 U6313 ( .A1(n5202), .A2(n3191), .B1(n5679), .B2(n5201), .ZN(U3459)
         );
  NOR3_X1 U6315 ( .A1(n5204), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5205), 
        .ZN(n5206) );
  AOI21_X1 U6316 ( .B1(n5207), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5206), 
        .ZN(n5208) );
  XNOR2_X1 U6317 ( .A(n5208), .B(n5518), .ZN(n5522) );
  NAND2_X1 U6318 ( .A1(n5261), .A2(n5209), .ZN(n5214) );
  AOI22_X1 U6319 ( .A1(n5211), .A2(EAX_REG_31__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n5210), .ZN(n5212) );
  INV_X1 U6320 ( .A(n5212), .ZN(n5213) );
  XNOR2_X2 U6321 ( .A(n5214), .B(n5213), .ZN(n5225) );
  INV_X1 U6322 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6918) );
  NOR2_X1 U6323 ( .A1(n5819), .A2(n6918), .ZN(n5516) );
  AOI21_X1 U6324 ( .B1(n6117), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5516), 
        .ZN(n5215) );
  OAI21_X1 U6325 ( .B1(n6111), .B2(n5216), .A(n5215), .ZN(n5217) );
  OAI21_X1 U6326 ( .B1(n5522), .B2(n5835), .A(n5218), .ZN(U2955) );
  NAND3_X1 U6327 ( .A1(n5225), .A2(n5220), .A3(n5219), .ZN(n5222) );
  AOI22_X1 U6328 ( .A1(n6029), .A2(DATAI_31_), .B1(n6025), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n5221) );
  NAND2_X1 U6329 ( .A1(n5222), .A2(n5221), .ZN(U2860) );
  INV_X1 U6330 ( .A(n5377), .ZN(n5224) );
  INV_X1 U6331 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5223) );
  OAI222_X1 U6332 ( .A1(n6012), .A2(n5224), .B1(n6022), .B2(n5223), .C1(n5257), 
        .C2(n6011), .ZN(U2829) );
  INV_X1 U6333 ( .A(n5225), .ZN(n5249) );
  NAND2_X1 U6334 ( .A1(n5226), .A2(n3174), .ZN(n5230) );
  NOR2_X1 U6335 ( .A1(n5227), .A2(EBX_REG_29__SCAN_IN), .ZN(n5264) );
  NAND2_X1 U6336 ( .A1(n5228), .A2(n5264), .ZN(n5229) );
  NAND2_X1 U6337 ( .A1(n5230), .A2(n5229), .ZN(n5268) );
  NAND2_X1 U6338 ( .A1(n5268), .A2(n5231), .ZN(n5233) );
  NAND2_X1 U6339 ( .A1(n5233), .A2(n5232), .ZN(n5238) );
  INV_X1 U6340 ( .A(n5234), .ZN(n5236) );
  NOR2_X1 U6341 ( .A1(n5168), .A2(EBX_REG_31__SCAN_IN), .ZN(n5235) );
  AOI21_X1 U6342 ( .B1(n5236), .B2(n5518), .A(n5235), .ZN(n5237) );
  XNOR2_X1 U6343 ( .A(n5238), .B(n5237), .ZN(n5517) );
  NAND3_X1 U6344 ( .A1(n5239), .A2(EBX_REG_31__SCAN_IN), .A3(n6725), .ZN(n5241) );
  NAND2_X1 U6345 ( .A1(n5997), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5240)
         );
  OAI21_X1 U6346 ( .B1(n6830), .B2(n5241), .A(n5240), .ZN(n5244) );
  INV_X1 U6347 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6786) );
  INV_X1 U6348 ( .A(REIP_REG_27__SCAN_IN), .ZN(n7012) );
  NOR2_X1 U6349 ( .A1(n6786), .A2(n7012), .ZN(n5242) );
  INV_X1 U6350 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6783) );
  INV_X1 U6351 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6967) );
  INV_X1 U6352 ( .A(REIP_REG_19__SCAN_IN), .ZN(n7043) );
  INV_X1 U6353 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6780) );
  INV_X1 U6354 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6779) );
  NOR3_X1 U6355 ( .A1(n6780), .A2(n6779), .A3(n5868), .ZN(n5245) );
  NAND3_X1 U6356 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5245), .A3(n5931), .ZN(
        n5746) );
  NOR4_X1 U6357 ( .A1(n6783), .A2(n6967), .A3(n7043), .A4(n5746), .ZN(n5302)
         );
  NAND4_X1 U6358 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5302), .ZN(n5282) );
  NAND3_X1 U6359 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n5246) );
  OAI21_X1 U6360 ( .B1(n5282), .B2(n5246), .A(n5989), .ZN(n5699) );
  OAI21_X1 U6361 ( .B1(n5242), .B2(n5934), .A(n5699), .ZN(n5681) );
  INV_X1 U6362 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6909) );
  NOR2_X1 U6363 ( .A1(n5681), .A2(n6909), .ZN(n5269) );
  AOI211_X1 U6364 ( .C1(n5269), .C2(REIP_REG_30__SCAN_IN), .A(n5303), .B(n6918), .ZN(n5243) );
  AOI211_X1 U6365 ( .C1(n5517), .C2(n5965), .A(n5244), .B(n5243), .ZN(n5248)
         );
  INV_X1 U6366 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6983) );
  NAND2_X1 U6367 ( .A1(n5977), .A2(n5245), .ZN(n5860) );
  NAND3_X1 U6368 ( .A1(n5747), .A2(REIP_REG_18__SCAN_IN), .A3(
        REIP_REG_19__SCAN_IN), .ZN(n5314) );
  NAND4_X1 U6369 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5297), .ZN(n5710) );
  NOR2_X1 U6370 ( .A1(n5710), .A2(n5246), .ZN(n5695) );
  NAND3_X1 U6371 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .A3(
        n5695), .ZN(n5270) );
  INV_X1 U6372 ( .A(n5270), .ZN(n5250) );
  NAND4_X1 U6373 ( .A1(n5250), .A2(REIP_REG_30__SCAN_IN), .A3(
        REIP_REG_29__SCAN_IN), .A4(n6918), .ZN(n5247) );
  OAI211_X1 U6374 ( .C1(n5249), .C2(n5937), .A(n5248), .B(n5247), .ZN(U2796)
         );
  INV_X1 U6375 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6930) );
  NAND3_X1 U6376 ( .A1(n5250), .A2(REIP_REG_29__SCAN_IN), .A3(n6930), .ZN(
        n5256) );
  NOR3_X1 U6377 ( .A1(n5303), .A2(n5269), .A3(n6930), .ZN(n5254) );
  OAI22_X1 U6378 ( .A1(n5252), .A2(n5872), .B1(n5251), .B2(n5988), .ZN(n5253)
         );
  AOI211_X1 U6379 ( .C1(n5980), .C2(EBX_REG_30__SCAN_IN), .A(n5254), .B(n5253), 
        .ZN(n5255) );
  OAI211_X1 U6380 ( .C1(n5992), .C2(n5257), .A(n5256), .B(n5255), .ZN(n5258)
         );
  AOI21_X1 U6381 ( .B1(n5377), .B2(n5951), .A(n5258), .ZN(n5259) );
  INV_X1 U6382 ( .A(n5259), .ZN(U2797) );
  INV_X1 U6383 ( .A(n5399), .ZN(n5322) );
  INV_X1 U6384 ( .A(n5263), .ZN(n5265) );
  AOI21_X1 U6385 ( .B1(n5265), .B2(n3174), .A(n5264), .ZN(n5266) );
  AND2_X1 U6386 ( .A1(n5328), .A2(n5266), .ZN(n5267) );
  NOR2_X1 U6387 ( .A1(n5268), .A2(n5267), .ZN(n5523) );
  AOI21_X1 U6388 ( .B1(n6909), .B2(n5270), .A(n5269), .ZN(n5271) );
  AOI21_X1 U6389 ( .B1(n5980), .B2(EBX_REG_29__SCAN_IN), .A(n5271), .ZN(n5272)
         );
  INV_X1 U6390 ( .A(n5272), .ZN(n5275) );
  INV_X1 U6391 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5273) );
  OAI22_X1 U6392 ( .A1(n5273), .A2(n5872), .B1(n5397), .B2(n5988), .ZN(n5274)
         );
  AOI211_X1 U6393 ( .C1(n5965), .C2(n5523), .A(n5275), .B(n5274), .ZN(n5276)
         );
  OAI21_X1 U6394 ( .B1(n5322), .B2(n5937), .A(n5276), .ZN(U2798) );
  NOR2_X1 U6395 ( .A1(n5279), .A2(n5280), .ZN(n5281) );
  OR2_X1 U6396 ( .A1(n5277), .A2(n5281), .ZN(n5450) );
  INV_X1 U6397 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6784) );
  NAND2_X1 U6398 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5297), .ZN(n5731) );
  INV_X1 U6399 ( .A(REIP_REG_23__SCAN_IN), .ZN(n7060) );
  OAI21_X1 U6400 ( .B1(n6784), .B2(n5731), .A(n7060), .ZN(n5290) );
  AND2_X1 U6401 ( .A1(n5989), .A2(n5282), .ZN(n5716) );
  NAND2_X1 U6402 ( .A1(n5283), .A2(n5284), .ZN(n5285) );
  NAND2_X1 U6403 ( .A1(n5350), .A2(n5285), .ZN(n5572) );
  INV_X1 U6404 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5286) );
  OAI22_X1 U6405 ( .A1(n5286), .A2(n6000), .B1(n5452), .B2(n5988), .ZN(n5287)
         );
  AOI21_X1 U6406 ( .B1(n5997), .B2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n5287), 
        .ZN(n5288) );
  OAI21_X1 U6407 ( .B1(n5572), .B2(n5992), .A(n5288), .ZN(n5289) );
  AOI21_X1 U6408 ( .B1(n5290), .B2(n5716), .A(n5289), .ZN(n5291) );
  OAI21_X1 U6409 ( .B1(n5450), .B2(n5937), .A(n5291), .ZN(U2804) );
  NAND2_X1 U6410 ( .A1(n5294), .A2(n5295), .ZN(n5296) );
  AND2_X1 U6411 ( .A1(n5293), .A2(n5296), .ZN(n5761) );
  INV_X1 U6412 ( .A(n5761), .ZN(n5360) );
  INV_X1 U6413 ( .A(REIP_REG_21__SCAN_IN), .ZN(n7026) );
  NAND2_X1 U6414 ( .A1(n5297), .A2(n7026), .ZN(n5737) );
  AND2_X1 U6415 ( .A1(n5299), .A2(n5298), .ZN(n5300) );
  OR2_X1 U6416 ( .A1(n5300), .A2(n5356), .ZN(n5588) );
  INV_X1 U6417 ( .A(n5588), .ZN(n5306) );
  INV_X1 U6418 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5361) );
  OAI22_X1 U6419 ( .A1(n5361), .A2(n6000), .B1(n5301), .B2(n5872), .ZN(n5305)
         );
  OR2_X1 U6420 ( .A1(n5303), .A2(n5302), .ZN(n5738) );
  OAI22_X1 U6421 ( .A1(n5467), .A2(n5988), .B1(n7026), .B2(n5738), .ZN(n5304)
         );
  AOI211_X1 U6422 ( .C1(n5306), .C2(n5965), .A(n5305), .B(n5304), .ZN(n5307)
         );
  OAI211_X1 U6423 ( .C1(n5360), .C2(n5937), .A(n5737), .B(n5307), .ZN(U2806)
         );
  XOR2_X1 U6424 ( .A(n5310), .B(n5309), .Z(n5764) );
  INV_X1 U6425 ( .A(n5764), .ZN(n5363) );
  MUX2_X1 U6426 ( .A(n3174), .B(n5366), .S(n5367), .Z(n5312) );
  XNOR2_X1 U6427 ( .A(n5312), .B(n5311), .ZN(n5600) );
  INV_X1 U6428 ( .A(n5600), .ZN(n5317) );
  INV_X1 U6429 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5474) );
  AOI22_X1 U6430 ( .A1(EBX_REG_20__SCAN_IN), .A2(n5980), .B1(n5472), .B2(n5996), .ZN(n5313) );
  OAI21_X1 U6431 ( .B1(n5474), .B2(n5872), .A(n5313), .ZN(n5316) );
  AOI21_X1 U6432 ( .B1(n6783), .B2(n5314), .A(n5738), .ZN(n5315) );
  AOI211_X1 U6433 ( .C1(n5317), .C2(n5965), .A(n5316), .B(n5315), .ZN(n5318)
         );
  OAI21_X1 U6434 ( .B1(n5363), .B2(n5937), .A(n5318), .ZN(U2807) );
  INV_X1 U6435 ( .A(n5517), .ZN(n5320) );
  INV_X1 U6436 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5319) );
  OAI22_X1 U6437 ( .A1(n5320), .A2(n6011), .B1(n5319), .B2(n6022), .ZN(U2828)
         );
  AOI22_X1 U6438 ( .A1(n5523), .A2(n6018), .B1(n5371), .B2(EBX_REG_29__SCAN_IN), .ZN(n5321) );
  OAI21_X1 U6439 ( .B1(n5322), .B2(n6012), .A(n5321), .ZN(U2830) );
  OR2_X1 U6440 ( .A1(n5417), .A2(n5324), .ZN(n5325) );
  INV_X1 U6441 ( .A(n6012), .ZN(n6019) );
  NAND2_X1 U6442 ( .A1(n5545), .A2(n5326), .ZN(n5327) );
  NAND2_X1 U6443 ( .A1(n5328), .A2(n5327), .ZN(n5683) );
  OAI22_X1 U6444 ( .A1(n5683), .A2(n6011), .B1(n5329), .B2(n6022), .ZN(n5330)
         );
  AOI21_X1 U6445 ( .B1(n5685), .B2(n6019), .A(n5330), .ZN(n5331) );
  INV_X1 U6446 ( .A(n5331), .ZN(U2831) );
  AOI21_X1 U6447 ( .B1(n5334), .B2(n5332), .A(n5333), .ZN(n5428) );
  OR2_X1 U6448 ( .A1(n5345), .A2(n5335), .ZN(n5336) );
  NAND2_X1 U6449 ( .A1(n5543), .A2(n5336), .ZN(n5700) );
  OAI22_X1 U6450 ( .A1(n5700), .A2(n6011), .B1(n5707), .B2(n6022), .ZN(n5337)
         );
  AOI21_X1 U6451 ( .B1(n5428), .B2(n6019), .A(n5337), .ZN(n5338) );
  INV_X1 U6452 ( .A(n5338), .ZN(U2833) );
  INV_X1 U6453 ( .A(n5332), .ZN(n5341) );
  AOI21_X1 U6454 ( .B1(n5342), .B2(n5340), .A(n5341), .ZN(n5770) );
  INV_X1 U6455 ( .A(n5770), .ZN(n5347) );
  INV_X1 U6456 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5346) );
  NOR2_X1 U6457 ( .A1(n5351), .A2(n5343), .ZN(n5344) );
  OR2_X1 U6458 ( .A1(n5345), .A2(n5344), .ZN(n5709) );
  OAI222_X1 U6459 ( .A1(n5347), .A2(n6012), .B1(n6022), .B2(n5346), .C1(n5709), 
        .C2(n6011), .ZN(U2834) );
  OAI21_X1 U6460 ( .B1(n5277), .B2(n5348), .A(n5340), .ZN(n5439) );
  AND2_X1 U6461 ( .A1(n5350), .A2(n5349), .ZN(n5352) );
  OR2_X1 U6462 ( .A1(n5352), .A2(n5351), .ZN(n5728) );
  OAI222_X1 U6463 ( .A1(n6012), .A2(n5439), .B1(n6022), .B2(n5721), .C1(n5728), 
        .C2(n6011), .ZN(U2835) );
  INV_X1 U6464 ( .A(n5572), .ZN(n5353) );
  AOI22_X1 U6465 ( .A1(n6018), .A2(n5353), .B1(n5371), .B2(EBX_REG_23__SCAN_IN), .ZN(n5354) );
  OAI21_X1 U6466 ( .B1(n5450), .B2(n6012), .A(n5354), .ZN(U2836) );
  OR2_X1 U6467 ( .A1(n5356), .A2(n5355), .ZN(n5357) );
  NAND2_X1 U6468 ( .A1(n5283), .A2(n5357), .ZN(n5732) );
  INV_X1 U6469 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5359) );
  AOI21_X1 U6470 ( .B1(n5358), .B2(n5293), .A(n5279), .ZN(n5461) );
  INV_X1 U6471 ( .A(n5461), .ZN(n5733) );
  OAI222_X1 U6472 ( .A1(n6011), .A2(n5732), .B1(n6022), .B2(n5359), .C1(n5733), 
        .C2(n6012), .ZN(U2837) );
  OAI222_X1 U6473 ( .A1(n5588), .A2(n6011), .B1(n6022), .B2(n5361), .C1(n6012), 
        .C2(n5360), .ZN(U2838) );
  OAI222_X1 U6474 ( .A1(n5363), .A2(n6012), .B1(n6022), .B2(n5362), .C1(n6011), 
        .C2(n5600), .ZN(U2839) );
  AOI21_X1 U6475 ( .B1(n5364), .B2(n4819), .A(n5309), .ZN(n5775) );
  INV_X1 U6476 ( .A(n5775), .ZN(n5374) );
  MUX2_X1 U6477 ( .A(n5366), .B(n5365), .S(n3475), .Z(n5376) );
  INV_X1 U6478 ( .A(n5367), .ZN(n5370) );
  INV_X1 U6479 ( .A(n5629), .ZN(n5375) );
  NOR2_X1 U6480 ( .A1(n5375), .A2(n5376), .ZN(n5369) );
  OAI22_X1 U6481 ( .A1(n5376), .A2(n5370), .B1(n5369), .B2(n5368), .ZN(n5750)
         );
  INV_X1 U6482 ( .A(n5750), .ZN(n5372) );
  AOI22_X1 U6483 ( .A1(n6018), .A2(n5372), .B1(n5371), .B2(EBX_REG_19__SCAN_IN), .ZN(n5373) );
  OAI21_X1 U6484 ( .B1(n5374), .B2(n6012), .A(n5373), .ZN(U2840) );
  XNOR2_X1 U6485 ( .A(n5376), .B(n5375), .ZN(n5859) );
  OAI222_X1 U6486 ( .A1(n5859), .A2(n6011), .B1(n6022), .B2(n5851), .C1(n6012), 
        .C2(n5855), .ZN(U2841) );
  NAND2_X1 U6487 ( .A1(n5377), .A2(n6030), .ZN(n5379) );
  AOI22_X1 U6488 ( .A1(n6029), .A2(DATAI_30_), .B1(n6025), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5378) );
  OAI211_X1 U6489 ( .C1(n6033), .C2(n6099), .A(n5379), .B(n5378), .ZN(U2861)
         );
  NAND2_X1 U6490 ( .A1(n5399), .A2(n6030), .ZN(n5381) );
  AOI22_X1 U6491 ( .A1(n6029), .A2(DATAI_29_), .B1(n6025), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5380) );
  OAI211_X1 U6492 ( .C1(n6033), .C2(n6993), .A(n5381), .B(n5380), .ZN(U2862)
         );
  INV_X1 U6493 ( .A(n5685), .ZN(n5384) );
  AOI22_X1 U6494 ( .A1(n6026), .A2(DATAI_12_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n6025), .ZN(n5383) );
  NAND2_X1 U6495 ( .A1(n6029), .A2(DATAI_28_), .ZN(n5382) );
  OAI211_X1 U6496 ( .C1(n5384), .C2(n5391), .A(n5383), .B(n5382), .ZN(U2863)
         );
  INV_X1 U6497 ( .A(n5428), .ZN(n5701) );
  AOI22_X1 U6498 ( .A1(n6026), .A2(DATAI_10_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n6025), .ZN(n5386) );
  NAND2_X1 U6499 ( .A1(n6029), .A2(DATAI_26_), .ZN(n5385) );
  OAI211_X1 U6500 ( .C1(n5701), .C2(n5391), .A(n5386), .B(n5385), .ZN(U2865)
         );
  AOI22_X1 U6501 ( .A1(n6026), .A2(DATAI_8_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n6025), .ZN(n5388) );
  NAND2_X1 U6502 ( .A1(n6029), .A2(DATAI_24_), .ZN(n5387) );
  OAI211_X1 U6503 ( .C1(n5439), .C2(n5391), .A(n5388), .B(n5387), .ZN(U2867)
         );
  AOI22_X1 U6504 ( .A1(n6026), .A2(DATAI_6_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n6025), .ZN(n5390) );
  NAND2_X1 U6505 ( .A1(n6029), .A2(DATAI_22_), .ZN(n5389) );
  OAI211_X1 U6506 ( .C1(n5733), .C2(n5391), .A(n5390), .B(n5389), .ZN(U2869)
         );
  NAND2_X1 U6507 ( .A1(n5401), .A2(n5393), .ZN(n5394) );
  NAND2_X1 U6508 ( .A1(n5392), .A2(n5394), .ZN(n5395) );
  XNOR2_X1 U6509 ( .A(n5395), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5533)
         );
  NOR2_X1 U6510 ( .A1(n5819), .A2(n6909), .ZN(n5526) );
  AOI21_X1 U6511 ( .B1(n6117), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5526), 
        .ZN(n5396) );
  OAI21_X1 U6512 ( .B1(n5397), .B2(n6111), .A(n5396), .ZN(n5398) );
  AOI21_X1 U6513 ( .B1(n5399), .B2(n6113), .A(n5398), .ZN(n5400) );
  OAI21_X1 U6514 ( .B1(n5533), .B2(n5835), .A(n5400), .ZN(U2957) );
  INV_X2 U6515 ( .A(n5401), .ZN(n5424) );
  NAND3_X1 U6516 ( .A1(n5424), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n3150), .ZN(n5405) );
  BUF_X1 U6517 ( .A(n5402), .Z(n5403) );
  NOR2_X1 U6518 ( .A1(n5422), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5404)
         );
  NAND2_X1 U6519 ( .A1(n5403), .A2(n5404), .ZN(n5411) );
  AOI22_X2 U6520 ( .A1(n5405), .A2(n5411), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5555), .ZN(n5406) );
  XNOR2_X1 U6521 ( .A(n5406), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5541)
         );
  NAND2_X1 U6522 ( .A1(n5781), .A2(n5682), .ZN(n5407) );
  NAND2_X1 U6523 ( .A1(n6176), .A2(REIP_REG_28__SCAN_IN), .ZN(n5534) );
  OAI211_X1 U6524 ( .C1(n5786), .C2(n5408), .A(n5407), .B(n5534), .ZN(n5409)
         );
  AOI21_X1 U6525 ( .B1(n5685), .B2(n6113), .A(n5409), .ZN(n5410) );
  OAI21_X1 U6526 ( .B1(n5835), .B2(n5541), .A(n5410), .ZN(U2958) );
  INV_X1 U6527 ( .A(n5411), .ZN(n5412) );
  OR2_X1 U6528 ( .A1(n5413), .A2(n5412), .ZN(n5414) );
  XNOR2_X1 U6529 ( .A(n5414), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5553)
         );
  NOR2_X1 U6530 ( .A1(n5333), .A2(n5415), .ZN(n5416) );
  NAND2_X1 U6531 ( .A1(n6176), .A2(REIP_REG_27__SCAN_IN), .ZN(n5547) );
  NAND2_X1 U6532 ( .A1(n6117), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5418)
         );
  OAI211_X1 U6533 ( .C1(n6111), .C2(n5690), .A(n5547), .B(n5418), .ZN(n5419)
         );
  AOI21_X1 U6534 ( .B1(n3183), .B2(n6113), .A(n5419), .ZN(n5420) );
  OAI21_X1 U6535 ( .B1(n5553), .B2(n5835), .A(n5420), .ZN(U2959) );
  NAND2_X1 U6536 ( .A1(n5422), .A2(n5421), .ZN(n5423) );
  XNOR2_X1 U6537 ( .A(n5424), .B(n5423), .ZN(n5561) );
  INV_X1 U6538 ( .A(n5698), .ZN(n5426) );
  NAND2_X1 U6539 ( .A1(n6117), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5425)
         );
  NAND2_X1 U6540 ( .A1(n5969), .A2(REIP_REG_26__SCAN_IN), .ZN(n5556) );
  OAI211_X1 U6541 ( .C1(n6111), .C2(n5426), .A(n5425), .B(n5556), .ZN(n5427)
         );
  AOI21_X1 U6542 ( .B1(n5428), .B2(n6113), .A(n5427), .ZN(n5429) );
  OAI21_X1 U6543 ( .B1(n5561), .B2(n5835), .A(n5429), .ZN(U2960) );
  NAND2_X1 U6544 ( .A1(n3150), .A2(n5609), .ZN(n5430) );
  AOI21_X2 U6545 ( .B1(n5443), .B2(n5430), .A(n3186), .ZN(n5470) );
  XNOR2_X1 U6546 ( .A(n5432), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5471)
         );
  INV_X1 U6547 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5431) );
  AOI21_X1 U6548 ( .B1(n5470), .B2(n5471), .A(n3184), .ZN(n5465) );
  XNOR2_X1 U6549 ( .A(n5489), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5464)
         );
  INV_X1 U6550 ( .A(n5435), .ZN(n5463) );
  NOR2_X1 U6551 ( .A1(n3150), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5455)
         );
  NAND2_X1 U6552 ( .A1(n5463), .A2(n5455), .ZN(n5448) );
  NAND2_X1 U6553 ( .A1(n5432), .A2(n5433), .ZN(n5434) );
  INV_X1 U6554 ( .A(n5457), .ZN(n5436) );
  NAND2_X1 U6555 ( .A1(n5436), .A2(n3180), .ZN(n5437) );
  XNOR2_X1 U6556 ( .A(n5438), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5568)
         );
  INV_X1 U6557 ( .A(n5439), .ZN(n5723) );
  NAND2_X1 U6558 ( .A1(n6176), .A2(REIP_REG_24__SCAN_IN), .ZN(n5564) );
  NAND2_X1 U6559 ( .A1(n6117), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5440)
         );
  OAI211_X1 U6560 ( .C1(n6111), .C2(n5717), .A(n5564), .B(n5440), .ZN(n5441)
         );
  AOI21_X1 U6561 ( .B1(n5723), .B2(n6113), .A(n5441), .ZN(n5442) );
  OAI21_X1 U6562 ( .B1(n5568), .B2(n5835), .A(n5442), .ZN(U2962) );
  INV_X1 U6563 ( .A(n5445), .ZN(n5446) );
  NAND3_X1 U6564 ( .A1(n5444), .A2(n5446), .A3(n3150), .ZN(n5447) );
  NAND2_X1 U6565 ( .A1(n5448), .A2(n5447), .ZN(n5449) );
  XNOR2_X1 U6566 ( .A(n5449), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5577)
         );
  INV_X1 U6567 ( .A(n5450), .ZN(n5758) );
  NAND2_X1 U6568 ( .A1(n6176), .A2(REIP_REG_23__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U6569 ( .A1(n6117), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5451)
         );
  OAI211_X1 U6570 ( .C1(n6111), .C2(n5452), .A(n5570), .B(n5451), .ZN(n5453)
         );
  AOI21_X1 U6571 ( .B1(n5758), .B2(n6113), .A(n5453), .ZN(n5454) );
  OAI21_X1 U6572 ( .B1(n5577), .B2(n5835), .A(n5454), .ZN(U2963) );
  AOI21_X1 U6573 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n3150), .A(n5455), 
        .ZN(n5456) );
  XNOR2_X1 U6574 ( .A(n5457), .B(n5456), .ZN(n5586) );
  NAND2_X1 U6575 ( .A1(n5781), .A2(n5729), .ZN(n5458) );
  NAND2_X1 U6576 ( .A1(n5969), .A2(REIP_REG_22__SCAN_IN), .ZN(n5579) );
  OAI211_X1 U6577 ( .C1(n5786), .C2(n5459), .A(n5458), .B(n5579), .ZN(n5460)
         );
  AOI21_X1 U6578 ( .B1(n5461), .B2(n6113), .A(n5460), .ZN(n5462) );
  OAI21_X1 U6579 ( .B1(n5586), .B2(n5835), .A(n5462), .ZN(U2964) );
  AOI21_X1 U6580 ( .B1(n5465), .B2(n5464), .A(n5463), .ZN(n5594) );
  NAND2_X1 U6581 ( .A1(n5969), .A2(REIP_REG_21__SCAN_IN), .ZN(n5587) );
  NAND2_X1 U6582 ( .A1(n6117), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5466)
         );
  OAI211_X1 U6583 ( .C1(n6111), .C2(n5467), .A(n5587), .B(n5466), .ZN(n5468)
         );
  AOI21_X1 U6584 ( .B1(n5761), .B2(n6113), .A(n5468), .ZN(n5469) );
  OAI21_X1 U6585 ( .B1(n5594), .B2(n5835), .A(n5469), .ZN(U2965) );
  XOR2_X1 U6586 ( .A(n5471), .B(n5470), .Z(n5608) );
  NAND2_X1 U6587 ( .A1(n5781), .A2(n5472), .ZN(n5473) );
  NAND2_X1 U6588 ( .A1(n5969), .A2(REIP_REG_20__SCAN_IN), .ZN(n5599) );
  OAI211_X1 U6589 ( .C1(n5786), .C2(n5474), .A(n5473), .B(n5599), .ZN(n5475)
         );
  AOI21_X1 U6590 ( .B1(n5764), .B2(n6113), .A(n5475), .ZN(n5476) );
  OAI21_X1 U6591 ( .B1(n5608), .B2(n5835), .A(n5476), .ZN(U2966) );
  NOR3_X1 U6592 ( .A1(n5478), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n3150), 
        .ZN(n5625) );
  NOR3_X1 U6593 ( .A1(n5479), .A2(n5489), .A3(n5481), .ZN(n5480) );
  AOI21_X1 U6594 ( .B1(n5625), .B2(n5481), .A(n5480), .ZN(n5483) );
  XNOR2_X1 U6595 ( .A(n5483), .B(n5482), .ZN(n5624) );
  INV_X1 U6596 ( .A(n5857), .ZN(n5485) );
  AOI22_X1 U6597 ( .A1(n6117), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .B1(n5969), 
        .B2(REIP_REG_18__SCAN_IN), .ZN(n5484) );
  OAI21_X1 U6598 ( .B1(n5485), .B2(n6111), .A(n5484), .ZN(n5486) );
  AOI21_X1 U6599 ( .B1(n5487), .B2(n6113), .A(n5486), .ZN(n5488) );
  OAI21_X1 U6600 ( .B1(n5624), .B2(n5835), .A(n5488), .ZN(U2968) );
  NOR2_X1 U6601 ( .A1(n5489), .A2(n4786), .ZN(n5491) );
  MUX2_X1 U6602 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .B(n4786), .S(n3150), 
        .Z(n5490) );
  MUX2_X1 U6603 ( .A(n5491), .B(n5490), .S(n5478), .Z(n5492) );
  NOR2_X1 U6604 ( .A1(n5625), .A2(n5492), .ZN(n5796) );
  AOI22_X1 U6605 ( .A1(n6117), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n5969), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n5493) );
  OAI21_X1 U6606 ( .B1(n5875), .B2(n6111), .A(n5493), .ZN(n5494) );
  AOI21_X1 U6607 ( .B1(n6031), .B2(n6113), .A(n5494), .ZN(n5495) );
  OAI21_X1 U6608 ( .B1(n5796), .B2(n5835), .A(n5495), .ZN(U2970) );
  XNOR2_X1 U6609 ( .A(n5432), .B(n5497), .ZN(n5498) );
  XNOR2_X1 U6610 ( .A(n5499), .B(n5498), .ZN(n5803) );
  INV_X1 U6611 ( .A(n6006), .ZN(n5503) );
  AOI22_X1 U6612 ( .A1(n6117), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n5969), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n5500) );
  OAI21_X1 U6613 ( .B1(n5501), .B2(n6111), .A(n5500), .ZN(n5502) );
  AOI21_X1 U6614 ( .B1(n5503), .B2(n6113), .A(n5502), .ZN(n5504) );
  OAI21_X1 U6615 ( .B1(n5803), .B2(n5835), .A(n5504), .ZN(U2971) );
  XNOR2_X1 U6616 ( .A(n5432), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5506)
         );
  XNOR2_X1 U6617 ( .A(n5505), .B(n5506), .ZN(n5638) );
  NAND2_X1 U6618 ( .A1(n5638), .A2(n6115), .ZN(n5510) );
  NOR2_X1 U6619 ( .A1(n5819), .A2(n6778), .ZN(n5657) );
  NOR2_X1 U6620 ( .A1(n6111), .A2(n5507), .ZN(n5508) );
  AOI211_X1 U6621 ( .C1(n6117), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n5657), 
        .B(n5508), .ZN(n5509) );
  OAI211_X1 U6622 ( .C1(n5512), .C2(n5511), .A(n5510), .B(n5509), .ZN(U2972)
         );
  NAND2_X1 U6623 ( .A1(n6170), .A2(n4797), .ZN(n5513) );
  AOI21_X1 U6624 ( .B1(n5514), .B2(n5513), .A(n5518), .ZN(n5515) );
  AOI211_X1 U6625 ( .C1(n5517), .C2(n6172), .A(n5516), .B(n5515), .ZN(n5521)
         );
  NAND3_X1 U6626 ( .A1(n5519), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5518), .ZN(n5520) );
  OAI211_X1 U6627 ( .C1(n5522), .C2(n6125), .A(n5521), .B(n5520), .ZN(U2987)
         );
  INV_X1 U6628 ( .A(n5523), .ZN(n5524) );
  NOR2_X1 U6629 ( .A1(n5524), .A2(n6163), .ZN(n5525) );
  INV_X1 U6630 ( .A(n5528), .ZN(n5551) );
  NAND3_X1 U6631 ( .A1(n5551), .A2(n5530), .A3(n5529), .ZN(n5531) );
  OAI211_X1 U6632 ( .C1(n5533), .C2(n6125), .A(n5532), .B(n5531), .ZN(U2989)
         );
  INV_X1 U6633 ( .A(n5548), .ZN(n5536) );
  OAI21_X1 U6634 ( .B1(n5683), .B2(n6163), .A(n5534), .ZN(n5535) );
  AOI21_X1 U6635 ( .B1(n5536), .B2(INSTADDRPOINTER_REG_28__SCAN_IN), .A(n5535), 
        .ZN(n5540) );
  NAND3_X1 U6636 ( .A1(n5551), .A2(n5538), .A3(n5537), .ZN(n5539) );
  OAI211_X1 U6637 ( .C1(n5541), .C2(n6125), .A(n5540), .B(n5539), .ZN(U2990)
         );
  NAND2_X1 U6638 ( .A1(n5543), .A2(n5542), .ZN(n5544) );
  AND2_X1 U6639 ( .A1(n5545), .A2(n5544), .ZN(n5751) );
  NAND2_X1 U6640 ( .A1(n5751), .A2(n6172), .ZN(n5546) );
  OAI211_X1 U6641 ( .C1(n5548), .C2(n5550), .A(n5547), .B(n5546), .ZN(n5549)
         );
  AOI21_X1 U6642 ( .B1(n5551), .B2(n5550), .A(n5549), .ZN(n5552) );
  OAI21_X1 U6643 ( .B1(n5553), .B2(n6125), .A(n5552), .ZN(U2991) );
  AOI21_X1 U6644 ( .B1(n5555), .B2(n5791), .A(n5554), .ZN(n5559) );
  NAND2_X1 U6645 ( .A1(n5790), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5557) );
  OAI211_X1 U6646 ( .C1(n6163), .C2(n5700), .A(n5557), .B(n5556), .ZN(n5558)
         );
  AOI21_X1 U6647 ( .B1(n5792), .B2(n5559), .A(n5558), .ZN(n5560) );
  OAI21_X1 U6648 ( .B1(n5561), .B2(n6125), .A(n5560), .ZN(U2992) );
  INV_X1 U6649 ( .A(n5575), .ZN(n5563) );
  OAI21_X1 U6650 ( .B1(n5563), .B2(n5574), .A(n5562), .ZN(n5566) );
  OAI21_X1 U6651 ( .B1(n6163), .B2(n5728), .A(n5564), .ZN(n5565) );
  AOI21_X1 U6652 ( .B1(n5566), .B2(n5790), .A(n5565), .ZN(n5567) );
  OAI21_X1 U6653 ( .B1(n5568), .B2(n6125), .A(n5567), .ZN(U2994) );
  NAND2_X1 U6654 ( .A1(n5569), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5571) );
  OAI211_X1 U6655 ( .C1(n6163), .C2(n5572), .A(n5571), .B(n5570), .ZN(n5573)
         );
  AOI21_X1 U6656 ( .B1(n5575), .B2(n5574), .A(n5573), .ZN(n5576) );
  OAI21_X1 U6657 ( .B1(n5577), .B2(n6125), .A(n5576), .ZN(U2995) );
  INV_X1 U6658 ( .A(n5578), .ZN(n5592) );
  OAI21_X1 U6659 ( .B1(n6163), .B2(n5732), .A(n5579), .ZN(n5584) );
  INV_X1 U6660 ( .A(n5580), .ZN(n5589) );
  NOR3_X1 U6661 ( .A1(n5589), .A2(n5582), .A3(n5581), .ZN(n5583) );
  AOI211_X1 U6662 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n5592), .A(n5584), .B(n5583), .ZN(n5585) );
  OAI21_X1 U6663 ( .B1(n5586), .B2(n6125), .A(n5585), .ZN(U2996) );
  OAI21_X1 U6664 ( .B1(n6163), .B2(n5588), .A(n5587), .ZN(n5591) );
  NOR2_X1 U6665 ( .A1(n5589), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5590)
         );
  AOI211_X1 U6666 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5592), .A(n5591), .B(n5590), .ZN(n5593) );
  OAI21_X1 U6667 ( .B1(n5594), .B2(n6125), .A(n5593), .ZN(U2997) );
  AOI221_X1 U6668 ( .B1(n5642), .B2(n5643), .C1(n5595), .C2(n5643), .A(n5641), 
        .ZN(n5596) );
  OAI221_X1 U6669 ( .B1(n5645), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .C1(
        n5645), .C2(n5597), .A(n5596), .ZN(n5632) );
  AOI21_X1 U6670 ( .B1(n6157), .B2(n5481), .A(n5632), .ZN(n5618) );
  OAI21_X1 U6671 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5598), .A(n5618), 
        .ZN(n5613) );
  INV_X1 U6672 ( .A(n5599), .ZN(n5602) );
  NOR2_X1 U6673 ( .A1(n6163), .A2(n5600), .ZN(n5601) );
  AOI211_X1 U6674 ( .C1(INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n5613), .A(n5602), .B(n5601), .ZN(n5607) );
  OR4_X1 U6675 ( .A1(n5634), .A2(n5605), .A3(n5604), .A4(n5603), .ZN(n5606) );
  OAI211_X1 U6676 ( .C1(n5608), .C2(n6125), .A(n5607), .B(n5606), .ZN(U2998)
         );
  XNOR2_X1 U6677 ( .A(n5432), .B(n5609), .ZN(n5610) );
  XNOR2_X1 U6678 ( .A(n5444), .B(n5610), .ZN(n5774) );
  INV_X1 U6679 ( .A(n5634), .ZN(n5612) );
  NAND3_X1 U6680 ( .A1(n5612), .A2(n5611), .A3(n5609), .ZN(n5615) );
  AOI22_X1 U6681 ( .A1(n5969), .A2(REIP_REG_19__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n5613), .ZN(n5614) );
  OAI211_X1 U6682 ( .C1(n6163), .C2(n5750), .A(n5615), .B(n5614), .ZN(n5616)
         );
  AOI21_X1 U6683 ( .B1(n5774), .B2(n6175), .A(n5616), .ZN(n5617) );
  INV_X1 U6684 ( .A(n5617), .ZN(U2999) );
  NOR3_X1 U6685 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n5481), .A3(n5634), 
        .ZN(n5620) );
  NOR2_X1 U6686 ( .A1(n5482), .A2(n5618), .ZN(n5619) );
  AOI211_X1 U6687 ( .C1(n6176), .C2(REIP_REG_18__SCAN_IN), .A(n5620), .B(n5619), .ZN(n5623) );
  INV_X1 U6688 ( .A(n5859), .ZN(n5621) );
  NAND2_X1 U6689 ( .A1(n6172), .A2(n5621), .ZN(n5622) );
  OAI211_X1 U6690 ( .C1(n5624), .C2(n6125), .A(n5623), .B(n5622), .ZN(U3000)
         );
  INV_X1 U6691 ( .A(n5625), .ZN(n5627) );
  NAND3_X1 U6692 ( .A1(n5478), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n3150), .ZN(n5626) );
  NAND2_X1 U6693 ( .A1(n5627), .A2(n5626), .ZN(n5628) );
  XNOR2_X1 U6694 ( .A(n5628), .B(n5481), .ZN(n5783) );
  INV_X1 U6695 ( .A(n5783), .ZN(n5637) );
  AOI21_X1 U6696 ( .B1(n5631), .B2(n5630), .A(n5629), .ZN(n6002) );
  INV_X1 U6697 ( .A(n5632), .ZN(n5633) );
  NAND2_X1 U6698 ( .A1(n6176), .A2(REIP_REG_17__SCAN_IN), .ZN(n5784) );
  OAI221_X1 U6699 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5634), .C1(
        n5481), .C2(n5633), .A(n5784), .ZN(n5635) );
  AOI21_X1 U6700 ( .B1(n6002), .B2(n6172), .A(n5635), .ZN(n5636) );
  OAI21_X1 U6701 ( .B1(n5637), .B2(n6125), .A(n5636), .ZN(U3001) );
  INV_X1 U6702 ( .A(n5638), .ZN(n5661) );
  NOR2_X1 U6703 ( .A1(n5813), .A2(n5639), .ZN(n5647) );
  INV_X1 U6704 ( .A(n5640), .ZN(n5646) );
  AOI21_X1 U6705 ( .B1(n5643), .B2(n5642), .A(n5641), .ZN(n5644) );
  OAI21_X1 U6706 ( .B1(n5646), .B2(n5645), .A(n5644), .ZN(n6134) );
  AOI211_X1 U6707 ( .C1(n5648), .C2(n5654), .A(n5647), .B(n6134), .ZN(n5815)
         );
  INV_X1 U6708 ( .A(n5649), .ZN(n5650) );
  OAI21_X1 U6709 ( .B1(n5651), .B2(n5650), .A(n5814), .ZN(n5653) );
  AOI21_X1 U6710 ( .B1(n5815), .B2(n5653), .A(n5652), .ZN(n5659) );
  NOR3_X1 U6711 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6138), .A3(n5654), 
        .ZN(n5658) );
  NOR2_X1 U6712 ( .A1(n6163), .A2(n5655), .ZN(n5656) );
  NOR4_X1 U6713 ( .A1(n5659), .A2(n5658), .A3(n5657), .A4(n5656), .ZN(n5660)
         );
  OAI21_X1 U6714 ( .B1(n5661), .B2(n6125), .A(n5660), .ZN(U3004) );
  NAND3_X1 U6715 ( .A1(n5664), .A2(n5663), .A3(n5662), .ZN(n5665) );
  OAI21_X1 U6716 ( .B1(n5666), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n5665), 
        .ZN(n5667) );
  AOI21_X1 U6717 ( .B1(n6181), .B2(n5668), .A(n5667), .ZN(n6699) );
  NOR3_X1 U6718 ( .A1(n5670), .A2(n5669), .A3(n6733), .ZN(n5671) );
  AOI21_X1 U6719 ( .B1(n5673), .B2(n5672), .A(n5671), .ZN(n5674) );
  OAI21_X1 U6720 ( .B1(n6699), .B2(n5677), .A(n5674), .ZN(n5675) );
  MUX2_X1 U6721 ( .A(n5675), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(n5679), 
        .Z(U3460) );
  OAI22_X1 U6722 ( .A1(n5678), .A2(n5677), .B1(n6733), .B2(n5676), .ZN(n5680)
         );
  MUX2_X1 U6723 ( .A(n5680), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n5679), 
        .Z(U3456) );
  AOI22_X1 U6724 ( .A1(EBX_REG_28__SCAN_IN), .A2(n5980), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n5997), .ZN(n5689) );
  AOI22_X1 U6725 ( .A1(n5682), .A2(n5996), .B1(REIP_REG_28__SCAN_IN), .B2(
        n5681), .ZN(n5688) );
  NOR2_X1 U6726 ( .A1(n5683), .A2(n5992), .ZN(n5684) );
  AOI21_X1 U6727 ( .B1(n5685), .B2(n5951), .A(n5684), .ZN(n5687) );
  NAND3_X1 U6728 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5695), .A3(n6786), .ZN(
        n5686) );
  NAND4_X1 U6729 ( .A1(n5689), .A2(n5688), .A3(n5687), .A4(n5686), .ZN(U2799)
         );
  INV_X1 U6730 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5691) );
  OAI22_X1 U6731 ( .A1(n5691), .A2(n5872), .B1(n5988), .B2(n5690), .ZN(n5692)
         );
  AOI21_X1 U6732 ( .B1(n5980), .B2(EBX_REG_27__SCAN_IN), .A(n5692), .ZN(n5693)
         );
  OAI21_X1 U6733 ( .B1(n5699), .B2(n7012), .A(n5693), .ZN(n5694) );
  AOI21_X1 U6734 ( .B1(n3183), .B2(n5951), .A(n5694), .ZN(n5697) );
  AOI22_X1 U6735 ( .A1(n5965), .A2(n5751), .B1(n5695), .B2(n7012), .ZN(n5696)
         );
  NAND2_X1 U6736 ( .A1(n5697), .A2(n5696), .ZN(U2800) );
  AOI22_X1 U6737 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n5997), .B1(n5698), 
        .B2(n5996), .ZN(n5706) );
  INV_X1 U6738 ( .A(n5699), .ZN(n5704) );
  NAND2_X1 U6739 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n5711) );
  INV_X1 U6740 ( .A(REIP_REG_26__SCAN_IN), .ZN(n7053) );
  OAI21_X1 U6741 ( .B1(n5710), .B2(n5711), .A(n7053), .ZN(n5703) );
  OAI22_X1 U6742 ( .A1(n5701), .A2(n5937), .B1(n5992), .B2(n5700), .ZN(n5702)
         );
  AOI21_X1 U6743 ( .B1(n5704), .B2(n5703), .A(n5702), .ZN(n5705) );
  OAI211_X1 U6744 ( .C1(n5707), .C2(n6000), .A(n5706), .B(n5705), .ZN(U2801)
         );
  AOI22_X1 U6745 ( .A1(EBX_REG_25__SCAN_IN), .A2(n5980), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n5997), .ZN(n5715) );
  INV_X1 U6746 ( .A(n5773), .ZN(n5708) );
  AOI22_X1 U6747 ( .A1(n5708), .A2(n5996), .B1(REIP_REG_25__SCAN_IN), .B2(
        n5716), .ZN(n5714) );
  INV_X1 U6748 ( .A(n5709), .ZN(n5787) );
  AOI22_X1 U6749 ( .A1(n5770), .A2(n5951), .B1(n5965), .B2(n5787), .ZN(n5713)
         );
  INV_X1 U6750 ( .A(n5710), .ZN(n5726) );
  OAI211_X1 U6751 ( .C1(REIP_REG_24__SCAN_IN), .C2(REIP_REG_25__SCAN_IN), .A(
        n5726), .B(n5711), .ZN(n5712) );
  NAND4_X1 U6752 ( .A1(n5715), .A2(n5714), .A3(n5713), .A4(n5712), .ZN(U2802)
         );
  INV_X1 U6753 ( .A(REIP_REG_24__SCAN_IN), .ZN(n7016) );
  AOI22_X1 U6754 ( .A1(n5997), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        REIP_REG_24__SCAN_IN), .B2(n5716), .ZN(n5720) );
  INV_X1 U6755 ( .A(n5717), .ZN(n5718) );
  NAND2_X1 U6756 ( .A1(n5996), .A2(n5718), .ZN(n5719) );
  OAI211_X1 U6757 ( .C1(n6000), .C2(n5721), .A(n5720), .B(n5719), .ZN(n5722)
         );
  AOI21_X1 U6758 ( .B1(n5723), .B2(n5951), .A(n5722), .ZN(n5724) );
  INV_X1 U6759 ( .A(n5724), .ZN(n5725) );
  AOI21_X1 U6760 ( .B1(n5726), .B2(n7016), .A(n5725), .ZN(n5727) );
  OAI21_X1 U6761 ( .B1(n5728), .B2(n5992), .A(n5727), .ZN(U2803) );
  AOI22_X1 U6762 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n5997), .B1(n5729), 
        .B2(n5996), .ZN(n5730) );
  OAI21_X1 U6763 ( .B1(REIP_REG_22__SCAN_IN), .B2(n5731), .A(n5730), .ZN(n5735) );
  OAI22_X1 U6764 ( .A1(n5733), .A2(n5937), .B1(n5732), .B2(n5992), .ZN(n5734)
         );
  AOI211_X1 U6765 ( .C1(EBX_REG_22__SCAN_IN), .C2(n5980), .A(n5735), .B(n5734), 
        .ZN(n5736) );
  OAI221_X1 U6766 ( .B1(n6784), .B2(n5738), .C1(n6784), .C2(n5737), .A(n5736), 
        .ZN(U2805) );
  NAND3_X1 U6767 ( .A1(REIP_REG_18__SCAN_IN), .A2(n5747), .A3(n7043), .ZN(
        n5743) );
  INV_X1 U6768 ( .A(n5778), .ZN(n5741) );
  INV_X1 U6769 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5739) );
  OAI21_X1 U6770 ( .B1(n5872), .B2(n5739), .A(n5819), .ZN(n5740) );
  AOI21_X1 U6771 ( .B1(n5741), .B2(n5996), .A(n5740), .ZN(n5742) );
  OAI211_X1 U6772 ( .C1(n5744), .C2(n6000), .A(n5743), .B(n5742), .ZN(n5745)
         );
  AOI21_X1 U6773 ( .B1(n5775), .B2(n5951), .A(n5745), .ZN(n5749) );
  AND2_X1 U6774 ( .A1(n5989), .A2(n5746), .ZN(n5864) );
  AND2_X1 U6775 ( .A1(n6967), .A2(n5747), .ZN(n5852) );
  OAI21_X1 U6776 ( .B1(n5864), .B2(n5852), .A(REIP_REG_19__SCAN_IN), .ZN(n5748) );
  OAI211_X1 U6777 ( .C1(n5750), .C2(n5992), .A(n5749), .B(n5748), .ZN(U2808)
         );
  INV_X1 U6778 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5753) );
  AOI22_X1 U6779 ( .A1(n3183), .A2(n6019), .B1(n5751), .B2(n6018), .ZN(n5752)
         );
  OAI21_X1 U6780 ( .B1(n5753), .B2(n6022), .A(n5752), .ZN(U2832) );
  AOI22_X1 U6781 ( .A1(n3183), .A2(n6030), .B1(n6029), .B2(DATAI_27_), .ZN(
        n5755) );
  AOI22_X1 U6782 ( .A1(n6026), .A2(DATAI_11_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n6025), .ZN(n5754) );
  NAND2_X1 U6783 ( .A1(n5755), .A2(n5754), .ZN(U2864) );
  AOI22_X1 U6784 ( .A1(n5770), .A2(n6030), .B1(n6029), .B2(DATAI_25_), .ZN(
        n5757) );
  AOI22_X1 U6785 ( .A1(n6026), .A2(DATAI_9_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n6025), .ZN(n5756) );
  NAND2_X1 U6786 ( .A1(n5757), .A2(n5756), .ZN(U2866) );
  AOI22_X1 U6787 ( .A1(n5758), .A2(n6030), .B1(n6029), .B2(DATAI_23_), .ZN(
        n5760) );
  AOI22_X1 U6788 ( .A1(n6026), .A2(DATAI_7_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n6025), .ZN(n5759) );
  NAND2_X1 U6789 ( .A1(n5760), .A2(n5759), .ZN(U2868) );
  AOI22_X1 U6790 ( .A1(n5761), .A2(n6030), .B1(n6029), .B2(DATAI_21_), .ZN(
        n5763) );
  AOI22_X1 U6791 ( .A1(n6026), .A2(DATAI_5_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n6025), .ZN(n5762) );
  NAND2_X1 U6792 ( .A1(n5763), .A2(n5762), .ZN(U2870) );
  AOI22_X1 U6793 ( .A1(n5764), .A2(n6030), .B1(n6029), .B2(DATAI_20_), .ZN(
        n5766) );
  AOI22_X1 U6794 ( .A1(n6026), .A2(DATAI_4_), .B1(EAX_REG_20__SCAN_IN), .B2(
        n6025), .ZN(n5765) );
  NAND2_X1 U6795 ( .A1(n5766), .A2(n5765), .ZN(U2871) );
  AOI22_X1 U6796 ( .A1(n5775), .A2(n6030), .B1(n6029), .B2(DATAI_19_), .ZN(
        n5768) );
  AOI22_X1 U6797 ( .A1(n6026), .A2(DATAI_3_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n6025), .ZN(n5767) );
  NAND2_X1 U6798 ( .A1(n5768), .A2(n5767), .ZN(U2872) );
  AOI22_X1 U6799 ( .A1(n6176), .A2(REIP_REG_25__SCAN_IN), .B1(n6117), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5772) );
  OAI21_X1 U6800 ( .B1(n5403), .B2(n5769), .A(n5204), .ZN(n5788) );
  AOI22_X1 U6801 ( .A1(n5770), .A2(n6113), .B1(n6115), .B2(n5788), .ZN(n5771)
         );
  OAI211_X1 U6802 ( .C1(n6111), .C2(n5773), .A(n5772), .B(n5771), .ZN(U2961)
         );
  AOI22_X1 U6803 ( .A1(n6176), .A2(REIP_REG_19__SCAN_IN), .B1(n6117), .B2(
        PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5777) );
  AOI22_X1 U6804 ( .A1(n6113), .A2(n5775), .B1(n5774), .B2(n6115), .ZN(n5776)
         );
  OAI211_X1 U6805 ( .C1(n6111), .C2(n5778), .A(n5777), .B(n5776), .ZN(U2967)
         );
  INV_X1 U6806 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5861) );
  INV_X1 U6807 ( .A(n5867), .ZN(n5782) );
  NAND2_X1 U6808 ( .A1(n4716), .A2(n5779), .ZN(n5780) );
  AND2_X1 U6809 ( .A1(n4766), .A2(n5780), .ZN(n6024) );
  AOI222_X1 U6810 ( .A1(n5783), .A2(n6115), .B1(n5782), .B2(n5781), .C1(n6113), 
        .C2(n6024), .ZN(n5785) );
  OAI211_X1 U6811 ( .C1(n5861), .C2(n5786), .A(n5785), .B(n5784), .ZN(U2969)
         );
  AOI22_X1 U6812 ( .A1(n5788), .A2(n6175), .B1(n6172), .B2(n5787), .ZN(n5794)
         );
  INV_X1 U6813 ( .A(REIP_REG_25__SCAN_IN), .ZN(n7164) );
  NOR2_X1 U6814 ( .A1(n5819), .A2(n7164), .ZN(n5789) );
  AOI221_X1 U6815 ( .B1(n5792), .B2(n5791), .C1(n5790), .C2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5789), .ZN(n5793) );
  NAND2_X1 U6816 ( .A1(n5794), .A2(n5793), .ZN(U2993) );
  INV_X1 U6817 ( .A(n5797), .ZN(n5795) );
  AOI21_X1 U6818 ( .B1(n5795), .B2(n6170), .A(n6134), .ZN(n5812) );
  INV_X1 U6819 ( .A(n5796), .ZN(n5801) );
  INV_X1 U6820 ( .A(n6138), .ZN(n6123) );
  NAND2_X1 U6821 ( .A1(n5797), .A2(n6123), .ZN(n5804) );
  AOI221_X1 U6822 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .C1(n5497), .C2(n4786), .A(n5804), 
        .ZN(n5798) );
  AOI21_X1 U6823 ( .B1(n5969), .B2(REIP_REG_16__SCAN_IN), .A(n5798), .ZN(n5799) );
  OAI21_X1 U6824 ( .B1(n6163), .B2(n5879), .A(n5799), .ZN(n5800) );
  AOI21_X1 U6825 ( .B1(n5801), .B2(n6175), .A(n5800), .ZN(n5802) );
  OAI21_X1 U6826 ( .B1(n5812), .B2(n4786), .A(n5802), .ZN(U3002) );
  INV_X1 U6827 ( .A(n5803), .ZN(n5810) );
  NOR2_X1 U6828 ( .A1(n5804), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5809)
         );
  AOI21_X1 U6829 ( .B1(n5807), .B2(n5806), .A(n5805), .ZN(n5885) );
  INV_X1 U6830 ( .A(n5885), .ZN(n6005) );
  OAI22_X1 U6831 ( .A1(n6163), .A2(n6005), .B1(n6779), .B2(n5819), .ZN(n5808)
         );
  AOI211_X1 U6832 ( .C1(n5810), .C2(n6175), .A(n5809), .B(n5808), .ZN(n5811)
         );
  OAI21_X1 U6833 ( .B1(n5812), .B2(n5497), .A(n5811), .ZN(U3003) );
  NAND2_X1 U6834 ( .A1(n5813), .A2(n5814), .ZN(n5824) );
  NOR2_X1 U6835 ( .A1(n5815), .A2(n5814), .ZN(n5821) );
  AOI21_X1 U6836 ( .B1(n5818), .B2(n5817), .A(n5816), .ZN(n5889) );
  INV_X1 U6837 ( .A(n5889), .ZN(n6010) );
  OAI22_X1 U6838 ( .A1(n6163), .A2(n6010), .B1(n5113), .B2(n5819), .ZN(n5820)
         );
  AOI211_X1 U6839 ( .C1(n5822), .C2(n6175), .A(n5821), .B(n5820), .ZN(n5823)
         );
  OAI21_X1 U6840 ( .B1(n6138), .B2(n5824), .A(n5823), .ZN(U3005) );
  INV_X1 U6841 ( .A(n5966), .ZN(n5829) );
  INV_X1 U6842 ( .A(n5825), .ZN(n5828) );
  NAND4_X1 U6843 ( .A1(n5829), .A2(n5828), .A3(n5827), .A4(n5826), .ZN(n5830)
         );
  OAI21_X1 U6844 ( .B1(n5832), .B2(n5831), .A(n5830), .ZN(U3455) );
  INV_X1 U6845 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6758) );
  NAND2_X1 U6846 ( .A1(n6758), .A2(STATE_REG_1__SCAN_IN), .ZN(n7220) );
  INV_X1 U6847 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6966) );
  INV_X1 U6848 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6959) );
  OAI221_X1 U6849 ( .B1(n6959), .B2(n6758), .C1(STATE_REG_1__SCAN_IN), .C2(
        n6758), .A(n7220), .ZN(n6748) );
  INV_X1 U6850 ( .A(n6748), .ZN(n6794) );
  INV_X1 U6851 ( .A(n6794), .ZN(n6791) );
  OAI21_X1 U6852 ( .B1(n7221), .B2(n6966), .A(n6791), .ZN(U2789) );
  INV_X1 U6853 ( .A(D_C_N_REG_SCAN_IN), .ZN(n6955) );
  NOR2_X1 U6854 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5834) );
  NOR2_X1 U6855 ( .A1(n7221), .A2(n5834), .ZN(n5833) );
  AOI22_X1 U6856 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(n7221), .B1(n6955), .B2(
        n5833), .ZN(U2791) );
  OAI21_X1 U6857 ( .B1(BS16_N), .B2(n5834), .A(n6794), .ZN(n6793) );
  OAI21_X1 U6858 ( .B1(n6794), .B2(n6912), .A(n6793), .ZN(U2792) );
  OAI21_X1 U6859 ( .B1(n5836), .B2(n6712), .A(n5835), .ZN(U2793) );
  NOR4_X1 U6860 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(DATAWIDTH_REG_6__SCAN_IN), .A3(DATAWIDTH_REG_17__SCAN_IN), .A4(DATAWIDTH_REG_2__SCAN_IN), .ZN(n5840) );
  NOR4_X1 U6861 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_9__SCAN_IN), .A4(DATAWIDTH_REG_3__SCAN_IN), .ZN(n5839) );
  NOR4_X1 U6862 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5838) );
  NOR4_X1 U6863 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n5837) );
  NAND4_X1 U6864 ( .A1(n5840), .A2(n5839), .A3(n5838), .A4(n5837), .ZN(n5846)
         );
  NOR4_X1 U6865 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_12__SCAN_IN), .A4(DATAWIDTH_REG_19__SCAN_IN), .ZN(
        n5844) );
  AOI211_X1 U6866 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_11__SCAN_IN), .B(
        DATAWIDTH_REG_16__SCAN_IN), .ZN(n5843) );
  NOR4_X1 U6867 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(
        DATAWIDTH_REG_18__SCAN_IN), .A3(DATAWIDTH_REG_13__SCAN_IN), .A4(
        DATAWIDTH_REG_7__SCAN_IN), .ZN(n5842) );
  NOR4_X1 U6868 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_23__SCAN_IN), .A3(DATAWIDTH_REG_10__SCAN_IN), .A4(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n5841) );
  NAND4_X1 U6869 ( .A1(n5844), .A2(n5843), .A3(n5842), .A4(n5841), .ZN(n5845)
         );
  NOR2_X1 U6870 ( .A1(n5846), .A2(n5845), .ZN(n6824) );
  INV_X1 U6871 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n7193) );
  NOR3_X1 U6872 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_0__SCAN_IN), 
        .A3(DATAWIDTH_REG_1__SCAN_IN), .ZN(n5848) );
  OAI21_X1 U6873 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5848), .A(n6824), .ZN(n5847)
         );
  OAI21_X1 U6874 ( .B1(n6824), .B2(n7193), .A(n5847), .ZN(U2794) );
  INV_X1 U6875 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6979) );
  AOI21_X1 U6876 ( .B1(n3739), .B2(n6979), .A(n5848), .ZN(n5849) );
  INV_X1 U6877 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n7192) );
  INV_X1 U6878 ( .A(n6824), .ZN(n6822) );
  AOI22_X1 U6879 ( .A1(n6824), .A2(n5849), .B1(n7192), .B2(n6822), .ZN(U2795)
         );
  AOI21_X1 U6880 ( .B1(n5997), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n5969), 
        .ZN(n5850) );
  OAI21_X1 U6881 ( .B1(n6000), .B2(n5851), .A(n5850), .ZN(n5853) );
  AOI211_X1 U6882 ( .C1(REIP_REG_18__SCAN_IN), .C2(n5864), .A(n5853), .B(n5852), .ZN(n5854) );
  OAI21_X1 U6883 ( .B1(n5855), .B2(n5937), .A(n5854), .ZN(n5856) );
  AOI21_X1 U6884 ( .B1(n5857), .B2(n5996), .A(n5856), .ZN(n5858) );
  OAI21_X1 U6885 ( .B1(n5992), .B2(n5859), .A(n5858), .ZN(U2809) );
  NAND2_X1 U6886 ( .A1(n6983), .A2(n5860), .ZN(n5863) );
  INV_X1 U6887 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6004) );
  OAI22_X1 U6888 ( .A1(n6004), .A2(n6000), .B1(n5861), .B2(n5872), .ZN(n5862)
         );
  AOI211_X1 U6889 ( .C1(n5864), .C2(n5863), .A(n5969), .B(n5862), .ZN(n5866)
         );
  AOI22_X1 U6890 ( .A1(n6024), .A2(n5951), .B1(n5965), .B2(n6002), .ZN(n5865)
         );
  OAI211_X1 U6891 ( .C1(n5867), .C2(n5988), .A(n5866), .B(n5865), .ZN(U2810)
         );
  OR2_X1 U6892 ( .A1(n5934), .A2(n5868), .ZN(n5869) );
  NOR3_X1 U6893 ( .A1(n5869), .A2(REIP_REG_16__SCAN_IN), .A3(n6779), .ZN(n5874) );
  NOR2_X1 U6894 ( .A1(n5869), .A2(REIP_REG_15__SCAN_IN), .ZN(n5881) );
  OAI21_X1 U6895 ( .B1(n5880), .B2(n5881), .A(REIP_REG_16__SCAN_IN), .ZN(n5870) );
  OAI211_X1 U6896 ( .C1(n5872), .C2(n5871), .A(n5819), .B(n5870), .ZN(n5873)
         );
  AOI211_X1 U6897 ( .C1(n5980), .C2(EBX_REG_16__SCAN_IN), .A(n5874), .B(n5873), 
        .ZN(n5878) );
  INV_X1 U6898 ( .A(n5875), .ZN(n5876) );
  AOI22_X1 U6899 ( .A1(n6031), .A2(n5951), .B1(n5876), .B2(n5996), .ZN(n5877)
         );
  OAI211_X1 U6900 ( .C1(n5992), .C2(n5879), .A(n5878), .B(n5877), .ZN(U2811)
         );
  AOI22_X1 U6901 ( .A1(EBX_REG_15__SCAN_IN), .A2(n5980), .B1(
        REIP_REG_15__SCAN_IN), .B2(n5880), .ZN(n5883) );
  AOI211_X1 U6902 ( .C1(n5997), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5969), 
        .B(n5881), .ZN(n5882) );
  OAI211_X1 U6903 ( .C1(n6006), .C2(n5937), .A(n5883), .B(n5882), .ZN(n5884)
         );
  INV_X1 U6904 ( .A(n5884), .ZN(n5888) );
  AOI22_X1 U6905 ( .A1(n5886), .A2(n5996), .B1(n5965), .B2(n5885), .ZN(n5887)
         );
  NAND2_X1 U6906 ( .A1(n5888), .A2(n5887), .ZN(U2812) );
  AOI22_X1 U6907 ( .A1(EBX_REG_13__SCAN_IN), .A2(n5980), .B1(n5965), .B2(n5889), .ZN(n5897) );
  NOR3_X1 U6908 ( .A1(REIP_REG_13__SCAN_IN), .A2(n4681), .A3(n5893), .ZN(n5890) );
  AOI211_X1 U6909 ( .C1(n5997), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5969), 
        .B(n5890), .ZN(n5896) );
  OAI22_X1 U6910 ( .A1(n6013), .A2(n5937), .B1(n5891), .B2(n5988), .ZN(n5892)
         );
  INV_X1 U6911 ( .A(n5892), .ZN(n5895) );
  NOR2_X1 U6912 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5893), .ZN(n5900) );
  OAI21_X1 U6913 ( .B1(n5900), .B2(n5898), .A(REIP_REG_13__SCAN_IN), .ZN(n5894) );
  NAND4_X1 U6914 ( .A1(n5897), .A2(n5896), .A3(n5895), .A4(n5894), .ZN(U2814)
         );
  INV_X1 U6915 ( .A(n6124), .ZN(n5899) );
  AOI22_X1 U6916 ( .A1(n5965), .A2(n5899), .B1(REIP_REG_12__SCAN_IN), .B2(
        n5898), .ZN(n5907) );
  AOI211_X1 U6917 ( .C1(n5997), .C2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n5969), 
        .B(n5900), .ZN(n5906) );
  INV_X1 U6918 ( .A(n5901), .ZN(n5903) );
  AOI22_X1 U6919 ( .A1(n5903), .A2(n5951), .B1(n5996), .B2(n5902), .ZN(n5905)
         );
  NAND2_X1 U6920 ( .A1(EBX_REG_12__SCAN_IN), .A2(n5980), .ZN(n5904) );
  NAND4_X1 U6921 ( .A1(n5907), .A2(n5906), .A3(n5905), .A4(n5904), .ZN(U2815)
         );
  OAI22_X1 U6922 ( .A1(n4542), .A2(n6000), .B1(n5992), .B2(n5908), .ZN(n5909)
         );
  AOI211_X1 U6923 ( .C1(n5997), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n5969), 
        .B(n5909), .ZN(n5919) );
  INV_X1 U6924 ( .A(n5910), .ZN(n5912) );
  AOI22_X1 U6925 ( .A1(n5912), .A2(n5951), .B1(n5996), .B2(n5911), .ZN(n5918)
         );
  OAI21_X1 U6926 ( .B1(n5913), .B2(n5920), .A(REIP_REG_10__SCAN_IN), .ZN(n5917) );
  INV_X1 U6927 ( .A(n5914), .ZN(n5915) );
  NAND3_X1 U6928 ( .A1(n5915), .A2(n6775), .A3(REIP_REG_9__SCAN_IN), .ZN(n5916) );
  NAND4_X1 U6929 ( .A1(n5919), .A2(n5918), .A3(n5917), .A4(n5916), .ZN(U2817)
         );
  AOI22_X1 U6930 ( .A1(n5965), .A2(n5921), .B1(REIP_REG_8__SCAN_IN), .B2(n5920), .ZN(n5930) );
  INV_X1 U6931 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5924) );
  OAI22_X1 U6932 ( .A1(n5924), .A2(n6000), .B1(n5923), .B2(n5922), .ZN(n5925)
         );
  AOI211_X1 U6933 ( .C1(n5997), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n5969), 
        .B(n5925), .ZN(n5929) );
  AOI22_X1 U6934 ( .A1(n5927), .A2(n5951), .B1(n5996), .B2(n5926), .ZN(n5928)
         );
  NAND3_X1 U6935 ( .A1(n5930), .A2(n5929), .A3(n5928), .ZN(U2819) );
  OAI21_X1 U6936 ( .B1(n5934), .B2(n5932), .A(n5931), .ZN(n5958) );
  INV_X1 U6937 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6772) );
  NOR2_X1 U6938 ( .A1(n5934), .A2(n5933), .ZN(n5959) );
  NAND2_X1 U6939 ( .A1(REIP_REG_5__SCAN_IN), .A2(n5959), .ZN(n5948) );
  AOI221_X1 U6940 ( .B1(REIP_REG_7__SCAN_IN), .B2(REIP_REG_6__SCAN_IN), .C1(
        n6772), .C2(n6770), .A(n5948), .ZN(n5943) );
  NAND2_X1 U6941 ( .A1(n5997), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5935)
         );
  OAI211_X1 U6942 ( .C1(n6000), .C2(n5936), .A(n5819), .B(n5935), .ZN(n5940)
         );
  NOR2_X1 U6943 ( .A1(n5938), .A2(n5937), .ZN(n5939) );
  AOI211_X1 U6944 ( .C1(n6148), .C2(n5965), .A(n5940), .B(n5939), .ZN(n5941)
         );
  INV_X1 U6945 ( .A(n5941), .ZN(n5942) );
  AOI211_X1 U6946 ( .C1(REIP_REG_7__SCAN_IN), .C2(n5958), .A(n5943), .B(n5942), 
        .ZN(n5944) );
  OAI21_X1 U6947 ( .B1(n5945), .B2(n5988), .A(n5944), .ZN(U2820) );
  INV_X1 U6948 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6023) );
  AOI22_X1 U6949 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n5997), .B1(n5965), 
        .B2(n6017), .ZN(n5946) );
  OAI211_X1 U6950 ( .C1(n6000), .C2(n6023), .A(n5819), .B(n5946), .ZN(n5950)
         );
  INV_X1 U6951 ( .A(n5958), .ZN(n5947) );
  AOI22_X1 U6952 ( .A1(n5948), .A2(n6770), .B1(REIP_REG_6__SCAN_IN), .B2(n5947), .ZN(n5949) );
  AOI211_X1 U6953 ( .C1(n6020), .C2(n5951), .A(n5950), .B(n5949), .ZN(n5952)
         );
  OAI21_X1 U6954 ( .B1(n5953), .B2(n5988), .A(n5952), .ZN(U2821) );
  AOI22_X1 U6955 ( .A1(EBX_REG_5__SCAN_IN), .A2(n5980), .B1(
        PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n5997), .ZN(n5962) );
  OAI22_X1 U6956 ( .A1(n5955), .A2(n5994), .B1(n5954), .B2(n5988), .ZN(n5956)
         );
  AOI21_X1 U6957 ( .B1(n5965), .B2(n5957), .A(n5956), .ZN(n5961) );
  OAI21_X1 U6958 ( .B1(REIP_REG_5__SCAN_IN), .B2(n5959), .A(n5958), .ZN(n5960)
         );
  NAND4_X1 U6959 ( .A1(n5962), .A2(n5961), .A3(n5819), .A4(n5960), .ZN(U2822)
         );
  AOI22_X1 U6960 ( .A1(n5965), .A2(n5964), .B1(REIP_REG_4__SCAN_IN), .B2(n5963), .ZN(n5976) );
  INV_X1 U6961 ( .A(EBX_REG_4__SCAN_IN), .ZN(n5967) );
  OAI22_X1 U6962 ( .A1(n5967), .A2(n6000), .B1(n5966), .B2(n5981), .ZN(n5968)
         );
  AOI211_X1 U6963 ( .C1(n5997), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n5969), 
        .B(n5968), .ZN(n5975) );
  INV_X1 U6964 ( .A(n5994), .ZN(n5986) );
  AOI22_X1 U6965 ( .A1(n5971), .A2(n5986), .B1(n5970), .B2(n5996), .ZN(n5974)
         );
  INV_X1 U6966 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6767) );
  NAND3_X1 U6967 ( .A1(n5977), .A2(n5972), .A3(n6767), .ZN(n5973) );
  NAND4_X1 U6968 ( .A1(n5976), .A2(n5975), .A3(n5974), .A4(n5973), .ZN(U2823)
         );
  AOI21_X1 U6969 ( .B1(n5977), .B2(REIP_REG_1__SCAN_IN), .A(
        REIP_REG_2__SCAN_IN), .ZN(n5978) );
  NOR2_X1 U6970 ( .A1(n5979), .A2(n5978), .ZN(n5985) );
  AOI22_X1 U6971 ( .A1(n5980), .A2(EBX_REG_2__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n5997), .ZN(n5983) );
  INV_X1 U6972 ( .A(n5981), .ZN(n5990) );
  NAND2_X1 U6973 ( .A1(n5990), .A2(n6182), .ZN(n5982) );
  OAI211_X1 U6974 ( .C1(n6164), .C2(n5992), .A(n5983), .B(n5982), .ZN(n5984)
         );
  AOI211_X1 U6975 ( .C1(n6107), .C2(n5986), .A(n5985), .B(n5984), .ZN(n5987)
         );
  OAI21_X1 U6976 ( .B1(n6110), .B2(n5988), .A(n5987), .ZN(U2825) );
  AOI22_X1 U6977 ( .A1(n6814), .A2(n5990), .B1(n5989), .B2(REIP_REG_0__SCAN_IN), .ZN(n5999) );
  OAI22_X1 U6978 ( .A1(n5994), .A2(n5993), .B1(n5992), .B2(n5991), .ZN(n5995)
         );
  AOI221_X1 U6979 ( .B1(n5997), .B2(PHYADDRPOINTER_REG_0__SCAN_IN), .C1(n5996), 
        .C2(PHYADDRPOINTER_REG_0__SCAN_IN), .A(n5995), .ZN(n5998) );
  OAI211_X1 U6980 ( .C1(n6001), .C2(n6000), .A(n5999), .B(n5998), .ZN(U2827)
         );
  AOI22_X1 U6981 ( .A1(n6024), .A2(n6019), .B1(n6018), .B2(n6002), .ZN(n6003)
         );
  OAI21_X1 U6982 ( .B1(n6004), .B2(n6022), .A(n6003), .ZN(U2842) );
  INV_X1 U6983 ( .A(EBX_REG_15__SCAN_IN), .ZN(n6009) );
  OAI22_X1 U6984 ( .A1(n6006), .A2(n6012), .B1(n6011), .B2(n6005), .ZN(n6007)
         );
  INV_X1 U6985 ( .A(n6007), .ZN(n6008) );
  OAI21_X1 U6986 ( .B1(n6009), .B2(n6022), .A(n6008), .ZN(U2844) );
  INV_X1 U6987 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6016) );
  OAI22_X1 U6988 ( .A1(n6013), .A2(n6012), .B1(n6011), .B2(n6010), .ZN(n6014)
         );
  INV_X1 U6989 ( .A(n6014), .ZN(n6015) );
  OAI21_X1 U6990 ( .B1(n6016), .B2(n6022), .A(n6015), .ZN(U2846) );
  AOI22_X1 U6991 ( .A1(n6020), .A2(n6019), .B1(n6018), .B2(n6017), .ZN(n6021)
         );
  OAI21_X1 U6992 ( .B1(n6023), .B2(n6022), .A(n6021), .ZN(U2853) );
  AOI22_X1 U6993 ( .A1(n6024), .A2(n6030), .B1(n6029), .B2(DATAI_17_), .ZN(
        n6028) );
  AOI22_X1 U6994 ( .A1(n6026), .A2(DATAI_1_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n6025), .ZN(n6027) );
  NAND2_X1 U6995 ( .A1(n6028), .A2(n6027), .ZN(U2874) );
  AOI22_X1 U6996 ( .A1(n6031), .A2(n6030), .B1(n6029), .B2(DATAI_16_), .ZN(
        n6036) );
  OAI22_X1 U6997 ( .A1(n6033), .A2(n6081), .B1(n4073), .B2(n6032), .ZN(n6034)
         );
  INV_X1 U6998 ( .A(n6034), .ZN(n6035) );
  NAND2_X1 U6999 ( .A1(n6036), .A2(n6035), .ZN(U2875) );
  AOI22_X1 U7000 ( .A1(n6059), .A2(LWORD_REG_15__SCAN_IN), .B1(n6058), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6038) );
  OAI21_X1 U7001 ( .B1(n6039), .B2(n6061), .A(n6038), .ZN(U2908) );
  AOI22_X1 U7002 ( .A1(n6059), .A2(LWORD_REG_14__SCAN_IN), .B1(n6058), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6040) );
  OAI21_X1 U7003 ( .B1(n4583), .B2(n6061), .A(n6040), .ZN(U2909) );
  AOI22_X1 U7004 ( .A1(n6059), .A2(LWORD_REG_13__SCAN_IN), .B1(n6058), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6041) );
  OAI21_X1 U7005 ( .B1(n4517), .B2(n6061), .A(n6041), .ZN(U2910) );
  AOI22_X1 U7006 ( .A1(n6059), .A2(LWORD_REG_12__SCAN_IN), .B1(n6058), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6042) );
  OAI21_X1 U7007 ( .B1(n4486), .B2(n6061), .A(n6042), .ZN(U2911) );
  AOI22_X1 U7008 ( .A1(n6059), .A2(LWORD_REG_11__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6043) );
  OAI21_X1 U7009 ( .B1(n6044), .B2(n6061), .A(n6043), .ZN(U2912) );
  AOI22_X1 U7010 ( .A1(n6059), .A2(LWORD_REG_10__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6045) );
  OAI21_X1 U7011 ( .B1(n4453), .B2(n6061), .A(n6045), .ZN(U2913) );
  AOI22_X1 U7012 ( .A1(n6059), .A2(LWORD_REG_9__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6046) );
  OAI21_X1 U7013 ( .B1(n4397), .B2(n6061), .A(n6046), .ZN(U2914) );
  AOI22_X1 U7014 ( .A1(n6059), .A2(LWORD_REG_8__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6048) );
  OAI21_X1 U7015 ( .B1(n4346), .B2(n6061), .A(n6048), .ZN(U2915) );
  AOI22_X1 U7016 ( .A1(n6059), .A2(LWORD_REG_7__SCAN_IN), .B1(n6058), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6049) );
  OAI21_X1 U7017 ( .B1(n4267), .B2(n6061), .A(n6049), .ZN(U2916) );
  AOI22_X1 U7018 ( .A1(n6059), .A2(LWORD_REG_6__SCAN_IN), .B1(n6058), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6050) );
  OAI21_X1 U7019 ( .B1(n4181), .B2(n6061), .A(n6050), .ZN(U2917) );
  AOI22_X1 U7020 ( .A1(n6059), .A2(LWORD_REG_5__SCAN_IN), .B1(n6058), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6051) );
  OAI21_X1 U7021 ( .B1(n4024), .B2(n6061), .A(n6051), .ZN(U2918) );
  AOI22_X1 U7022 ( .A1(n6059), .A2(LWORD_REG_4__SCAN_IN), .B1(n6058), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6052) );
  OAI21_X1 U7023 ( .B1(n6053), .B2(n6061), .A(n6052), .ZN(U2919) );
  AOI22_X1 U7024 ( .A1(n6059), .A2(LWORD_REG_3__SCAN_IN), .B1(n6058), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6054) );
  OAI21_X1 U7025 ( .B1(n3837), .B2(n6061), .A(n6054), .ZN(U2920) );
  AOI22_X1 U7026 ( .A1(n6059), .A2(LWORD_REG_2__SCAN_IN), .B1(n6058), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6055) );
  OAI21_X1 U7027 ( .B1(n6056), .B2(n6061), .A(n6055), .ZN(U2921) );
  AOI22_X1 U7028 ( .A1(n6059), .A2(LWORD_REG_1__SCAN_IN), .B1(n6058), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6057) );
  OAI21_X1 U7029 ( .B1(n3621), .B2(n6061), .A(n6057), .ZN(U2922) );
  AOI22_X1 U7030 ( .A1(n6059), .A2(LWORD_REG_0__SCAN_IN), .B1(n6058), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6060) );
  OAI21_X1 U7031 ( .B1(n3524), .B2(n6061), .A(n6060), .ZN(U2923) );
  INV_X1 U7032 ( .A(n6062), .ZN(n6063) );
  OAI21_X1 U7033 ( .B1(n5239), .B2(n7199), .A(n6063), .ZN(n6093) );
  INV_X2 U7034 ( .A(n6064), .ZN(n6100) );
  AOI22_X1 U7035 ( .A1(UWORD_REG_0__SCAN_IN), .A2(n6097), .B1(n6100), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6065) );
  OAI21_X1 U7036 ( .B1(n6102), .B2(n6081), .A(n6065), .ZN(U2924) );
  AOI22_X1 U7037 ( .A1(UWORD_REG_1__SCAN_IN), .A2(n6097), .B1(n6100), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6066) );
  OAI21_X1 U7038 ( .B1(n6102), .B2(n7170), .A(n6066), .ZN(U2925) );
  AOI22_X1 U7039 ( .A1(UWORD_REG_2__SCAN_IN), .A2(n6097), .B1(n6100), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6067) );
  OAI21_X1 U7040 ( .B1(n6102), .B2(n7145), .A(n6067), .ZN(U2926) );
  AOI22_X1 U7041 ( .A1(UWORD_REG_3__SCAN_IN), .A2(n6097), .B1(n6100), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n6068) );
  OAI21_X1 U7042 ( .B1(n6102), .B2(n6934), .A(n6068), .ZN(U2927) );
  AOI22_X1 U7043 ( .A1(UWORD_REG_4__SCAN_IN), .A2(n6097), .B1(n6100), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n6069) );
  OAI21_X1 U7044 ( .B1(n6102), .B2(n6972), .A(n6069), .ZN(U2928) );
  AOI22_X1 U7045 ( .A1(UWORD_REG_5__SCAN_IN), .A2(n6097), .B1(n6100), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n6070) );
  OAI21_X1 U7046 ( .B1(n6102), .B2(n7161), .A(n6070), .ZN(U2929) );
  AOI22_X1 U7047 ( .A1(UWORD_REG_6__SCAN_IN), .A2(n6097), .B1(n6100), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n6071) );
  OAI21_X1 U7048 ( .B1(n6102), .B2(n6995), .A(n6071), .ZN(U2930) );
  AOI22_X1 U7049 ( .A1(UWORD_REG_7__SCAN_IN), .A2(n6097), .B1(n6100), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n6072) );
  OAI21_X1 U7050 ( .B1(n6102), .B2(n6991), .A(n6072), .ZN(U2931) );
  AOI22_X1 U7051 ( .A1(UWORD_REG_8__SCAN_IN), .A2(n6097), .B1(n6100), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n6073) );
  OAI21_X1 U7052 ( .B1(n6102), .B2(n7196), .A(n6073), .ZN(U2932) );
  AOI22_X1 U7053 ( .A1(UWORD_REG_9__SCAN_IN), .A2(n6097), .B1(n6100), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n6074) );
  OAI21_X1 U7054 ( .B1(n6102), .B2(n6091), .A(n6074), .ZN(U2933) );
  AOI22_X1 U7055 ( .A1(UWORD_REG_10__SCAN_IN), .A2(n6097), .B1(n6100), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n6075) );
  OAI21_X1 U7056 ( .B1(n6102), .B2(n6921), .A(n6075), .ZN(U2934) );
  AOI22_X1 U7057 ( .A1(UWORD_REG_11__SCAN_IN), .A2(n6097), .B1(n6100), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n6076) );
  OAI21_X1 U7058 ( .B1(n6102), .B2(n7040), .A(n6076), .ZN(U2935) );
  AOI22_X1 U7059 ( .A1(UWORD_REG_12__SCAN_IN), .A2(n6093), .B1(n6100), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n6077) );
  OAI21_X1 U7060 ( .B1(n6102), .B2(n7186), .A(n6077), .ZN(U2936) );
  AOI22_X1 U7061 ( .A1(UWORD_REG_13__SCAN_IN), .A2(n6093), .B1(n6100), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n6078) );
  OAI21_X1 U7062 ( .B1(n6102), .B2(n6993), .A(n6078), .ZN(U2937) );
  AOI22_X1 U7063 ( .A1(UWORD_REG_14__SCAN_IN), .A2(n6093), .B1(n6100), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n6079) );
  OAI21_X1 U7064 ( .B1(n6102), .B2(n6099), .A(n6079), .ZN(U2938) );
  AOI22_X1 U7065 ( .A1(LWORD_REG_0__SCAN_IN), .A2(n6093), .B1(n6100), .B2(
        EAX_REG_0__SCAN_IN), .ZN(n6080) );
  OAI21_X1 U7066 ( .B1(n6102), .B2(n6081), .A(n6080), .ZN(U2939) );
  AOI22_X1 U7067 ( .A1(LWORD_REG_1__SCAN_IN), .A2(n6093), .B1(n6100), .B2(
        EAX_REG_1__SCAN_IN), .ZN(n6082) );
  OAI21_X1 U7068 ( .B1(n6102), .B2(n7170), .A(n6082), .ZN(U2940) );
  AOI22_X1 U7069 ( .A1(LWORD_REG_2__SCAN_IN), .A2(n6093), .B1(n6100), .B2(
        EAX_REG_2__SCAN_IN), .ZN(n6083) );
  OAI21_X1 U7070 ( .B1(n6102), .B2(n7145), .A(n6083), .ZN(U2941) );
  AOI22_X1 U7071 ( .A1(LWORD_REG_3__SCAN_IN), .A2(n6093), .B1(n6100), .B2(
        EAX_REG_3__SCAN_IN), .ZN(n6084) );
  OAI21_X1 U7072 ( .B1(n6102), .B2(n6934), .A(n6084), .ZN(U2942) );
  AOI22_X1 U7073 ( .A1(LWORD_REG_4__SCAN_IN), .A2(n6097), .B1(n6100), .B2(
        EAX_REG_4__SCAN_IN), .ZN(n6085) );
  OAI21_X1 U7074 ( .B1(n6102), .B2(n6972), .A(n6085), .ZN(U2943) );
  AOI22_X1 U7075 ( .A1(LWORD_REG_5__SCAN_IN), .A2(n6097), .B1(n6100), .B2(
        EAX_REG_5__SCAN_IN), .ZN(n6086) );
  OAI21_X1 U7076 ( .B1(n6102), .B2(n7161), .A(n6086), .ZN(U2944) );
  AOI22_X1 U7077 ( .A1(LWORD_REG_6__SCAN_IN), .A2(n6097), .B1(n6100), .B2(
        EAX_REG_6__SCAN_IN), .ZN(n6087) );
  OAI21_X1 U7078 ( .B1(n6102), .B2(n6995), .A(n6087), .ZN(U2945) );
  AOI22_X1 U7079 ( .A1(LWORD_REG_7__SCAN_IN), .A2(n6097), .B1(n6100), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n6088) );
  OAI21_X1 U7080 ( .B1(n6102), .B2(n6991), .A(n6088), .ZN(U2946) );
  AOI22_X1 U7081 ( .A1(LWORD_REG_8__SCAN_IN), .A2(n6097), .B1(n6100), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n6089) );
  OAI21_X1 U7082 ( .B1(n6102), .B2(n7196), .A(n6089), .ZN(U2947) );
  AOI22_X1 U7083 ( .A1(LWORD_REG_9__SCAN_IN), .A2(n6093), .B1(n6100), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n6090) );
  OAI21_X1 U7084 ( .B1(n6102), .B2(n6091), .A(n6090), .ZN(U2948) );
  AOI22_X1 U7085 ( .A1(LWORD_REG_10__SCAN_IN), .A2(n6093), .B1(n6100), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n6092) );
  OAI21_X1 U7086 ( .B1(n6102), .B2(n6921), .A(n6092), .ZN(U2949) );
  AOI22_X1 U7087 ( .A1(LWORD_REG_11__SCAN_IN), .A2(n6093), .B1(n6100), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n6094) );
  OAI21_X1 U7088 ( .B1(n6102), .B2(n7040), .A(n6094), .ZN(U2950) );
  AOI22_X1 U7089 ( .A1(LWORD_REG_12__SCAN_IN), .A2(n6097), .B1(n6100), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n6095) );
  OAI21_X1 U7090 ( .B1(n6102), .B2(n7186), .A(n6095), .ZN(U2951) );
  AOI22_X1 U7091 ( .A1(LWORD_REG_13__SCAN_IN), .A2(n6097), .B1(n6100), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n6096) );
  OAI21_X1 U7092 ( .B1(n6102), .B2(n6993), .A(n6096), .ZN(U2952) );
  AOI22_X1 U7093 ( .A1(LWORD_REG_14__SCAN_IN), .A2(n6097), .B1(n6100), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n6098) );
  OAI21_X1 U7094 ( .B1(n6102), .B2(n6099), .A(n6098), .ZN(U2953) );
  AOI22_X1 U7095 ( .A1(LWORD_REG_15__SCAN_IN), .A2(n6097), .B1(n6100), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n6101) );
  OAI21_X1 U7096 ( .B1(n6102), .B2(n7028), .A(n6101), .ZN(U2954) );
  AOI22_X1 U7097 ( .A1(n6176), .A2(REIP_REG_2__SCAN_IN), .B1(n6117), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6109) );
  NAND2_X1 U7098 ( .A1(n6104), .A2(n6103), .ZN(n6105) );
  XOR2_X1 U7099 ( .A(n6106), .B(n6105), .Z(n6166) );
  AOI22_X1 U7100 ( .A1(n6166), .A2(n6115), .B1(n6107), .B2(n6113), .ZN(n6108)
         );
  OAI211_X1 U7101 ( .C1(n6111), .C2(n6110), .A(n6109), .B(n6108), .ZN(U2984)
         );
  AOI22_X1 U7102 ( .A1(n6115), .A2(n6114), .B1(n6113), .B2(n6112), .ZN(n6120)
         );
  OAI21_X1 U7103 ( .B1(n6117), .B2(n6116), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n6118) );
  NAND3_X1 U7104 ( .A1(n6120), .A2(n6119), .A3(n6118), .ZN(U2986) );
  AOI221_X1 U7105 ( .B1(n6161), .B2(n6122), .C1(n6121), .C2(n6122), .A(n6134), 
        .ZN(n6130) );
  AOI21_X1 U7106 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6123), .A(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6129) );
  OAI22_X1 U7107 ( .A1(n6126), .A2(n6125), .B1(n6163), .B2(n6124), .ZN(n6127)
         );
  AOI21_X1 U7108 ( .B1(n6176), .B2(REIP_REG_12__SCAN_IN), .A(n6127), .ZN(n6128) );
  OAI21_X1 U7109 ( .B1(n6130), .B2(n6129), .A(n6128), .ZN(U3006) );
  INV_X1 U7110 ( .A(n6131), .ZN(n6132) );
  AOI21_X1 U7111 ( .B1(n6172), .B2(n6133), .A(n6132), .ZN(n6137) );
  AOI22_X1 U7112 ( .A1(n6135), .A2(n6175), .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6134), .ZN(n6136) );
  OAI211_X1 U7113 ( .C1(INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n6138), .A(n6137), .B(n6136), .ZN(U3007) );
  INV_X1 U7114 ( .A(n6139), .ZN(n6147) );
  AOI21_X1 U7115 ( .B1(n6172), .B2(n6141), .A(n6140), .ZN(n6145) );
  AOI22_X1 U7116 ( .A1(n6143), .A2(n6175), .B1(n6142), .B2(n6146), .ZN(n6144)
         );
  OAI211_X1 U7117 ( .C1(n6147), .C2(n6146), .A(n6145), .B(n6144), .ZN(U3009)
         );
  NAND2_X1 U7118 ( .A1(n6172), .A2(n6148), .ZN(n6150) );
  OAI211_X1 U7119 ( .C1(n6151), .C2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n6150), 
        .B(n6149), .ZN(n6152) );
  AOI21_X1 U7120 ( .B1(n6153), .B2(n6175), .A(n6152), .ZN(n6154) );
  OAI21_X1 U7121 ( .B1(n6156), .B2(n6155), .A(n6154), .ZN(U3011) );
  NAND2_X1 U7122 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6157), .ZN(n6169)
         );
  OAI21_X1 U7123 ( .B1(n6159), .B2(n3881), .A(n6158), .ZN(n6160) );
  AOI22_X1 U7124 ( .A1(n6161), .A2(n6160), .B1(n5969), .B2(REIP_REG_2__SCAN_IN), .ZN(n6162) );
  OAI21_X1 U7125 ( .B1(n6164), .B2(n6163), .A(n6162), .ZN(n6165) );
  AOI21_X1 U7126 ( .B1(n6166), .B2(n6175), .A(n6165), .ZN(n6167) );
  OAI221_X1 U7127 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6169), .C1(n3881), .C2(n6168), .A(n6167), .ZN(U3016) );
  NAND2_X1 U7128 ( .A1(n6171), .A2(n6170), .ZN(n6179) );
  AOI222_X1 U7129 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6176), .B1(n6175), .B2(
        n6174), .C1(n6173), .C2(n6172), .ZN(n6177) );
  OAI221_X1 U7130 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n6179), .C1(n3876), .C2(n6178), .A(n6177), .ZN(U3017) );
  AND2_X1 U7131 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n6818), .ZN(U3019)
         );
  NAND3_X1 U7132 ( .A1(n6806), .A2(n6180), .A3(n6394), .ZN(n6216) );
  NOR2_X1 U7133 ( .A1(n6182), .A2(n6181), .ZN(n6432) );
  NAND2_X1 U7134 ( .A1(n6432), .A2(n6804), .ZN(n6213) );
  INV_X1 U7135 ( .A(n6324), .ZN(n6538) );
  INV_X1 U7136 ( .A(n6183), .ZN(n6184) );
  OAI22_X1 U7137 ( .A1(n6213), .A2(n6802), .B1(n6538), .B2(n6184), .ZN(n6208)
         );
  INV_X1 U7138 ( .A(n6471), .ZN(n6638) );
  NAND3_X1 U7139 ( .A1(n6810), .A2(n6704), .A3(n6400), .ZN(n6220) );
  NOR2_X1 U7140 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6220), .ZN(n6207)
         );
  AOI22_X1 U7141 ( .A1(n6639), .A2(n6208), .B1(n6638), .B2(n6207), .ZN(n6194)
         );
  INV_X1 U7142 ( .A(n6207), .ZN(n6186) );
  AOI211_X1 U7143 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6186), .A(n6317), .B(
        n6185), .ZN(n6192) );
  INV_X1 U7144 ( .A(n6243), .ZN(n6189) );
  AND2_X1 U7145 ( .A1(n6187), .A2(n3935), .ZN(n6188) );
  OAI21_X1 U7146 ( .B1(n6189), .B2(n6690), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6190) );
  NAND3_X1 U7147 ( .A1(n6190), .A2(n6812), .A3(n6213), .ZN(n6191) );
  NAND2_X1 U7148 ( .A1(n6192), .A2(n6191), .ZN(n6209) );
  AOI22_X1 U7149 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n6209), .B1(n6598), 
        .B2(n6690), .ZN(n6193) );
  OAI211_X1 U7150 ( .C1(n6601), .C2(n6243), .A(n6194), .B(n6193), .ZN(U3020)
         );
  INV_X1 U7151 ( .A(n6485), .ZN(n6650) );
  AOI22_X1 U7152 ( .A1(n6651), .A2(n6208), .B1(n6650), .B2(n6207), .ZN(n6196)
         );
  AOI22_X1 U7153 ( .A1(INSTQUEUE_REG_0__1__SCAN_IN), .A2(n6209), .B1(n6602), 
        .B2(n6690), .ZN(n6195) );
  OAI211_X1 U7154 ( .C1(n6605), .C2(n6243), .A(n6196), .B(n6195), .ZN(U3021)
         );
  INV_X1 U7155 ( .A(n6489), .ZN(n6656) );
  AOI22_X1 U7156 ( .A1(n6657), .A2(n6208), .B1(n6656), .B2(n6207), .ZN(n6198)
         );
  AOI22_X1 U7157 ( .A1(INSTQUEUE_REG_0__2__SCAN_IN), .A2(n6209), .B1(n6606), 
        .B2(n6690), .ZN(n6197) );
  OAI211_X1 U7158 ( .C1(n6609), .C2(n6243), .A(n6198), .B(n6197), .ZN(U3022)
         );
  INV_X1 U7159 ( .A(n6493), .ZN(n6662) );
  AOI22_X1 U7160 ( .A1(n6663), .A2(n6208), .B1(n6662), .B2(n6207), .ZN(n6200)
         );
  AOI22_X1 U7161 ( .A1(INSTQUEUE_REG_0__3__SCAN_IN), .A2(n6209), .B1(n6610), 
        .B2(n6690), .ZN(n6199) );
  OAI211_X1 U7162 ( .C1(n6613), .C2(n6243), .A(n6200), .B(n6199), .ZN(U3023)
         );
  INV_X1 U7163 ( .A(n6497), .ZN(n6668) );
  AOI22_X1 U7164 ( .A1(n6669), .A2(n6208), .B1(n6668), .B2(n6207), .ZN(n6202)
         );
  AOI22_X1 U7165 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n6209), .B1(n6614), 
        .B2(n6690), .ZN(n6201) );
  OAI211_X1 U7166 ( .C1(n6617), .C2(n6243), .A(n6202), .B(n6201), .ZN(U3024)
         );
  AOI22_X1 U7167 ( .A1(n6675), .A2(n6208), .B1(n6674), .B2(n6207), .ZN(n6204)
         );
  AOI22_X1 U7168 ( .A1(INSTQUEUE_REG_0__5__SCAN_IN), .A2(n6209), .B1(n6618), 
        .B2(n6690), .ZN(n6203) );
  OAI211_X1 U7169 ( .C1(n6621), .C2(n6243), .A(n6204), .B(n6203), .ZN(U3025)
         );
  AOI22_X1 U7170 ( .A1(n6681), .A2(n6208), .B1(n6680), .B2(n6207), .ZN(n6206)
         );
  AOI22_X1 U7171 ( .A1(INSTQUEUE_REG_0__6__SCAN_IN), .A2(n6209), .B1(n6622), 
        .B2(n6690), .ZN(n6205) );
  OAI211_X1 U7172 ( .C1(n6625), .C2(n6243), .A(n6206), .B(n6205), .ZN(U3026)
         );
  AOI22_X1 U7173 ( .A1(n6689), .A2(n6208), .B1(n6686), .B2(n6207), .ZN(n6211)
         );
  AOI22_X1 U7174 ( .A1(INSTQUEUE_REG_0__7__SCAN_IN), .A2(n6209), .B1(n6629), 
        .B2(n6690), .ZN(n6210) );
  OAI211_X1 U7175 ( .C1(n6633), .C2(n6243), .A(n6211), .B(n6210), .ZN(U3027)
         );
  NOR2_X1 U7176 ( .A1(n6819), .A2(n6220), .ZN(n6214) );
  INV_X1 U7177 ( .A(n6214), .ZN(n6244) );
  OAI22_X1 U7178 ( .A1(n6471), .A2(n6244), .B1(n6243), .B2(n6649), .ZN(n6212)
         );
  INV_X1 U7179 ( .A(n6212), .ZN(n6224) );
  INV_X1 U7180 ( .A(n6284), .ZN(n6645) );
  INV_X1 U7181 ( .A(n6213), .ZN(n6215) );
  AOI21_X1 U7182 ( .B1(n6215), .B2(n6814), .A(n6214), .ZN(n6222) );
  OR2_X1 U7183 ( .A1(n6216), .A2(n6912), .ZN(n6217) );
  AOI22_X1 U7184 ( .A1(n6222), .A2(n6219), .B1(n6802), .B2(n6220), .ZN(n6218)
         );
  NAND2_X1 U7185 ( .A1(n6645), .A2(n6218), .ZN(n6247) );
  INV_X1 U7186 ( .A(n6219), .ZN(n6221) );
  OAI22_X1 U7187 ( .A1(n6222), .A2(n6221), .B1(n6478), .B2(n6220), .ZN(n6246)
         );
  AOI22_X1 U7188 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n6247), .B1(n6639), 
        .B2(n6246), .ZN(n6223) );
  OAI211_X1 U7189 ( .C1(n6278), .C2(n6601), .A(n6224), .B(n6223), .ZN(U3028)
         );
  OAI22_X1 U7190 ( .A1(n6485), .A2(n6244), .B1(n6278), .B2(n6605), .ZN(n6225)
         );
  INV_X1 U7191 ( .A(n6225), .ZN(n6227) );
  AOI22_X1 U7192 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n6247), .B1(n6651), 
        .B2(n6246), .ZN(n6226) );
  OAI211_X1 U7193 ( .C1(n6655), .C2(n6243), .A(n6227), .B(n6226), .ZN(U3029)
         );
  OAI22_X1 U7194 ( .A1(n6489), .A2(n6244), .B1(n6278), .B2(n6609), .ZN(n6228)
         );
  INV_X1 U7195 ( .A(n6228), .ZN(n6230) );
  AOI22_X1 U7196 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n6247), .B1(n6657), 
        .B2(n6246), .ZN(n6229) );
  OAI211_X1 U7197 ( .C1(n6661), .C2(n6243), .A(n6230), .B(n6229), .ZN(U3030)
         );
  OAI22_X1 U7198 ( .A1(n6493), .A2(n6244), .B1(n6243), .B2(n6667), .ZN(n6231)
         );
  INV_X1 U7199 ( .A(n6231), .ZN(n6233) );
  AOI22_X1 U7200 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n6247), .B1(n6663), 
        .B2(n6246), .ZN(n6232) );
  OAI211_X1 U7201 ( .C1(n6278), .C2(n6613), .A(n6233), .B(n6232), .ZN(U3031)
         );
  OAI22_X1 U7202 ( .A1(n6497), .A2(n6244), .B1(n6278), .B2(n6617), .ZN(n6234)
         );
  INV_X1 U7203 ( .A(n6234), .ZN(n6236) );
  AOI22_X1 U7204 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n6247), .B1(n6669), 
        .B2(n6246), .ZN(n6235) );
  OAI211_X1 U7205 ( .C1(n6673), .C2(n6243), .A(n6236), .B(n6235), .ZN(U3032)
         );
  OAI22_X1 U7206 ( .A1(n6501), .A2(n6244), .B1(n6278), .B2(n6621), .ZN(n6237)
         );
  INV_X1 U7207 ( .A(n6237), .ZN(n6239) );
  AOI22_X1 U7208 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n6247), .B1(n6675), 
        .B2(n6246), .ZN(n6238) );
  OAI211_X1 U7209 ( .C1(n6679), .C2(n6243), .A(n6239), .B(n6238), .ZN(U3033)
         );
  OAI22_X1 U7210 ( .A1(n6505), .A2(n6244), .B1(n6278), .B2(n6625), .ZN(n6240)
         );
  INV_X1 U7211 ( .A(n6240), .ZN(n6242) );
  AOI22_X1 U7212 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n6247), .B1(n6681), 
        .B2(n6246), .ZN(n6241) );
  OAI211_X1 U7213 ( .C1(n6685), .C2(n6243), .A(n6242), .B(n6241), .ZN(U3034)
         );
  OAI22_X1 U7214 ( .A1(n6510), .A2(n6244), .B1(n6243), .B2(n6696), .ZN(n6245)
         );
  INV_X1 U7215 ( .A(n6245), .ZN(n6249) );
  AOI22_X1 U7216 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n6247), .B1(n6689), 
        .B2(n6246), .ZN(n6248) );
  OAI211_X1 U7217 ( .C1(n6278), .C2(n6633), .A(n6249), .B(n6248), .ZN(U3035)
         );
  NAND2_X1 U7218 ( .A1(n6480), .A2(n6810), .ZN(n6318) );
  OAI22_X1 U7219 ( .A1(n6254), .A2(n6802), .B1(n6538), .B2(n6318), .ZN(n6273)
         );
  NOR2_X1 U7220 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6250), .ZN(n6272)
         );
  AOI22_X1 U7221 ( .A1(n6639), .A2(n6273), .B1(n6638), .B2(n6272), .ZN(n6259)
         );
  INV_X1 U7222 ( .A(n6278), .ZN(n6253) );
  INV_X1 U7223 ( .A(n6252), .ZN(n6805) );
  OAI21_X1 U7224 ( .B1(n6253), .B2(n6274), .A(n6805), .ZN(n6255) );
  AOI21_X1 U7225 ( .B1(n6255), .B2(n6254), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n6257) );
  OAI21_X1 U7226 ( .B1(n6480), .B2(n6637), .A(n6256), .ZN(n6323) );
  NOR2_X1 U7227 ( .A1(n6317), .A2(n6323), .ZN(n6477) );
  OAI21_X1 U7228 ( .B1(n6257), .B2(n6272), .A(n6477), .ZN(n6275) );
  AOI22_X1 U7229 ( .A1(n6275), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n6646), 
        .B2(n6274), .ZN(n6258) );
  OAI211_X1 U7230 ( .C1(n6649), .C2(n6278), .A(n6259), .B(n6258), .ZN(U3036)
         );
  AOI22_X1 U7231 ( .A1(n6651), .A2(n6273), .B1(n6650), .B2(n6272), .ZN(n6261)
         );
  AOI22_X1 U7232 ( .A1(n6275), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n6274), 
        .B2(n6652), .ZN(n6260) );
  OAI211_X1 U7233 ( .C1(n6278), .C2(n6655), .A(n6261), .B(n6260), .ZN(U3037)
         );
  AOI22_X1 U7234 ( .A1(n6657), .A2(n6273), .B1(n6656), .B2(n6272), .ZN(n6263)
         );
  AOI22_X1 U7235 ( .A1(n6275), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n6274), 
        .B2(n6658), .ZN(n6262) );
  OAI211_X1 U7236 ( .C1(n6278), .C2(n6661), .A(n6263), .B(n6262), .ZN(U3038)
         );
  AOI22_X1 U7237 ( .A1(n6663), .A2(n6273), .B1(n6662), .B2(n6272), .ZN(n6265)
         );
  AOI22_X1 U7238 ( .A1(n6275), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n6274), 
        .B2(n6664), .ZN(n6264) );
  OAI211_X1 U7239 ( .C1(n6278), .C2(n6667), .A(n6265), .B(n6264), .ZN(U3039)
         );
  AOI22_X1 U7240 ( .A1(n6669), .A2(n6273), .B1(n6668), .B2(n6272), .ZN(n6267)
         );
  AOI22_X1 U7241 ( .A1(n6275), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n6274), 
        .B2(n6670), .ZN(n6266) );
  OAI211_X1 U7242 ( .C1(n6278), .C2(n6673), .A(n6267), .B(n6266), .ZN(U3040)
         );
  AOI22_X1 U7243 ( .A1(n6675), .A2(n6273), .B1(n6674), .B2(n6272), .ZN(n6269)
         );
  AOI22_X1 U7244 ( .A1(n6275), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n6274), 
        .B2(n6676), .ZN(n6268) );
  OAI211_X1 U7245 ( .C1(n6278), .C2(n6679), .A(n6269), .B(n6268), .ZN(U3041)
         );
  AOI22_X1 U7246 ( .A1(n6681), .A2(n6273), .B1(n6680), .B2(n6272), .ZN(n6271)
         );
  AOI22_X1 U7247 ( .A1(n6275), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n6274), 
        .B2(n6682), .ZN(n6270) );
  OAI211_X1 U7248 ( .C1(n6278), .C2(n6685), .A(n6271), .B(n6270), .ZN(U3042)
         );
  AOI22_X1 U7249 ( .A1(n6689), .A2(n6273), .B1(n6686), .B2(n6272), .ZN(n6277)
         );
  AOI22_X1 U7250 ( .A1(n6275), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n6274), 
        .B2(n6691), .ZN(n6276) );
  OAI211_X1 U7251 ( .C1(n6278), .C2(n6696), .A(n6277), .B(n6276), .ZN(U3043)
         );
  NOR2_X1 U7252 ( .A1(n6819), .A2(n6287), .ZN(n6282) );
  INV_X1 U7253 ( .A(n6282), .ZN(n6310) );
  OAI22_X1 U7254 ( .A1(n6471), .A2(n6310), .B1(n6326), .B2(n6601), .ZN(n6280)
         );
  INV_X1 U7255 ( .A(n6280), .ZN(n6291) );
  INV_X1 U7256 ( .A(n6281), .ZN(n6561) );
  OR2_X1 U7257 ( .A1(n6430), .A2(n6536), .ZN(n6348) );
  INV_X1 U7258 ( .A(n6348), .ZN(n6283) );
  AOI21_X1 U7259 ( .B1(n6561), .B2(n6283), .A(n6282), .ZN(n6289) );
  INV_X1 U7260 ( .A(n6289), .ZN(n6286) );
  AOI21_X1 U7261 ( .B1(n6802), .B2(n6287), .A(n6284), .ZN(n6285) );
  OAI21_X1 U7262 ( .B1(n6288), .B2(n6286), .A(n6285), .ZN(n6313) );
  OAI22_X1 U7263 ( .A1(n6289), .A2(n6288), .B1(n6478), .B2(n6287), .ZN(n6312)
         );
  AOI22_X1 U7264 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n6313), .B1(n6639), 
        .B2(n6312), .ZN(n6290) );
  OAI211_X1 U7265 ( .C1(n6649), .C2(n6316), .A(n6291), .B(n6290), .ZN(U3060)
         );
  OAI22_X1 U7266 ( .A1(n6485), .A2(n6310), .B1(n6326), .B2(n6605), .ZN(n6292)
         );
  INV_X1 U7267 ( .A(n6292), .ZN(n6294) );
  AOI22_X1 U7268 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n6313), .B1(n6651), 
        .B2(n6312), .ZN(n6293) );
  OAI211_X1 U7269 ( .C1(n6655), .C2(n6316), .A(n6294), .B(n6293), .ZN(U3061)
         );
  OAI22_X1 U7270 ( .A1(n6489), .A2(n6310), .B1(n6326), .B2(n6609), .ZN(n6295)
         );
  INV_X1 U7271 ( .A(n6295), .ZN(n6297) );
  AOI22_X1 U7272 ( .A1(INSTQUEUE_REG_5__2__SCAN_IN), .A2(n6313), .B1(n6657), 
        .B2(n6312), .ZN(n6296) );
  OAI211_X1 U7273 ( .C1(n6661), .C2(n6316), .A(n6297), .B(n6296), .ZN(U3062)
         );
  OAI22_X1 U7274 ( .A1(n6493), .A2(n6310), .B1(n6326), .B2(n6613), .ZN(n6298)
         );
  INV_X1 U7275 ( .A(n6298), .ZN(n6300) );
  AOI22_X1 U7276 ( .A1(INSTQUEUE_REG_5__3__SCAN_IN), .A2(n6313), .B1(n6663), 
        .B2(n6312), .ZN(n6299) );
  OAI211_X1 U7277 ( .C1(n6667), .C2(n6316), .A(n6300), .B(n6299), .ZN(U3063)
         );
  OAI22_X1 U7278 ( .A1(n6497), .A2(n6310), .B1(n6326), .B2(n6617), .ZN(n6301)
         );
  INV_X1 U7279 ( .A(n6301), .ZN(n6303) );
  AOI22_X1 U7280 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n6313), .B1(n6669), 
        .B2(n6312), .ZN(n6302) );
  OAI211_X1 U7281 ( .C1(n6673), .C2(n6316), .A(n6303), .B(n6302), .ZN(U3064)
         );
  OAI22_X1 U7282 ( .A1(n6501), .A2(n6310), .B1(n6326), .B2(n6621), .ZN(n6304)
         );
  INV_X1 U7283 ( .A(n6304), .ZN(n6306) );
  AOI22_X1 U7284 ( .A1(INSTQUEUE_REG_5__5__SCAN_IN), .A2(n6313), .B1(n6675), 
        .B2(n6312), .ZN(n6305) );
  OAI211_X1 U7285 ( .C1(n6679), .C2(n6316), .A(n6306), .B(n6305), .ZN(U3065)
         );
  OAI22_X1 U7286 ( .A1(n6505), .A2(n6310), .B1(n6326), .B2(n6625), .ZN(n6307)
         );
  INV_X1 U7287 ( .A(n6307), .ZN(n6309) );
  AOI22_X1 U7288 ( .A1(INSTQUEUE_REG_5__6__SCAN_IN), .A2(n6313), .B1(n6681), 
        .B2(n6312), .ZN(n6308) );
  OAI211_X1 U7289 ( .C1(n6685), .C2(n6316), .A(n6309), .B(n6308), .ZN(U3066)
         );
  OAI22_X1 U7290 ( .A1(n6510), .A2(n6310), .B1(n6326), .B2(n6633), .ZN(n6311)
         );
  INV_X1 U7291 ( .A(n6311), .ZN(n6315) );
  AOI22_X1 U7292 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n6313), .B1(n6689), 
        .B2(n6312), .ZN(n6314) );
  OAI211_X1 U7293 ( .C1(n6696), .C2(n6316), .A(n6315), .B(n6314), .ZN(U3067)
         );
  OR2_X1 U7294 ( .A1(n3907), .A2(n3940), .ZN(n6349) );
  INV_X1 U7295 ( .A(n6349), .ZN(n6635) );
  NAND2_X1 U7296 ( .A1(n6635), .A2(n6812), .ZN(n6592) );
  INV_X1 U7297 ( .A(n6317), .ZN(n6591) );
  OAI22_X1 U7298 ( .A1(n6592), .A2(n6319), .B1(n6591), .B2(n6318), .ZN(n6342)
         );
  NAND2_X1 U7299 ( .A1(n6819), .A2(n6357), .ZN(n6322) );
  INV_X1 U7300 ( .A(n6322), .ZN(n6341) );
  AOI22_X1 U7301 ( .A1(n6639), .A2(n6342), .B1(n6638), .B2(n6341), .ZN(n6328)
         );
  NAND3_X1 U7302 ( .A1(n6326), .A2(n6812), .A3(n6386), .ZN(n6320) );
  AOI21_X1 U7303 ( .B1(n6805), .B2(n6320), .A(n6635), .ZN(n6321) );
  AOI21_X1 U7304 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6322), .A(n6321), .ZN(
        n6325) );
  NOR2_X1 U7305 ( .A1(n6324), .A2(n6323), .ZN(n6597) );
  NAND3_X1 U7306 ( .A1(n6810), .A2(n6325), .A3(n6597), .ZN(n6344) );
  AOI22_X1 U7307 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n6344), .B1(n6598), 
        .B2(n6343), .ZN(n6327) );
  OAI211_X1 U7308 ( .C1(n6601), .C2(n6386), .A(n6328), .B(n6327), .ZN(U3068)
         );
  AOI22_X1 U7309 ( .A1(n6651), .A2(n6342), .B1(n6650), .B2(n6341), .ZN(n6330)
         );
  AOI22_X1 U7310 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(n6344), .B1(n6602), 
        .B2(n6343), .ZN(n6329) );
  OAI211_X1 U7311 ( .C1(n6605), .C2(n6386), .A(n6330), .B(n6329), .ZN(U3069)
         );
  AOI22_X1 U7312 ( .A1(n6657), .A2(n6342), .B1(n6656), .B2(n6341), .ZN(n6332)
         );
  AOI22_X1 U7313 ( .A1(INSTQUEUE_REG_6__2__SCAN_IN), .A2(n6344), .B1(n6606), 
        .B2(n6343), .ZN(n6331) );
  OAI211_X1 U7314 ( .C1(n6609), .C2(n6386), .A(n6332), .B(n6331), .ZN(U3070)
         );
  AOI22_X1 U7315 ( .A1(n6663), .A2(n6342), .B1(n6662), .B2(n6341), .ZN(n6334)
         );
  AOI22_X1 U7316 ( .A1(INSTQUEUE_REG_6__3__SCAN_IN), .A2(n6344), .B1(n6610), 
        .B2(n6343), .ZN(n6333) );
  OAI211_X1 U7317 ( .C1(n6613), .C2(n6386), .A(n6334), .B(n6333), .ZN(U3071)
         );
  AOI22_X1 U7318 ( .A1(n6669), .A2(n6342), .B1(n6668), .B2(n6341), .ZN(n6336)
         );
  AOI22_X1 U7319 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n6344), .B1(n6614), 
        .B2(n6343), .ZN(n6335) );
  OAI211_X1 U7320 ( .C1(n6617), .C2(n6386), .A(n6336), .B(n6335), .ZN(U3072)
         );
  AOI22_X1 U7321 ( .A1(n6675), .A2(n6342), .B1(n6674), .B2(n6341), .ZN(n6338)
         );
  AOI22_X1 U7322 ( .A1(INSTQUEUE_REG_6__5__SCAN_IN), .A2(n6344), .B1(n6618), 
        .B2(n6343), .ZN(n6337) );
  OAI211_X1 U7323 ( .C1(n6621), .C2(n6386), .A(n6338), .B(n6337), .ZN(U3073)
         );
  AOI22_X1 U7324 ( .A1(n6681), .A2(n6342), .B1(n6680), .B2(n6341), .ZN(n6340)
         );
  AOI22_X1 U7325 ( .A1(INSTQUEUE_REG_6__6__SCAN_IN), .A2(n6344), .B1(n6622), 
        .B2(n6343), .ZN(n6339) );
  OAI211_X1 U7326 ( .C1(n6625), .C2(n6386), .A(n6340), .B(n6339), .ZN(U3074)
         );
  AOI22_X1 U7327 ( .A1(n6689), .A2(n6342), .B1(n6686), .B2(n6341), .ZN(n6346)
         );
  AOI22_X1 U7328 ( .A1(INSTQUEUE_REG_6__7__SCAN_IN), .A2(n6344), .B1(n6629), 
        .B2(n6343), .ZN(n6345) );
  OAI211_X1 U7329 ( .C1(n6633), .C2(n6386), .A(n6346), .B(n6345), .ZN(U3075)
         );
  NOR2_X1 U7330 ( .A1(n6351), .A2(n6347), .ZN(n6799) );
  NOR2_X1 U7331 ( .A1(n6799), .A2(n6802), .ZN(n6355) );
  OAI21_X1 U7332 ( .B1(n6349), .B2(n6348), .A(n6387), .ZN(n6353) );
  AOI22_X1 U7333 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6357), .B1(n6355), .B2(
        n6353), .ZN(n6393) );
  OR2_X1 U7334 ( .A1(n6351), .A2(n6350), .ZN(n6401) );
  OAI22_X1 U7335 ( .A1(n6471), .A2(n6387), .B1(n6601), .B2(n6401), .ZN(n6352)
         );
  INV_X1 U7336 ( .A(n6352), .ZN(n6359) );
  INV_X1 U7337 ( .A(n6353), .ZN(n6354) );
  NAND2_X1 U7338 ( .A1(n6355), .A2(n6354), .ZN(n6356) );
  OAI211_X1 U7339 ( .C1(n6357), .C2(n6812), .A(n6645), .B(n6356), .ZN(n6389)
         );
  INV_X1 U7340 ( .A(n6386), .ZN(n6362) );
  AOI22_X1 U7341 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6389), .B1(n6598), 
        .B2(n6362), .ZN(n6358) );
  OAI211_X1 U7342 ( .C1(n6393), .C2(n6360), .A(n6359), .B(n6358), .ZN(U3076)
         );
  OAI22_X1 U7343 ( .A1(n6485), .A2(n6387), .B1(n6605), .B2(n6401), .ZN(n6361)
         );
  INV_X1 U7344 ( .A(n6361), .ZN(n6364) );
  AOI22_X1 U7345 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6389), .B1(n6602), 
        .B2(n6362), .ZN(n6363) );
  OAI211_X1 U7346 ( .C1(n6393), .C2(n6365), .A(n6364), .B(n6363), .ZN(U3077)
         );
  OAI22_X1 U7347 ( .A1(n6489), .A2(n6387), .B1(n6661), .B2(n6386), .ZN(n6366)
         );
  INV_X1 U7348 ( .A(n6366), .ZN(n6368) );
  AOI22_X1 U7349 ( .A1(n6389), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n6658), 
        .B2(n6423), .ZN(n6367) );
  OAI211_X1 U7350 ( .C1(n6393), .C2(n6369), .A(n6368), .B(n6367), .ZN(U3078)
         );
  OAI22_X1 U7351 ( .A1(n6493), .A2(n6387), .B1(n6667), .B2(n6386), .ZN(n6370)
         );
  INV_X1 U7352 ( .A(n6370), .ZN(n6372) );
  AOI22_X1 U7353 ( .A1(n6389), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n6664), 
        .B2(n6423), .ZN(n6371) );
  OAI211_X1 U7354 ( .C1(n6393), .C2(n6373), .A(n6372), .B(n6371), .ZN(U3079)
         );
  OAI22_X1 U7355 ( .A1(n6497), .A2(n6387), .B1(n6673), .B2(n6386), .ZN(n6374)
         );
  INV_X1 U7356 ( .A(n6374), .ZN(n6376) );
  AOI22_X1 U7357 ( .A1(n6389), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n6670), 
        .B2(n6423), .ZN(n6375) );
  OAI211_X1 U7358 ( .C1(n6393), .C2(n6377), .A(n6376), .B(n6375), .ZN(U3080)
         );
  OAI22_X1 U7359 ( .A1(n6501), .A2(n6387), .B1(n6679), .B2(n6386), .ZN(n6378)
         );
  INV_X1 U7360 ( .A(n6378), .ZN(n6380) );
  AOI22_X1 U7361 ( .A1(n6389), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n6676), 
        .B2(n6423), .ZN(n6379) );
  OAI211_X1 U7362 ( .C1(n6393), .C2(n6381), .A(n6380), .B(n6379), .ZN(U3081)
         );
  OAI22_X1 U7363 ( .A1(n6505), .A2(n6387), .B1(n6685), .B2(n6386), .ZN(n6382)
         );
  INV_X1 U7364 ( .A(n6382), .ZN(n6384) );
  AOI22_X1 U7365 ( .A1(n6389), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n6682), 
        .B2(n6423), .ZN(n6383) );
  OAI211_X1 U7366 ( .C1(n6393), .C2(n6385), .A(n6384), .B(n6383), .ZN(U3082)
         );
  OAI22_X1 U7367 ( .A1(n6510), .A2(n6387), .B1(n6696), .B2(n6386), .ZN(n6388)
         );
  INV_X1 U7368 ( .A(n6388), .ZN(n6391) );
  AOI22_X1 U7369 ( .A1(n6389), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n6691), 
        .B2(n6423), .ZN(n6390) );
  OAI211_X1 U7370 ( .C1(n6393), .C2(n6392), .A(n6391), .B(n6390), .ZN(U3083)
         );
  INV_X1 U7371 ( .A(n6432), .ZN(n6396) );
  NOR2_X1 U7372 ( .A1(n6396), .A2(n6804), .ZN(n6402) );
  INV_X1 U7373 ( .A(n6402), .ZN(n6399) );
  INV_X1 U7374 ( .A(n6480), .ZN(n6398) );
  NAND2_X1 U7375 ( .A1(n6398), .A2(n6397), .ZN(n6532) );
  OAI22_X1 U7376 ( .A1(n6399), .A2(n6802), .B1(n6538), .B2(n6532), .ZN(n6422)
         );
  NAND3_X1 U7377 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6704), .A3(n6400), .ZN(n6437) );
  NOR2_X1 U7378 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6437), .ZN(n6421)
         );
  AOI22_X1 U7379 ( .A1(n6639), .A2(n6422), .B1(n6638), .B2(n6421), .ZN(n6408)
         );
  AOI21_X1 U7380 ( .B1(n6464), .B2(n6401), .A(n6912), .ZN(n6403) );
  NOR3_X1 U7381 ( .A1(n6403), .A2(n6402), .A3(n6802), .ZN(n6406) );
  AOI21_X1 U7382 ( .B1(n6532), .B2(STATE2_REG_2__SCAN_IN), .A(n6404), .ZN(
        n6537) );
  OAI211_X1 U7383 ( .C1(n6798), .C2(n6421), .A(n6591), .B(n6537), .ZN(n6405)
         );
  AOI22_X1 U7384 ( .A1(n6424), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n6598), 
        .B2(n6423), .ZN(n6407) );
  OAI211_X1 U7385 ( .C1(n6601), .C2(n6464), .A(n6408), .B(n6407), .ZN(U3084)
         );
  AOI22_X1 U7386 ( .A1(n6651), .A2(n6422), .B1(n6650), .B2(n6421), .ZN(n6410)
         );
  AOI22_X1 U7387 ( .A1(n6424), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n6602), 
        .B2(n6423), .ZN(n6409) );
  OAI211_X1 U7388 ( .C1(n6605), .C2(n6464), .A(n6410), .B(n6409), .ZN(U3085)
         );
  AOI22_X1 U7389 ( .A1(n6657), .A2(n6422), .B1(n6656), .B2(n6421), .ZN(n6412)
         );
  AOI22_X1 U7390 ( .A1(n6424), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n6606), 
        .B2(n6423), .ZN(n6411) );
  OAI211_X1 U7391 ( .C1(n6609), .C2(n6464), .A(n6412), .B(n6411), .ZN(U3086)
         );
  AOI22_X1 U7392 ( .A1(n6663), .A2(n6422), .B1(n6662), .B2(n6421), .ZN(n6414)
         );
  AOI22_X1 U7393 ( .A1(n6424), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n6610), 
        .B2(n6423), .ZN(n6413) );
  OAI211_X1 U7394 ( .C1(n6613), .C2(n6464), .A(n6414), .B(n6413), .ZN(U3087)
         );
  AOI22_X1 U7395 ( .A1(n6669), .A2(n6422), .B1(n6668), .B2(n6421), .ZN(n6416)
         );
  AOI22_X1 U7396 ( .A1(n6424), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n6614), 
        .B2(n6423), .ZN(n6415) );
  OAI211_X1 U7397 ( .C1(n6617), .C2(n6464), .A(n6416), .B(n6415), .ZN(U3088)
         );
  AOI22_X1 U7398 ( .A1(n6675), .A2(n6422), .B1(n6674), .B2(n6421), .ZN(n6418)
         );
  AOI22_X1 U7399 ( .A1(n6424), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n6618), 
        .B2(n6423), .ZN(n6417) );
  OAI211_X1 U7400 ( .C1(n6621), .C2(n6464), .A(n6418), .B(n6417), .ZN(U3089)
         );
  AOI22_X1 U7401 ( .A1(n6681), .A2(n6422), .B1(n6680), .B2(n6421), .ZN(n6420)
         );
  AOI22_X1 U7402 ( .A1(n6424), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n6622), 
        .B2(n6423), .ZN(n6419) );
  OAI211_X1 U7403 ( .C1(n6625), .C2(n6464), .A(n6420), .B(n6419), .ZN(U3090)
         );
  AOI22_X1 U7404 ( .A1(n6689), .A2(n6422), .B1(n6686), .B2(n6421), .ZN(n6426)
         );
  AOI22_X1 U7405 ( .A1(n6424), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n6629), 
        .B2(n6423), .ZN(n6425) );
  OAI211_X1 U7406 ( .C1(n6633), .C2(n6464), .A(n6426), .B(n6425), .ZN(U3091)
         );
  INV_X1 U7407 ( .A(n6427), .ZN(n6434) );
  NOR2_X1 U7408 ( .A1(n3935), .A2(n6589), .ZN(n6428) );
  NOR2_X1 U7409 ( .A1(n6819), .A2(n6437), .ZN(n6431) );
  INV_X1 U7410 ( .A(n6431), .ZN(n6463) );
  OAI22_X1 U7411 ( .A1(n6464), .A2(n6649), .B1(n6471), .B2(n6463), .ZN(n6429)
         );
  INV_X1 U7412 ( .A(n6429), .ZN(n6441) );
  NOR2_X1 U7413 ( .A1(n6804), .A2(n6430), .ZN(n6636) );
  AOI21_X1 U7414 ( .B1(n6636), .B2(n6432), .A(n6431), .ZN(n6439) );
  NOR2_X1 U7415 ( .A1(n3935), .A2(n6912), .ZN(n6433) );
  AOI21_X1 U7416 ( .B1(n6434), .B2(n6433), .A(n6802), .ZN(n6436) );
  AOI22_X1 U7417 ( .A1(n6439), .A2(n6436), .B1(n6802), .B2(n6437), .ZN(n6435)
         );
  NAND2_X1 U7418 ( .A1(n6645), .A2(n6435), .ZN(n6467) );
  INV_X1 U7419 ( .A(n6436), .ZN(n6438) );
  OAI22_X1 U7420 ( .A1(n6439), .A2(n6438), .B1(n6478), .B2(n6437), .ZN(n6466)
         );
  AOI22_X1 U7421 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n6467), .B1(n6639), 
        .B2(n6466), .ZN(n6440) );
  OAI211_X1 U7422 ( .C1(n6601), .C2(n6516), .A(n6441), .B(n6440), .ZN(U3092)
         );
  OR2_X1 U7423 ( .A1(n6485), .A2(n6463), .ZN(n6442) );
  OAI21_X1 U7424 ( .B1(n6516), .B2(n6605), .A(n6442), .ZN(n6443) );
  INV_X1 U7425 ( .A(n6443), .ZN(n6445) );
  AOI22_X1 U7426 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n6467), .B1(n6651), 
        .B2(n6466), .ZN(n6444) );
  OAI211_X1 U7427 ( .C1(n6655), .C2(n6464), .A(n6445), .B(n6444), .ZN(U3093)
         );
  OR2_X1 U7428 ( .A1(n6489), .A2(n6463), .ZN(n6446) );
  OAI21_X1 U7429 ( .B1(n6516), .B2(n6609), .A(n6446), .ZN(n6447) );
  INV_X1 U7430 ( .A(n6447), .ZN(n6449) );
  AOI22_X1 U7431 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n6467), .B1(n6657), 
        .B2(n6466), .ZN(n6448) );
  OAI211_X1 U7432 ( .C1(n6661), .C2(n6464), .A(n6449), .B(n6448), .ZN(U3094)
         );
  OAI22_X1 U7433 ( .A1(n6464), .A2(n6667), .B1(n6493), .B2(n6463), .ZN(n6450)
         );
  INV_X1 U7434 ( .A(n6450), .ZN(n6452) );
  AOI22_X1 U7435 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n6467), .B1(n6663), 
        .B2(n6466), .ZN(n6451) );
  OAI211_X1 U7436 ( .C1(n6613), .C2(n6516), .A(n6452), .B(n6451), .ZN(U3095)
         );
  OAI22_X1 U7437 ( .A1(n6464), .A2(n6673), .B1(n6497), .B2(n6463), .ZN(n6453)
         );
  INV_X1 U7438 ( .A(n6453), .ZN(n6455) );
  AOI22_X1 U7439 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n6467), .B1(n6669), 
        .B2(n6466), .ZN(n6454) );
  OAI211_X1 U7440 ( .C1(n6617), .C2(n6516), .A(n6455), .B(n6454), .ZN(U3096)
         );
  OAI22_X1 U7441 ( .A1(n6464), .A2(n6679), .B1(n6501), .B2(n6463), .ZN(n6456)
         );
  INV_X1 U7442 ( .A(n6456), .ZN(n6458) );
  AOI22_X1 U7443 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n6467), .B1(n6675), 
        .B2(n6466), .ZN(n6457) );
  OAI211_X1 U7444 ( .C1(n6621), .C2(n6516), .A(n6458), .B(n6457), .ZN(U3097)
         );
  OR2_X1 U7445 ( .A1(n6505), .A2(n6463), .ZN(n6459) );
  OAI21_X1 U7446 ( .B1(n6516), .B2(n6625), .A(n6459), .ZN(n6460) );
  INV_X1 U7447 ( .A(n6460), .ZN(n6462) );
  AOI22_X1 U7448 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n6467), .B1(n6681), 
        .B2(n6466), .ZN(n6461) );
  OAI211_X1 U7449 ( .C1(n6685), .C2(n6464), .A(n6462), .B(n6461), .ZN(U3098)
         );
  OAI22_X1 U7450 ( .A1(n6464), .A2(n6696), .B1(n6510), .B2(n6463), .ZN(n6465)
         );
  INV_X1 U7451 ( .A(n6465), .ZN(n6469) );
  AOI22_X1 U7452 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n6467), .B1(n6689), 
        .B2(n6466), .ZN(n6468) );
  OAI211_X1 U7453 ( .C1(n6633), .C2(n6516), .A(n6469), .B(n6468), .ZN(U3099)
         );
  NOR2_X1 U7454 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6470), .ZN(n6474)
         );
  INV_X1 U7455 ( .A(n6474), .ZN(n6509) );
  OAI22_X1 U7456 ( .A1(n6530), .A2(n6601), .B1(n6471), .B2(n6509), .ZN(n6472)
         );
  INV_X1 U7457 ( .A(n6472), .ZN(n6484) );
  NAND2_X1 U7458 ( .A1(n6530), .A2(n6516), .ZN(n6473) );
  AOI21_X1 U7459 ( .B1(n6473), .B2(STATEBS16_REG_SCAN_IN), .A(n6802), .ZN(
        n6479) );
  NOR2_X1 U7460 ( .A1(n6474), .A2(n6798), .ZN(n6475) );
  AOI21_X1 U7461 ( .B1(n6479), .B2(n6481), .A(n6475), .ZN(n6476) );
  OAI211_X1 U7462 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6478), .A(n6477), .B(n6476), .ZN(n6513) );
  INV_X1 U7463 ( .A(n6479), .ZN(n6482) );
  NAND2_X1 U7464 ( .A1(n6480), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6590) );
  OAI22_X1 U7465 ( .A1(n6482), .A2(n6481), .B1(n6538), .B2(n6590), .ZN(n6512)
         );
  AOI22_X1 U7466 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n6513), .B1(n6639), 
        .B2(n6512), .ZN(n6483) );
  OAI211_X1 U7467 ( .C1(n6649), .C2(n6516), .A(n6484), .B(n6483), .ZN(U3100)
         );
  OAI22_X1 U7468 ( .A1(n6530), .A2(n6605), .B1(n6485), .B2(n6509), .ZN(n6486)
         );
  INV_X1 U7469 ( .A(n6486), .ZN(n6488) );
  AOI22_X1 U7470 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(n6513), .B1(n6651), 
        .B2(n6512), .ZN(n6487) );
  OAI211_X1 U7471 ( .C1(n6655), .C2(n6516), .A(n6488), .B(n6487), .ZN(U3101)
         );
  OAI22_X1 U7472 ( .A1(n6530), .A2(n6609), .B1(n6489), .B2(n6509), .ZN(n6490)
         );
  INV_X1 U7473 ( .A(n6490), .ZN(n6492) );
  AOI22_X1 U7474 ( .A1(INSTQUEUE_REG_10__2__SCAN_IN), .A2(n6513), .B1(n6657), 
        .B2(n6512), .ZN(n6491) );
  OAI211_X1 U7475 ( .C1(n6661), .C2(n6516), .A(n6492), .B(n6491), .ZN(U3102)
         );
  OAI22_X1 U7476 ( .A1(n6530), .A2(n6613), .B1(n6493), .B2(n6509), .ZN(n6494)
         );
  INV_X1 U7477 ( .A(n6494), .ZN(n6496) );
  AOI22_X1 U7478 ( .A1(INSTQUEUE_REG_10__3__SCAN_IN), .A2(n6513), .B1(n6663), 
        .B2(n6512), .ZN(n6495) );
  OAI211_X1 U7479 ( .C1(n6667), .C2(n6516), .A(n6496), .B(n6495), .ZN(U3103)
         );
  OAI22_X1 U7480 ( .A1(n6530), .A2(n6617), .B1(n6497), .B2(n6509), .ZN(n6498)
         );
  INV_X1 U7481 ( .A(n6498), .ZN(n6500) );
  AOI22_X1 U7482 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n6513), .B1(n6669), 
        .B2(n6512), .ZN(n6499) );
  OAI211_X1 U7483 ( .C1(n6673), .C2(n6516), .A(n6500), .B(n6499), .ZN(U3104)
         );
  OAI22_X1 U7484 ( .A1(n6530), .A2(n6621), .B1(n6501), .B2(n6509), .ZN(n6502)
         );
  INV_X1 U7485 ( .A(n6502), .ZN(n6504) );
  AOI22_X1 U7486 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(n6513), .B1(n6675), 
        .B2(n6512), .ZN(n6503) );
  OAI211_X1 U7487 ( .C1(n6679), .C2(n6516), .A(n6504), .B(n6503), .ZN(U3105)
         );
  OAI22_X1 U7488 ( .A1(n6530), .A2(n6625), .B1(n6505), .B2(n6509), .ZN(n6506)
         );
  INV_X1 U7489 ( .A(n6506), .ZN(n6508) );
  AOI22_X1 U7490 ( .A1(INSTQUEUE_REG_10__6__SCAN_IN), .A2(n6513), .B1(n6681), 
        .B2(n6512), .ZN(n6507) );
  OAI211_X1 U7491 ( .C1(n6685), .C2(n6516), .A(n6508), .B(n6507), .ZN(U3106)
         );
  OAI22_X1 U7492 ( .A1(n6530), .A2(n6633), .B1(n6510), .B2(n6509), .ZN(n6511)
         );
  INV_X1 U7493 ( .A(n6511), .ZN(n6515) );
  AOI22_X1 U7494 ( .A1(INSTQUEUE_REG_10__7__SCAN_IN), .A2(n6513), .B1(n6689), 
        .B2(n6512), .ZN(n6514) );
  OAI211_X1 U7495 ( .C1(n6696), .C2(n6516), .A(n6515), .B(n6514), .ZN(U3107)
         );
  AOI22_X1 U7496 ( .A1(n6638), .A2(n6525), .B1(n6557), .B2(n6646), .ZN(n6518)
         );
  AOI22_X1 U7497 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6527), .B1(n6639), 
        .B2(n6526), .ZN(n6517) );
  OAI211_X1 U7498 ( .C1(n6649), .C2(n6530), .A(n6518), .B(n6517), .ZN(U3108)
         );
  AOI22_X1 U7499 ( .A1(n6650), .A2(n6525), .B1(n6557), .B2(n6652), .ZN(n6520)
         );
  AOI22_X1 U7500 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6527), .B1(n6651), 
        .B2(n6526), .ZN(n6519) );
  OAI211_X1 U7501 ( .C1(n6655), .C2(n6530), .A(n6520), .B(n6519), .ZN(U3109)
         );
  AOI22_X1 U7502 ( .A1(n6656), .A2(n6525), .B1(n6557), .B2(n6658), .ZN(n6522)
         );
  AOI22_X1 U7503 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6527), .B1(n6657), 
        .B2(n6526), .ZN(n6521) );
  OAI211_X1 U7504 ( .C1(n6661), .C2(n6530), .A(n6522), .B(n6521), .ZN(U3110)
         );
  AOI22_X1 U7505 ( .A1(n6662), .A2(n6525), .B1(n6557), .B2(n6664), .ZN(n6524)
         );
  AOI22_X1 U7506 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6527), .B1(n6663), 
        .B2(n6526), .ZN(n6523) );
  OAI211_X1 U7507 ( .C1(n6667), .C2(n6530), .A(n6524), .B(n6523), .ZN(U3111)
         );
  AOI22_X1 U7508 ( .A1(n6668), .A2(n6525), .B1(n6557), .B2(n6670), .ZN(n6529)
         );
  AOI22_X1 U7509 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6527), .B1(n6669), 
        .B2(n6526), .ZN(n6528) );
  OAI211_X1 U7510 ( .C1(n6673), .C2(n6530), .A(n6529), .B(n6528), .ZN(U3112)
         );
  INV_X1 U7511 ( .A(n6531), .ZN(n6533) );
  OAI22_X1 U7512 ( .A1(n6533), .A2(n6804), .B1(n6532), .B2(n6591), .ZN(n6556)
         );
  NOR2_X1 U7513 ( .A1(n6810), .A2(n6562), .ZN(n6567) );
  AND2_X1 U7514 ( .A1(n6819), .A2(n6567), .ZN(n6555) );
  AOI22_X1 U7515 ( .A1(n6639), .A2(n6556), .B1(n6638), .B2(n6555), .ZN(n6542)
         );
  INV_X1 U7516 ( .A(n6557), .ZN(n6534) );
  AOI21_X1 U7517 ( .B1(n6534), .B2(n6588), .A(n6912), .ZN(n6535) );
  AOI211_X1 U7518 ( .C1(n6561), .C2(n6536), .A(n6802), .B(n6535), .ZN(n6540)
         );
  OAI211_X1 U7519 ( .C1(n6798), .C2(n6555), .A(n6538), .B(n6537), .ZN(n6539)
         );
  AOI22_X1 U7520 ( .A1(n6558), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n6598), 
        .B2(n6557), .ZN(n6541) );
  OAI211_X1 U7521 ( .C1(n6601), .C2(n6588), .A(n6542), .B(n6541), .ZN(U3116)
         );
  AOI22_X1 U7522 ( .A1(n6651), .A2(n6556), .B1(n6650), .B2(n6555), .ZN(n6544)
         );
  AOI22_X1 U7523 ( .A1(n6558), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n6602), 
        .B2(n6557), .ZN(n6543) );
  OAI211_X1 U7524 ( .C1(n6605), .C2(n6588), .A(n6544), .B(n6543), .ZN(U3117)
         );
  AOI22_X1 U7525 ( .A1(n6657), .A2(n6556), .B1(n6656), .B2(n6555), .ZN(n6546)
         );
  AOI22_X1 U7526 ( .A1(n6558), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n6606), 
        .B2(n6557), .ZN(n6545) );
  OAI211_X1 U7527 ( .C1(n6609), .C2(n6588), .A(n6546), .B(n6545), .ZN(U3118)
         );
  AOI22_X1 U7528 ( .A1(n6663), .A2(n6556), .B1(n6662), .B2(n6555), .ZN(n6548)
         );
  AOI22_X1 U7529 ( .A1(n6558), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n6610), 
        .B2(n6557), .ZN(n6547) );
  OAI211_X1 U7530 ( .C1(n6613), .C2(n6588), .A(n6548), .B(n6547), .ZN(U3119)
         );
  AOI22_X1 U7531 ( .A1(n6669), .A2(n6556), .B1(n6668), .B2(n6555), .ZN(n6550)
         );
  AOI22_X1 U7532 ( .A1(n6558), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n6614), 
        .B2(n6557), .ZN(n6549) );
  OAI211_X1 U7533 ( .C1(n6617), .C2(n6588), .A(n6550), .B(n6549), .ZN(U3120)
         );
  AOI22_X1 U7534 ( .A1(n6675), .A2(n6556), .B1(n6674), .B2(n6555), .ZN(n6552)
         );
  AOI22_X1 U7535 ( .A1(n6558), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n6618), 
        .B2(n6557), .ZN(n6551) );
  OAI211_X1 U7536 ( .C1(n6621), .C2(n6588), .A(n6552), .B(n6551), .ZN(U3121)
         );
  AOI22_X1 U7537 ( .A1(n6681), .A2(n6556), .B1(n6680), .B2(n6555), .ZN(n6554)
         );
  AOI22_X1 U7538 ( .A1(n6558), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n6622), 
        .B2(n6557), .ZN(n6553) );
  OAI211_X1 U7539 ( .C1(n6625), .C2(n6588), .A(n6554), .B(n6553), .ZN(U3122)
         );
  AOI22_X1 U7540 ( .A1(n6689), .A2(n6556), .B1(n6686), .B2(n6555), .ZN(n6560)
         );
  AOI22_X1 U7541 ( .A1(n6558), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n6629), 
        .B2(n6557), .ZN(n6559) );
  OAI211_X1 U7542 ( .C1(n6633), .C2(n6588), .A(n6560), .B(n6559), .ZN(U3123)
         );
  AND2_X1 U7543 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6567), .ZN(n6583)
         );
  AOI21_X1 U7544 ( .B1(n6636), .B2(n6561), .A(n6583), .ZN(n6565) );
  NAND2_X1 U7545 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6563) );
  OAI22_X1 U7546 ( .A1(n6565), .A2(n6802), .B1(n6563), .B2(n6562), .ZN(n6584)
         );
  AOI22_X1 U7547 ( .A1(n6639), .A2(n6584), .B1(n6638), .B2(n6583), .ZN(n6570)
         );
  NAND2_X1 U7548 ( .A1(n6565), .A2(n6564), .ZN(n6566) );
  OAI221_X1 U7549 ( .B1(n6812), .B2(n6567), .C1(n6802), .C2(n6566), .A(n6645), 
        .ZN(n6585) );
  OR2_X1 U7550 ( .A1(n6568), .A2(n6589), .ZN(n6593) );
  AOI22_X1 U7551 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n6585), .B1(n6646), 
        .B2(n6628), .ZN(n6569) );
  OAI211_X1 U7552 ( .C1(n6649), .C2(n6588), .A(n6570), .B(n6569), .ZN(U3124)
         );
  AOI22_X1 U7553 ( .A1(n6651), .A2(n6584), .B1(n6650), .B2(n6583), .ZN(n6572)
         );
  AOI22_X1 U7554 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n6585), .B1(n6652), 
        .B2(n6628), .ZN(n6571) );
  OAI211_X1 U7555 ( .C1(n6655), .C2(n6588), .A(n6572), .B(n6571), .ZN(U3125)
         );
  AOI22_X1 U7556 ( .A1(n6657), .A2(n6584), .B1(n6656), .B2(n6583), .ZN(n6574)
         );
  AOI22_X1 U7557 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n6585), .B1(n6658), 
        .B2(n6628), .ZN(n6573) );
  OAI211_X1 U7558 ( .C1(n6661), .C2(n6588), .A(n6574), .B(n6573), .ZN(U3126)
         );
  AOI22_X1 U7559 ( .A1(n6663), .A2(n6584), .B1(n6662), .B2(n6583), .ZN(n6576)
         );
  AOI22_X1 U7560 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n6585), .B1(n6664), 
        .B2(n6628), .ZN(n6575) );
  OAI211_X1 U7561 ( .C1(n6667), .C2(n6588), .A(n6576), .B(n6575), .ZN(U3127)
         );
  AOI22_X1 U7562 ( .A1(n6669), .A2(n6584), .B1(n6668), .B2(n6583), .ZN(n6578)
         );
  AOI22_X1 U7563 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n6585), .B1(n6670), 
        .B2(n6628), .ZN(n6577) );
  OAI211_X1 U7564 ( .C1(n6673), .C2(n6588), .A(n6578), .B(n6577), .ZN(U3128)
         );
  AOI22_X1 U7565 ( .A1(n6675), .A2(n6584), .B1(n6674), .B2(n6583), .ZN(n6580)
         );
  AOI22_X1 U7566 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n6585), .B1(n6676), 
        .B2(n6628), .ZN(n6579) );
  OAI211_X1 U7567 ( .C1(n6679), .C2(n6588), .A(n6580), .B(n6579), .ZN(U3129)
         );
  AOI22_X1 U7568 ( .A1(n6681), .A2(n6584), .B1(n6680), .B2(n6583), .ZN(n6582)
         );
  AOI22_X1 U7569 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n6585), .B1(n6682), 
        .B2(n6628), .ZN(n6581) );
  OAI211_X1 U7570 ( .C1(n6685), .C2(n6588), .A(n6582), .B(n6581), .ZN(U3130)
         );
  AOI22_X1 U7571 ( .A1(n6689), .A2(n6584), .B1(n6686), .B2(n6583), .ZN(n6587)
         );
  AOI22_X1 U7572 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n6585), .B1(n6691), 
        .B2(n6628), .ZN(n6586) );
  OAI211_X1 U7573 ( .C1(n6696), .C2(n6588), .A(n6587), .B(n6586), .ZN(U3131)
         );
  OAI22_X1 U7574 ( .A1(n6592), .A2(n6804), .B1(n6591), .B2(n6590), .ZN(n6627)
         );
  NOR2_X1 U7575 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6641), .ZN(n6626)
         );
  AOI22_X1 U7576 ( .A1(n6639), .A2(n6627), .B1(n6638), .B2(n6626), .ZN(n6600)
         );
  AOI21_X1 U7577 ( .B1(n6695), .B2(n6593), .A(n6912), .ZN(n6594) );
  NOR3_X1 U7578 ( .A1(n6594), .A2(n6635), .A3(n6802), .ZN(n6595) );
  NOR2_X1 U7579 ( .A1(n6810), .A2(n6595), .ZN(n6596) );
  OAI211_X1 U7580 ( .C1(n6626), .C2(n6798), .A(n6597), .B(n6596), .ZN(n6630)
         );
  AOI22_X1 U7581 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n6630), .B1(n6598), 
        .B2(n6628), .ZN(n6599) );
  OAI211_X1 U7582 ( .C1(n6601), .C2(n6695), .A(n6600), .B(n6599), .ZN(U3132)
         );
  AOI22_X1 U7583 ( .A1(n6651), .A2(n6627), .B1(n6650), .B2(n6626), .ZN(n6604)
         );
  AOI22_X1 U7584 ( .A1(INSTQUEUE_REG_14__1__SCAN_IN), .A2(n6630), .B1(n6602), 
        .B2(n6628), .ZN(n6603) );
  OAI211_X1 U7585 ( .C1(n6605), .C2(n6695), .A(n6604), .B(n6603), .ZN(U3133)
         );
  AOI22_X1 U7586 ( .A1(n6657), .A2(n6627), .B1(n6656), .B2(n6626), .ZN(n6608)
         );
  AOI22_X1 U7587 ( .A1(INSTQUEUE_REG_14__2__SCAN_IN), .A2(n6630), .B1(n6606), 
        .B2(n6628), .ZN(n6607) );
  OAI211_X1 U7588 ( .C1(n6609), .C2(n6695), .A(n6608), .B(n6607), .ZN(U3134)
         );
  AOI22_X1 U7589 ( .A1(n6663), .A2(n6627), .B1(n6662), .B2(n6626), .ZN(n6612)
         );
  AOI22_X1 U7590 ( .A1(INSTQUEUE_REG_14__3__SCAN_IN), .A2(n6630), .B1(n6610), 
        .B2(n6628), .ZN(n6611) );
  OAI211_X1 U7591 ( .C1(n6613), .C2(n6695), .A(n6612), .B(n6611), .ZN(U3135)
         );
  AOI22_X1 U7592 ( .A1(n6669), .A2(n6627), .B1(n6668), .B2(n6626), .ZN(n6616)
         );
  AOI22_X1 U7593 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n6630), .B1(n6614), 
        .B2(n6628), .ZN(n6615) );
  OAI211_X1 U7594 ( .C1(n6617), .C2(n6695), .A(n6616), .B(n6615), .ZN(U3136)
         );
  AOI22_X1 U7595 ( .A1(n6675), .A2(n6627), .B1(n6674), .B2(n6626), .ZN(n6620)
         );
  AOI22_X1 U7596 ( .A1(INSTQUEUE_REG_14__5__SCAN_IN), .A2(n6630), .B1(n6618), 
        .B2(n6628), .ZN(n6619) );
  OAI211_X1 U7597 ( .C1(n6621), .C2(n6695), .A(n6620), .B(n6619), .ZN(U3137)
         );
  AOI22_X1 U7598 ( .A1(n6681), .A2(n6627), .B1(n6680), .B2(n6626), .ZN(n6624)
         );
  AOI22_X1 U7599 ( .A1(INSTQUEUE_REG_14__6__SCAN_IN), .A2(n6630), .B1(n6622), 
        .B2(n6628), .ZN(n6623) );
  OAI211_X1 U7600 ( .C1(n6625), .C2(n6695), .A(n6624), .B(n6623), .ZN(U3138)
         );
  AOI22_X1 U7601 ( .A1(n6689), .A2(n6627), .B1(n6686), .B2(n6626), .ZN(n6632)
         );
  AOI22_X1 U7602 ( .A1(INSTQUEUE_REG_14__7__SCAN_IN), .A2(n6630), .B1(n6629), 
        .B2(n6628), .ZN(n6631) );
  OAI211_X1 U7603 ( .C1(n6633), .C2(n6695), .A(n6632), .B(n6631), .ZN(U3139)
         );
  INV_X1 U7604 ( .A(n6634), .ZN(n6687) );
  AOI21_X1 U7605 ( .B1(n6636), .B2(n6635), .A(n6687), .ZN(n6643) );
  OAI22_X1 U7606 ( .A1(n6643), .A2(n6802), .B1(n6641), .B2(n6637), .ZN(n6688)
         );
  AOI22_X1 U7607 ( .A1(n6639), .A2(n6688), .B1(n6687), .B2(n6638), .ZN(n6648)
         );
  OAI21_X1 U7608 ( .B1(n6640), .B2(n5512), .A(n6805), .ZN(n6642) );
  AOI22_X1 U7609 ( .A1(n6643), .A2(n6642), .B1(n6641), .B2(n6802), .ZN(n6644)
         );
  NAND2_X1 U7610 ( .A1(n6645), .A2(n6644), .ZN(n6692) );
  AOI22_X1 U7611 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n6692), .B1(n6646), 
        .B2(n6690), .ZN(n6647) );
  OAI211_X1 U7612 ( .C1(n6649), .C2(n6695), .A(n6648), .B(n6647), .ZN(U3140)
         );
  AOI22_X1 U7613 ( .A1(n6651), .A2(n6688), .B1(n6687), .B2(n6650), .ZN(n6654)
         );
  AOI22_X1 U7614 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n6692), .B1(n6652), 
        .B2(n6690), .ZN(n6653) );
  OAI211_X1 U7615 ( .C1(n6655), .C2(n6695), .A(n6654), .B(n6653), .ZN(U3141)
         );
  AOI22_X1 U7616 ( .A1(n6657), .A2(n6688), .B1(n6687), .B2(n6656), .ZN(n6660)
         );
  AOI22_X1 U7617 ( .A1(INSTQUEUE_REG_15__2__SCAN_IN), .A2(n6692), .B1(n6658), 
        .B2(n6690), .ZN(n6659) );
  OAI211_X1 U7618 ( .C1(n6661), .C2(n6695), .A(n6660), .B(n6659), .ZN(U3142)
         );
  AOI22_X1 U7619 ( .A1(n6663), .A2(n6688), .B1(n6687), .B2(n6662), .ZN(n6666)
         );
  AOI22_X1 U7620 ( .A1(INSTQUEUE_REG_15__3__SCAN_IN), .A2(n6692), .B1(n6664), 
        .B2(n6690), .ZN(n6665) );
  OAI211_X1 U7621 ( .C1(n6667), .C2(n6695), .A(n6666), .B(n6665), .ZN(U3143)
         );
  AOI22_X1 U7622 ( .A1(n6669), .A2(n6688), .B1(n6687), .B2(n6668), .ZN(n6672)
         );
  AOI22_X1 U7623 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n6692), .B1(n6670), 
        .B2(n6690), .ZN(n6671) );
  OAI211_X1 U7624 ( .C1(n6673), .C2(n6695), .A(n6672), .B(n6671), .ZN(U3144)
         );
  AOI22_X1 U7625 ( .A1(n6675), .A2(n6688), .B1(n6687), .B2(n6674), .ZN(n6678)
         );
  AOI22_X1 U7626 ( .A1(INSTQUEUE_REG_15__5__SCAN_IN), .A2(n6692), .B1(n6676), 
        .B2(n6690), .ZN(n6677) );
  OAI211_X1 U7627 ( .C1(n6679), .C2(n6695), .A(n6678), .B(n6677), .ZN(U3145)
         );
  AOI22_X1 U7628 ( .A1(n6681), .A2(n6688), .B1(n6687), .B2(n6680), .ZN(n6684)
         );
  AOI22_X1 U7629 ( .A1(INSTQUEUE_REG_15__6__SCAN_IN), .A2(n6692), .B1(n6682), 
        .B2(n6690), .ZN(n6683) );
  OAI211_X1 U7630 ( .C1(n6685), .C2(n6695), .A(n6684), .B(n6683), .ZN(U3146)
         );
  AOI22_X1 U7631 ( .A1(n6689), .A2(n6688), .B1(n6687), .B2(n6686), .ZN(n6694)
         );
  AOI22_X1 U7632 ( .A1(INSTQUEUE_REG_15__7__SCAN_IN), .A2(n6692), .B1(n6691), 
        .B2(n6690), .ZN(n6693) );
  OAI211_X1 U7633 ( .C1(n6696), .C2(n6695), .A(n6694), .B(n6693), .ZN(U3147)
         );
  INV_X1 U7634 ( .A(n6711), .ZN(n6709) );
  INV_X1 U7635 ( .A(n6707), .ZN(n6705) );
  NOR3_X1 U7636 ( .A1(n6698), .A2(n6697), .A3(n6819), .ZN(n6701) );
  NAND2_X1 U7637 ( .A1(n6701), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6703) );
  OAI22_X1 U7638 ( .A1(n6701), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n6700), .B2(n6699), .ZN(n6702) );
  OAI211_X1 U7639 ( .C1(n6705), .C2(n6704), .A(n6703), .B(n6702), .ZN(n6706)
         );
  OAI21_X1 U7640 ( .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6707), .A(n6706), 
        .ZN(n6708) );
  OAI21_X1 U7641 ( .B1(n6709), .B2(n6810), .A(n6708), .ZN(n6710) );
  OAI21_X1 U7642 ( .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n6711), .A(n6710), 
        .ZN(n6722) );
  INV_X1 U7643 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6721) );
  NAND2_X1 U7644 ( .A1(n7029), .A2(n6712), .ZN(n6715) );
  AOI211_X1 U7645 ( .C1(n6716), .C2(n6715), .A(n6714), .B(n6713), .ZN(n6717)
         );
  NAND2_X1 U7646 ( .A1(n6718), .A2(n6717), .ZN(n6719) );
  AOI211_X1 U7647 ( .C1(n6722), .C2(n6721), .A(n6720), .B(n6719), .ZN(n6737)
         );
  NOR2_X1 U7648 ( .A1(n6724), .A2(n6723), .ZN(n6815) );
  OAI21_X1 U7649 ( .B1(n6726), .B2(n6725), .A(STATE2_REG_2__SCAN_IN), .ZN(
        n6727) );
  AOI221_X1 U7650 ( .B1(n6728), .B2(n6828), .C1(n7199), .C2(n6828), .A(n6727), 
        .ZN(n6731) );
  OAI221_X1 U7651 ( .B1(n6828), .B2(n6737), .C1(n6828), .C2(n6728), .A(n6731), 
        .ZN(n6797) );
  OAI21_X1 U7652 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n7199), .A(n6797), .ZN(
        n6740) );
  INV_X1 U7653 ( .A(n6729), .ZN(n6730) );
  AOI221_X1 U7654 ( .B1(n6815), .B2(STATE2_REG_0__SCAN_IN), .C1(n6740), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6730), .ZN(n6735) );
  INV_X1 U7655 ( .A(n6731), .ZN(n6732) );
  OAI211_X1 U7656 ( .C1(n6827), .C2(n6733), .A(n6828), .B(n6732), .ZN(n6734)
         );
  OAI211_X1 U7657 ( .C1(n6737), .C2(n6736), .A(n6735), .B(n6734), .ZN(U3148)
         );
  INV_X1 U7658 ( .A(n6797), .ZN(n6744) );
  AOI21_X1 U7659 ( .B1(n6739), .B2(n7199), .A(n6738), .ZN(n6743) );
  OAI211_X1 U7660 ( .C1(STATE2_REG_0__SCAN_IN), .C2(STATE2_REG_2__SCAN_IN), 
        .A(STATE2_REG_1__SCAN_IN), .B(n6740), .ZN(n6741) );
  OAI211_X1 U7661 ( .C1(n6744), .C2(n6743), .A(n6742), .B(n6741), .ZN(U3149)
         );
  OAI221_X1 U7662 ( .B1(STATE2_REG_2__SCAN_IN), .B2(STATE2_REG_0__SCAN_IN), 
        .C1(STATE2_REG_2__SCAN_IN), .C2(n7199), .A(n6795), .ZN(n6746) );
  OAI21_X1 U7663 ( .B1(n6747), .B2(n6746), .A(n6745), .ZN(U3150) );
  AND2_X1 U7664 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6791), .ZN(U3151) );
  AND2_X1 U7665 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6791), .ZN(U3152) );
  AND2_X1 U7666 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6791), .ZN(U3153) );
  AND2_X1 U7667 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6791), .ZN(U3154) );
  AND2_X1 U7668 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6791), .ZN(U3155) );
  AND2_X1 U7669 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6791), .ZN(U3156) );
  AND2_X1 U7670 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6791), .ZN(U3157) );
  AND2_X1 U7671 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6791), .ZN(U3158) );
  AND2_X1 U7672 ( .A1(n6791), .A2(DATAWIDTH_REG_23__SCAN_IN), .ZN(U3159) );
  AND2_X1 U7673 ( .A1(n6791), .A2(DATAWIDTH_REG_22__SCAN_IN), .ZN(U3160) );
  AND2_X1 U7674 ( .A1(n6791), .A2(DATAWIDTH_REG_21__SCAN_IN), .ZN(U3161) );
  INV_X1 U7675 ( .A(DATAWIDTH_REG_20__SCAN_IN), .ZN(n6945) );
  NOR2_X1 U7676 ( .A1(n6794), .A2(n6945), .ZN(U3162) );
  AND2_X1 U7677 ( .A1(n6791), .A2(DATAWIDTH_REG_19__SCAN_IN), .ZN(U3163) );
  AND2_X1 U7678 ( .A1(n6791), .A2(DATAWIDTH_REG_18__SCAN_IN), .ZN(U3164) );
  AND2_X1 U7679 ( .A1(n6791), .A2(DATAWIDTH_REG_17__SCAN_IN), .ZN(U3165) );
  INV_X1 U7680 ( .A(DATAWIDTH_REG_16__SCAN_IN), .ZN(n6998) );
  NOR2_X1 U7681 ( .A1(n6794), .A2(n6998), .ZN(U3166) );
  AND2_X1 U7682 ( .A1(n6791), .A2(DATAWIDTH_REG_15__SCAN_IN), .ZN(U3167) );
  AND2_X1 U7683 ( .A1(n6748), .A2(DATAWIDTH_REG_14__SCAN_IN), .ZN(U3168) );
  AND2_X1 U7684 ( .A1(n6748), .A2(DATAWIDTH_REG_13__SCAN_IN), .ZN(U3169) );
  AND2_X1 U7685 ( .A1(n6748), .A2(DATAWIDTH_REG_12__SCAN_IN), .ZN(U3170) );
  INV_X1 U7686 ( .A(DATAWIDTH_REG_11__SCAN_IN), .ZN(n6942) );
  NOR2_X1 U7687 ( .A1(n6794), .A2(n6942), .ZN(U3171) );
  AND2_X1 U7688 ( .A1(n6748), .A2(DATAWIDTH_REG_10__SCAN_IN), .ZN(U3172) );
  AND2_X1 U7689 ( .A1(n6791), .A2(DATAWIDTH_REG_9__SCAN_IN), .ZN(U3173) );
  AND2_X1 U7690 ( .A1(n6791), .A2(DATAWIDTH_REG_8__SCAN_IN), .ZN(U3174) );
  INV_X1 U7691 ( .A(DATAWIDTH_REG_7__SCAN_IN), .ZN(n7135) );
  NOR2_X1 U7692 ( .A1(n6794), .A2(n7135), .ZN(U3175) );
  INV_X1 U7693 ( .A(DATAWIDTH_REG_6__SCAN_IN), .ZN(n7177) );
  NOR2_X1 U7694 ( .A1(n6794), .A2(n7177), .ZN(U3176) );
  AND2_X1 U7695 ( .A1(n6791), .A2(DATAWIDTH_REG_5__SCAN_IN), .ZN(U3177) );
  AND2_X1 U7696 ( .A1(n6791), .A2(DATAWIDTH_REG_4__SCAN_IN), .ZN(U3178) );
  INV_X1 U7697 ( .A(DATAWIDTH_REG_3__SCAN_IN), .ZN(n7163) );
  NOR2_X1 U7698 ( .A1(n6794), .A2(n7163), .ZN(U3179) );
  INV_X1 U7699 ( .A(DATAWIDTH_REG_2__SCAN_IN), .ZN(n6931) );
  NOR2_X1 U7700 ( .A1(n6794), .A2(n6931), .ZN(U3180) );
  INV_X1 U7701 ( .A(n6749), .ZN(n6752) );
  NAND2_X1 U7702 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .ZN(n6754) );
  INV_X1 U7703 ( .A(n6754), .ZN(n6760) );
  AOI21_X1 U7704 ( .B1(HOLD), .B2(STATE_REG_2__SCAN_IN), .A(n6760), .ZN(n6751)
         );
  AND2_X1 U7705 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6753) );
  INV_X1 U7706 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n7154) );
  INV_X1 U7707 ( .A(NA_N), .ZN(n7160) );
  AOI211_X1 U7708 ( .C1(STATE_REG_2__SCAN_IN), .C2(n7160), .A(
        STATE_REG_0__SCAN_IN), .B(n6752), .ZN(n6764) );
  AOI221_X1 U7709 ( .B1(n6753), .B2(n7220), .C1(n7154), .C2(n7220), .A(n6764), 
        .ZN(n6750) );
  OAI21_X1 U7710 ( .B1(n6752), .B2(n6751), .A(n6750), .ZN(U3181) );
  AND2_X1 U7711 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6757) );
  AOI21_X1 U7712 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(STATE_REG_0__SCAN_IN), 
        .A(n6753), .ZN(n6756) );
  OAI211_X1 U7713 ( .C1(n6757), .C2(n6756), .A(n6755), .B(n6754), .ZN(U3182)
         );
  AOI221_X1 U7714 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n7199), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6759) );
  AOI221_X1 U7715 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6759), .C2(HOLD), .A(n6758), .ZN(n6763) );
  NAND3_X1 U7716 ( .A1(READY_N), .A2(STATE_REG_2__SCAN_IN), .A3(
        STATE_REG_1__SCAN_IN), .ZN(n6762) );
  NAND4_X1 U7717 ( .A1(REQUESTPENDING_REG_SCAN_IN), .A2(STATE_REG_0__SCAN_IN), 
        .A3(n6760), .A4(n7160), .ZN(n6761) );
  OAI211_X1 U7718 ( .C1(n6764), .C2(n6763), .A(n6762), .B(n6761), .ZN(U3183)
         );
  NAND2_X1 U7719 ( .A1(n7221), .A2(n6959), .ZN(n6789) );
  INV_X1 U7720 ( .A(ADDRESS_REG_0__SCAN_IN), .ZN(n7054) );
  OAI222_X1 U7721 ( .A1(n6789), .A2(n6765), .B1(n7054), .B2(n7221), .C1(n3739), 
        .C2(n6787), .ZN(U3184) );
  INV_X1 U7722 ( .A(ADDRESS_REG_1__SCAN_IN), .ZN(n7169) );
  OAI222_X1 U7723 ( .A1(n6787), .A2(n6765), .B1(n7169), .B2(n7221), .C1(n6766), 
        .C2(n6788), .ZN(U3185) );
  INV_X1 U7724 ( .A(ADDRESS_REG_2__SCAN_IN), .ZN(n7166) );
  OAI222_X1 U7725 ( .A1(n6787), .A2(n6766), .B1(n7166), .B2(n7221), .C1(n6767), 
        .C2(n6788), .ZN(U3186) );
  INV_X1 U7726 ( .A(ADDRESS_REG_3__SCAN_IN), .ZN(n6923) );
  OAI222_X1 U7727 ( .A1(n6787), .A2(n6767), .B1(n6923), .B2(n7221), .C1(n6768), 
        .C2(n6788), .ZN(U3187) );
  INV_X1 U7728 ( .A(ADDRESS_REG_4__SCAN_IN), .ZN(n7063) );
  OAI222_X1 U7729 ( .A1(n6789), .A2(n6770), .B1(n7063), .B2(n7221), .C1(n6768), 
        .C2(n6787), .ZN(U3188) );
  INV_X1 U7730 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n6769) );
  OAI222_X1 U7731 ( .A1(n6787), .A2(n6770), .B1(n6769), .B2(n7221), .C1(n6772), 
        .C2(n6788), .ZN(U3189) );
  INV_X1 U7732 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n6771) );
  OAI222_X1 U7733 ( .A1(n6787), .A2(n6772), .B1(n6771), .B2(n7221), .C1(n6773), 
        .C2(n6789), .ZN(U3190) );
  INV_X1 U7734 ( .A(ADDRESS_REG_7__SCAN_IN), .ZN(n6970) );
  INV_X1 U7735 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6774) );
  OAI222_X1 U7736 ( .A1(n6787), .A2(n6773), .B1(n6970), .B2(n7221), .C1(n6774), 
        .C2(n6788), .ZN(U3191) );
  INV_X1 U7737 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n7018) );
  OAI222_X1 U7738 ( .A1(n6787), .A2(n6774), .B1(n7018), .B2(n7221), .C1(n6775), 
        .C2(n6789), .ZN(U3192) );
  INV_X1 U7739 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n7183) );
  OAI222_X1 U7740 ( .A1(n6787), .A2(n6775), .B1(n7183), .B2(n7221), .C1(n6776), 
        .C2(n6789), .ZN(U3193) );
  INV_X1 U7741 ( .A(ADDRESS_REG_10__SCAN_IN), .ZN(n7046) );
  OAI222_X1 U7742 ( .A1(n6788), .A2(n4681), .B1(n7046), .B2(n7221), .C1(n6776), 
        .C2(n6787), .ZN(U3194) );
  INV_X1 U7743 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n7148) );
  OAI222_X1 U7744 ( .A1(n6787), .A2(n4681), .B1(n7148), .B2(n7221), .C1(n5113), 
        .C2(n6789), .ZN(U3195) );
  INV_X1 U7745 ( .A(ADDRESS_REG_12__SCAN_IN), .ZN(n6777) );
  OAI222_X1 U7746 ( .A1(n6787), .A2(n5113), .B1(n6777), .B2(n7221), .C1(n6778), 
        .C2(n6789), .ZN(U3196) );
  INV_X1 U7747 ( .A(ADDRESS_REG_13__SCAN_IN), .ZN(n6969) );
  OAI222_X1 U7748 ( .A1(n6787), .A2(n6778), .B1(n6969), .B2(n7221), .C1(n6779), 
        .C2(n6789), .ZN(U3197) );
  INV_X1 U7749 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n7180) );
  OAI222_X1 U7750 ( .A1(n6787), .A2(n6779), .B1(n7180), .B2(n7221), .C1(n6780), 
        .C2(n6788), .ZN(U3198) );
  INV_X1 U7751 ( .A(ADDRESS_REG_15__SCAN_IN), .ZN(n7150) );
  OAI222_X1 U7752 ( .A1(n6787), .A2(n6780), .B1(n7150), .B2(n7221), .C1(n6983), 
        .C2(n6788), .ZN(U3199) );
  INV_X1 U7753 ( .A(ADDRESS_REG_16__SCAN_IN), .ZN(n6781) );
  OAI222_X1 U7754 ( .A1(n6789), .A2(n6967), .B1(n6781), .B2(n7221), .C1(n6983), 
        .C2(n6787), .ZN(U3200) );
  INV_X1 U7755 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n6782) );
  OAI222_X1 U7756 ( .A1(n6788), .A2(n7043), .B1(n6782), .B2(n7221), .C1(n6967), 
        .C2(n6787), .ZN(U3201) );
  INV_X1 U7757 ( .A(ADDRESS_REG_18__SCAN_IN), .ZN(n6981) );
  OAI222_X1 U7758 ( .A1(n6787), .A2(n7043), .B1(n6981), .B2(n7221), .C1(n6783), 
        .C2(n6788), .ZN(U3202) );
  INV_X1 U7759 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n7013) );
  OAI222_X1 U7760 ( .A1(n6787), .A2(n6783), .B1(n7013), .B2(n7221), .C1(n7026), 
        .C2(n6788), .ZN(U3203) );
  INV_X1 U7761 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n6933) );
  OAI222_X1 U7762 ( .A1(n6787), .A2(n7026), .B1(n6933), .B2(n7221), .C1(n6784), 
        .C2(n6788), .ZN(U3204) );
  INV_X1 U7763 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n7179) );
  OAI222_X1 U7764 ( .A1(n6787), .A2(n6784), .B1(n7179), .B2(n7221), .C1(n7060), 
        .C2(n6788), .ZN(U3205) );
  INV_X1 U7765 ( .A(ADDRESS_REG_22__SCAN_IN), .ZN(n6984) );
  OAI222_X1 U7766 ( .A1(n6787), .A2(n7060), .B1(n6984), .B2(n7221), .C1(n7016), 
        .C2(n6788), .ZN(U3206) );
  INV_X1 U7767 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n7015) );
  OAI222_X1 U7768 ( .A1(n6788), .A2(n7164), .B1(n7015), .B2(n7221), .C1(n7016), 
        .C2(n6787), .ZN(U3207) );
  INV_X1 U7769 ( .A(ADDRESS_REG_24__SCAN_IN), .ZN(n7167) );
  OAI222_X1 U7770 ( .A1(n6787), .A2(n7164), .B1(n7167), .B2(n7221), .C1(n7053), 
        .C2(n6788), .ZN(U3208) );
  INV_X1 U7771 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n6785) );
  OAI222_X1 U7772 ( .A1(n6787), .A2(n7053), .B1(n6785), .B2(n7221), .C1(n7012), 
        .C2(n6788), .ZN(U3209) );
  INV_X1 U7773 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n7038) );
  OAI222_X1 U7774 ( .A1(n6787), .A2(n7012), .B1(n7038), .B2(n7221), .C1(n6786), 
        .C2(n6788), .ZN(U3210) );
  INV_X1 U7775 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n7031) );
  OAI222_X1 U7776 ( .A1(n6787), .A2(n6786), .B1(n7031), .B2(n7221), .C1(n6909), 
        .C2(n6788), .ZN(U3211) );
  INV_X1 U7777 ( .A(ADDRESS_REG_28__SCAN_IN), .ZN(n7182) );
  OAI222_X1 U7778 ( .A1(n6787), .A2(n6909), .B1(n7182), .B2(n7221), .C1(n6930), 
        .C2(n6788), .ZN(U3212) );
  INV_X1 U7779 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n7176) );
  OAI222_X1 U7780 ( .A1(n6789), .A2(n6918), .B1(n7176), .B2(n7221), .C1(n6930), 
        .C2(n6787), .ZN(U3213) );
  INV_X1 U7781 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n7025) );
  INV_X1 U7782 ( .A(BE_N_REG_2__SCAN_IN), .ZN(n7019) );
  AOI22_X1 U7783 ( .A1(n7221), .A2(n7025), .B1(n7019), .B2(n7220), .ZN(U3446)
         );
  INV_X1 U7784 ( .A(BE_N_REG_1__SCAN_IN), .ZN(n6997) );
  AOI22_X1 U7785 ( .A1(n7221), .A2(n7193), .B1(n6997), .B2(n7220), .ZN(U3447)
         );
  INV_X1 U7786 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6990) );
  INV_X1 U7787 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n7041) );
  AOI22_X1 U7788 ( .A1(n7221), .A2(n6990), .B1(n7041), .B2(n7220), .ZN(U3448)
         );
  INV_X1 U7789 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6792) );
  INV_X1 U7790 ( .A(n6793), .ZN(n6790) );
  AOI21_X1 U7791 ( .B1(n6792), .B2(n6791), .A(n6790), .ZN(U3451) );
  OAI21_X1 U7792 ( .B1(n6794), .B2(n6979), .A(n6793), .ZN(U3452) );
  OAI211_X1 U7793 ( .C1(n6798), .C2(n6797), .A(n6796), .B(n6795), .ZN(U3453)
         );
  NOR2_X1 U7794 ( .A1(n6800), .A2(n6799), .ZN(n6801) );
  OAI222_X1 U7795 ( .A1(n6806), .A2(n6805), .B1(n6804), .B2(n6803), .C1(n6802), 
        .C2(n6801), .ZN(n6807) );
  INV_X1 U7796 ( .A(n6807), .ZN(n6809) );
  AOI22_X1 U7797 ( .A1(n6818), .A2(n6810), .B1(n6809), .B2(n6808), .ZN(U3462)
         );
  AOI22_X1 U7798 ( .A1(n6814), .A2(n6813), .B1(n6812), .B2(n6811), .ZN(n6817)
         );
  NOR2_X1 U7799 ( .A1(n6818), .A2(n6815), .ZN(n6816) );
  AOI22_X1 U7800 ( .A1(n6819), .A2(n6818), .B1(n6817), .B2(n6816), .ZN(U3465)
         );
  AOI211_X1 U7801 ( .C1(REIP_REG_0__SCAN_IN), .C2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(REIP_REG_1__SCAN_IN), .B(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6820) );
  AOI21_X1 U7802 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6820), .ZN(n6821) );
  AOI22_X1 U7803 ( .A1(n6824), .A2(n6821), .B1(n7025), .B2(n6822), .ZN(U3468)
         );
  NOR2_X1 U7804 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .ZN(
        n6823) );
  AOI22_X1 U7805 ( .A1(n6824), .A2(n6823), .B1(n6990), .B2(n6822), .ZN(U3469)
         );
  INV_X1 U7806 ( .A(W_R_N_REG_SCAN_IN), .ZN(n7195) );
  AOI22_X1 U7807 ( .A1(n7221), .A2(READREQUEST_REG_SCAN_IN), .B1(n7195), .B2(
        n7220), .ZN(U3470) );
  AOI211_X1 U7808 ( .C1(n5239), .C2(n6912), .A(n6637), .B(READY_N), .ZN(n6825)
         );
  AND2_X1 U7809 ( .A1(n6826), .A2(n6825), .ZN(n6829) );
  OAI21_X1 U7810 ( .B1(n6829), .B2(n6828), .A(n6827), .ZN(n6834) );
  OAI211_X1 U7811 ( .C1(READY_N), .C2(n6832), .A(n6831), .B(n6830), .ZN(n6833)
         );
  MUX2_X1 U7812 ( .A(REQUESTPENDING_REG_SCAN_IN), .B(n6834), .S(n6833), .Z(
        U3472) );
  INV_X1 U7813 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n6835) );
  AOI22_X1 U7814 ( .A1(n7221), .A2(n7062), .B1(n6835), .B2(n7220), .ZN(U3473)
         );
  XOR2_X1 U7815 ( .A(DATAWIDTH_REG_13__SCAN_IN), .B(keyinput_g117), .Z(n6842)
         );
  AOI22_X1 U7816 ( .A1(ADDRESS_REG_23__SCAN_IN), .A2(keyinput_g77), .B1(
        REIP_REG_22__SCAN_IN), .B2(keyinput_g60), .ZN(n6836) );
  OAI221_X1 U7817 ( .B1(ADDRESS_REG_23__SCAN_IN), .B2(keyinput_g77), .C1(
        REIP_REG_22__SCAN_IN), .C2(keyinput_g60), .A(n6836), .ZN(n6841) );
  AOI22_X1 U7818 ( .A1(ADDRESS_REG_12__SCAN_IN), .A2(keyinput_g88), .B1(
        REIP_REG_26__SCAN_IN), .B2(keyinput_g56), .ZN(n6837) );
  OAI221_X1 U7819 ( .B1(ADDRESS_REG_12__SCAN_IN), .B2(keyinput_g88), .C1(
        REIP_REG_26__SCAN_IN), .C2(keyinput_g56), .A(n6837), .ZN(n6840) );
  AOI22_X1 U7820 ( .A1(REIP_REG_16__SCAN_IN), .A2(keyinput_g66), .B1(
        REIP_REG_20__SCAN_IN), .B2(keyinput_g62), .ZN(n6838) );
  OAI221_X1 U7821 ( .B1(REIP_REG_16__SCAN_IN), .B2(keyinput_g66), .C1(
        REIP_REG_20__SCAN_IN), .C2(keyinput_g62), .A(n6838), .ZN(n6839) );
  NOR4_X1 U7822 ( .A1(n6842), .A2(n6841), .A3(n6840), .A4(n6839), .ZN(n6870)
         );
  AOI22_X1 U7823 ( .A1(BE_N_REG_3__SCAN_IN), .A2(keyinput_g67), .B1(
        DATAWIDTH_REG_21__SCAN_IN), .B2(keyinput_g125), .ZN(n6843) );
  OAI221_X1 U7824 ( .B1(BE_N_REG_3__SCAN_IN), .B2(keyinput_g67), .C1(
        DATAWIDTH_REG_21__SCAN_IN), .C2(keyinput_g125), .A(n6843), .ZN(n6850)
         );
  AOI22_X1 U7825 ( .A1(DATAI_29_), .A2(keyinput_g2), .B1(REIP_REG_27__SCAN_IN), 
        .B2(keyinput_g55), .ZN(n6844) );
  OAI221_X1 U7826 ( .B1(DATAI_29_), .B2(keyinput_g2), .C1(REIP_REG_27__SCAN_IN), .C2(keyinput_g55), .A(n6844), .ZN(n6849) );
  AOI22_X1 U7827 ( .A1(ADDRESS_REG_19__SCAN_IN), .A2(keyinput_g81), .B1(
        STATE_REG_1__SCAN_IN), .B2(keyinput_g102), .ZN(n6845) );
  OAI221_X1 U7828 ( .B1(ADDRESS_REG_19__SCAN_IN), .B2(keyinput_g81), .C1(
        STATE_REG_1__SCAN_IN), .C2(keyinput_g102), .A(n6845), .ZN(n6848) );
  AOI22_X1 U7829 ( .A1(DATAI_16_), .A2(keyinput_g15), .B1(DATAI_31_), .B2(
        keyinput_g0), .ZN(n6846) );
  OAI221_X1 U7830 ( .B1(DATAI_16_), .B2(keyinput_g15), .C1(DATAI_31_), .C2(
        keyinput_g0), .A(n6846), .ZN(n6847) );
  NOR4_X1 U7831 ( .A1(n6850), .A2(n6849), .A3(n6848), .A4(n6847), .ZN(n6869)
         );
  AOI22_X1 U7832 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(keyinput_g123), .B1(
        DATAI_26_), .B2(keyinput_g5), .ZN(n6851) );
  OAI221_X1 U7833 ( .B1(DATAWIDTH_REG_19__SCAN_IN), .B2(keyinput_g123), .C1(
        DATAI_26_), .C2(keyinput_g5), .A(n6851), .ZN(n6858) );
  AOI22_X1 U7834 ( .A1(MORE_REG_SCAN_IN), .A2(keyinput_g44), .B1(DATAI_25_), 
        .B2(keyinput_g6), .ZN(n6852) );
  OAI221_X1 U7835 ( .B1(MORE_REG_SCAN_IN), .B2(keyinput_g44), .C1(DATAI_25_), 
        .C2(keyinput_g6), .A(n6852), .ZN(n6857) );
  AOI22_X1 U7836 ( .A1(DATAI_0_), .A2(keyinput_g31), .B1(REIP_REG_19__SCAN_IN), 
        .B2(keyinput_g63), .ZN(n6853) );
  OAI221_X1 U7837 ( .B1(DATAI_0_), .B2(keyinput_g31), .C1(REIP_REG_19__SCAN_IN), .C2(keyinput_g63), .A(n6853), .ZN(n6856) );
  AOI22_X1 U7838 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(keyinput_g108), .B1(
        CODEFETCH_REG_SCAN_IN), .B2(keyinput_g39), .ZN(n6854) );
  OAI221_X1 U7839 ( .B1(DATAWIDTH_REG_4__SCAN_IN), .B2(keyinput_g108), .C1(
        CODEFETCH_REG_SCAN_IN), .C2(keyinput_g39), .A(n6854), .ZN(n6855) );
  NOR4_X1 U7840 ( .A1(n6858), .A2(n6857), .A3(n6856), .A4(n6855), .ZN(n6868)
         );
  AOI22_X1 U7841 ( .A1(ADDRESS_REG_17__SCAN_IN), .A2(keyinput_g83), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(keyinput_g94), .ZN(n6859) );
  OAI221_X1 U7842 ( .B1(ADDRESS_REG_17__SCAN_IN), .B2(keyinput_g83), .C1(
        ADDRESS_REG_6__SCAN_IN), .C2(keyinput_g94), .A(n6859), .ZN(n6866) );
  AOI22_X1 U7843 ( .A1(ADDRESS_REG_16__SCAN_IN), .A2(keyinput_g84), .B1(
        DATAI_2_), .B2(keyinput_g29), .ZN(n6860) );
  OAI221_X1 U7844 ( .B1(ADDRESS_REG_16__SCAN_IN), .B2(keyinput_g84), .C1(
        DATAI_2_), .C2(keyinput_g29), .A(n6860), .ZN(n6865) );
  AOI22_X1 U7845 ( .A1(FLUSH_REG_SCAN_IN), .A2(keyinput_g45), .B1(DATAI_27_), 
        .B2(keyinput_g4), .ZN(n6861) );
  OAI221_X1 U7846 ( .B1(FLUSH_REG_SCAN_IN), .B2(keyinput_g45), .C1(DATAI_27_), 
        .C2(keyinput_g4), .A(n6861), .ZN(n6864) );
  AOI22_X1 U7847 ( .A1(HOLD), .A2(keyinput_g36), .B1(DATAI_18_), .B2(
        keyinput_g13), .ZN(n6862) );
  OAI221_X1 U7848 ( .B1(HOLD), .B2(keyinput_g36), .C1(DATAI_18_), .C2(
        keyinput_g13), .A(n6862), .ZN(n6863) );
  NOR4_X1 U7849 ( .A1(n6866), .A2(n6865), .A3(n6864), .A4(n6863), .ZN(n6867)
         );
  NAND4_X1 U7850 ( .A1(n6870), .A2(n6869), .A3(n6868), .A4(n6867), .ZN(n7010)
         );
  AOI22_X1 U7851 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(keyinput_g118), .B1(
        DATAWIDTH_REG_15__SCAN_IN), .B2(keyinput_g119), .ZN(n6871) );
  OAI221_X1 U7852 ( .B1(DATAWIDTH_REG_14__SCAN_IN), .B2(keyinput_g118), .C1(
        DATAWIDTH_REG_15__SCAN_IN), .C2(keyinput_g119), .A(n6871), .ZN(n6878)
         );
  AOI22_X1 U7853 ( .A1(BS16_N), .A2(keyinput_g34), .B1(
        DATAWIDTH_REG_22__SCAN_IN), .B2(keyinput_g126), .ZN(n6872) );
  OAI221_X1 U7854 ( .B1(BS16_N), .B2(keyinput_g34), .C1(
        DATAWIDTH_REG_22__SCAN_IN), .C2(keyinput_g126), .A(n6872), .ZN(n6877)
         );
  AOI22_X1 U7855 ( .A1(DATAI_20_), .A2(keyinput_g11), .B1(DATAI_23_), .B2(
        keyinput_g8), .ZN(n6873) );
  OAI221_X1 U7856 ( .B1(DATAI_20_), .B2(keyinput_g11), .C1(DATAI_23_), .C2(
        keyinput_g8), .A(n6873), .ZN(n6876) );
  AOI22_X1 U7857 ( .A1(ADDRESS_REG_25__SCAN_IN), .A2(keyinput_g75), .B1(
        DATAI_14_), .B2(keyinput_g17), .ZN(n6874) );
  OAI221_X1 U7858 ( .B1(ADDRESS_REG_25__SCAN_IN), .B2(keyinput_g75), .C1(
        DATAI_14_), .C2(keyinput_g17), .A(n6874), .ZN(n6875) );
  NOR4_X1 U7859 ( .A1(n6878), .A2(n6877), .A3(n6876), .A4(n6875), .ZN(n6906)
         );
  AOI22_X1 U7860 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(keyinput_g121), .B1(
        DATAI_24_), .B2(keyinput_g7), .ZN(n6879) );
  OAI221_X1 U7861 ( .B1(DATAWIDTH_REG_17__SCAN_IN), .B2(keyinput_g121), .C1(
        DATAI_24_), .C2(keyinput_g7), .A(n6879), .ZN(n6886) );
  AOI22_X1 U7862 ( .A1(READREQUEST_REG_SCAN_IN), .A2(keyinput_g37), .B1(
        DATAI_28_), .B2(keyinput_g3), .ZN(n6880) );
  OAI221_X1 U7863 ( .B1(READREQUEST_REG_SCAN_IN), .B2(keyinput_g37), .C1(
        DATAI_28_), .C2(keyinput_g3), .A(n6880), .ZN(n6885) );
  AOI22_X1 U7864 ( .A1(ADDRESS_REG_14__SCAN_IN), .A2(keyinput_g86), .B1(NA_N), 
        .B2(keyinput_g33), .ZN(n6881) );
  OAI221_X1 U7865 ( .B1(ADDRESS_REG_14__SCAN_IN), .B2(keyinput_g86), .C1(NA_N), 
        .C2(keyinput_g33), .A(n6881), .ZN(n6884) );
  AOI22_X1 U7866 ( .A1(ADDRESS_REG_21__SCAN_IN), .A2(keyinput_g79), .B1(
        DATAWIDTH_REG_0__SCAN_IN), .B2(keyinput_g104), .ZN(n6882) );
  OAI221_X1 U7867 ( .B1(ADDRESS_REG_21__SCAN_IN), .B2(keyinput_g79), .C1(
        DATAWIDTH_REG_0__SCAN_IN), .C2(keyinput_g104), .A(n6882), .ZN(n6883)
         );
  NOR4_X1 U7868 ( .A1(n6886), .A2(n6885), .A3(n6884), .A4(n6883), .ZN(n6905)
         );
  AOI22_X1 U7869 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(keyinput_g127), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(keyinput_g95), .ZN(n6887) );
  OAI221_X1 U7870 ( .B1(DATAWIDTH_REG_23__SCAN_IN), .B2(keyinput_g127), .C1(
        ADDRESS_REG_5__SCAN_IN), .C2(keyinput_g95), .A(n6887), .ZN(n6894) );
  AOI22_X1 U7871 ( .A1(BYTEENABLE_REG_1__SCAN_IN), .A2(keyinput_g48), .B1(
        STATE_REG_0__SCAN_IN), .B2(keyinput_g103), .ZN(n6888) );
  OAI221_X1 U7872 ( .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_g48), .C1(
        STATE_REG_0__SCAN_IN), .C2(keyinput_g103), .A(n6888), .ZN(n6893) );
  AOI22_X1 U7873 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(keyinput_g112), .B1(
        DATAWIDTH_REG_10__SCAN_IN), .B2(keyinput_g114), .ZN(n6889) );
  OAI221_X1 U7874 ( .B1(DATAWIDTH_REG_8__SCAN_IN), .B2(keyinput_g112), .C1(
        DATAWIDTH_REG_10__SCAN_IN), .C2(keyinput_g114), .A(n6889), .ZN(n6892)
         );
  AOI22_X1 U7875 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(keyinput_g109), .B1(
        MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_g32), .ZN(n6890) );
  OAI221_X1 U7876 ( .B1(DATAWIDTH_REG_5__SCAN_IN), .B2(keyinput_g109), .C1(
        MEMORYFETCH_REG_SCAN_IN), .C2(keyinput_g32), .A(n6890), .ZN(n6891) );
  NOR4_X1 U7877 ( .A1(n6894), .A2(n6893), .A3(n6892), .A4(n6891), .ZN(n6904)
         );
  AOI22_X1 U7878 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(keyinput_g122), .B1(
        DATAI_19_), .B2(keyinput_g12), .ZN(n6895) );
  OAI221_X1 U7879 ( .B1(DATAWIDTH_REG_18__SCAN_IN), .B2(keyinput_g122), .C1(
        DATAI_19_), .C2(keyinput_g12), .A(n6895), .ZN(n6902) );
  AOI22_X1 U7880 ( .A1(ADDRESS_REG_15__SCAN_IN), .A2(keyinput_g85), .B1(
        DATAI_1_), .B2(keyinput_g30), .ZN(n6896) );
  OAI221_X1 U7881 ( .B1(ADDRESS_REG_15__SCAN_IN), .B2(keyinput_g85), .C1(
        DATAI_1_), .C2(keyinput_g30), .A(n6896), .ZN(n6901) );
  AOI22_X1 U7882 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(keyinput_g50), .B1(
        M_IO_N_REG_SCAN_IN), .B2(keyinput_g40), .ZN(n6897) );
  OAI221_X1 U7883 ( .B1(BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_g50), .C1(
        M_IO_N_REG_SCAN_IN), .C2(keyinput_g40), .A(n6897), .ZN(n6900) );
  AOI22_X1 U7884 ( .A1(ADDRESS_REG_10__SCAN_IN), .A2(keyinput_g90), .B1(
        REIP_REG_28__SCAN_IN), .B2(keyinput_g54), .ZN(n6898) );
  OAI221_X1 U7885 ( .B1(ADDRESS_REG_10__SCAN_IN), .B2(keyinput_g90), .C1(
        REIP_REG_28__SCAN_IN), .C2(keyinput_g54), .A(n6898), .ZN(n6899) );
  NOR4_X1 U7886 ( .A1(n6902), .A2(n6901), .A3(n6900), .A4(n6899), .ZN(n6903)
         );
  NAND4_X1 U7887 ( .A1(n6906), .A2(n6905), .A3(n6904), .A4(n6903), .ZN(n7009)
         );
  AOI22_X1 U7888 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(keyinput_g113), .B1(
        DATAWIDTH_REG_12__SCAN_IN), .B2(keyinput_g116), .ZN(n6907) );
  OAI221_X1 U7889 ( .B1(DATAWIDTH_REG_9__SCAN_IN), .B2(keyinput_g113), .C1(
        DATAWIDTH_REG_12__SCAN_IN), .C2(keyinput_g116), .A(n6907), .ZN(n6916)
         );
  AOI22_X1 U7890 ( .A1(n6909), .A2(keyinput_g53), .B1(keyinput_g72), .B2(n7182), .ZN(n6908) );
  OAI221_X1 U7891 ( .B1(n6909), .B2(keyinput_g53), .C1(n7182), .C2(
        keyinput_g72), .A(n6908), .ZN(n6915) );
  AOI22_X1 U7892 ( .A1(n7016), .A2(keyinput_g58), .B1(keyinput_g42), .B2(n7154), .ZN(n6910) );
  OAI221_X1 U7893 ( .B1(n7016), .B2(keyinput_g58), .C1(n7154), .C2(
        keyinput_g42), .A(n6910), .ZN(n6914) );
  AOI22_X1 U7894 ( .A1(n7186), .A2(keyinput_g19), .B1(n6912), .B2(keyinput_g43), .ZN(n6911) );
  OAI221_X1 U7895 ( .B1(n7186), .B2(keyinput_g19), .C1(n6912), .C2(
        keyinput_g43), .A(n6911), .ZN(n6913) );
  NOR4_X1 U7896 ( .A1(n6916), .A2(n6915), .A3(n6914), .A4(n6913), .ZN(n6953)
         );
  AOI22_X1 U7897 ( .A1(n6918), .A2(keyinput_g51), .B1(keyinput_g74), .B2(n7038), .ZN(n6917) );
  OAI221_X1 U7898 ( .B1(n6918), .B2(keyinput_g51), .C1(n7038), .C2(
        keyinput_g74), .A(n6917), .ZN(n6927) );
  AOI22_X1 U7899 ( .A1(n7040), .A2(keyinput_g20), .B1(n7164), .B2(keyinput_g57), .ZN(n6919) );
  OAI221_X1 U7900 ( .B1(n7040), .B2(keyinput_g20), .C1(n7164), .C2(
        keyinput_g57), .A(n6919), .ZN(n6926) );
  AOI22_X1 U7901 ( .A1(n7054), .A2(keyinput_g100), .B1(n6921), .B2(
        keyinput_g21), .ZN(n6920) );
  OAI221_X1 U7902 ( .B1(n7054), .B2(keyinput_g100), .C1(n6921), .C2(
        keyinput_g21), .A(n6920), .ZN(n6925) );
  AOI22_X1 U7903 ( .A1(n6923), .A2(keyinput_g97), .B1(keyinput_g91), .B2(n7183), .ZN(n6922) );
  OAI221_X1 U7904 ( .B1(n6923), .B2(keyinput_g97), .C1(n7183), .C2(
        keyinput_g91), .A(n6922), .ZN(n6924) );
  NOR4_X1 U7905 ( .A1(n6927), .A2(n6926), .A3(n6925), .A4(n6924), .ZN(n6952)
         );
  AOI22_X1 U7906 ( .A1(n7028), .A2(keyinput_g16), .B1(keyinput_g89), .B2(n7148), .ZN(n6928) );
  OAI221_X1 U7907 ( .B1(n7028), .B2(keyinput_g16), .C1(n7148), .C2(
        keyinput_g89), .A(n6928), .ZN(n6939) );
  AOI22_X1 U7908 ( .A1(n6931), .A2(keyinput_g106), .B1(n6930), .B2(
        keyinput_g52), .ZN(n6929) );
  OAI221_X1 U7909 ( .B1(n6931), .B2(keyinput_g106), .C1(n6930), .C2(
        keyinput_g52), .A(n6929), .ZN(n6938) );
  AOI22_X1 U7910 ( .A1(n6934), .A2(keyinput_g28), .B1(keyinput_g80), .B2(n6933), .ZN(n6932) );
  OAI221_X1 U7911 ( .B1(n6934), .B2(keyinput_g28), .C1(n6933), .C2(
        keyinput_g80), .A(n6932), .ZN(n6937) );
  AOI22_X1 U7912 ( .A1(n7198), .A2(keyinput_g14), .B1(keyinput_g92), .B2(n7018), .ZN(n6935) );
  OAI221_X1 U7913 ( .B1(n7198), .B2(keyinput_g14), .C1(n7018), .C2(
        keyinput_g92), .A(n6935), .ZN(n6936) );
  NOR4_X1 U7914 ( .A1(n6939), .A2(n6938), .A3(n6937), .A4(n6936), .ZN(n6951)
         );
  AOI22_X1 U7915 ( .A1(n7163), .A2(keyinput_g107), .B1(n7060), .B2(
        keyinput_g59), .ZN(n6940) );
  OAI221_X1 U7916 ( .B1(n7163), .B2(keyinput_g107), .C1(n7060), .C2(
        keyinput_g59), .A(n6940), .ZN(n6949) );
  AOI22_X1 U7917 ( .A1(n7026), .A2(keyinput_g61), .B1(keyinput_g115), .B2(
        n6942), .ZN(n6941) );
  OAI221_X1 U7918 ( .B1(n7026), .B2(keyinput_g61), .C1(n6942), .C2(
        keyinput_g115), .A(n6941), .ZN(n6948) );
  AOI22_X1 U7919 ( .A1(n7151), .A2(keyinput_g10), .B1(keyinput_g46), .B2(n7195), .ZN(n6943) );
  OAI221_X1 U7920 ( .B1(n7151), .B2(keyinput_g10), .C1(n7195), .C2(
        keyinput_g46), .A(n6943), .ZN(n6947) );
  AOI22_X1 U7921 ( .A1(n6945), .A2(keyinput_g124), .B1(n7153), .B2(keyinput_g9), .ZN(n6944) );
  OAI221_X1 U7922 ( .B1(n6945), .B2(keyinput_g124), .C1(n7153), .C2(
        keyinput_g9), .A(n6944), .ZN(n6946) );
  NOR4_X1 U7923 ( .A1(n6949), .A2(n6948), .A3(n6947), .A4(n6946), .ZN(n6950)
         );
  NAND4_X1 U7924 ( .A1(n6953), .A2(n6952), .A3(n6951), .A4(n6950), .ZN(n7008)
         );
  AOI22_X1 U7925 ( .A1(n7025), .A2(keyinput_g49), .B1(n6955), .B2(keyinput_g41), .ZN(n6954) );
  OAI221_X1 U7926 ( .B1(n7025), .B2(keyinput_g49), .C1(n6955), .C2(
        keyinput_g41), .A(n6954), .ZN(n6963) );
  AOI22_X1 U7927 ( .A1(n4099), .A2(keyinput_g1), .B1(keyinput_g99), .B2(n7169), 
        .ZN(n6956) );
  OAI221_X1 U7928 ( .B1(n4099), .B2(keyinput_g1), .C1(n7169), .C2(keyinput_g99), .A(n6956), .ZN(n6962) );
  AOI22_X1 U7929 ( .A1(n7019), .A2(keyinput_g68), .B1(n7199), .B2(keyinput_g35), .ZN(n6957) );
  OAI221_X1 U7930 ( .B1(n7019), .B2(keyinput_g68), .C1(n7199), .C2(
        keyinput_g35), .A(n6957), .ZN(n6961) );
  AOI22_X1 U7931 ( .A1(n6959), .A2(keyinput_g101), .B1(keyinput_g111), .B2(
        n7135), .ZN(n6958) );
  OAI221_X1 U7932 ( .B1(n6959), .B2(keyinput_g101), .C1(n7135), .C2(
        keyinput_g111), .A(n6958), .ZN(n6960) );
  NOR4_X1 U7933 ( .A1(n6963), .A2(n6962), .A3(n6961), .A4(n6960), .ZN(n7006)
         );
  AOI22_X1 U7934 ( .A1(n7167), .A2(keyinput_g76), .B1(n7161), .B2(keyinput_g26), .ZN(n6964) );
  OAI221_X1 U7935 ( .B1(n7167), .B2(keyinput_g76), .C1(n7161), .C2(
        keyinput_g26), .A(n6964), .ZN(n6976) );
  AOI22_X1 U7936 ( .A1(n6967), .A2(keyinput_g64), .B1(keyinput_g38), .B2(n6966), .ZN(n6965) );
  OAI221_X1 U7937 ( .B1(n6967), .B2(keyinput_g64), .C1(n6966), .C2(
        keyinput_g38), .A(n6965), .ZN(n6975) );
  AOI22_X1 U7938 ( .A1(n6970), .A2(keyinput_g93), .B1(keyinput_g87), .B2(n6969), .ZN(n6968) );
  OAI221_X1 U7939 ( .B1(n6970), .B2(keyinput_g93), .C1(n6969), .C2(
        keyinput_g87), .A(n6968), .ZN(n6974) );
  AOI22_X1 U7940 ( .A1(n6972), .A2(keyinput_g27), .B1(keyinput_g73), .B2(n7031), .ZN(n6971) );
  OAI221_X1 U7941 ( .B1(n6972), .B2(keyinput_g27), .C1(n7031), .C2(
        keyinput_g73), .A(n6971), .ZN(n6973) );
  NOR4_X1 U7942 ( .A1(n6976), .A2(n6975), .A3(n6974), .A4(n6973), .ZN(n7005)
         );
  AOI22_X1 U7943 ( .A1(n7063), .A2(keyinput_g96), .B1(keyinput_g110), .B2(
        n7177), .ZN(n6977) );
  OAI221_X1 U7944 ( .B1(n7063), .B2(keyinput_g96), .C1(n7177), .C2(
        keyinput_g110), .A(n6977), .ZN(n6988) );
  AOI22_X1 U7945 ( .A1(n7196), .A2(keyinput_g23), .B1(keyinput_g105), .B2(
        n6979), .ZN(n6978) );
  OAI221_X1 U7946 ( .B1(n7196), .B2(keyinput_g23), .C1(n6979), .C2(
        keyinput_g105), .A(n6978), .ZN(n6987) );
  AOI22_X1 U7947 ( .A1(n7166), .A2(keyinput_g98), .B1(n6981), .B2(keyinput_g82), .ZN(n6980) );
  OAI221_X1 U7948 ( .B1(n7166), .B2(keyinput_g98), .C1(n6981), .C2(
        keyinput_g82), .A(n6980), .ZN(n6986) );
  AOI22_X1 U7949 ( .A1(n6984), .A2(keyinput_g78), .B1(n6983), .B2(keyinput_g65), .ZN(n6982) );
  OAI221_X1 U7950 ( .B1(n6984), .B2(keyinput_g78), .C1(n6983), .C2(
        keyinput_g65), .A(n6982), .ZN(n6985) );
  NOR4_X1 U7951 ( .A1(n6988), .A2(n6987), .A3(n6986), .A4(n6985), .ZN(n7004)
         );
  AOI22_X1 U7952 ( .A1(n6991), .A2(keyinput_g24), .B1(keyinput_g47), .B2(n6990), .ZN(n6989) );
  OAI221_X1 U7953 ( .B1(n6991), .B2(keyinput_g24), .C1(n6990), .C2(
        keyinput_g47), .A(n6989), .ZN(n7002) );
  AOI22_X1 U7954 ( .A1(n7176), .A2(keyinput_g71), .B1(n6993), .B2(keyinput_g18), .ZN(n6992) );
  OAI221_X1 U7955 ( .B1(n7176), .B2(keyinput_g71), .C1(n6993), .C2(
        keyinput_g18), .A(n6992), .ZN(n7001) );
  AOI22_X1 U7956 ( .A1(n7041), .A2(keyinput_g70), .B1(n6995), .B2(keyinput_g25), .ZN(n6994) );
  OAI221_X1 U7957 ( .B1(n7041), .B2(keyinput_g70), .C1(n6995), .C2(
        keyinput_g25), .A(n6994), .ZN(n7000) );
  AOI22_X1 U7958 ( .A1(n6998), .A2(keyinput_g120), .B1(keyinput_g69), .B2(
        n6997), .ZN(n6996) );
  OAI221_X1 U7959 ( .B1(n6998), .B2(keyinput_g120), .C1(n6997), .C2(
        keyinput_g69), .A(n6996), .ZN(n6999) );
  NOR4_X1 U7960 ( .A1(n7002), .A2(n7001), .A3(n7000), .A4(n6999), .ZN(n7003)
         );
  NAND4_X1 U7961 ( .A1(n7006), .A2(n7005), .A3(n7004), .A4(n7003), .ZN(n7007)
         );
  NOR4_X1 U7962 ( .A1(n7010), .A2(n7009), .A3(n7008), .A4(n7007), .ZN(n7219)
         );
  AOI22_X1 U7963 ( .A1(n7013), .A2(keyinput_f81), .B1(n7012), .B2(keyinput_f55), .ZN(n7011) );
  OAI221_X1 U7964 ( .B1(n7013), .B2(keyinput_f81), .C1(n7012), .C2(
        keyinput_f55), .A(n7011), .ZN(n7215) );
  OAI22_X1 U7965 ( .A1(n7016), .A2(keyinput_f58), .B1(n7015), .B2(keyinput_f77), .ZN(n7014) );
  AOI221_X1 U7966 ( .B1(n7016), .B2(keyinput_f58), .C1(keyinput_f77), .C2(
        n7015), .A(n7014), .ZN(n7023) );
  OAI22_X1 U7967 ( .A1(n7019), .A2(keyinput_f68), .B1(n7018), .B2(keyinput_f92), .ZN(n7017) );
  AOI221_X1 U7968 ( .B1(n7019), .B2(keyinput_f68), .C1(keyinput_f92), .C2(
        n7018), .A(n7017), .ZN(n7022) );
  XNOR2_X1 U7969 ( .A(keyinput_f113), .B(DATAWIDTH_REG_9__SCAN_IN), .ZN(n7021)
         );
  XNOR2_X1 U7970 ( .A(keyinput_f124), .B(DATAWIDTH_REG_20__SCAN_IN), .ZN(n7020) );
  NAND4_X1 U7971 ( .A1(n7023), .A2(n7022), .A3(n7021), .A4(n7020), .ZN(n7214)
         );
  OAI22_X1 U7972 ( .A1(n7026), .A2(keyinput_f61), .B1(n7025), .B2(keyinput_f49), .ZN(n7024) );
  AOI221_X1 U7973 ( .B1(n7026), .B2(keyinput_f61), .C1(keyinput_f49), .C2(
        n7025), .A(n7024), .ZN(n7071) );
  XOR2_X1 U7974 ( .A(ADDRESS_REG_3__SCAN_IN), .B(keyinput_f97), .Z(n7035) );
  XOR2_X1 U7975 ( .A(keyinput_f112), .B(DATAWIDTH_REG_8__SCAN_IN), .Z(n7034)
         );
  AOI22_X1 U7976 ( .A1(n7029), .A2(keyinput_f44), .B1(n7028), .B2(keyinput_f16), .ZN(n7027) );
  OAI221_X1 U7977 ( .B1(n7029), .B2(keyinput_f44), .C1(n7028), .C2(
        keyinput_f16), .A(n7027), .ZN(n7033) );
  AOI22_X1 U7978 ( .A1(n7031), .A2(keyinput_f73), .B1(n4077), .B2(keyinput_f4), 
        .ZN(n7030) );
  OAI221_X1 U7979 ( .B1(n7031), .B2(keyinput_f73), .C1(n4077), .C2(keyinput_f4), .A(n7030), .ZN(n7032) );
  NOR4_X1 U7980 ( .A1(n7035), .A2(n7034), .A3(n7033), .A4(n7032), .ZN(n7070)
         );
  INV_X1 U7981 ( .A(DATAI_26_), .ZN(n7037) );
  AOI22_X1 U7982 ( .A1(n7038), .A2(keyinput_f74), .B1(n7037), .B2(keyinput_f5), 
        .ZN(n7036) );
  OAI221_X1 U7983 ( .B1(n7038), .B2(keyinput_f74), .C1(n7037), .C2(keyinput_f5), .A(n7036), .ZN(n7051) );
  AOI22_X1 U7984 ( .A1(n7041), .A2(keyinput_f70), .B1(n7040), .B2(keyinput_f20), .ZN(n7039) );
  OAI221_X1 U7985 ( .B1(n7041), .B2(keyinput_f70), .C1(n7040), .C2(
        keyinput_f20), .A(n7039), .ZN(n7050) );
  AOI22_X1 U7986 ( .A1(n7044), .A2(keyinput_f15), .B1(n7043), .B2(keyinput_f63), .ZN(n7042) );
  OAI221_X1 U7987 ( .B1(n7044), .B2(keyinput_f15), .C1(n7043), .C2(
        keyinput_f63), .A(n7042), .ZN(n7049) );
  AOI22_X1 U7988 ( .A1(n7047), .A2(keyinput_f12), .B1(keyinput_f90), .B2(n7046), .ZN(n7045) );
  OAI221_X1 U7989 ( .B1(n7047), .B2(keyinput_f12), .C1(n7046), .C2(
        keyinput_f90), .A(n7045), .ZN(n7048) );
  NOR4_X1 U7990 ( .A1(n7051), .A2(n7050), .A3(n7049), .A4(n7048), .ZN(n7069)
         );
  AOI22_X1 U7991 ( .A1(n7054), .A2(keyinput_f100), .B1(n7053), .B2(
        keyinput_f56), .ZN(n7052) );
  OAI221_X1 U7992 ( .B1(n7054), .B2(keyinput_f100), .C1(n7053), .C2(
        keyinput_f56), .A(n7052), .ZN(n7067) );
  INV_X1 U7993 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n7057) );
  INV_X1 U7994 ( .A(keyinput_f105), .ZN(n7056) );
  AOI22_X1 U7995 ( .A1(n7057), .A2(keyinput_f37), .B1(DATAWIDTH_REG_1__SCAN_IN), .B2(n7056), .ZN(n7055) );
  OAI221_X1 U7996 ( .B1(n7057), .B2(keyinput_f37), .C1(n7056), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(n7055), .ZN(n7066) );
  AOI22_X1 U7997 ( .A1(n7060), .A2(keyinput_f59), .B1(keyinput_f11), .B2(n7059), .ZN(n7058) );
  OAI221_X1 U7998 ( .B1(n7060), .B2(keyinput_f59), .C1(n7059), .C2(
        keyinput_f11), .A(n7058), .ZN(n7065) );
  AOI22_X1 U7999 ( .A1(n7063), .A2(keyinput_f96), .B1(n7062), .B2(keyinput_f32), .ZN(n7061) );
  OAI221_X1 U8000 ( .B1(n7063), .B2(keyinput_f96), .C1(n7062), .C2(
        keyinput_f32), .A(n7061), .ZN(n7064) );
  NOR4_X1 U8001 ( .A1(n7067), .A2(n7066), .A3(n7065), .A4(n7064), .ZN(n7068)
         );
  NAND4_X1 U8002 ( .A1(n7071), .A2(n7070), .A3(n7069), .A4(n7068), .ZN(n7213)
         );
  OAI22_X1 U8003 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(keyinput_f39), .B1(
        keyinput_f94), .B2(ADDRESS_REG_6__SCAN_IN), .ZN(n7072) );
  AOI221_X1 U8004 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(keyinput_f39), .C1(
        ADDRESS_REG_6__SCAN_IN), .C2(keyinput_f94), .A(n7072), .ZN(n7078) );
  OAI22_X1 U8005 ( .A1(DATAI_31_), .A2(keyinput_f0), .B1(DATAI_29_), .B2(
        keyinput_f2), .ZN(n7073) );
  AOI221_X1 U8006 ( .B1(DATAI_31_), .B2(keyinput_f0), .C1(keyinput_f2), .C2(
        DATAI_29_), .A(n7073), .ZN(n7077) );
  OAI22_X1 U8007 ( .A1(REIP_REG_17__SCAN_IN), .A2(keyinput_f65), .B1(
        keyinput_f83), .B2(ADDRESS_REG_17__SCAN_IN), .ZN(n7074) );
  AOI221_X1 U8008 ( .B1(REIP_REG_17__SCAN_IN), .B2(keyinput_f65), .C1(
        ADDRESS_REG_17__SCAN_IN), .C2(keyinput_f83), .A(n7074), .ZN(n7076) );
  XNOR2_X1 U8009 ( .A(keyinput_f125), .B(DATAWIDTH_REG_21__SCAN_IN), .ZN(n7075) );
  NAND4_X1 U8010 ( .A1(n7078), .A2(n7077), .A3(n7076), .A4(n7075), .ZN(n7106)
         );
  OAI22_X1 U8011 ( .A1(keyinput_f115), .A2(DATAWIDTH_REG_11__SCAN_IN), .B1(
        keyinput_f95), .B2(ADDRESS_REG_5__SCAN_IN), .ZN(n7079) );
  AOI221_X1 U8012 ( .B1(keyinput_f115), .B2(DATAWIDTH_REG_11__SCAN_IN), .C1(
        ADDRESS_REG_5__SCAN_IN), .C2(keyinput_f95), .A(n7079), .ZN(n7086) );
  OAI22_X1 U8013 ( .A1(REIP_REG_16__SCAN_IN), .A2(keyinput_f66), .B1(
        keyinput_f27), .B2(DATAI_4_), .ZN(n7080) );
  AOI221_X1 U8014 ( .B1(REIP_REG_16__SCAN_IN), .B2(keyinput_f66), .C1(DATAI_4_), .C2(keyinput_f27), .A(n7080), .ZN(n7085) );
  OAI22_X1 U8015 ( .A1(REIP_REG_29__SCAN_IN), .A2(keyinput_f53), .B1(
        keyinput_f45), .B2(FLUSH_REG_SCAN_IN), .ZN(n7081) );
  AOI221_X1 U8016 ( .B1(REIP_REG_29__SCAN_IN), .B2(keyinput_f53), .C1(
        FLUSH_REG_SCAN_IN), .C2(keyinput_f45), .A(n7081), .ZN(n7084) );
  OAI22_X1 U8017 ( .A1(DATAI_24_), .A2(keyinput_f7), .B1(
        DATAWIDTH_REG_16__SCAN_IN), .B2(keyinput_f120), .ZN(n7082) );
  AOI221_X1 U8018 ( .B1(DATAI_24_), .B2(keyinput_f7), .C1(keyinput_f120), .C2(
        DATAWIDTH_REG_16__SCAN_IN), .A(n7082), .ZN(n7083) );
  NAND4_X1 U8019 ( .A1(n7086), .A2(n7085), .A3(n7084), .A4(n7083), .ZN(n7105)
         );
  OAI22_X1 U8020 ( .A1(DATAI_14_), .A2(keyinput_f17), .B1(keyinput_f80), .B2(
        ADDRESS_REG_20__SCAN_IN), .ZN(n7087) );
  AOI221_X1 U8021 ( .B1(DATAI_14_), .B2(keyinput_f17), .C1(
        ADDRESS_REG_20__SCAN_IN), .C2(keyinput_f80), .A(n7087), .ZN(n7094) );
  OAI22_X1 U8022 ( .A1(REIP_REG_22__SCAN_IN), .A2(keyinput_f60), .B1(
        DATAWIDTH_REG_4__SCAN_IN), .B2(keyinput_f108), .ZN(n7088) );
  AOI221_X1 U8023 ( .B1(REIP_REG_22__SCAN_IN), .B2(keyinput_f60), .C1(
        keyinput_f108), .C2(DATAWIDTH_REG_4__SCAN_IN), .A(n7088), .ZN(n7093)
         );
  OAI22_X1 U8024 ( .A1(DATAI_3_), .A2(keyinput_f28), .B1(
        DATAWIDTH_REG_0__SCAN_IN), .B2(keyinput_f104), .ZN(n7089) );
  AOI221_X1 U8025 ( .B1(DATAI_3_), .B2(keyinput_f28), .C1(keyinput_f104), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(n7089), .ZN(n7092) );
  OAI22_X1 U8026 ( .A1(DATAI_6_), .A2(keyinput_f25), .B1(keyinput_f47), .B2(
        BYTEENABLE_REG_0__SCAN_IN), .ZN(n7090) );
  AOI221_X1 U8027 ( .B1(DATAI_6_), .B2(keyinput_f25), .C1(
        BYTEENABLE_REG_0__SCAN_IN), .C2(keyinput_f47), .A(n7090), .ZN(n7091)
         );
  NAND4_X1 U8028 ( .A1(n7094), .A2(n7093), .A3(n7092), .A4(n7091), .ZN(n7104)
         );
  OAI22_X1 U8029 ( .A1(DATAI_10_), .A2(keyinput_f21), .B1(
        DATAWIDTH_REG_5__SCAN_IN), .B2(keyinput_f109), .ZN(n7095) );
  AOI221_X1 U8030 ( .B1(DATAI_10_), .B2(keyinput_f21), .C1(keyinput_f109), 
        .C2(DATAWIDTH_REG_5__SCAN_IN), .A(n7095), .ZN(n7102) );
  OAI22_X1 U8031 ( .A1(keyinput_f116), .A2(DATAWIDTH_REG_12__SCAN_IN), .B1(
        keyinput_f40), .B2(M_IO_N_REG_SCAN_IN), .ZN(n7096) );
  AOI221_X1 U8032 ( .B1(keyinput_f116), .B2(DATAWIDTH_REG_12__SCAN_IN), .C1(
        M_IO_N_REG_SCAN_IN), .C2(keyinput_f40), .A(n7096), .ZN(n7101) );
  OAI22_X1 U8033 ( .A1(REIP_REG_30__SCAN_IN), .A2(keyinput_f52), .B1(
        BE_N_REG_3__SCAN_IN), .B2(keyinput_f67), .ZN(n7097) );
  AOI221_X1 U8034 ( .B1(REIP_REG_30__SCAN_IN), .B2(keyinput_f52), .C1(
        keyinput_f67), .C2(BE_N_REG_3__SCAN_IN), .A(n7097), .ZN(n7100) );
  OAI22_X1 U8035 ( .A1(STATE_REG_1__SCAN_IN), .A2(keyinput_f102), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(keyinput_f88), .ZN(n7098) );
  AOI221_X1 U8036 ( .B1(STATE_REG_1__SCAN_IN), .B2(keyinput_f102), .C1(
        keyinput_f88), .C2(ADDRESS_REG_12__SCAN_IN), .A(n7098), .ZN(n7099) );
  NAND4_X1 U8037 ( .A1(n7102), .A2(n7101), .A3(n7100), .A4(n7099), .ZN(n7103)
         );
  NOR4_X1 U8038 ( .A1(n7106), .A2(n7105), .A3(n7104), .A4(n7103), .ZN(n7211)
         );
  OAI22_X1 U8039 ( .A1(DATAI_25_), .A2(keyinput_f6), .B1(keyinput_f69), .B2(
        BE_N_REG_1__SCAN_IN), .ZN(n7107) );
  AOI221_X1 U8040 ( .B1(DATAI_25_), .B2(keyinput_f6), .C1(BE_N_REG_1__SCAN_IN), 
        .C2(keyinput_f69), .A(n7107), .ZN(n7114) );
  OAI22_X1 U8041 ( .A1(keyinput_f123), .A2(DATAWIDTH_REG_19__SCAN_IN), .B1(
        keyinput_f78), .B2(ADDRESS_REG_22__SCAN_IN), .ZN(n7108) );
  AOI221_X1 U8042 ( .B1(keyinput_f123), .B2(DATAWIDTH_REG_19__SCAN_IN), .C1(
        ADDRESS_REG_22__SCAN_IN), .C2(keyinput_f78), .A(n7108), .ZN(n7113) );
  OAI22_X1 U8043 ( .A1(STATEBS16_REG_SCAN_IN), .A2(keyinput_f43), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(keyinput_f82), .ZN(n7109) );
  AOI221_X1 U8044 ( .B1(STATEBS16_REG_SCAN_IN), .B2(keyinput_f43), .C1(
        keyinput_f82), .C2(ADDRESS_REG_18__SCAN_IN), .A(n7109), .ZN(n7112) );
  OAI22_X1 U8045 ( .A1(D_C_N_REG_SCAN_IN), .A2(keyinput_f41), .B1(
        keyinput_f126), .B2(DATAWIDTH_REG_22__SCAN_IN), .ZN(n7110) );
  AOI221_X1 U8046 ( .B1(D_C_N_REG_SCAN_IN), .B2(keyinput_f41), .C1(
        DATAWIDTH_REG_22__SCAN_IN), .C2(keyinput_f126), .A(n7110), .ZN(n7111)
         );
  NAND4_X1 U8047 ( .A1(n7114), .A2(n7113), .A3(n7112), .A4(n7111), .ZN(n7143)
         );
  OAI22_X1 U8048 ( .A1(keyinput_f75), .A2(ADDRESS_REG_25__SCAN_IN), .B1(
        keyinput_f38), .B2(ADS_N_REG_SCAN_IN), .ZN(n7115) );
  AOI221_X1 U8049 ( .B1(keyinput_f75), .B2(ADDRESS_REG_25__SCAN_IN), .C1(
        ADS_N_REG_SCAN_IN), .C2(keyinput_f38), .A(n7115), .ZN(n7122) );
  OAI22_X1 U8050 ( .A1(STATE_REG_0__SCAN_IN), .A2(keyinput_f103), .B1(
        DATAWIDTH_REG_23__SCAN_IN), .B2(keyinput_f127), .ZN(n7116) );
  AOI221_X1 U8051 ( .B1(STATE_REG_0__SCAN_IN), .B2(keyinput_f103), .C1(
        keyinput_f127), .C2(DATAWIDTH_REG_23__SCAN_IN), .A(n7116), .ZN(n7121)
         );
  OAI22_X1 U8052 ( .A1(REIP_REG_28__SCAN_IN), .A2(keyinput_f54), .B1(
        keyinput_f13), .B2(DATAI_18_), .ZN(n7117) );
  AOI221_X1 U8053 ( .B1(REIP_REG_28__SCAN_IN), .B2(keyinput_f54), .C1(
        DATAI_18_), .C2(keyinput_f13), .A(n7117), .ZN(n7120) );
  OAI22_X1 U8054 ( .A1(keyinput_f114), .A2(DATAWIDTH_REG_10__SCAN_IN), .B1(
        keyinput_f36), .B2(HOLD), .ZN(n7118) );
  AOI221_X1 U8055 ( .B1(keyinput_f114), .B2(DATAWIDTH_REG_10__SCAN_IN), .C1(
        HOLD), .C2(keyinput_f36), .A(n7118), .ZN(n7119) );
  NAND4_X1 U8056 ( .A1(n7122), .A2(n7121), .A3(n7120), .A4(n7119), .ZN(n7142)
         );
  OAI22_X1 U8057 ( .A1(keyinput_f119), .A2(DATAWIDTH_REG_15__SCAN_IN), .B1(
        keyinput_f118), .B2(DATAWIDTH_REG_14__SCAN_IN), .ZN(n7123) );
  AOI221_X1 U8058 ( .B1(keyinput_f119), .B2(DATAWIDTH_REG_15__SCAN_IN), .C1(
        DATAWIDTH_REG_14__SCAN_IN), .C2(keyinput_f118), .A(n7123), .ZN(n7130)
         );
  OAI22_X1 U8059 ( .A1(REIP_REG_20__SCAN_IN), .A2(keyinput_f62), .B1(
        DATAWIDTH_REG_18__SCAN_IN), .B2(keyinput_f122), .ZN(n7124) );
  AOI221_X1 U8060 ( .B1(REIP_REG_20__SCAN_IN), .B2(keyinput_f62), .C1(
        keyinput_f122), .C2(DATAWIDTH_REG_18__SCAN_IN), .A(n7124), .ZN(n7129)
         );
  OAI22_X1 U8061 ( .A1(REIP_REG_18__SCAN_IN), .A2(keyinput_f64), .B1(
        keyinput_f24), .B2(DATAI_7_), .ZN(n7125) );
  AOI221_X1 U8062 ( .B1(REIP_REG_18__SCAN_IN), .B2(keyinput_f64), .C1(DATAI_7_), .C2(keyinput_f24), .A(n7125), .ZN(n7128) );
  OAI22_X1 U8063 ( .A1(REIP_REG_31__SCAN_IN), .A2(keyinput_f51), .B1(
        keyinput_f93), .B2(ADDRESS_REG_7__SCAN_IN), .ZN(n7126) );
  AOI221_X1 U8064 ( .B1(REIP_REG_31__SCAN_IN), .B2(keyinput_f51), .C1(
        ADDRESS_REG_7__SCAN_IN), .C2(keyinput_f93), .A(n7126), .ZN(n7127) );
  NAND4_X1 U8065 ( .A1(n7130), .A2(n7129), .A3(n7128), .A4(n7127), .ZN(n7141)
         );
  OAI22_X1 U8066 ( .A1(DATAI_0_), .A2(keyinput_f31), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(keyinput_f84), .ZN(n7131) );
  AOI221_X1 U8067 ( .B1(DATAI_0_), .B2(keyinput_f31), .C1(keyinput_f84), .C2(
        ADDRESS_REG_16__SCAN_IN), .A(n7131), .ZN(n7139) );
  OAI22_X1 U8068 ( .A1(keyinput_f87), .A2(ADDRESS_REG_13__SCAN_IN), .B1(
        keyinput_f117), .B2(DATAWIDTH_REG_13__SCAN_IN), .ZN(n7132) );
  AOI221_X1 U8069 ( .B1(keyinput_f87), .B2(ADDRESS_REG_13__SCAN_IN), .C1(
        DATAWIDTH_REG_13__SCAN_IN), .C2(keyinput_f117), .A(n7132), .ZN(n7138)
         );
  OAI22_X1 U8070 ( .A1(DATAI_30_), .A2(keyinput_f1), .B1(keyinput_f18), .B2(
        DATAI_13_), .ZN(n7133) );
  AOI221_X1 U8071 ( .B1(DATAI_30_), .B2(keyinput_f1), .C1(DATAI_13_), .C2(
        keyinput_f18), .A(n7133), .ZN(n7137) );
  OAI22_X1 U8072 ( .A1(keyinput_f111), .A2(n7135), .B1(STATE_REG_2__SCAN_IN), 
        .B2(keyinput_f101), .ZN(n7134) );
  AOI221_X1 U8073 ( .B1(n7135), .B2(keyinput_f111), .C1(STATE_REG_2__SCAN_IN), 
        .C2(keyinput_f101), .A(n7134), .ZN(n7136) );
  NAND4_X1 U8074 ( .A1(n7139), .A2(n7138), .A3(n7137), .A4(n7136), .ZN(n7140)
         );
  NOR4_X1 U8075 ( .A1(n7143), .A2(n7142), .A3(n7141), .A4(n7140), .ZN(n7210)
         );
  AOI22_X1 U8076 ( .A1(n7145), .A2(keyinput_f29), .B1(n4090), .B2(keyinput_f3), 
        .ZN(n7144) );
  OAI221_X1 U8077 ( .B1(n7145), .B2(keyinput_f29), .C1(n4090), .C2(keyinput_f3), .A(n7144), .ZN(n7158) );
  AOI22_X1 U8078 ( .A1(n7148), .A2(keyinput_f89), .B1(n7147), .B2(keyinput_f8), 
        .ZN(n7146) );
  OAI221_X1 U8079 ( .B1(n7148), .B2(keyinput_f89), .C1(n7147), .C2(keyinput_f8), .A(n7146), .ZN(n7157) );
  AOI22_X1 U8080 ( .A1(n7151), .A2(keyinput_f10), .B1(keyinput_f85), .B2(n7150), .ZN(n7149) );
  OAI221_X1 U8081 ( .B1(n7151), .B2(keyinput_f10), .C1(n7150), .C2(
        keyinput_f85), .A(n7149), .ZN(n7156) );
  AOI22_X1 U8082 ( .A1(n7154), .A2(keyinput_f42), .B1(n7153), .B2(keyinput_f9), 
        .ZN(n7152) );
  OAI221_X1 U8083 ( .B1(n7154), .B2(keyinput_f42), .C1(n7153), .C2(keyinput_f9), .A(n7152), .ZN(n7155) );
  NOR4_X1 U8084 ( .A1(n7158), .A2(n7157), .A3(n7156), .A4(n7155), .ZN(n7209)
         );
  OAI22_X1 U8085 ( .A1(n7161), .A2(keyinput_f26), .B1(n7160), .B2(keyinput_f33), .ZN(n7159) );
  AOI221_X1 U8086 ( .B1(n7161), .B2(keyinput_f26), .C1(keyinput_f33), .C2(
        n7160), .A(n7159), .ZN(n7174) );
  OAI22_X1 U8087 ( .A1(n7164), .A2(keyinput_f57), .B1(n7163), .B2(
        keyinput_f107), .ZN(n7162) );
  AOI221_X1 U8088 ( .B1(n7164), .B2(keyinput_f57), .C1(keyinput_f107), .C2(
        n7163), .A(n7162), .ZN(n7173) );
  OAI22_X1 U8089 ( .A1(n7167), .A2(keyinput_f76), .B1(n7166), .B2(keyinput_f98), .ZN(n7165) );
  AOI221_X1 U8090 ( .B1(n7167), .B2(keyinput_f76), .C1(keyinput_f98), .C2(
        n7166), .A(n7165), .ZN(n7172) );
  OAI22_X1 U8091 ( .A1(n7170), .A2(keyinput_f30), .B1(n7169), .B2(keyinput_f99), .ZN(n7168) );
  AOI221_X1 U8092 ( .B1(n7170), .B2(keyinput_f30), .C1(keyinput_f99), .C2(
        n7169), .A(n7168), .ZN(n7171) );
  NAND4_X1 U8093 ( .A1(n7174), .A2(n7173), .A3(n7172), .A4(n7171), .ZN(n7207)
         );
  OAI22_X1 U8094 ( .A1(keyinput_f110), .A2(n7177), .B1(n7176), .B2(
        keyinput_f71), .ZN(n7175) );
  AOI221_X1 U8095 ( .B1(n7177), .B2(keyinput_f110), .C1(n7176), .C2(
        keyinput_f71), .A(n7175), .ZN(n7190) );
  OAI22_X1 U8096 ( .A1(n7180), .A2(keyinput_f86), .B1(n7179), .B2(keyinput_f79), .ZN(n7178) );
  AOI221_X1 U8097 ( .B1(n7180), .B2(keyinput_f86), .C1(keyinput_f79), .C2(
        n7179), .A(n7178), .ZN(n7189) );
  OAI22_X1 U8098 ( .A1(n7183), .A2(keyinput_f91), .B1(n7182), .B2(keyinput_f72), .ZN(n7181) );
  AOI221_X1 U8099 ( .B1(n7183), .B2(keyinput_f91), .C1(keyinput_f72), .C2(
        n7182), .A(n7181), .ZN(n7188) );
  INV_X1 U8100 ( .A(keyinput_f121), .ZN(n7185) );
  OAI22_X1 U8101 ( .A1(n7186), .A2(keyinput_f19), .B1(n7185), .B2(
        DATAWIDTH_REG_17__SCAN_IN), .ZN(n7184) );
  AOI221_X1 U8102 ( .B1(n7186), .B2(keyinput_f19), .C1(
        DATAWIDTH_REG_17__SCAN_IN), .C2(n7185), .A(n7184), .ZN(n7187) );
  NAND4_X1 U8103 ( .A1(n7190), .A2(n7189), .A3(n7188), .A4(n7187), .ZN(n7206)
         );
  AOI22_X1 U8104 ( .A1(n7193), .A2(keyinput_f48), .B1(keyinput_f50), .B2(n7192), .ZN(n7191) );
  OAI221_X1 U8105 ( .B1(n7193), .B2(keyinput_f48), .C1(n7192), .C2(
        keyinput_f50), .A(n7191), .ZN(n7205) );
  OAI22_X1 U8106 ( .A1(n7196), .A2(keyinput_f23), .B1(n7195), .B2(keyinput_f46), .ZN(n7194) );
  AOI221_X1 U8107 ( .B1(n7196), .B2(keyinput_f23), .C1(keyinput_f46), .C2(
        n7195), .A(n7194), .ZN(n7203) );
  OAI22_X1 U8108 ( .A1(n7199), .A2(keyinput_f35), .B1(n7198), .B2(keyinput_f14), .ZN(n7197) );
  AOI221_X1 U8109 ( .B1(n7199), .B2(keyinput_f35), .C1(keyinput_f14), .C2(
        n7198), .A(n7197), .ZN(n7202) );
  XNOR2_X1 U8110 ( .A(keyinput_f106), .B(DATAWIDTH_REG_2__SCAN_IN), .ZN(n7201)
         );
  XNOR2_X1 U8111 ( .A(keyinput_f34), .B(BS16_N), .ZN(n7200) );
  NAND4_X1 U8112 ( .A1(n7203), .A2(n7202), .A3(n7201), .A4(n7200), .ZN(n7204)
         );
  NOR4_X1 U8113 ( .A1(n7207), .A2(n7206), .A3(n7205), .A4(n7204), .ZN(n7208)
         );
  NAND4_X1 U8114 ( .A1(n7211), .A2(n7210), .A3(n7209), .A4(n7208), .ZN(n7212)
         );
  NOR4_X1 U8115 ( .A1(n7215), .A2(n7214), .A3(n7213), .A4(n7212), .ZN(n7217)
         );
  XNOR2_X1 U8116 ( .A(DATAI_9_), .B(keyinput_f22), .ZN(n7216) );
  OAI22_X1 U8117 ( .A1(n7217), .A2(n7216), .B1(DATAI_9_), .B2(keyinput_g22), 
        .ZN(n7218) );
  AOI211_X1 U8118 ( .C1(DATAI_9_), .C2(keyinput_g22), .A(n7219), .B(n7218), 
        .ZN(n7223) );
  AOI22_X1 U8119 ( .A1(n7221), .A2(BYTEENABLE_REG_3__SCAN_IN), .B1(
        BE_N_REG_3__SCAN_IN), .B2(n7220), .ZN(n7222) );
  XNOR2_X1 U8120 ( .A(n7223), .B(n7222), .ZN(U3445) );
  AND2_X2 U4089 ( .A1(n3219), .A2(n3217), .ZN(n3776) );
  INV_X1 U4275 ( .A(n3460), .ZN(n5220) );
  AND2_X1 U4215 ( .A1(n3455), .A2(n3361), .ZN(n3438) );
  BUF_X2 U3632 ( .A(n3457), .Z(n4091) );
  AND2_X1 U3722 ( .A1(n3574), .A2(n3631), .ZN(n3151) );
  CLKBUF_X1 U3685 ( .A(n3361), .Z(n3717) );
  CLKBUF_X2 U3604 ( .A(n3776), .Z(n3534) );
  CLKBUF_X2 U4407 ( .A(n3407), .Z(n3599) );
  CLKBUF_X1 U3621 ( .A(n3597), .Z(n3538) );
  AND4_X1 U3631 ( .A1(n3234), .A2(n3233), .A3(n3232), .A4(n3231), .ZN(n3235)
         );
  AND4_X1 U3643 ( .A1(n3230), .A2(n3229), .A3(n3228), .A4(n3227), .ZN(n3236)
         );
  AND2_X2 U3645 ( .A1(n3894), .A2(n3220), .ZN(n5087) );
  AND2_X1 U3653 ( .A1(n3643), .A2(n4385), .ZN(n3428) );
  NAND2_X1 U3674 ( .A1(n3151), .A2(n4772), .ZN(n3716) );
  CLKBUF_X3 U3723 ( .A(n3159), .Z(n4773) );
  AND2_X2 U3739 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5669) );
  CLKBUF_X1 U3898 ( .A(n3868), .Z(n6806) );
  CLKBUF_X1 U4085 ( .A(n6047), .Z(n6058) );
  CLKBUF_X1 U4100 ( .A(n5203), .Z(n5204) );
  AND2_X2 U4107 ( .A1(n4604), .A2(n3166), .ZN(n4715) );
  AOI21_X2 U4112 ( .B1(n5225), .B2(n6113), .A(n5217), .ZN(n5218) );
  CLKBUF_X1 U4269 ( .A(n5111), .Z(n3152) );
  CLKBUF_X1 U4406 ( .A(n5051), .Z(n5085) );
endmodule

