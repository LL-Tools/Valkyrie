

module b15_C_SARLock_k_128_8 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3445, 
        U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208, U3207, 
        U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198, U3197, 
        U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188, U3187, 
        U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180, U3179, 
        U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170, U3169, 
        U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160, U3159, 
        U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453, U3150, 
        U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141, U3140, 
        U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131, U3130, 
        U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121, U3120, 
        U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111, U3110, 
        U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101, U3100, 
        U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091, U3090, 
        U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081, U3080, 
        U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071, U3070, 
        U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061, U3060, 
        U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051, U3050, 
        U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041, U3040, 
        U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031, U3030, 
        U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021, U3020, 
        U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464, U3465, 
        U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010, U3009, 
        U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000, U2999, 
        U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990, U2989, 
        U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980, U2979, 
        U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970, U2969, 
        U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960, U2959, 
        U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950, U2949, 
        U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940, U2939, 
        U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930, U2929, 
        U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920, U2919, 
        U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910, U2909, 
        U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900, U2899, 
        U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890, U2889, 
        U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880, U2879, 
        U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870, U2869, 
        U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860, U2859, 
        U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850, U2849, 
        U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840, U2839, 
        U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830, U2829, 
        U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820, U2819, 
        U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810, U2809, 
        U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800, U2799, 
        U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793, U3471, 
        U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3129, n3130, n3132, n3133, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3656, n3657, n3658, n3659, n3660, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121;

  AOI21_X1 U3567 ( .B1(n5497), .B2(n5496), .A(n5485), .ZN(n5706) );
  OR2_X1 U3568 ( .A1(n5495), .A2(n3213), .ZN(n4071) );
  NOR2_X1 U3569 ( .A1(n3915), .A2(n3850), .ZN(n3851) );
  CLKBUF_X1 U3570 ( .A(n3476), .Z(n3975) );
  CLKBUF_X2 U3571 ( .A(n4001), .Z(n3140) );
  INV_X2 U3572 ( .A(n3492), .ZN(n4585) );
  AND2_X2 U3573 ( .A1(n3259), .A2(n4604), .ZN(n3470) );
  NAND2_X2 U3574 ( .A1(n3259), .A2(n3258), .ZN(n3455) );
  AND2_X1 U3575 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4621) );
  NOR2_X1 U3576 ( .A1(n3915), .A2(n6934), .ZN(n3916) );
  CLKBUF_X2 U3577 ( .A(n3462), .Z(n4430) );
  CLKBUF_X2 U3578 ( .A(n3404), .Z(n4421) );
  NAND2_X1 U3579 ( .A1(n4495), .A2(n4621), .ZN(n3436) );
  OAI22_X1 U3580 ( .A1(n6934), .A2(keyinput119), .B1(n6933), .B2(
        ADDRESS_REG_11__SCAN_IN), .ZN(n6932) );
  AOI221_X1 U3581 ( .B1(n6934), .B2(keyinput119), .C1(ADDRESS_REG_11__SCAN_IN), 
        .C2(n6933), .A(n6932), .ZN(n6947) );
  NAND2_X1 U3582 ( .A1(n3488), .A2(n3392), .ZN(n3425) );
  NAND2_X1 U3583 ( .A1(n3492), .A2(n4656), .ZN(n3174) );
  NOR2_X1 U3584 ( .A1(n5513), .A2(n5498), .ZN(n4237) );
  INV_X1 U3585 ( .A(n4578), .ZN(n4574) );
  INV_X4 U3586 ( .A(n6133), .ZN(n6222) );
  INV_X1 U3587 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6937) );
  INV_X1 U3588 ( .A(n3510), .ZN(n3392) );
  AND2_X4 U3589 ( .A1(n3618), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3259)
         );
  OAI22_X2 U3590 ( .A1(n4133), .A2(n4132), .B1(n4136), .B2(n4363), .ZN(n4141)
         );
  XNOR2_X1 U3591 ( .A(n5423), .B(n5422), .ZN(n5429) );
  OR2_X1 U3592 ( .A1(n5495), .A2(n3211), .ZN(n4449) );
  CLKBUF_X1 U3593 ( .A(n5495), .Z(n5496) );
  NAND2_X1 U3594 ( .A1(n5508), .A2(n5509), .ZN(n5495) );
  AOI21_X1 U3595 ( .B1(n5754), .B2(n5721), .A(n5720), .ZN(n5747) );
  NOR2_X2 U3596 ( .A1(n5522), .A2(n5628), .ZN(n5508) );
  NOR2_X1 U3597 ( .A1(n5535), .A2(n5663), .ZN(n5654) );
  CLKBUF_X1 U3598 ( .A(n5383), .Z(n5557) );
  NAND2_X1 U3599 ( .A1(n5772), .A2(n5773), .ZN(n5758) );
  OAI21_X1 U3600 ( .B1(n5772), .B2(n3239), .A(n3236), .ZN(n5996) );
  INV_X2 U3601 ( .A(n6156), .ZN(n6110) );
  NAND2_X1 U3602 ( .A1(n3160), .A2(n3152), .ZN(n4316) );
  INV_X1 U3603 ( .A(n6206), .ZN(n6171) );
  NOR3_X2 U3604 ( .A1(n5648), .A2(n5629), .A3(n3175), .ZN(n5512) );
  CLKBUF_X2 U3605 ( .A(n6283), .Z(n6346) );
  AND2_X1 U3606 ( .A1(n5394), .A2(n3184), .ZN(n5658) );
  BUF_X1 U3607 ( .A(n3617), .Z(n3133) );
  NAND2_X1 U3609 ( .A1(n3507), .A2(n3506), .ZN(n4372) );
  AND2_X1 U3610 ( .A1(n3495), .A2(n4084), .ZN(n3534) );
  INV_X2 U3611 ( .A(n6782), .ZN(n4309) );
  NAND2_X1 U3612 ( .A1(n3500), .A2(n3487), .ZN(n3555) );
  NAND2_X1 U3613 ( .A1(n3493), .A2(n3392), .ZN(n3536) );
  CLKBUF_X2 U3614 ( .A(n3489), .Z(n4848) );
  NAND2_X2 U3615 ( .A1(n3356), .A2(n3355), .ZN(n3510) );
  INV_X2 U3616 ( .A(n5400), .ZN(n3118) );
  AND4_X1 U3617 ( .A1(n3373), .A2(n3372), .A3(n3371), .A4(n3370), .ZN(n3385)
         );
  AND4_X1 U3618 ( .A1(n3382), .A2(n3381), .A3(n3380), .A4(n3379), .ZN(n3383)
         );
  AND4_X1 U3619 ( .A1(n3444), .A2(n3443), .A3(n3442), .A4(n3441), .ZN(n3450)
         );
  BUF_X2 U3620 ( .A(n4428), .Z(n4015) );
  CLKBUF_X2 U3621 ( .A(n3471), .Z(n3920) );
  CLKBUF_X2 U3622 ( .A(n3453), .Z(n4423) );
  CLKBUF_X2 U3623 ( .A(n3470), .Z(n4429) );
  BUF_X2 U3624 ( .A(n3461), .Z(n4431) );
  CLKBUF_X2 U3625 ( .A(n3477), .Z(n3996) );
  INV_X2 U3626 ( .A(n3455), .ZN(n4428) );
  NOR2_X1 U3627 ( .A1(n7021), .A2(n6211), .ZN(n3691) );
  INV_X2 U3628 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3166) );
  AND2_X2 U3629 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4491) );
  NOR2_X1 U3630 ( .A1(n5427), .A2(n3242), .ZN(n5428) );
  AOI21_X1 U3631 ( .B1(n3194), .B2(n6356), .A(n4458), .ZN(n4459) );
  AOI21_X1 U3632 ( .B1(n3194), .B2(n6110), .A(n3191), .ZN(n3190) );
  INV_X1 U3633 ( .A(n5466), .ZN(n3194) );
  NOR2_X1 U3634 ( .A1(n5745), .A2(n3240), .ZN(n5739) );
  NAND2_X1 U3636 ( .A1(n5974), .A2(n5709), .ZN(n5701) );
  AND2_X1 U3637 ( .A1(n5654), .A2(n3202), .ZN(n5521) );
  NAND2_X1 U3638 ( .A1(n5717), .A2(n5718), .ZN(n5983) );
  CLKBUF_X1 U3639 ( .A(n5535), .Z(n5536) );
  INV_X1 U3640 ( .A(n5383), .ZN(n3199) );
  OAI21_X1 U3641 ( .B1(n5996), .B2(n3159), .A(n5994), .ZN(n3158) );
  NAND2_X1 U3642 ( .A1(n3223), .A2(n3226), .ZN(n4337) );
  NAND2_X1 U3643 ( .A1(n4329), .A2(n3229), .ZN(n3162) );
  NAND2_X1 U3644 ( .A1(n4326), .A2(n4325), .ZN(n5299) );
  INV_X1 U3645 ( .A(n4677), .ZN(n3767) );
  AND2_X1 U3646 ( .A1(n4247), .A2(n4246), .ZN(n4248) );
  AND2_X1 U3647 ( .A1(n3230), .A2(n4331), .ZN(n3161) );
  OR2_X1 U3648 ( .A1(n5809), .A2(n5671), .ZN(n4247) );
  AND2_X1 U3649 ( .A1(n3234), .A2(n5319), .ZN(n3229) );
  INV_X1 U3650 ( .A(n3231), .ZN(n3230) );
  OR2_X1 U3651 ( .A1(n5462), .A2(n4244), .ZN(n5809) );
  NAND2_X1 U3652 ( .A1(n5422), .A2(n3212), .ZN(n3211) );
  AND2_X2 U3653 ( .A1(n6193), .A2(n5391), .ZN(n6133) );
  XNOR2_X1 U3654 ( .A(n4303), .B(n4302), .ZN(n4788) );
  NAND2_X1 U3655 ( .A1(n4517), .A2(n4532), .ZN(n4555) );
  INV_X1 U3656 ( .A(n5446), .ZN(n5444) );
  AND2_X1 U3657 ( .A1(n4552), .A2(n3125), .ZN(n3126) );
  NAND2_X1 U3658 ( .A1(n3766), .A2(n3765), .ZN(n4798) );
  OAI211_X1 U3659 ( .C1(n4294), .C2(n3883), .A(n3736), .B(n3735), .ZN(n4552)
         );
  NAND2_X1 U3660 ( .A1(n7121), .A2(n3656), .ZN(n3196) );
  OAI21_X1 U3661 ( .B1(n4276), .B2(n4091), .A(n4275), .ZN(n4277) );
  NAND2_X1 U3662 ( .A1(n3160), .A2(n3730), .ZN(n3756) );
  NOR2_X1 U3663 ( .A1(n4068), .A2(n5488), .ZN(n3249) );
  NAND2_X2 U3664 ( .A1(n3689), .A2(n3715), .ZN(n4276) );
  OR2_X1 U3665 ( .A1(n4055), .A2(n7097), .ZN(n4068) );
  CLKBUF_X1 U3666 ( .A(n4573), .Z(n5030) );
  NAND2_X1 U3667 ( .A1(n6362), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4260)
         );
  NAND2_X1 U3668 ( .A1(n3627), .A2(n3605), .ZN(n4573) );
  NOR2_X1 U3669 ( .A1(n4735), .A2(n4819), .ZN(n6437) );
  NOR2_X1 U3670 ( .A1(n4700), .A2(n4819), .ZN(n6454) );
  OR2_X1 U3671 ( .A1(n4040), .A2(n3247), .ZN(n4052) );
  OR2_X2 U3672 ( .A1(n6776), .A2(n5387), .ZN(n6193) );
  NAND2_X1 U3673 ( .A1(n3687), .A2(n3686), .ZN(n4743) );
  NAND2_X1 U3674 ( .A1(n3602), .A2(n3601), .ZN(n3627) );
  NAND2_X2 U3675 ( .A1(n3615), .A2(n3614), .ZN(n4578) );
  NAND2_X1 U3676 ( .A1(n3669), .A2(n3668), .ZN(n4625) );
  NOR2_X2 U3677 ( .A1(n6645), .A2(n6660), .ZN(n4703) );
  NAND2_X1 U3678 ( .A1(n3599), .A2(n3611), .ZN(n3615) );
  AND2_X2 U3679 ( .A1(n4146), .A2(n4145), .ZN(n6645) );
  NOR2_X1 U3680 ( .A1(n3994), .A2(n3993), .ZN(n4023) );
  AND2_X1 U3681 ( .A1(n4899), .A2(n3148), .ZN(n5347) );
  NOR2_X2 U3682 ( .A1(n4799), .A2(n4800), .ZN(n4899) );
  NAND2_X1 U3683 ( .A1(n3577), .A2(n3576), .ZN(n3628) );
  NAND3_X1 U3684 ( .A1(n3178), .A2(n3179), .A3(n3181), .ZN(n4799) );
  INV_X1 U3685 ( .A(n3576), .ZN(n3578) );
  NAND2_X1 U3686 ( .A1(n3639), .A2(n3638), .ZN(n3668) );
  NAND2_X1 U3687 ( .A1(n3527), .A2(n3526), .ZN(n3577) );
  NOR2_X1 U3688 ( .A1(n6934), .A2(n3902), .ZN(n3935) );
  NOR2_X1 U3689 ( .A1(n4163), .A2(n4162), .ZN(n4546) );
  NOR2_X1 U3690 ( .A1(n4553), .A2(n3183), .ZN(n3179) );
  NOR2_X1 U3691 ( .A1(n3850), .A2(n3847), .ZN(n3879) );
  XNOR2_X1 U3692 ( .A(n4161), .B(n4469), .ZN(n4539) );
  AND3_X1 U3693 ( .A1(n3570), .A2(n3579), .A3(n3569), .ZN(n3573) );
  NAND2_X1 U3694 ( .A1(n4158), .A2(n4157), .ZN(n4161) );
  CLKBUF_X1 U3695 ( .A(n3501), .Z(n4076) );
  OR2_X1 U3696 ( .A1(n4147), .A2(n4319), .ZN(n3579) );
  AND2_X1 U3697 ( .A1(n4147), .A2(n3674), .ZN(n4138) );
  AND3_X1 U3698 ( .A1(n3596), .A2(n3595), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n3597) );
  NAND2_X1 U3699 ( .A1(n4848), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4147) );
  NOR2_X4 U3700 ( .A1(n4168), .A2(n3174), .ZN(n4164) );
  NAND2_X2 U3701 ( .A1(n3118), .A2(n3492), .ZN(n4168) );
  OR2_X1 U3702 ( .A1(n3567), .A2(n3566), .ZN(n4319) );
  NOR2_X1 U3703 ( .A1(n5400), .A2(n6872), .ZN(n3500) );
  NOR2_X1 U3704 ( .A1(n6889), .A2(n3768), .ZN(n3784) );
  NAND2_X1 U3705 ( .A1(n5400), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3674) );
  OR2_X1 U3706 ( .A1(n3590), .A2(n3589), .ZN(n4254) );
  OR2_X1 U3707 ( .A1(n3553), .A2(n3552), .ZN(n4253) );
  NAND2_X1 U3708 ( .A1(n4656), .A2(n4599), .ZN(n4354) );
  AND3_X2 U3709 ( .A1(n3485), .A2(n3484), .A3(n3483), .ZN(n5400) );
  AND4_X2 U3710 ( .A1(n3145), .A2(n3423), .A3(n3422), .A4(n3421), .ZN(n4599)
         );
  NAND2_X1 U3711 ( .A1(n3365), .A2(n3245), .ZN(n3487) );
  AND4_X1 U3712 ( .A1(n3350), .A2(n3349), .A3(n3348), .A4(n3347), .ZN(n3356)
         );
  AND4_X1 U3713 ( .A1(n3354), .A2(n3353), .A3(n3352), .A4(n3351), .ZN(n3355)
         );
  AND2_X1 U3714 ( .A1(n3241), .A2(n3475), .ZN(n3484) );
  AND2_X1 U3715 ( .A1(n3468), .A2(n3467), .ZN(n3485) );
  NOR2_X1 U3716 ( .A1(n3750), .A2(n5278), .ZN(n3761) );
  AND4_X1 U3717 ( .A1(n3360), .A2(n3359), .A3(n3358), .A4(n3357), .ZN(n3365)
         );
  NAND2_X1 U3718 ( .A1(n3734), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3750)
         );
  AND4_X1 U3719 ( .A1(n3412), .A2(n3411), .A3(n3410), .A4(n3409), .ZN(n3423)
         );
  AND4_X1 U3720 ( .A1(n3448), .A2(n3447), .A3(n3446), .A4(n3445), .ZN(n3449)
         );
  AND4_X1 U3721 ( .A1(n3440), .A2(n3439), .A3(n3438), .A4(n3437), .ZN(n3451)
         );
  AND4_X1 U3722 ( .A1(n3433), .A2(n3432), .A3(n3431), .A4(n3430), .ZN(n3452)
         );
  AND4_X1 U3723 ( .A1(n3466), .A2(n3465), .A3(n3464), .A4(n3463), .ZN(n3467)
         );
  AND4_X1 U3724 ( .A1(n3459), .A2(n3458), .A3(n3457), .A4(n3456), .ZN(n3468)
         );
  AND4_X1 U3725 ( .A1(n3378), .A2(n3377), .A3(n3376), .A4(n3375), .ZN(n3384)
         );
  AND4_X1 U3726 ( .A1(n3369), .A2(n3368), .A3(n3367), .A4(n3366), .ZN(n3386)
         );
  AND4_X1 U3727 ( .A1(n3416), .A2(n3415), .A3(n3414), .A4(n3413), .ZN(n3422)
         );
  AND4_X1 U3728 ( .A1(n3420), .A2(n3419), .A3(n3418), .A4(n3417), .ZN(n3421)
         );
  BUF_X1 U3729 ( .A(n3460), .Z(n3644) );
  BUF_X2 U3730 ( .A(n3469), .Z(n3257) );
  BUF_X2 U3731 ( .A(n3478), .Z(n4610) );
  NOR2_X1 U3732 ( .A1(n3711), .A2(n6180), .ZN(n3734) );
  INV_X1 U3733 ( .A(n4450), .ZN(n3637) );
  AND2_X2 U3734 ( .A1(n4495), .A2(n4608), .ZN(n3471) );
  AND2_X2 U3735 ( .A1(n4490), .A2(n4621), .ZN(n3143) );
  AND2_X1 U3736 ( .A1(n4604), .A2(n4491), .ZN(n3462) );
  AND2_X2 U3737 ( .A1(n3166), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4495)
         );
  AND2_X2 U3738 ( .A1(n3215), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4608)
         );
  AND2_X4 U3739 ( .A1(n4621), .A2(n4491), .ZN(n3561) );
  INV_X1 U3740 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3215) );
  NOR2_X2 U3741 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4490) );
  CLKBUF_X1 U3742 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n6925) );
  INV_X2 U3743 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6872) );
  NAND2_X1 U3744 ( .A1(n3162), .A2(n3161), .ZN(n3119) );
  CLKBUF_X1 U3745 ( .A(n4662), .Z(n3120) );
  NAND2_X1 U3746 ( .A1(n3162), .A2(n3161), .ZN(n4333) );
  NAND2_X1 U3747 ( .A1(n4288), .A2(n4287), .ZN(n4662) );
  OAI21_X1 U3748 ( .B1(n4276), .B2(n3883), .A(n3695), .ZN(n4532) );
  NAND2_X1 U3749 ( .A1(n5758), .A2(n3238), .ZN(n3246) );
  XNOR2_X1 U3750 ( .A(n3653), .B(n3652), .ZN(n3664) );
  NAND2_X2 U3751 ( .A1(n5983), .A2(n5981), .ZN(n5754) );
  NOR2_X1 U3752 ( .A1(n5535), .A2(n5663), .ZN(n3121) );
  NAND2_X1 U3753 ( .A1(n3121), .A2(n3122), .ZN(n5522) );
  AND2_X1 U3754 ( .A1(n5523), .A2(n3202), .ZN(n3122) );
  INV_X1 U3755 ( .A(n4555), .ZN(n3124) );
  NAND2_X2 U3756 ( .A1(n4337), .A2(n4336), .ZN(n5772) );
  NAND2_X4 U3757 ( .A1(n4316), .A2(n4318), .ZN(n4327) );
  CLKBUF_X1 U3758 ( .A(n5352), .Z(n3123) );
  INV_X1 U3759 ( .A(n4556), .ZN(n3125) );
  AND2_X1 U3760 ( .A1(n3124), .A2(n3125), .ZN(n4550) );
  INV_X1 U3761 ( .A(n7121), .ZN(n3127) );
  AND2_X1 U3762 ( .A1(n4978), .A2(n3207), .ZN(n3129) );
  OAI211_X1 U3763 ( .C1(n6641), .C2(n3514), .A(n4381), .B(n4378), .ZN(n3130)
         );
  OAI211_X1 U3764 ( .C1(n6641), .C2(n3514), .A(n4381), .B(n4378), .ZN(n3519)
         );
  AND2_X1 U3765 ( .A1(n3489), .A2(n3488), .ZN(n3490) );
  AND2_X2 U3766 ( .A1(n3498), .A2(n3497), .ZN(n4073) );
  AND2_X1 U3767 ( .A1(n4495), .A2(n4608), .ZN(n3132) );
  XNOR2_X1 U3768 ( .A(n3578), .B(n3577), .ZN(n3617) );
  AND2_X2 U3769 ( .A1(n4490), .A2(n4604), .ZN(n4001) );
  NAND2_X2 U3770 ( .A1(n3505), .A2(n3504), .ZN(n3632) );
  AOI21_X2 U3771 ( .B1(n3503), .B2(STATE2_REG_0__SCAN_IN), .A(n3502), .ZN(
        n3504) );
  NAND2_X2 U3772 ( .A1(n3663), .A2(n3662), .ZN(n4517) );
  OAI222_X1 U3773 ( .A1(n5670), .A2(n5429), .B1(n6231), .B2(n5459), .C1(n5799), 
        .C2(n5671), .ZN(U2829) );
  AND2_X2 U3774 ( .A1(n4896), .A2(n4979), .ZN(n4978) );
  NOR2_X2 U3775 ( .A1(n4796), .A2(n4897), .ZN(n4896) );
  NAND4_X4 U3776 ( .A1(n3386), .A2(n3385), .A3(n3384), .A4(n3383), .ZN(n3493)
         );
  AND2_X1 U3777 ( .A1(n4604), .A2(n4491), .ZN(n3135) );
  AND2_X1 U3778 ( .A1(n4604), .A2(n4491), .ZN(n3136) );
  INV_X2 U3779 ( .A(n3487), .ZN(n3489) );
  XNOR2_X2 U3780 ( .A(n3865), .B(n3866), .ZN(n5357) );
  AND2_X4 U3781 ( .A1(n4490), .A2(n4608), .ZN(n3460) );
  AND2_X2 U3782 ( .A1(n3259), .A2(n4608), .ZN(n3137) );
  INV_X1 U3783 ( .A(n3137), .ZN(n3138) );
  AND2_X1 U3784 ( .A1(n3259), .A2(n4608), .ZN(n3560) );
  AND2_X1 U3785 ( .A1(n3259), .A2(n4608), .ZN(n3139) );
  AND2_X4 U3786 ( .A1(n4495), .A2(n4604), .ZN(n3476) );
  NOR2_X2 U3787 ( .A1(n5495), .A2(n3210), .ZN(n5423) );
  AND2_X4 U3788 ( .A1(n4608), .A2(n4491), .ZN(n3477) );
  INV_X1 U3789 ( .A(n3732), .ZN(n3160) );
  INV_X1 U3790 ( .A(n4334), .ZN(n3228) );
  NOR2_X1 U3791 ( .A1(n5647), .A2(n3206), .ZN(n3205) );
  INV_X1 U3792 ( .A(n5655), .ZN(n3206) );
  OAI22_X1 U3793 ( .A1(n4138), .A2(n3759), .B1(n3555), .B2(n5235), .ZN(n3760)
         );
  NOR2_X2 U3794 ( .A1(n3510), .A2(n6937), .ZN(n3893) );
  NAND2_X1 U3795 ( .A1(n5879), .A2(n6909), .ZN(n3159) );
  INV_X1 U3796 ( .A(n4230), .ZN(n4238) );
  NAND2_X1 U3797 ( .A1(n4301), .A2(n4300), .ZN(n4303) );
  OAI21_X1 U3798 ( .B1(n4294), .B2(n4091), .A(n4293), .ZN(n4295) );
  INV_X1 U3799 ( .A(n4234), .ZN(n4201) );
  OR2_X1 U3800 ( .A1(n4656), .A2(n5400), .ZN(n4230) );
  NAND2_X1 U3801 ( .A1(n4099), .A2(n4134), .ZN(n4365) );
  OR2_X1 U3802 ( .A1(n4135), .A2(n4098), .ZN(n4099) );
  AND2_X1 U3803 ( .A1(n3535), .A2(n3488), .ZN(n3429) );
  AND2_X1 U3804 ( .A1(n6193), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5607) );
  INV_X1 U3805 ( .A(n4281), .ZN(n4289) );
  INV_X1 U3806 ( .A(n4106), .ZN(n4102) );
  AOI21_X1 U3807 ( .B1(n4486), .B2(n6872), .A(n3554), .ZN(n3574) );
  NOR2_X1 U3808 ( .A1(n3650), .A2(n3649), .ZN(n4264) );
  AND2_X2 U3809 ( .A1(n3690), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3258)
         );
  INV_X1 U3810 ( .A(n4077), .ZN(n3532) );
  NOR2_X1 U3811 ( .A1(n3555), .A2(n4076), .ZN(n3502) );
  NAND2_X1 U3812 ( .A1(n5486), .A2(n3214), .ZN(n3213) );
  INV_X1 U3813 ( .A(n5497), .ZN(n3214) );
  INV_X1 U3814 ( .A(n4061), .ZN(n4440) );
  NAND2_X1 U3815 ( .A1(n4492), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4061) );
  NAND2_X1 U3816 ( .A1(n4978), .A2(n3207), .ZN(n3865) );
  NOR2_X1 U3817 ( .A1(n5316), .A2(n3208), .ZN(n3207) );
  INV_X1 U3818 ( .A(n3209), .ZN(n3208) );
  INV_X1 U3819 ( .A(n3757), .ZN(n3758) );
  AND2_X1 U3820 ( .A1(n3182), .A2(n4559), .ZN(n3181) );
  INV_X1 U3821 ( .A(n4534), .ZN(n3182) );
  OR2_X1 U3822 ( .A1(n3685), .A2(n3684), .ZN(n4274) );
  INV_X1 U3823 ( .A(n4138), .ZN(n4129) );
  INV_X1 U3824 ( .A(n3555), .ZN(n4136) );
  OR2_X1 U3825 ( .A1(n6763), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4450) );
  AND2_X1 U3826 ( .A1(n4352), .A2(n4353), .ZN(n6644) );
  AND2_X1 U3827 ( .A1(n3151), .A2(n3185), .ZN(n3184) );
  INV_X1 U3828 ( .A(n5665), .ZN(n3185) );
  NOR2_X1 U3829 ( .A1(n4072), .A2(n3213), .ZN(n3212) );
  INV_X1 U3830 ( .A(n3915), .ZN(n4447) );
  NAND2_X1 U3831 ( .A1(n4703), .A2(n4521), .ZN(n6302) );
  NOR2_X1 U3832 ( .A1(n5635), .A2(n3203), .ZN(n3202) );
  INV_X1 U3833 ( .A(n3204), .ZN(n3203) );
  NAND2_X1 U3834 ( .A1(n5654), .A2(n3204), .ZN(n5634) );
  AOI21_X1 U3835 ( .B1(n4298), .B2(n3893), .A(n3753), .ZN(n4678) );
  AND2_X1 U3836 ( .A1(n3220), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3219)
         );
  AND2_X1 U3837 ( .A1(n5708), .A2(n3156), .ZN(n3220) );
  AND2_X1 U3838 ( .A1(n4221), .A2(n4220), .ZN(n5644) );
  INV_X1 U3839 ( .A(n3227), .ZN(n3226) );
  NAND2_X1 U3840 ( .A1(n3119), .A2(n5328), .ZN(n5364) );
  NAND2_X1 U3841 ( .A1(n5364), .A2(n5363), .ZN(n5362) );
  NOR2_X1 U3842 ( .A1(n5283), .A2(n3235), .ZN(n3234) );
  INV_X1 U3843 ( .A(n4328), .ZN(n3235) );
  INV_X1 U3844 ( .A(n5275), .ZN(n3187) );
  OR2_X1 U3845 ( .A1(n4327), .A2(n5291), .ZN(n5284) );
  AND2_X1 U3846 ( .A1(n4384), .A2(n4359), .ZN(n6640) );
  AND2_X1 U3847 ( .A1(n4377), .A2(n4376), .ZN(n4403) );
  NOR2_X1 U3848 ( .A1(n4450), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6368) );
  OR2_X1 U3849 ( .A1(n4114), .A2(n4365), .ZN(n4146) );
  NAND2_X1 U3850 ( .A1(n4144), .A2(n4143), .ZN(n4145) );
  OR2_X1 U3851 ( .A1(n4138), .A2(n4365), .ZN(n4144) );
  OR2_X1 U3852 ( .A1(n4276), .A2(n4572), .ZN(n5031) );
  INV_X1 U3853 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n7081) );
  NOR2_X1 U3854 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4584), .ZN(n4860) );
  AND2_X1 U3855 ( .A1(n5389), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4149) );
  INV_X1 U3856 ( .A(n6672), .ZN(n6660) );
  AND2_X1 U3857 ( .A1(n5476), .A2(REIP_REG_31__SCAN_IN), .ZN(n3193) );
  AND2_X1 U3858 ( .A1(n6193), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U3859 ( .A1(n5607), .A2(n5393), .ZN(n6095) );
  INV_X1 U3860 ( .A(n6166), .ZN(n6220) );
  INV_X1 U3861 ( .A(n5464), .ZN(n3195) );
  INV_X1 U3862 ( .A(n6413), .ZN(n6389) );
  INV_X1 U3863 ( .A(n6520), .ZN(n6564) );
  CLKBUF_X1 U3864 ( .A(n4571), .Z(n4572) );
  NAND2_X1 U3865 ( .A1(n5400), .A2(n4599), .ZN(n4077) );
  OR2_X1 U3866 ( .A1(n4138), .A2(n4289), .ZN(n3707) );
  INV_X1 U3867 ( .A(n3731), .ZN(n3730) );
  OR2_X1 U3868 ( .A1(n3746), .A2(n3745), .ZN(n4307) );
  OR2_X1 U3869 ( .A1(n3705), .A2(n3704), .ZN(n4281) );
  NAND2_X1 U3870 ( .A1(n4090), .A2(n3489), .ZN(n3528) );
  OR2_X1 U3871 ( .A1(n3455), .A2(n3374), .ZN(n3377) );
  OR2_X1 U3872 ( .A1(n3455), .A2(n3434), .ZN(n3438) );
  INV_X1 U3873 ( .A(n5644), .ZN(n3176) );
  AND2_X1 U3874 ( .A1(n3205), .A2(n5643), .ZN(n3204) );
  NOR2_X1 U3875 ( .A1(n3951), .A2(n5760), .ZN(n3968) );
  NOR2_X1 U3876 ( .A1(n5538), .A2(n3198), .ZN(n3197) );
  INV_X1 U3877 ( .A(n3200), .ZN(n3198) );
  AND2_X1 U3878 ( .A1(n6001), .A2(n3201), .ZN(n3200) );
  INV_X1 U3879 ( .A(n5556), .ZN(n3201) );
  AND2_X1 U3880 ( .A1(n5272), .A2(n5215), .ZN(n3209) );
  INV_X1 U3881 ( .A(n3893), .ZN(n3883) );
  INV_X1 U3882 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n7021) );
  NOR2_X1 U3883 ( .A1(n4168), .A2(n5540), .ZN(n4234) );
  INV_X1 U3884 ( .A(n6021), .ZN(n3186) );
  OAI21_X1 U3885 ( .B1(n5363), .B2(n3228), .A(n4335), .ZN(n3227) );
  NOR2_X1 U3886 ( .A1(n3228), .A2(n3225), .ZN(n3224) );
  NOR2_X1 U3887 ( .A1(n5178), .A2(n3189), .ZN(n3188) );
  INV_X1 U3888 ( .A(n4900), .ZN(n3189) );
  NAND2_X1 U3889 ( .A1(n4268), .A2(n4267), .ZN(n4269) );
  INV_X1 U3890 ( .A(n4149), .ZN(n3636) );
  NAND2_X1 U3891 ( .A1(n3627), .A2(n3626), .ZN(n3665) );
  OR2_X1 U3892 ( .A1(n3555), .A2(n4091), .ZN(n4114) );
  AOI22_X1 U3893 ( .A1(n4137), .A2(n4136), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6872), .ZN(n4140) );
  AOI21_X1 U3894 ( .B1(n4138), .B2(n4090), .A(n4366), .ZN(n4139) );
  AND2_X1 U3895 ( .A1(n4807), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6555) );
  AOI21_X1 U3896 ( .B1(n6677), .B2(n4707), .A(n4576), .ZN(n4584) );
  AND2_X1 U3897 ( .A1(n4367), .A2(n4366), .ZN(n6643) );
  INV_X1 U3898 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6211) );
  NAND2_X1 U3899 ( .A1(n4083), .A2(n3543), .ZN(n3576) );
  AND4_X1 U3900 ( .A1(n3542), .A2(n3534), .A3(n3541), .A4(n3540), .ZN(n3543)
         );
  NAND2_X1 U3901 ( .A1(n3535), .A2(n4309), .ZN(n3541) );
  AND2_X1 U3902 ( .A1(n4213), .A2(n5539), .ZN(n5656) );
  OAI21_X1 U3903 ( .B1(n5930), .B2(n3150), .A(n4010), .ZN(n5647) );
  AND2_X1 U3904 ( .A1(n4706), .A2(n4705), .ZN(n6245) );
  NAND2_X1 U3905 ( .A1(n3249), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4454)
         );
  INV_X1 U3906 ( .A(n3212), .ZN(n3210) );
  NAND2_X1 U3907 ( .A1(n3248), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4055)
         );
  INV_X1 U3908 ( .A(n4052), .ZN(n3248) );
  NAND2_X1 U3909 ( .A1(n4036), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4040)
         );
  OAI21_X1 U3910 ( .B1(n3150), .B2(n5980), .A(n4047), .ZN(n5628) );
  OAI21_X1 U3911 ( .B1(n3150), .B2(n5918), .A(n4033), .ZN(n5635) );
  NAND2_X1 U3912 ( .A1(n3990), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3994)
         );
  AND2_X1 U3913 ( .A1(n3992), .A2(n3991), .ZN(n5655) );
  AND2_X1 U3914 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n3968), .ZN(n3990)
         );
  OR2_X1 U3915 ( .A1(n5993), .A2(n3150), .ZN(n3973) );
  NAND2_X1 U3916 ( .A1(n3199), .A2(n3200), .ZN(n5534) );
  NAND2_X1 U3917 ( .A1(n3884), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3902)
         );
  AND2_X1 U3918 ( .A1(n3879), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3884)
         );
  NAND2_X1 U3919 ( .A1(n3129), .A2(n3866), .ZN(n3867) );
  CLKBUF_X1 U3920 ( .A(n5353), .Z(n5354) );
  NAND2_X1 U3921 ( .A1(n3831), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3847)
         );
  NAND2_X1 U3922 ( .A1(n3800), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3814)
         );
  INV_X1 U3923 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3827) );
  AND2_X1 U3924 ( .A1(n3783), .A2(n3782), .ZN(n4897) );
  NAND2_X1 U3925 ( .A1(n3761), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3768)
         );
  INV_X1 U3926 ( .A(n3764), .ZN(n3765) );
  NAND2_X1 U3927 ( .A1(n4305), .A2(n3893), .ZN(n3766) );
  CLKBUF_X1 U3928 ( .A(n4796), .Z(n4797) );
  NAND2_X1 U3929 ( .A1(n3222), .A2(n7006), .ZN(n3221) );
  INV_X1 U3930 ( .A(n4470), .ZN(n5460) );
  NAND2_X1 U3931 ( .A1(n3173), .A2(n3172), .ZN(n5446) );
  INV_X1 U3932 ( .A(n4242), .ZN(n3172) );
  NAND2_X1 U3933 ( .A1(n5416), .A2(n5708), .ZN(n4417) );
  NAND2_X1 U3934 ( .A1(n5717), .A2(n4341), .ZN(n3216) );
  OR2_X1 U3935 ( .A1(n3240), .A2(n3168), .ZN(n3167) );
  NAND2_X1 U3936 ( .A1(n4327), .A2(n3157), .ZN(n3168) );
  NAND2_X1 U3937 ( .A1(n5745), .A2(n5738), .ZN(n5732) );
  AND2_X1 U3938 ( .A1(n4211), .A2(n4210), .ZN(n5665) );
  AOI21_X1 U3939 ( .B1(n3237), .B2(n3238), .A(INSTADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n3236) );
  INV_X1 U3940 ( .A(n5773), .ZN(n3237) );
  NAND2_X1 U3941 ( .A1(n5394), .A2(n5560), .ZN(n6020) );
  NAND2_X1 U3942 ( .A1(n5377), .A2(n5378), .ZN(n5395) );
  OAI21_X1 U3943 ( .B1(n5284), .B2(n3232), .A(n5320), .ZN(n3231) );
  NAND2_X1 U3944 ( .A1(n4899), .A2(n3144), .ZN(n5274) );
  AND2_X1 U3945 ( .A1(n4899), .A2(n3188), .ZN(n5267) );
  NAND2_X1 U3946 ( .A1(n4899), .A2(n4900), .ZN(n5177) );
  INV_X1 U3947 ( .A(n4296), .ZN(n3170) );
  INV_X1 U3948 ( .A(n4788), .ZN(n3171) );
  INV_X1 U3949 ( .A(n4680), .ZN(n3183) );
  NAND2_X1 U3950 ( .A1(n3178), .A2(n3181), .ZN(n4557) );
  NOR2_X1 U3951 ( .A1(n4533), .A2(n4534), .ZN(n4558) );
  INV_X1 U3952 ( .A(n4168), .ZN(n4540) );
  XNOR2_X1 U3953 ( .A(n4260), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4563)
         );
  OR2_X1 U3954 ( .A1(n5338), .A2(n4391), .ZN(n5370) );
  AND2_X1 U3955 ( .A1(n4230), .A2(n3174), .ZN(n4470) );
  INV_X1 U3956 ( .A(n3522), .ZN(n3523) );
  OAI21_X1 U3957 ( .B1(n3521), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        STATE2_REG_0__SCAN_IN), .ZN(n3522) );
  NAND2_X1 U3958 ( .A1(n5074), .A2(n6872), .ZN(n3687) );
  OR2_X1 U3959 ( .A1(n3425), .A2(n3387), .ZN(n6619) );
  INV_X1 U3960 ( .A(n6619), .ZN(n4492) );
  INV_X1 U3961 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n6889) );
  OR2_X1 U3962 ( .A1(n4584), .A2(n6754), .ZN(n4862) );
  INV_X1 U3963 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n5389) );
  NOR2_X1 U3964 ( .A1(n5924), .A2(n5432), .ZN(n5906) );
  NOR2_X1 U3965 ( .A1(n5878), .A2(n5947), .ZN(n5950) );
  INV_X1 U3966 ( .A(n6163), .ZN(n6182) );
  AND2_X1 U3967 ( .A1(n5607), .A2(n5407), .ZN(n6209) );
  AND2_X1 U3968 ( .A1(n5608), .A2(n6156), .ZN(n6166) );
  NAND2_X2 U3969 ( .A1(n4154), .A2(n4153), .ZN(n6231) );
  OR2_X1 U3970 ( .A1(n4523), .A2(n4168), .ZN(n4153) );
  AND2_X1 U3971 ( .A1(n5467), .A2(n3511), .ZN(n6238) );
  AND2_X1 U3972 ( .A1(n5467), .A2(n5456), .ZN(n6242) );
  AND2_X1 U3973 ( .A1(n5467), .A2(n4530), .ZN(n5414) );
  INV_X1 U3974 ( .A(n5414), .ZN(n5381) );
  NOR2_X1 U3975 ( .A1(n6779), .A2(n6245), .ZN(n6260) );
  INV_X1 U3976 ( .A(n6659), .ZN(n6779) );
  INV_X1 U3978 ( .A(n4701), .ZN(n4702) );
  INV_X1 U3979 ( .A(n4457), .ZN(n4458) );
  INV_X1 U3980 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n5278) );
  INV_X1 U3981 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6180) );
  OR2_X1 U3982 ( .A1(n6350), .A2(n6364), .ZN(n6361) );
  AND2_X1 U3983 ( .A1(n6068), .A2(n4451), .ZN(n6350) );
  INV_X1 U3984 ( .A(n6350), .ZN(n6365) );
  OAI21_X1 U3985 ( .B1(n5701), .B2(n3155), .A(n3218), .ZN(n3217) );
  NOR2_X1 U3986 ( .A1(n5648), .A2(n5644), .ZN(n5637) );
  NAND2_X1 U3987 ( .A1(n5758), .A2(n4338), .ZN(n5765) );
  NAND2_X1 U3988 ( .A1(n5362), .A2(n4334), .ZN(n5782) );
  NAND2_X1 U3989 ( .A1(n3233), .A2(n5284), .ZN(n5322) );
  NAND2_X1 U3990 ( .A1(n4329), .A2(n3234), .ZN(n3233) );
  NAND2_X1 U3991 ( .A1(n4329), .A2(n4328), .ZN(n5287) );
  NAND2_X1 U3992 ( .A1(n6640), .A2(n4385), .ZN(n6403) );
  OR2_X1 U3993 ( .A1(n4403), .A2(n4402), .ZN(n6413) );
  INV_X1 U3994 ( .A(n6014), .ZN(n6415) );
  INV_X1 U3995 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6556) );
  INV_X1 U3996 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n7064) );
  INV_X1 U3997 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6631) );
  INV_X1 U3998 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6637) );
  NOR2_X1 U3999 ( .A1(n3515), .A2(n6645), .ZN(n4576) );
  AND2_X1 U4000 ( .A1(n4582), .A2(n4581), .ZN(n4934) );
  OR2_X1 U4001 ( .A1(n4642), .A2(n4578), .ZN(n6796) );
  OAI211_X1 U4002 ( .C1(n6458), .C2(n3515), .A(n6433), .B(n7081), .ZN(n6462)
         );
  OR3_X1 U4003 ( .A1(n5079), .A2(n5078), .A3(n5077), .ZN(n5114) );
  INV_X1 U4004 ( .A(n5063), .ZN(n6502) );
  INV_X1 U4005 ( .A(n6601), .ZN(n6503) );
  OR2_X1 U4006 ( .A1(n5031), .A2(n4714), .ZN(n6547) );
  INV_X1 U4007 ( .A(n6572), .ZN(n6498) );
  INV_X1 U4008 ( .A(n6595), .ZN(n6447) );
  AND2_X1 U4009 ( .A1(n4807), .A2(n4578), .ZN(n6612) );
  INV_X1 U4010 ( .A(n6589), .ZN(n6444) );
  OR3_X1 U4011 ( .A1(n4749), .A2(n4748), .A3(n4747), .ZN(n4972) );
  AND2_X1 U4012 ( .A1(n4149), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6672) );
  AND2_X1 U4013 ( .A1(n6663), .A2(n6662), .ZN(n6752) );
  OAI21_X1 U4014 ( .B1(n5793), .B2(n6095), .A(n3190), .ZN(U2796) );
  OR3_X1 U4015 ( .A1(n5475), .A2(n3193), .A3(n3192), .ZN(n3191) );
  NAND2_X1 U4016 ( .A1(n5472), .A2(n5471), .ZN(n3192) );
  INV_X1 U4017 ( .A(n4327), .ZN(n5994) );
  INV_X2 U4018 ( .A(n3174), .ZN(n5540) );
  NAND2_X1 U4019 ( .A1(n4978), .A2(n3209), .ZN(n5271) );
  NAND2_X1 U4020 ( .A1(n5654), .A2(n5655), .ZN(n5646) );
  NAND2_X1 U4021 ( .A1(n3536), .A2(n4656), .ZN(n3535) );
  OR2_X1 U4022 ( .A1(n5648), .A2(n3175), .ZN(n3141) );
  AND2_X1 U4023 ( .A1(n3154), .A2(n3178), .ZN(n3142) );
  AND2_X1 U4024 ( .A1(n5654), .A2(n3205), .ZN(n5642) );
  NAND2_X1 U4025 ( .A1(n6193), .A2(n5388), .ZN(n6156) );
  AND2_X1 U4026 ( .A1(n3188), .A2(n5268), .ZN(n3144) );
  AND4_X1 U4027 ( .A1(n3408), .A2(n3407), .A3(n3406), .A4(n3405), .ZN(n3145)
         );
  NOR2_X1 U4028 ( .A1(n5383), .A2(n5556), .ZN(n5558) );
  NAND2_X1 U4029 ( .A1(n3216), .A2(n4343), .ZN(n5973) );
  INV_X1 U4030 ( .A(n4553), .ZN(n3180) );
  OR2_X1 U4031 ( .A1(n5745), .A2(n3167), .ZN(n3146) );
  INV_X1 U4032 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n6906) );
  INV_X1 U4033 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3690) );
  AND2_X1 U4034 ( .A1(n4536), .A2(n4537), .ZN(n3660) );
  INV_X1 U4035 ( .A(n5319), .ZN(n3232) );
  NOR2_X1 U4036 ( .A1(n4327), .A2(n5300), .ZN(n3147) );
  AND2_X1 U4037 ( .A1(n3144), .A2(n3187), .ZN(n3148) );
  NAND2_X1 U4038 ( .A1(n3707), .A2(n3706), .ZN(n3716) );
  NAND2_X1 U4039 ( .A1(n4327), .A2(n5893), .ZN(n3149) );
  OR2_X1 U4040 ( .A1(n3488), .A2(n6937), .ZN(n3244) );
  OR2_X1 U4041 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3150) );
  INV_X1 U4042 ( .A(n4373), .ZN(n3511) );
  AND2_X1 U4043 ( .A1(n4978), .A2(n5215), .ZN(n5214) );
  AND2_X1 U4044 ( .A1(n5560), .A2(n3186), .ZN(n3151) );
  NAND2_X1 U4045 ( .A1(n3162), .A2(n3230), .ZN(n5327) );
  AOI21_X1 U4046 ( .B1(n4788), .B2(n3170), .A(n3165), .ZN(n3169) );
  NAND2_X1 U4047 ( .A1(n5394), .A2(n3151), .ZN(n5544) );
  AND2_X1 U4048 ( .A1(n3429), .A2(n3428), .ZN(n4352) );
  INV_X1 U4049 ( .A(n3173), .ZN(n5445) );
  NOR2_X1 U4050 ( .A1(n5500), .A2(n4404), .ZN(n3173) );
  AND2_X1 U4051 ( .A1(n3730), .A2(n3758), .ZN(n3152) );
  INV_X1 U4052 ( .A(n3239), .ZN(n3238) );
  NAND2_X1 U4053 ( .A1(n3149), .A2(n4338), .ZN(n3239) );
  NOR3_X1 U4054 ( .A1(n5648), .A2(n5644), .A3(n3177), .ZN(n5524) );
  AND2_X1 U4055 ( .A1(n4344), .A2(n4343), .ZN(n3153) );
  NAND2_X1 U4056 ( .A1(n6231), .A2(n4148), .ZN(n5671) );
  NAND2_X1 U4057 ( .A1(n4703), .A2(n6649), .ZN(n6068) );
  NAND2_X1 U4058 ( .A1(n4297), .A2(n4296), .ZN(n4787) );
  INV_X1 U4059 ( .A(n5328), .ZN(n3225) );
  NOR2_X1 U4060 ( .A1(n5395), .A2(n5396), .ZN(n5394) );
  INV_X1 U4061 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3618) );
  AND2_X1 U4062 ( .A1(n3181), .A2(n3180), .ZN(n3154) );
  INV_X1 U4063 ( .A(n5636), .ZN(n3177) );
  OR2_X2 U4064 ( .A1(n3402), .A2(n3401), .ZN(n4656) );
  OR2_X1 U4065 ( .A1(n5417), .A2(n3221), .ZN(n3155) );
  INV_X1 U4066 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3222) );
  AND2_X1 U4067 ( .A1(n5805), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3156)
         );
  AND2_X1 U4068 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3157) );
  NOR2_X2 U4069 ( .A1(n6370), .A2(n4590), .ZN(n6604) );
  OR2_X1 U4070 ( .A1(n6679), .A2(n6564), .ZN(n6370) );
  NAND2_X2 U4071 ( .A1(n4339), .A2(n3158), .ZN(n5717) );
  AND2_X2 U4072 ( .A1(n5747), .A2(n5748), .ZN(n5745) );
  NAND3_X1 U4073 ( .A1(n3164), .A2(n5262), .A3(n3163), .ZN(n4315) );
  NAND2_X1 U4074 ( .A1(n3171), .A2(n4304), .ZN(n3163) );
  NAND2_X1 U4075 ( .A1(n4297), .A2(n3169), .ZN(n3164) );
  INV_X1 U4076 ( .A(n4304), .ZN(n3165) );
  NAND2_X1 U4077 ( .A1(n5724), .A2(n3146), .ZN(n5725) );
  OAI21_X1 U4078 ( .B1(n4297), .B2(n3171), .A(n3169), .ZN(n5263) );
  OR2_X2 U4079 ( .A1(n3246), .A2(n4393), .ZN(n4339) );
  OR2_X2 U4080 ( .A1(n5299), .A2(n3147), .ZN(n4329) );
  NAND2_X2 U4081 ( .A1(n3118), .A2(n4585), .ZN(n6782) );
  NAND3_X1 U4082 ( .A1(n3176), .A2(n5525), .A3(n5636), .ZN(n3175) );
  INV_X1 U4083 ( .A(n4533), .ZN(n3178) );
  XNOR2_X2 U4084 ( .A(n3195), .B(n5465), .ZN(n5793) );
  NAND2_X1 U4085 ( .A1(n3469), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3446) );
  AND2_X2 U4086 ( .A1(n3258), .A2(n4490), .ZN(n3469) );
  NAND2_X1 U4087 ( .A1(n3196), .A2(n4518), .ZN(n3663) );
  NOR2_X1 U4088 ( .A1(n3196), .A2(n4518), .ZN(n4519) );
  NAND2_X1 U4089 ( .A1(n3199), .A2(n3197), .ZN(n5535) );
  NOR2_X1 U4090 ( .A1(n5495), .A2(n5497), .ZN(n5485) );
  NAND2_X1 U4091 ( .A1(n3688), .A2(n4743), .ZN(n3715) );
  NAND3_X1 U4092 ( .A1(n3688), .A2(n4743), .A3(n3716), .ZN(n3732) );
  INV_X1 U4093 ( .A(n4074), .ZN(n3507) );
  NAND2_X1 U4094 ( .A1(n3491), .A2(n4074), .ZN(n3495) );
  NAND2_X1 U4095 ( .A1(n3490), .A2(n3496), .ZN(n4074) );
  NAND2_X1 U4096 ( .A1(n3216), .A2(n3153), .ZN(n4346) );
  AND2_X1 U4097 ( .A1(n5416), .A2(n3220), .ZN(n5420) );
  NAND2_X1 U4098 ( .A1(n5416), .A2(n3219), .ZN(n3218) );
  XNOR2_X1 U4099 ( .A(n3217), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5796)
         );
  NAND2_X1 U4100 ( .A1(n4333), .A2(n3224), .ZN(n3223) );
  NAND2_X1 U4101 ( .A1(n5723), .A2(n5722), .ZN(n5724) );
  XNOR2_X1 U4102 ( .A(n5725), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5838)
         );
  NAND2_X1 U4103 ( .A1(n3868), .A2(n3867), .ZN(n5352) );
  NAND2_X1 U4104 ( .A1(n3615), .A2(n4317), .ZN(n3604) );
  NAND2_X1 U4105 ( .A1(n5352), .A2(n5355), .ZN(n5353) );
  NAND2_X1 U4106 ( .A1(n4352), .A2(n3513), .ZN(n4378) );
  AOI21_X1 U4107 ( .B1(n4499), .B2(n6872), .A(n3651), .ZN(n3653) );
  INV_X1 U4108 ( .A(n5353), .ZN(n3901) );
  NAND2_X1 U4109 ( .A1(n3901), .A2(n3900), .ZN(n5383) );
  XNOR2_X1 U4110 ( .A(n3715), .B(n3716), .ZN(n4280) );
  AOI21_X1 U4111 ( .B1(n4072), .B2(n4071), .A(n5423), .ZN(n5691) );
  INV_X1 U4112 ( .A(n5684), .ZN(n6239) );
  NAND2_X1 U4113 ( .A1(n5467), .A2(n4529), .ZN(n5684) );
  AND2_X1 U4114 ( .A1(n4327), .A2(n5860), .ZN(n3240) );
  AND3_X1 U4115 ( .A1(n3474), .A2(n3473), .A3(n3472), .ZN(n3241) );
  NAND2_X1 U4116 ( .A1(n3610), .A2(n3609), .ZN(n4536) );
  OR2_X1 U4117 ( .A1(n5426), .A2(n5425), .ZN(n3242) );
  AND2_X1 U4118 ( .A1(n3529), .A2(n3528), .ZN(n3243) );
  INV_X1 U4119 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4270) );
  AND4_X1 U4120 ( .A1(n3364), .A2(n3363), .A3(n3362), .A4(n3361), .ZN(n3245)
         );
  INV_X1 U4121 ( .A(n4253), .ZN(n3568) );
  NAND2_X1 U4122 ( .A1(n4327), .A2(n4340), .ZN(n4341) );
  INV_X1 U4123 ( .A(n4656), .ZN(n3531) );
  NAND2_X1 U4124 ( .A1(n5455), .A2(n3510), .ZN(n3496) );
  OR2_X1 U4125 ( .A1(n4138), .A2(n3727), .ZN(n3729) );
  INV_X1 U4126 ( .A(n4319), .ZN(n3759) );
  NAND2_X1 U4127 ( .A1(n3118), .A2(n4599), .ZN(n3530) );
  NAND2_X1 U4128 ( .A1(n3532), .A2(n3531), .ZN(n4085) );
  AND2_X1 U4129 ( .A1(n3729), .A2(n3728), .ZN(n3731) );
  OR2_X1 U4130 ( .A1(n3726), .A2(n3725), .ZN(n4291) );
  AND4_X1 U4131 ( .A1(n4081), .A2(n4356), .A3(n4080), .A4(n4079), .ZN(n4082)
         );
  OR2_X1 U4132 ( .A1(n3436), .A2(n3435), .ZN(n3437) );
  AND2_X1 U4133 ( .A1(n3749), .A2(n3748), .ZN(n3757) );
  OR2_X1 U4134 ( .A1(n3688), .A2(n4743), .ZN(n3689) );
  INV_X1 U4135 ( .A(n5382), .ZN(n3900) );
  INV_X1 U4136 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3850) );
  AND2_X1 U4137 ( .A1(n3784), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3800)
         );
  INV_X1 U4138 ( .A(n4269), .ZN(n4271) );
  NAND2_X1 U4139 ( .A1(n3631), .A2(n3630), .ZN(n3667) );
  NAND2_X1 U4140 ( .A1(n3404), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3475)
         );
  OR2_X1 U4141 ( .A1(n4135), .A2(n4134), .ZN(n4366) );
  NOR2_X1 U4142 ( .A1(n5563), .A2(n5566), .ZN(n6085) );
  OR2_X1 U4143 ( .A1(n4454), .A2(n6923), .ZN(n4455) );
  NAND2_X1 U4144 ( .A1(n5400), .A2(n4585), .ZN(n4522) );
  AND2_X1 U4145 ( .A1(n5449), .A2(n4443), .ZN(n4444) );
  AND2_X1 U4146 ( .A1(n3937), .A2(n3936), .ZN(n6001) );
  INV_X1 U4147 ( .A(n6403), .ZN(n4391) );
  INV_X1 U4148 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4627) );
  INV_X1 U4149 ( .A(n5227), .ZN(n5082) );
  AND4_X1 U4150 ( .A1(n3482), .A2(n3481), .A3(n3480), .A4(n3479), .ZN(n3483)
         );
  NAND2_X1 U4151 ( .A1(n3613), .A2(n3612), .ZN(n3614) );
  AND2_X1 U4152 ( .A1(n4023), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4026)
         );
  NOR2_X1 U4153 ( .A1(n3814), .A2(n3827), .ZN(n3831) );
  XNOR2_X1 U4154 ( .A(n4455), .B(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5390)
         );
  OR2_X1 U4155 ( .A1(n6351), .A2(n5386), .ZN(n5387) );
  INV_X1 U4156 ( .A(n4522), .ZN(n5606) );
  AND2_X1 U4157 ( .A1(n4160), .A2(n4159), .ZN(n4469) );
  AOI21_X1 U4158 ( .B1(n5776), .B2(n5390), .A(n4456), .ZN(n4457) );
  OAI21_X1 U4159 ( .B1(n3150), .B2(n5704), .A(n4063), .ZN(n5497) );
  INV_X1 U4160 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6934) );
  NAND2_X1 U4161 ( .A1(n3691), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3711)
         );
  INV_X1 U4162 ( .A(n4105), .ZN(n4379) );
  AND2_X1 U4163 ( .A1(n4406), .A2(n6397), .ZN(n5868) );
  INV_X1 U4164 ( .A(n5887), .ZN(n5288) );
  OR2_X1 U4165 ( .A1(n5009), .A2(n4574), .ZN(n5248) );
  OR2_X1 U4166 ( .A1(n4642), .A2(n4574), .ZN(n6792) );
  AND2_X1 U4167 ( .A1(n4572), .A2(n4715), .ZN(n6423) );
  OR2_X1 U4168 ( .A1(n5031), .A2(n6421), .ZN(n6541) );
  AND2_X1 U4169 ( .A1(n5030), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6508) );
  NAND2_X1 U4170 ( .A1(n3673), .A2(n3672), .ZN(n4717) );
  AND2_X1 U4171 ( .A1(n4572), .A2(n4716), .ZN(n4807) );
  INV_X1 U4172 ( .A(n4860), .ZN(n4819) );
  AOI21_X1 U4173 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6556), .A(n4819), .ZN(
        n6568) );
  NAND2_X1 U4174 ( .A1(n6265), .A2(n4465), .ZN(n6776) );
  OR2_X1 U4175 ( .A1(n5911), .A2(n5436), .ZN(n5517) );
  AND2_X1 U4176 ( .A1(n4026), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4036)
         );
  AND2_X1 U4177 ( .A1(n5390), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5388) );
  INV_X1 U4178 ( .A(n6095), .ZN(n6214) );
  OR2_X1 U4179 ( .A1(n6231), .A2(n4245), .ZN(n4246) );
  INV_X1 U4180 ( .A(n5671), .ZN(n6227) );
  INV_X1 U4181 ( .A(n5467), .ZN(n6241) );
  OAI21_X1 U4182 ( .B1(n4309), .B2(n6778), .A(n6266), .ZN(n6283) );
  NAND2_X1 U4183 ( .A1(n3935), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3951)
         );
  INV_X1 U4184 ( .A(n6361), .ZN(n5776) );
  AND2_X1 U4185 ( .A1(n4417), .A2(n5805), .ZN(n4350) );
  INV_X1 U4186 ( .A(n6401), .ZN(n6351) );
  AND2_X1 U4187 ( .A1(n5890), .A2(n5889), .ZN(n6043) );
  OR2_X1 U4188 ( .A1(n4392), .A2(n4666), .ZN(n5341) );
  XNOR2_X1 U4189 ( .A(n4286), .B(n4285), .ZN(n4778) );
  INV_X1 U4190 ( .A(n6368), .ZN(n6401) );
  NOR2_X1 U4191 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6520) );
  INV_X1 U4192 ( .A(n4647), .ZN(n5201) );
  INV_X1 U4193 ( .A(n6796), .ZN(n5175) );
  AND2_X1 U4194 ( .A1(n6423), .A2(n6422), .ZN(n6491) );
  AND2_X1 U4195 ( .A1(n6423), .A2(n5072), .ZN(n6493) );
  NOR2_X1 U4196 ( .A1(n5031), .A2(n5030), .ZN(n4876) );
  INV_X1 U4197 ( .A(n6583), .ZN(n6440) );
  INV_X1 U4198 ( .A(n6617), .ZN(n6460) );
  INV_X1 U4199 ( .A(n6541), .ZN(n6550) );
  INV_X1 U4200 ( .A(n6547), .ZN(n6543) );
  INV_X1 U4201 ( .A(n6370), .ZN(n6356) );
  AND2_X1 U4202 ( .A1(n4807), .A2(n4574), .ZN(n6608) );
  NAND2_X1 U4203 ( .A1(n4703), .A2(n4462), .ZN(n6265) );
  OR3_X1 U4204 ( .A1(n5507), .A2(n6737), .A3(n5437), .ZN(n5484) );
  INV_X1 U4205 ( .A(n6148), .ZN(n6212) );
  INV_X1 U4206 ( .A(n6209), .ZN(n6150) );
  NAND4_X1 U4207 ( .A1(n6302), .A2(n4528), .A3(n4527), .A4(n4526), .ZN(n5467)
         );
  NAND2_X1 U4208 ( .A1(n6245), .A2(n3118), .ZN(n5130) );
  INV_X1 U4209 ( .A(n6245), .ZN(n6264) );
  NAND2_X2 U4210 ( .A1(n4703), .A2(n4702), .ZN(n6348) );
  INV_X1 U4211 ( .A(n6356), .ZN(n5989) );
  AND2_X1 U4212 ( .A1(n4397), .A2(n5865), .ZN(n5861) );
  OR2_X1 U4213 ( .A1(n4403), .A2(n4383), .ZN(n6014) );
  OR2_X1 U4214 ( .A1(n4403), .A2(n6622), .ZN(n6419) );
  OR2_X1 U4215 ( .A1(n4860), .A2(n4633), .ZN(n6420) );
  AND2_X1 U4216 ( .A1(n5224), .A2(n5223), .ZN(n5261) );
  AOI21_X1 U4217 ( .B1(n4646), .B2(n4645), .A(n4644), .ZN(n4941) );
  OR2_X1 U4218 ( .A1(n4827), .A2(n4574), .ZN(n4865) );
  AOI21_X1 U4219 ( .B1(n4821), .B2(n4822), .A(n4820), .ZN(n4870) );
  INV_X1 U4220 ( .A(n6491), .ZN(n6465) );
  NAND2_X1 U4221 ( .A1(n4876), .A2(n4578), .ZN(n5121) );
  AOI21_X1 U4222 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5041), .A(n5038), .ZN(
        n6507) );
  AOI21_X1 U4223 ( .B1(n4721), .B2(n4720), .A(n4719), .ZN(n4949) );
  NAND2_X1 U4224 ( .A1(n4950), .A2(n4578), .ZN(n5003) );
  AND2_X1 U4225 ( .A1(n6683), .A2(STATE_REG_1__SCAN_IN), .ZN(n6788) );
  OAI21_X1 U4226 ( .B1(n5674), .B2(n5670), .A(n4248), .ZN(U2830) );
  OAI21_X1 U4227 ( .B1(n5700), .B2(n6014), .A(n4416), .ZN(U2990) );
  INV_X1 U4228 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5760) );
  INV_X1 U4229 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3993) );
  INV_X1 U4230 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3247) );
  INV_X1 U4231 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n7097) );
  INV_X1 U4232 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5488) );
  INV_X1 U4233 ( .A(n3249), .ZN(n3251) );
  INV_X1 U4234 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n3250) );
  NAND2_X1 U4235 ( .A1(n3251), .A2(n3250), .ZN(n3252) );
  NAND2_X1 U4236 ( .A1(n4454), .A2(n3252), .ZN(n5689) );
  AND2_X2 U4237 ( .A1(n3258), .A2(n4495), .ZN(n3453) );
  AOI22_X1 U4238 ( .A1(n3560), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4423), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3256) );
  AND2_X2 U4239 ( .A1(n3259), .A2(n4621), .ZN(n3461) );
  AOI22_X1 U4240 ( .A1(n3460), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3255) );
  INV_X2 U4241 ( .A(n3436), .ZN(n3404) );
  NOR2_X4 U4242 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4604) );
  AOI22_X1 U4243 ( .A1(n4421), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3254) );
  AND2_X2 U4244 ( .A1(n3258), .A2(n4491), .ZN(n3478) );
  AOI22_X1 U4245 ( .A1(n3477), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4610), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3253) );
  NAND4_X1 U4246 ( .A1(n3256), .A2(n3255), .A3(n3254), .A4(n3253), .ZN(n3266)
         );
  AOI22_X1 U4247 ( .A1(n3920), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3257), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3264) );
  AOI22_X1 U4248 ( .A1(n3476), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3263) );
  INV_X1 U4249 ( .A(n3143), .ZN(n3260) );
  INV_X2 U4250 ( .A(n3260), .ZN(n4422) );
  AOI22_X1 U4251 ( .A1(n4015), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4422), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3262) );
  AOI22_X1 U4252 ( .A1(n4430), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3261) );
  NAND4_X1 U4253 ( .A1(n3264), .A2(n3263), .A3(n3262), .A4(n3261), .ZN(n3265)
         );
  NOR2_X1 U4254 ( .A1(n3266), .A2(n3265), .ZN(n4420) );
  AOI22_X1 U4255 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n3920), .B1(n4431), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3270) );
  AOI22_X1 U4256 ( .A1(n4423), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4610), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3269) );
  AOI22_X1 U4257 ( .A1(n3996), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3268) );
  AOI22_X1 U4258 ( .A1(n3137), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3267) );
  NAND4_X1 U4259 ( .A1(n3270), .A2(n3269), .A3(n3268), .A4(n3267), .ZN(n3276)
         );
  AOI22_X1 U4260 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n3460), .B1(n4015), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3274) );
  AOI22_X1 U4261 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n3470), .B1(n3257), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3273) );
  AOI22_X1 U4262 ( .A1(n3975), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4422), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3272) );
  AOI22_X1 U4263 ( .A1(n4421), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3584), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3271) );
  NAND4_X1 U4264 ( .A1(n3274), .A2(n3273), .A3(n3272), .A4(n3271), .ZN(n3275)
         );
  NOR2_X1 U4265 ( .A1(n3276), .A2(n3275), .ZN(n4058) );
  AOI22_X1 U4266 ( .A1(n4431), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4421), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3280) );
  AOI22_X1 U4267 ( .A1(n3137), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4610), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3279) );
  AOI22_X1 U4268 ( .A1(n3975), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3278) );
  AOI22_X1 U4269 ( .A1(n4430), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3277) );
  NAND4_X1 U4270 ( .A1(n3280), .A2(n3279), .A3(n3278), .A4(n3277), .ZN(n3286)
         );
  AOI22_X1 U4271 ( .A1(n4423), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4015), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3284) );
  AOI22_X1 U4272 ( .A1(n3920), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3644), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3283) );
  AOI22_X1 U4273 ( .A1(n3470), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3257), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3282) );
  AOI22_X1 U4274 ( .A1(n3996), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4422), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3281) );
  NAND4_X1 U4275 ( .A1(n3284), .A2(n3283), .A3(n3282), .A4(n3281), .ZN(n3285)
         );
  NOR2_X1 U4276 ( .A1(n3286), .A2(n3285), .ZN(n4043) );
  AOI22_X1 U4277 ( .A1(n3996), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4610), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3290) );
  AOI22_X1 U4278 ( .A1(n4423), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4015), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3289) );
  AOI22_X1 U4279 ( .A1(n4421), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3257), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3288) );
  AOI22_X1 U4280 ( .A1(n4431), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3584), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3287) );
  NAND4_X1 U4281 ( .A1(n3290), .A2(n3289), .A3(n3288), .A4(n3287), .ZN(n3296)
         );
  AOI22_X1 U4282 ( .A1(n3920), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4429), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3294) );
  AOI22_X1 U4283 ( .A1(n3476), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3293) );
  AOI22_X1 U4284 ( .A1(n3137), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4422), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3292) );
  AOI22_X1 U4285 ( .A1(n3644), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3291) );
  NAND4_X1 U4286 ( .A1(n3294), .A2(n3293), .A3(n3292), .A4(n3291), .ZN(n3295)
         );
  NOR2_X1 U4287 ( .A1(n3296), .A2(n3295), .ZN(n4028) );
  AOI22_X1 U4288 ( .A1(n3477), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3476), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3300) );
  AOI22_X1 U4289 ( .A1(n3920), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3257), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3299) );
  AOI22_X1 U4290 ( .A1(n4610), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4422), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3298) );
  AOI22_X1 U4291 ( .A1(n4431), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3297) );
  NAND4_X1 U4292 ( .A1(n3300), .A2(n3299), .A3(n3298), .A4(n3297), .ZN(n3306)
         );
  AOI22_X1 U4293 ( .A1(n3137), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4015), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3304) );
  AOI22_X1 U4294 ( .A1(n4421), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4429), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3303) );
  AOI22_X1 U4295 ( .A1(n4423), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3302) );
  AOI22_X1 U4296 ( .A1(n3644), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3584), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3301) );
  NAND4_X1 U4297 ( .A1(n3304), .A2(n3303), .A3(n3302), .A4(n3301), .ZN(n3305)
         );
  NOR2_X1 U4298 ( .A1(n3306), .A2(n3305), .ZN(n4029) );
  OR2_X1 U4299 ( .A1(n4028), .A2(n4029), .ZN(n4035) );
  AOI22_X1 U4300 ( .A1(n3920), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3310) );
  AOI22_X1 U4301 ( .A1(n3477), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3476), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3309) );
  AOI22_X1 U4302 ( .A1(n4423), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3644), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3308) );
  AOI22_X1 U4303 ( .A1(n4610), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4422), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3307) );
  NAND4_X1 U4304 ( .A1(n3310), .A2(n3309), .A3(n3308), .A4(n3307), .ZN(n3316)
         );
  AOI22_X1 U4305 ( .A1(n3137), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4421), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3314) );
  AOI22_X1 U4306 ( .A1(n3257), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3313) );
  AOI22_X1 U4307 ( .A1(n4015), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3312) );
  AOI22_X1 U4308 ( .A1(n4429), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3311) );
  NAND4_X1 U4309 ( .A1(n3314), .A2(n3313), .A3(n3312), .A4(n3311), .ZN(n3315)
         );
  NOR2_X1 U4310 ( .A1(n3316), .A2(n3315), .ZN(n4034) );
  OR2_X1 U4311 ( .A1(n4035), .A2(n4034), .ZN(n4042) );
  NOR2_X1 U4312 ( .A1(n4043), .A2(n4042), .ZN(n4048) );
  INV_X1 U4313 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3679) );
  NOR2_X1 U4314 ( .A1(n3260), .A2(n3679), .ZN(n3318) );
  INV_X1 U4315 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4761) );
  INV_X1 U4316 ( .A(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5049) );
  OAI22_X1 U4317 ( .A1(n3138), .A2(n4761), .B1(n3455), .B2(n5049), .ZN(n3317)
         );
  AOI211_X1 U4318 ( .C1(INSTQUEUE_REG_9__3__SCAN_IN), .C2(n4423), .A(n3318), 
        .B(n3317), .ZN(n3326) );
  AOI22_X1 U4319 ( .A1(n3996), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3325) );
  AOI22_X1 U4320 ( .A1(n3975), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4610), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3324) );
  AOI22_X1 U4321 ( .A1(n3920), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4421), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3322) );
  AOI22_X1 U4322 ( .A1(n4429), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3257), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3321) );
  AOI22_X1 U4323 ( .A1(n3644), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3320) );
  AOI22_X1 U4324 ( .A1(n4431), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3319) );
  AND4_X1 U4325 ( .A1(n3322), .A2(n3321), .A3(n3320), .A4(n3319), .ZN(n3323)
         );
  NAND4_X1 U4326 ( .A1(n3326), .A2(n3325), .A3(n3324), .A4(n3323), .ZN(n4049)
         );
  NAND2_X1 U4327 ( .A1(n4048), .A2(n4049), .ZN(n4057) );
  NOR2_X1 U4328 ( .A1(n4058), .A2(n4057), .ZN(n4064) );
  AOI22_X1 U4329 ( .A1(n3137), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4428), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3330) );
  AOI22_X1 U4330 ( .A1(n3476), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4610), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3329) );
  AOI22_X1 U4331 ( .A1(n3996), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3328) );
  INV_X1 U4332 ( .A(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n7078) );
  AOI22_X1 U4333 ( .A1(n4423), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4422), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3327) );
  NAND4_X1 U4334 ( .A1(n3330), .A2(n3329), .A3(n3328), .A4(n3327), .ZN(n3336)
         );
  AOI22_X1 U4335 ( .A1(n3920), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4421), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3334) );
  AOI22_X1 U4336 ( .A1(n4429), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3257), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3333) );
  AOI22_X1 U4337 ( .A1(n3460), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3332) );
  AOI22_X1 U4338 ( .A1(n4431), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3331) );
  NAND4_X1 U4339 ( .A1(n3334), .A2(n3333), .A3(n3332), .A4(n3331), .ZN(n3335)
         );
  OR2_X1 U4340 ( .A1(n3336), .A2(n3335), .ZN(n4065) );
  NAND2_X1 U4341 ( .A1(n4064), .A2(n4065), .ZN(n4419) );
  XNOR2_X1 U4342 ( .A(n4420), .B(n4419), .ZN(n3390) );
  AOI22_X1 U4343 ( .A1(n4428), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3340) );
  AOI22_X1 U4344 ( .A1(n3476), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3478), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3339) );
  AOI22_X1 U4345 ( .A1(n3404), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3338) );
  AOI22_X1 U4346 ( .A1(n3560), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3453), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3337) );
  NAND4_X1 U4347 ( .A1(n3340), .A2(n3339), .A3(n3338), .A4(n3337), .ZN(n3346)
         );
  AOI22_X1 U4348 ( .A1(n3471), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3344) );
  AOI22_X1 U4349 ( .A1(n3477), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4001), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3343) );
  AOI22_X1 U4350 ( .A1(n3143), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3136), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3342) );
  AOI22_X1 U4351 ( .A1(n3461), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3341) );
  NAND4_X1 U4352 ( .A1(n3344), .A2(n3343), .A3(n3342), .A4(n3341), .ZN(n3345)
         );
  OR2_X2 U4353 ( .A1(n3346), .A2(n3345), .ZN(n3488) );
  AOI22_X1 U4354 ( .A1(n3471), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3404), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3350) );
  AOI22_X1 U4355 ( .A1(n3460), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3349) );
  AOI22_X1 U4356 ( .A1(n3470), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3348) );
  AOI22_X1 U4357 ( .A1(n3461), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3347) );
  AOI22_X1 U4358 ( .A1(n3560), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4428), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3354) );
  AOI22_X1 U4359 ( .A1(n3476), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3478), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3353) );
  AOI22_X1 U4360 ( .A1(n3477), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4001), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3352) );
  AOI22_X1 U4361 ( .A1(n3453), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3143), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3351) );
  AOI22_X1 U4362 ( .A1(n4428), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3139), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3360) );
  AOI22_X1 U4363 ( .A1(n3476), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3478), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3359) );
  AOI22_X1 U4364 ( .A1(n3477), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4001), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3358) );
  AOI22_X1 U4365 ( .A1(n3453), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3143), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3357) );
  AOI22_X1 U4366 ( .A1(n3460), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3136), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3364) );
  AOI22_X1 U4367 ( .A1(n3470), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3363) );
  AOI22_X1 U4368 ( .A1(n3404), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3132), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3362) );
  AOI22_X1 U4369 ( .A1(n3461), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3361) );
  NAND2_X1 U4370 ( .A1(n3139), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3369)
         );
  NAND2_X1 U4371 ( .A1(n3477), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3368)
         );
  NAND2_X1 U4372 ( .A1(n3461), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3367)
         );
  NAND2_X1 U4373 ( .A1(n3460), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3366) );
  NAND2_X1 U4374 ( .A1(n3404), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3373)
         );
  NAND2_X1 U4375 ( .A1(n3471), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3372) );
  NAND2_X1 U4376 ( .A1(n3470), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3371) );
  NAND2_X1 U4377 ( .A1(n3469), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3370) );
  NAND2_X1 U4378 ( .A1(n3453), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3378) );
  INV_X1 U4379 ( .A(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3374) );
  NAND2_X1 U4380 ( .A1(n3561), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3376)
         );
  NAND2_X1 U4381 ( .A1(n3135), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3375) );
  NAND2_X1 U4382 ( .A1(n3478), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3382) );
  NAND2_X1 U4383 ( .A1(n3476), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3381) );
  NAND2_X1 U4384 ( .A1(n4001), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3380) );
  NAND2_X1 U4385 ( .A1(n3143), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3379)
         );
  NAND2_X1 U4386 ( .A1(n3487), .A2(n3493), .ZN(n3387) );
  INV_X2 U4387 ( .A(n3150), .ZN(n4443) );
  AOI21_X1 U4388 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6937), .A(n4443), 
        .ZN(n3389) );
  NAND2_X1 U4389 ( .A1(n3987), .A2(EAX_REG_29__SCAN_IN), .ZN(n3388) );
  OAI211_X1 U4390 ( .C1(n3390), .C2(n4061), .A(n3389), .B(n3388), .ZN(n3391)
         );
  OAI21_X1 U4391 ( .B1(n3150), .B2(n5689), .A(n3391), .ZN(n4072) );
  AOI22_X1 U4392 ( .A1(n3471), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3396) );
  AOI22_X1 U4393 ( .A1(n3404), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3395) );
  AOI22_X1 U4394 ( .A1(n3477), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4001), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3394) );
  AOI22_X1 U4395 ( .A1(n3460), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3393) );
  NAND4_X1 U4396 ( .A1(n3396), .A2(n3395), .A3(n3394), .A4(n3393), .ZN(n3402)
         );
  AOI22_X1 U4397 ( .A1(n4428), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        INSTQUEUE_REG_10__3__SCAN_IN), .B2(n3560), .ZN(n3400) );
  AOI22_X1 U4398 ( .A1(n3476), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3478), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3399) );
  AOI22_X1 U4399 ( .A1(n3453), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3143), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3398) );
  AOI22_X1 U4400 ( .A1(n3469), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3136), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3397) );
  NAND4_X1 U4401 ( .A1(n3400), .A2(n3399), .A3(n3398), .A4(n3397), .ZN(n3401)
         );
  OAI21_X1 U4402 ( .B1(n3489), .B2(n3510), .A(n3493), .ZN(n3424) );
  NAND2_X1 U4403 ( .A1(n3461), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3408)
         );
  INV_X1 U4404 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3403) );
  OR2_X1 U4405 ( .A1(n3455), .A2(n3403), .ZN(n3407) );
  NAND2_X1 U4406 ( .A1(n3470), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3406) );
  NAND2_X1 U4407 ( .A1(n3404), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3405)
         );
  NAND2_X1 U4408 ( .A1(n3460), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3412) );
  NAND2_X1 U4409 ( .A1(n3471), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3411) );
  NAND2_X1 U4410 ( .A1(n3469), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3410) );
  NAND2_X1 U4411 ( .A1(n3561), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3409)
         );
  NAND2_X1 U4412 ( .A1(n3560), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3416)
         );
  NAND2_X1 U4413 ( .A1(n3453), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3415) );
  NAND2_X1 U4414 ( .A1(n3478), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3414) );
  NAND2_X1 U4415 ( .A1(n4001), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3413) );
  NAND2_X1 U4416 ( .A1(n3476), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3420) );
  NAND2_X1 U4417 ( .A1(n3477), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3419)
         );
  NAND2_X1 U4418 ( .A1(n3136), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3418) );
  NAND2_X1 U4419 ( .A1(n3143), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3417)
         );
  NAND2_X1 U4420 ( .A1(n3424), .A2(n4599), .ZN(n3427) );
  INV_X1 U4421 ( .A(n4599), .ZN(n4368) );
  NAND4_X1 U4422 ( .A1(n3425), .A2(n3489), .A3(n3496), .A4(n4368), .ZN(n3426)
         );
  NAND2_X1 U4423 ( .A1(n3427), .A2(n3426), .ZN(n3428) );
  NAND2_X1 U4424 ( .A1(n3477), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3433)
         );
  NAND2_X1 U4425 ( .A1(n3453), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3432) );
  NAND2_X1 U4426 ( .A1(n3478), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3431) );
  NAND2_X1 U4427 ( .A1(n3143), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3430)
         );
  NAND2_X1 U4428 ( .A1(n3471), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3440) );
  NAND2_X1 U4429 ( .A1(n3461), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3439)
         );
  INV_X1 U4430 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3434) );
  INV_X1 U4431 ( .A(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3435) );
  NAND2_X1 U4432 ( .A1(n3560), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3444)
         );
  NAND2_X1 U4433 ( .A1(n3462), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3443) );
  NAND2_X1 U4434 ( .A1(n4001), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3442) );
  NAND2_X1 U4435 ( .A1(n3476), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3441) );
  NAND2_X1 U4436 ( .A1(n3460), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3448) );
  NAND2_X1 U4437 ( .A1(n3470), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3447) );
  NAND2_X1 U4438 ( .A1(n3561), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3445)
         );
  NAND4_X4 U4439 ( .A1(n3452), .A2(n3451), .A3(n3450), .A4(n3449), .ZN(n3492)
         );
  NAND2_X1 U4440 ( .A1(n4352), .A2(n4585), .ZN(n3529) );
  NAND2_X1 U4441 ( .A1(n3453), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3459) );
  NAND2_X1 U4442 ( .A1(n3560), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3458)
         );
  INV_X1 U4443 ( .A(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3454) );
  OR2_X1 U4444 ( .A1(n3455), .A2(n3454), .ZN(n3457) );
  NAND2_X1 U4445 ( .A1(n3143), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3456)
         );
  NAND2_X1 U4446 ( .A1(n3460), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3466) );
  NAND2_X1 U4447 ( .A1(n3461), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3465)
         );
  NAND2_X1 U4448 ( .A1(n3462), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3464) );
  NAND2_X1 U4449 ( .A1(n3561), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3463)
         );
  NAND2_X1 U4450 ( .A1(n3469), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3474) );
  NAND2_X1 U4451 ( .A1(n3470), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3473) );
  NAND2_X1 U4452 ( .A1(n3471), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3472) );
  NAND2_X1 U4453 ( .A1(n3476), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3482) );
  NAND2_X1 U4454 ( .A1(n4001), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3481) );
  NAND2_X1 U4455 ( .A1(n3477), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3480)
         );
  NAND2_X1 U4456 ( .A1(n3478), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3479) );
  INV_X1 U4457 ( .A(n3674), .ZN(n3486) );
  NAND2_X1 U4458 ( .A1(n3529), .A2(n3486), .ZN(n3505) );
  NOR2_X1 U4459 ( .A1(n5400), .A2(n3492), .ZN(n3491) );
  AND2_X4 U4460 ( .A1(n3493), .A2(n3492), .ZN(n4090) );
  INV_X1 U4461 ( .A(n3528), .ZN(n3494) );
  NAND2_X1 U4462 ( .A1(n3494), .A2(n4656), .ZN(n4084) );
  INV_X1 U4463 ( .A(n3536), .ZN(n3501) );
  NAND2_X1 U4464 ( .A1(n3501), .A2(n3489), .ZN(n3498) );
  AND2_X1 U4465 ( .A1(n3496), .A2(n3488), .ZN(n3497) );
  INV_X1 U4466 ( .A(n3493), .ZN(n5455) );
  NAND2_X1 U4467 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6694) );
  OAI21_X1 U4468 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .A(
        n6694), .ZN(n4360) );
  NAND2_X1 U4469 ( .A1(n4585), .A2(n4360), .ZN(n3508) );
  AOI21_X1 U4470 ( .B1(n5455), .B2(n3508), .A(n4354), .ZN(n3499) );
  NAND3_X1 U4471 ( .A1(n3534), .A2(n4073), .A3(n3499), .ZN(n3503) );
  NAND2_X1 U4472 ( .A1(n3632), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3518) );
  NOR2_X1 U4473 ( .A1(n4354), .A2(n3493), .ZN(n3506) );
  OR2_X2 U4474 ( .A1(n4372), .A2(n5400), .ZN(n6641) );
  INV_X1 U4475 ( .A(n3508), .ZN(n3514) );
  NOR2_X1 U4476 ( .A1(n4656), .A2(n3493), .ZN(n3509) );
  AND2_X1 U4477 ( .A1(n4599), .A2(n3509), .ZN(n4151) );
  NAND2_X1 U4478 ( .A1(n5606), .A2(n4151), .ZN(n4087) );
  INV_X1 U4479 ( .A(n4087), .ZN(n3512) );
  NAND2_X1 U4480 ( .A1(n3510), .A2(n3488), .ZN(n4373) );
  NAND2_X1 U4481 ( .A1(n3512), .A2(n3511), .ZN(n4381) );
  NAND2_X1 U4482 ( .A1(n3493), .A2(n3489), .ZN(n4105) );
  NOR2_X1 U4483 ( .A1(n4522), .A2(n4105), .ZN(n3513) );
  NAND2_X1 U4484 ( .A1(n3519), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3517) );
  INV_X1 U4485 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n3515) );
  NAND2_X1 U4486 ( .A1(n3515), .A2(n5389), .ZN(n6763) );
  XNOR2_X1 U4487 ( .A(n6556), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6424)
         );
  AND2_X1 U4488 ( .A1(n3636), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3516)
         );
  AOI21_X1 U4489 ( .B1(n3637), .B2(n6424), .A(n3516), .ZN(n3520) );
  NAND3_X1 U4490 ( .A1(n3518), .A2(n3517), .A3(n3520), .ZN(n3630) );
  INV_X1 U4491 ( .A(n3520), .ZN(n3521) );
  NAND2_X1 U4492 ( .A1(n3130), .A2(n3523), .ZN(n3524) );
  AND2_X2 U4493 ( .A1(n3630), .A2(n3524), .ZN(n3629) );
  NAND2_X1 U4494 ( .A1(n3632), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3527) );
  MUX2_X1 U4495 ( .A(n3636), .B(n3637), .S(n6556), .Z(n3525) );
  INV_X1 U4496 ( .A(n3525), .ZN(n3526) );
  NAND2_X1 U4497 ( .A1(n3243), .A2(n3530), .ZN(n4083) );
  INV_X1 U4498 ( .A(n6763), .ZN(n6050) );
  OAI211_X1 U4499 ( .C1(n4085), .C2(n3425), .A(STATE2_REG_0__SCAN_IN), .B(
        n6050), .ZN(n3533) );
  INV_X1 U4500 ( .A(n3533), .ZN(n3542) );
  INV_X1 U4501 ( .A(n4073), .ZN(n3539) );
  NAND2_X1 U4502 ( .A1(n3536), .A2(n3487), .ZN(n3537) );
  NAND2_X1 U4503 ( .A1(n3537), .A2(n4656), .ZN(n3538) );
  OAI21_X1 U4504 ( .B1(n3539), .B2(n3538), .A(n3492), .ZN(n3540) );
  XNOR2_X2 U4505 ( .A(n3629), .B(n3628), .ZN(n4486) );
  AOI22_X1 U4506 ( .A1(n3137), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4423), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3547) );
  AOI22_X1 U4507 ( .A1(n4015), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4421), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3546) );
  AOI22_X1 U4508 ( .A1(n4429), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3257), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3545) );
  AOI22_X1 U4509 ( .A1(n3975), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3544) );
  NAND4_X1 U4510 ( .A1(n3547), .A2(n3546), .A3(n3545), .A4(n3544), .ZN(n3553)
         );
  AOI22_X1 U4511 ( .A1(n3471), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3551) );
  AOI22_X1 U4512 ( .A1(n3996), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4610), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3550) );
  AOI22_X1 U4513 ( .A1(n4422), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3549) );
  BUF_X1 U4514 ( .A(n3561), .Z(n3584) );
  AOI22_X1 U4515 ( .A1(n3460), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3584), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3548) );
  NAND4_X1 U4516 ( .A1(n3551), .A2(n3550), .A3(n3549), .A4(n3548), .ZN(n3552)
         );
  NOR2_X1 U4517 ( .A1(n4147), .A2(n3568), .ZN(n3554) );
  INV_X1 U4518 ( .A(n3574), .ZN(n3572) );
  INV_X1 U4519 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5260) );
  OR2_X1 U4520 ( .A1(n3555), .A2(n5260), .ZN(n3570) );
  AOI22_X1 U4521 ( .A1(n3996), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3476), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3559) );
  AOI22_X1 U4522 ( .A1(n3453), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3558) );
  AOI22_X1 U4523 ( .A1(n4431), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4421), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3557) );
  AOI22_X1 U4524 ( .A1(n3470), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3257), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3556) );
  NAND4_X1 U4525 ( .A1(n3559), .A2(n3558), .A3(n3557), .A4(n3556), .ZN(n3567)
         );
  AOI22_X1 U4526 ( .A1(n4610), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3565) );
  AOI22_X1 U4527 ( .A1(n3137), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4422), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3564) );
  AOI22_X1 U4528 ( .A1(n4015), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3563) );
  AOI22_X1 U4529 ( .A1(n3471), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3562) );
  NAND4_X1 U4530 ( .A1(n3565), .A2(n3564), .A3(n3563), .A4(n3562), .ZN(n3566)
         );
  OR2_X1 U4531 ( .A1(n3568), .A2(n3674), .ZN(n3569) );
  INV_X1 U4532 ( .A(n3573), .ZN(n3571) );
  NAND2_X1 U4533 ( .A1(n3572), .A2(n3571), .ZN(n3575) );
  NAND2_X1 U4534 ( .A1(n3574), .A2(n3573), .ZN(n3626) );
  NAND2_X1 U4535 ( .A1(n3575), .A2(n3626), .ZN(n3603) );
  INV_X1 U4536 ( .A(n3603), .ZN(n3602) );
  NAND2_X1 U4537 ( .A1(n3617), .A2(n6872), .ZN(n3594) );
  INV_X1 U4538 ( .A(n3579), .ZN(n3592) );
  NOR2_X1 U4539 ( .A1(n4147), .A2(n3759), .ZN(n3600) );
  AOI22_X1 U4540 ( .A1(n3975), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3453), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3583) );
  AOI22_X1 U4541 ( .A1(n3471), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4421), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3582) );
  AOI22_X1 U4542 ( .A1(n3996), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3581) );
  AOI22_X1 U4543 ( .A1(n4015), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3580) );
  NAND4_X1 U4544 ( .A1(n3583), .A2(n3582), .A3(n3581), .A4(n3580), .ZN(n3590)
         );
  AOI22_X1 U4545 ( .A1(n3137), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3588) );
  AOI22_X1 U4546 ( .A1(n4429), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3257), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3587) );
  AOI22_X1 U4547 ( .A1(n4610), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4422), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3586) );
  AOI22_X1 U4548 ( .A1(n4431), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3584), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3585) );
  NAND4_X1 U4549 ( .A1(n3588), .A2(n3587), .A3(n3586), .A4(n3585), .ZN(n3589)
         );
  INV_X1 U4550 ( .A(n4254), .ZN(n3591) );
  MUX2_X1 U4551 ( .A(n3592), .B(n3600), .S(n3591), .Z(n3593) );
  INV_X1 U4552 ( .A(n3593), .ZN(n3613) );
  NAND2_X1 U4553 ( .A1(n3594), .A2(n3613), .ZN(n3599) );
  INV_X1 U4554 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n6902) );
  OR2_X1 U4555 ( .A1(n3555), .A2(n6902), .ZN(n3598) );
  NAND2_X1 U4556 ( .A1(n4848), .A2(n4319), .ZN(n3596) );
  NAND2_X1 U4557 ( .A1(n5400), .A2(n4254), .ZN(n3595) );
  NAND2_X1 U4558 ( .A1(n3598), .A2(n3597), .ZN(n3611) );
  INV_X1 U4559 ( .A(n3600), .ZN(n4317) );
  INV_X1 U4560 ( .A(n3604), .ZN(n3601) );
  NAND2_X1 U4561 ( .A1(n3603), .A2(n3604), .ZN(n3605) );
  NAND2_X1 U4562 ( .A1(n4573), .A2(n3893), .ZN(n3610) );
  NAND2_X1 U4563 ( .A1(n3511), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3710) );
  NAND2_X1 U4564 ( .A1(n3987), .A2(EAX_REG_1__SCAN_IN), .ZN(n3607) );
  NAND2_X1 U4565 ( .A1(n6937), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3606)
         );
  OAI211_X1 U4566 ( .C1(n3710), .C2(n3166), .A(n3607), .B(n3606), .ZN(n3608)
         );
  INV_X1 U4567 ( .A(n3608), .ZN(n3609) );
  INV_X1 U4568 ( .A(n3611), .ZN(n3612) );
  INV_X1 U4569 ( .A(n3425), .ZN(n3616) );
  AOI21_X1 U4570 ( .B1(n4578), .B2(n3616), .A(n6937), .ZN(n4475) );
  NAND2_X1 U4571 ( .A1(n3133), .A2(n3893), .ZN(n3623) );
  INV_X2 U4572 ( .A(n3244), .ZN(n3987) );
  NAND2_X1 U4573 ( .A1(n3987), .A2(EAX_REG_0__SCAN_IN), .ZN(n3620) );
  NAND2_X1 U4574 ( .A1(n6937), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n3619)
         );
  OAI211_X1 U4575 ( .C1(n3710), .C2(n3618), .A(n3620), .B(n3619), .ZN(n3621)
         );
  INV_X1 U4576 ( .A(n3621), .ZN(n3622) );
  NAND2_X1 U4577 ( .A1(n3623), .A2(n3622), .ZN(n4474) );
  NAND2_X1 U4578 ( .A1(n4475), .A2(n4474), .ZN(n4473) );
  INV_X1 U4579 ( .A(n4474), .ZN(n3624) );
  NAND2_X1 U4580 ( .A1(n3624), .A2(n4443), .ZN(n3625) );
  NAND2_X1 U4581 ( .A1(n4473), .A2(n3625), .ZN(n4537) );
  INV_X1 U4582 ( .A(n3660), .ZN(n3656) );
  NAND2_X1 U4583 ( .A1(n3629), .A2(n3628), .ZN(n3631) );
  NAND2_X1 U4584 ( .A1(n3632), .A2(n6925), .ZN(n3639) );
  AND2_X1 U4585 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3633) );
  NAND2_X1 U4586 ( .A1(n3633), .A2(n6631), .ZN(n6512) );
  INV_X1 U4587 ( .A(n3633), .ZN(n3634) );
  NAND2_X1 U4588 ( .A1(n3634), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3635) );
  NAND2_X1 U4589 ( .A1(n6512), .A2(n3635), .ZN(n4583) );
  AOI22_X1 U4590 ( .A1(n3637), .A2(n4583), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3636), .ZN(n3638) );
  XNOR2_X2 U4591 ( .A(n3667), .B(n3668), .ZN(n4499) );
  AOI22_X1 U4592 ( .A1(n3137), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4015), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3643) );
  INV_X1 U4593 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n6924) );
  AOI22_X1 U4594 ( .A1(n3975), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4610), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3642) );
  AOI22_X1 U4595 ( .A1(n3996), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3641) );
  AOI22_X1 U4596 ( .A1(n4423), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4422), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3640) );
  NAND4_X1 U4597 ( .A1(n3643), .A2(n3642), .A3(n3641), .A4(n3640), .ZN(n3650)
         );
  AOI22_X1 U4598 ( .A1(n3471), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4421), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3648) );
  AOI22_X1 U4599 ( .A1(n4429), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3257), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3647) );
  AOI22_X1 U4600 ( .A1(n3644), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3646) );
  AOI22_X1 U4601 ( .A1(n4431), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3584), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3645) );
  NAND4_X1 U4602 ( .A1(n3648), .A2(n3647), .A3(n3646), .A4(n3645), .ZN(n3649)
         );
  NOR2_X1 U4603 ( .A1(n4147), .A2(n4264), .ZN(n3651) );
  INV_X1 U4604 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5242) );
  OAI22_X1 U4605 ( .A1(n3555), .A2(n5242), .B1(n4264), .B2(n3674), .ZN(n3652)
         );
  XNOR2_X1 U4606 ( .A(n3665), .B(n3664), .ZN(n4571) );
  NAND2_X1 U4607 ( .A1(n4571), .A2(n3893), .ZN(n3654) );
  NAND2_X1 U4608 ( .A1(n6937), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3915) );
  INV_X1 U4611 ( .A(n6925), .ZN(n4515) );
  INV_X1 U4612 ( .A(n3691), .ZN(n3657) );
  OAI21_X1 U4613 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3657), .ZN(n6360) );
  AOI22_X1 U4614 ( .A1(n4443), .A2(n6360), .B1(n4447), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3659) );
  NAND2_X1 U4615 ( .A1(n3987), .A2(EAX_REG_2__SCAN_IN), .ZN(n3658) );
  OAI211_X1 U4616 ( .C1(n3710), .C2(n4515), .A(n3659), .B(n3658), .ZN(n4518)
         );
  NAND2_X1 U4617 ( .A1(n3127), .A2(n3660), .ZN(n3662) );
  INV_X1 U4618 ( .A(n3664), .ZN(n3666) );
  NOR2_X2 U4619 ( .A1(n3666), .A2(n3665), .ZN(n3688) );
  INV_X1 U4620 ( .A(n3667), .ZN(n3669) );
  NAND2_X1 U4621 ( .A1(n3632), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3673) );
  NAND3_X1 U4622 ( .A1(n7081), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6473) );
  INV_X1 U4623 ( .A(n6473), .ZN(n6471) );
  NAND2_X1 U4624 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6471), .ZN(n6472) );
  NAND2_X1 U4625 ( .A1(n7081), .A2(n6472), .ZN(n3670) );
  NOR3_X1 U4626 ( .A1(n7081), .A2(n6631), .A3(n7064), .ZN(n4955) );
  NAND2_X1 U4627 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4955), .ZN(n4998) );
  NAND2_X1 U4628 ( .A1(n3670), .A2(n4998), .ZN(n4718) );
  OAI22_X1 U4629 ( .A1(n4450), .A2(n4718), .B1(n4149), .B2(n7081), .ZN(n3671)
         );
  INV_X1 U4630 ( .A(n3671), .ZN(n3672) );
  XNOR2_X2 U4631 ( .A(n4625), .B(n4717), .ZN(n5074) );
  AOI22_X1 U4632 ( .A1(n3137), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4015), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3678) );
  AOI22_X1 U4633 ( .A1(n3975), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4610), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3677) );
  AOI22_X1 U4634 ( .A1(n3996), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3676) );
  AOI22_X1 U4635 ( .A1(n4423), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4422), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3675) );
  NAND4_X1 U4636 ( .A1(n3678), .A2(n3677), .A3(n3676), .A4(n3675), .ZN(n3685)
         );
  AOI22_X1 U4637 ( .A1(n3132), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4421), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3683) );
  AOI22_X1 U4638 ( .A1(n4429), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3257), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3682) );
  AOI22_X1 U4639 ( .A1(n3644), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3681) );
  AOI22_X1 U4640 ( .A1(n4431), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3584), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3680) );
  NAND4_X1 U4641 ( .A1(n3683), .A2(n3682), .A3(n3681), .A4(n3680), .ZN(n3684)
         );
  AOI22_X1 U4642 ( .A1(n4129), .A2(n4274), .B1(INSTQUEUE_REG_0__3__SCAN_IN), 
        .B2(n4136), .ZN(n3686) );
  OAI21_X1 U4643 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3691), .A(n3711), 
        .ZN(n6194) );
  AOI22_X1 U4644 ( .A1(n4443), .A2(n6194), .B1(n4447), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3693) );
  NAND2_X1 U4645 ( .A1(n3987), .A2(EAX_REG_3__SCAN_IN), .ZN(n3692) );
  OAI211_X1 U4646 ( .C1(n3710), .C2(n3690), .A(n3693), .B(n3692), .ZN(n3694)
         );
  INV_X1 U4647 ( .A(n3694), .ZN(n3695) );
  AOI22_X1 U4648 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n3137), .B1(n4423), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3699) );
  AOI22_X1 U4649 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n3132), .B1(n4429), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3698) );
  AOI22_X1 U4650 ( .A1(n3975), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4422), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3697) );
  AOI22_X1 U4651 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n4015), .B1(n4430), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3696) );
  NAND4_X1 U4652 ( .A1(n3699), .A2(n3698), .A3(n3697), .A4(n3696), .ZN(n3705)
         );
  AOI22_X1 U4653 ( .A1(n3644), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4610), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3703) );
  AOI22_X1 U4654 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n4421), .B1(n3257), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3702) );
  AOI22_X1 U4655 ( .A1(n3996), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3701) );
  AOI22_X1 U4656 ( .A1(n4431), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3584), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3700) );
  NAND4_X1 U4657 ( .A1(n3703), .A2(n3702), .A3(n3701), .A4(n3700), .ZN(n3704)
         );
  INV_X1 U4658 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5246) );
  OR2_X1 U4659 ( .A1(n3555), .A2(n5246), .ZN(n3706) );
  NAND2_X1 U4660 ( .A1(n3987), .A2(EAX_REG_4__SCAN_IN), .ZN(n3709) );
  INV_X1 U4661 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6064) );
  OAI21_X1 U4662 ( .B1(n6064), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6937), 
        .ZN(n3708) );
  OAI211_X1 U4663 ( .C1(n3710), .C2(n4627), .A(n3709), .B(n3708), .ZN(n3713)
         );
  AOI21_X1 U4664 ( .B1(n6180), .B2(n3711), .A(n3734), .ZN(n6177) );
  NAND2_X1 U4665 ( .A1(n6177), .A2(n4443), .ZN(n3712) );
  AND2_X1 U4666 ( .A1(n3713), .A2(n3712), .ZN(n3714) );
  AOI21_X1 U4667 ( .B1(n4280), .B2(n3893), .A(n3714), .ZN(n4556) );
  AOI22_X1 U4668 ( .A1(n3137), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4015), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3720) );
  AOI22_X1 U4669 ( .A1(n3975), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4610), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3719) );
  AOI22_X1 U4670 ( .A1(n3996), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3718) );
  AOI22_X1 U4671 ( .A1(n4423), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4422), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3717) );
  NAND4_X1 U4672 ( .A1(n3720), .A2(n3719), .A3(n3718), .A4(n3717), .ZN(n3726)
         );
  AOI22_X1 U4673 ( .A1(n3471), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4421), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3724) );
  AOI22_X1 U4674 ( .A1(n4429), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3257), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3723) );
  AOI22_X1 U4675 ( .A1(n3644), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3722) );
  AOI22_X1 U4676 ( .A1(n4431), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3584), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3721) );
  NAND4_X1 U4677 ( .A1(n3724), .A2(n3723), .A3(n3722), .A4(n3721), .ZN(n3725)
         );
  INV_X1 U4678 ( .A(n4291), .ZN(n3727) );
  INV_X1 U4679 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5231) );
  OR2_X1 U4680 ( .A1(n3555), .A2(n5231), .ZN(n3728) );
  NAND2_X1 U4681 ( .A1(n3732), .A2(n3731), .ZN(n3733) );
  NAND2_X1 U4682 ( .A1(n3756), .A2(n3733), .ZN(n4294) );
  OAI21_X1 U4683 ( .B1(PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n3734), .A(n3750), 
        .ZN(n6176) );
  AOI22_X1 U4684 ( .A1(n4443), .A2(n6176), .B1(n4447), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3736) );
  NAND2_X1 U4685 ( .A1(n3987), .A2(EAX_REG_5__SCAN_IN), .ZN(n3735) );
  NAND2_X1 U4686 ( .A1(n3126), .A2(n3124), .ZN(n4551) );
  INV_X1 U4687 ( .A(n4551), .ZN(n3755) );
  AOI22_X1 U4688 ( .A1(n3137), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3740) );
  AOI22_X1 U4689 ( .A1(n3920), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4421), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3739) );
  AOI22_X1 U4690 ( .A1(n3644), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3738) );
  AOI22_X1 U4691 ( .A1(n4431), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3584), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3737) );
  NAND4_X1 U4692 ( .A1(n3740), .A2(n3739), .A3(n3738), .A4(n3737), .ZN(n3746)
         );
  AOI22_X1 U4693 ( .A1(n4423), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4015), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3744) );
  AOI22_X1 U4694 ( .A1(n4429), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3257), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3743) );
  AOI22_X1 U4695 ( .A1(n3996), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3742) );
  AOI22_X1 U4696 ( .A1(n4610), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4422), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3741) );
  NAND4_X1 U4697 ( .A1(n3744), .A2(n3743), .A3(n3742), .A4(n3741), .ZN(n3745)
         );
  INV_X1 U4698 ( .A(n4307), .ZN(n3747) );
  OR2_X1 U4699 ( .A1(n4138), .A2(n3747), .ZN(n3749) );
  INV_X1 U4700 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5253) );
  OR2_X1 U4701 ( .A1(n3555), .A2(n5253), .ZN(n3748) );
  NAND2_X1 U4702 ( .A1(n3756), .A2(n3757), .ZN(n4298) );
  NAND2_X1 U4703 ( .A1(n3987), .A2(EAX_REG_6__SCAN_IN), .ZN(n3752) );
  OAI21_X1 U4704 ( .B1(n6064), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6937), 
        .ZN(n3751) );
  XNOR2_X1 U4705 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .B(n3750), .ZN(n6154) );
  AOI22_X1 U4706 ( .A1(n3752), .A2(n3751), .B1(n4443), .B2(n6154), .ZN(n3753)
         );
  INV_X1 U4707 ( .A(n4678), .ZN(n3754) );
  NAND2_X1 U4708 ( .A1(n3755), .A2(n3754), .ZN(n4677) );
  INV_X1 U4709 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5235) );
  XNOR2_X1 U4710 ( .A(n4316), .B(n3760), .ZN(n4305) );
  INV_X1 U4711 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3763) );
  OAI21_X1 U4712 ( .B1(PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n3761), .A(n3768), 
        .ZN(n6140) );
  AOI22_X1 U4713 ( .A1(n4443), .A2(n6140), .B1(n4447), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3762) );
  OAI21_X1 U4714 ( .B1(n3244), .B2(n3763), .A(n3762), .ZN(n3764) );
  NAND2_X1 U4715 ( .A1(n3767), .A2(n4798), .ZN(n4796) );
  AOI21_X1 U4716 ( .B1(n6889), .B2(n3768), .A(n3784), .ZN(n5592) );
  OR2_X1 U4717 ( .A1(n5592), .A2(n3150), .ZN(n3783) );
  NAND2_X1 U4718 ( .A1(n3987), .A2(EAX_REG_8__SCAN_IN), .ZN(n3781) );
  AOI22_X1 U4719 ( .A1(n3137), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4423), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3772) );
  AOI22_X1 U4720 ( .A1(n4429), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3257), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3771) );
  AOI22_X1 U4721 ( .A1(n3975), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4422), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3770) );
  AOI22_X1 U4722 ( .A1(n4430), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3584), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3769) );
  NAND4_X1 U4723 ( .A1(n3772), .A2(n3771), .A3(n3770), .A4(n3769), .ZN(n3778)
         );
  AOI22_X1 U4724 ( .A1(n3644), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3776) );
  AOI22_X1 U4725 ( .A1(n3920), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4421), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3775) );
  AOI22_X1 U4726 ( .A1(n4015), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4610), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3774) );
  AOI22_X1 U4727 ( .A1(n3996), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3773) );
  NAND4_X1 U4728 ( .A1(n3776), .A2(n3775), .A3(n3774), .A4(n3773), .ZN(n3777)
         );
  OAI21_X1 U4729 ( .B1(n3778), .B2(n3777), .A(n3893), .ZN(n3780) );
  NAND2_X1 U4730 ( .A1(n4447), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3779)
         );
  AND3_X1 U4731 ( .A1(n3781), .A2(n3780), .A3(n3779), .ZN(n3782) );
  INV_X1 U4732 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6128) );
  XNOR2_X1 U4733 ( .A(n3784), .B(n6128), .ZN(n6134) );
  OR2_X1 U4734 ( .A1(n6134), .A2(n3150), .ZN(n3799) );
  AOI22_X1 U4735 ( .A1(n4431), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3257), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3788) );
  AOI22_X1 U4736 ( .A1(n3996), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4422), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4737 ( .A1(n4015), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3786) );
  AOI22_X1 U4738 ( .A1(n3644), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3584), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3785) );
  NAND4_X1 U4739 ( .A1(n3788), .A2(n3787), .A3(n3786), .A4(n3785), .ZN(n3794)
         );
  AOI22_X1 U4740 ( .A1(n3137), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4741 ( .A1(n4421), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4429), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3791) );
  AOI22_X1 U4742 ( .A1(n4423), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4610), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3790) );
  AOI22_X1 U4743 ( .A1(n3975), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3789) );
  NAND4_X1 U4744 ( .A1(n3792), .A2(n3791), .A3(n3790), .A4(n3789), .ZN(n3793)
         );
  OAI21_X1 U4745 ( .B1(n3794), .B2(n3793), .A(n3893), .ZN(n3796) );
  NAND2_X1 U4746 ( .A1(n3987), .A2(EAX_REG_9__SCAN_IN), .ZN(n3795) );
  OAI211_X1 U4747 ( .C1(n3915), .C2(n6128), .A(n3796), .B(n3795), .ZN(n3797)
         );
  INV_X1 U4748 ( .A(n3797), .ZN(n3798) );
  NAND2_X1 U4749 ( .A1(n3799), .A2(n3798), .ZN(n4979) );
  XOR2_X1 U4750 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3800), .Z(n5310) );
  AOI22_X1 U4751 ( .A1(n3137), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3644), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3804) );
  AOI22_X1 U4752 ( .A1(n3920), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3803) );
  AOI22_X1 U4753 ( .A1(n4421), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4429), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3802) );
  AOI22_X1 U4754 ( .A1(n4610), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4422), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3801) );
  NAND4_X1 U4755 ( .A1(n3804), .A2(n3803), .A3(n3802), .A4(n3801), .ZN(n3810)
         );
  AOI22_X1 U4756 ( .A1(n3975), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4423), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3808) );
  AOI22_X1 U4757 ( .A1(n3996), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4758 ( .A1(n4015), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4759 ( .A1(n3257), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3584), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3805) );
  NAND4_X1 U4760 ( .A1(n3808), .A2(n3807), .A3(n3806), .A4(n3805), .ZN(n3809)
         );
  OR2_X1 U4761 ( .A1(n3810), .A2(n3809), .ZN(n3811) );
  AOI22_X1 U4762 ( .A1(n3893), .A2(n3811), .B1(n4447), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3813) );
  NAND2_X1 U4763 ( .A1(n3987), .A2(EAX_REG_10__SCAN_IN), .ZN(n3812) );
  OAI211_X1 U4764 ( .C1(n5310), .C2(n3150), .A(n3813), .B(n3812), .ZN(n5215)
         );
  XNOR2_X1 U4765 ( .A(n3814), .B(n3827), .ZN(n5582) );
  NAND2_X1 U4766 ( .A1(n5582), .A2(n4443), .ZN(n3830) );
  AOI22_X1 U4767 ( .A1(n3975), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4423), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3818) );
  AOI22_X1 U4768 ( .A1(n3137), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4015), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3817) );
  AOI22_X1 U4769 ( .A1(n3920), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3257), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3816) );
  AOI22_X1 U4770 ( .A1(n4430), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3584), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3815) );
  NAND4_X1 U4771 ( .A1(n3818), .A2(n3817), .A3(n3816), .A4(n3815), .ZN(n3824)
         );
  AOI22_X1 U4772 ( .A1(n3644), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4773 ( .A1(n4421), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4429), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4774 ( .A1(n3996), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3820) );
  AOI22_X1 U4775 ( .A1(n4610), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4422), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3819) );
  NAND4_X1 U4776 ( .A1(n3822), .A2(n3821), .A3(n3820), .A4(n3819), .ZN(n3823)
         );
  OAI21_X1 U4777 ( .B1(n3824), .B2(n3823), .A(n3893), .ZN(n3826) );
  NAND2_X1 U4778 ( .A1(n3987), .A2(EAX_REG_11__SCAN_IN), .ZN(n3825) );
  OAI211_X1 U4779 ( .C1(n3915), .C2(n3827), .A(n3826), .B(n3825), .ZN(n3828)
         );
  INV_X1 U4780 ( .A(n3828), .ZN(n3829) );
  NAND2_X1 U4781 ( .A1(n3830), .A2(n3829), .ZN(n5272) );
  XOR2_X1 U4782 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3831), .Z(n6109) );
  NAND2_X1 U4783 ( .A1(n6109), .A2(n4443), .ZN(n3846) );
  INV_X1 U4784 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5317) );
  OAI21_X1 U4785 ( .B1(PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n6064), .A(n6937), 
        .ZN(n3832) );
  OAI21_X1 U4786 ( .B1(n3244), .B2(n5317), .A(n3832), .ZN(n3845) );
  AOI22_X1 U4787 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n3920), .B1(n3644), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3836) );
  AOI22_X1 U4788 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n4421), .B1(n4429), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3835) );
  AOI22_X1 U4789 ( .A1(n3996), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4610), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3834) );
  AOI22_X1 U4790 ( .A1(n3137), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4422), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3833) );
  NAND4_X1 U4791 ( .A1(n3836), .A2(n3835), .A3(n3834), .A4(n3833), .ZN(n3842)
         );
  AOI22_X1 U4792 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n4423), .B1(n4015), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4793 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n4431), .B1(n3257), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3839) );
  AOI22_X1 U4794 ( .A1(n3975), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3838) );
  AOI22_X1 U4795 ( .A1(n4430), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3584), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3837) );
  NAND4_X1 U4796 ( .A1(n3840), .A2(n3839), .A3(n3838), .A4(n3837), .ZN(n3841)
         );
  NOR2_X1 U4797 ( .A1(n3842), .A2(n3841), .ZN(n3843) );
  NOR2_X1 U4798 ( .A1(n3883), .A2(n3843), .ZN(n3844) );
  AOI21_X1 U4799 ( .B1(n3846), .B2(n3845), .A(n3844), .ZN(n5316) );
  NAND2_X1 U4800 ( .A1(n3847), .A2(n3850), .ZN(n3849) );
  INV_X1 U4801 ( .A(n3879), .ZN(n3848) );
  NAND2_X1 U4802 ( .A1(n3849), .A2(n3848), .ZN(n6097) );
  NAND2_X1 U4803 ( .A1(n6097), .A2(n4443), .ZN(n3853) );
  AOI21_X1 U4804 ( .B1(n3987), .B2(EAX_REG_13__SCAN_IN), .A(n3851), .ZN(n3852)
         );
  NAND2_X1 U4805 ( .A1(n3853), .A2(n3852), .ZN(n3866) );
  AOI22_X1 U4806 ( .A1(n3137), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4015), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3857) );
  AOI22_X1 U4807 ( .A1(n3975), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4610), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3856) );
  AOI22_X1 U4808 ( .A1(n3477), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4809 ( .A1(n4423), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4422), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3854) );
  NAND4_X1 U4810 ( .A1(n3857), .A2(n3856), .A3(n3855), .A4(n3854), .ZN(n3863)
         );
  AOI22_X1 U4811 ( .A1(n3920), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4421), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3861) );
  AOI22_X1 U4812 ( .A1(n4429), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3257), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4813 ( .A1(n3644), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4814 ( .A1(n4431), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3858) );
  NAND4_X1 U4815 ( .A1(n3861), .A2(n3860), .A3(n3859), .A4(n3858), .ZN(n3862)
         );
  OR2_X1 U4816 ( .A1(n3863), .A2(n3862), .ZN(n3864) );
  AND2_X1 U4817 ( .A1(n3893), .A2(n3864), .ZN(n5358) );
  NAND2_X1 U4818 ( .A1(n5357), .A2(n5358), .ZN(n3868) );
  AOI22_X1 U4819 ( .A1(n3137), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4015), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3872) );
  AOI22_X1 U4820 ( .A1(n4421), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4429), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3871) );
  AOI22_X1 U4821 ( .A1(n4423), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4422), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3870) );
  AOI22_X1 U4822 ( .A1(n4431), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3584), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3869) );
  NAND4_X1 U4823 ( .A1(n3872), .A2(n3871), .A3(n3870), .A4(n3869), .ZN(n3878)
         );
  AOI22_X1 U4824 ( .A1(n3975), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4610), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3876) );
  AOI22_X1 U4825 ( .A1(n3920), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3257), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3875) );
  AOI22_X1 U4826 ( .A1(n3996), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3874) );
  AOI22_X1 U4827 ( .A1(n3644), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3873) );
  NAND4_X1 U4828 ( .A1(n3876), .A2(n3875), .A3(n3874), .A4(n3873), .ZN(n3877)
         );
  NOR2_X1 U4829 ( .A1(n3878), .A2(n3877), .ZN(n3882) );
  NAND2_X1 U4830 ( .A1(n3987), .A2(EAX_REG_14__SCAN_IN), .ZN(n3881) );
  XNOR2_X1 U4831 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3879), .ZN(n5783)
         );
  AOI22_X1 U4832 ( .A1(n4443), .A2(n5783), .B1(n4447), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3880) );
  OAI211_X1 U4833 ( .C1(n3883), .C2(n3882), .A(n3881), .B(n3880), .ZN(n5355)
         );
  XOR2_X1 U4834 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n3884), .Z(n5777) );
  INV_X1 U4835 ( .A(n5777), .ZN(n3899) );
  INV_X1 U4836 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5774) );
  AOI22_X1 U4837 ( .A1(n3920), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3888) );
  AOI22_X1 U4838 ( .A1(n4421), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4429), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3887) );
  AOI22_X1 U4839 ( .A1(n3137), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4422), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3886) );
  AOI22_X1 U4840 ( .A1(n4430), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3584), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3885) );
  NAND4_X1 U4841 ( .A1(n3888), .A2(n3887), .A3(n3886), .A4(n3885), .ZN(n3895)
         );
  AOI22_X1 U4842 ( .A1(n3975), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4610), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4843 ( .A1(n4423), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4015), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4844 ( .A1(n3644), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3257), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4845 ( .A1(n3996), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3889) );
  NAND4_X1 U4846 ( .A1(n3892), .A2(n3891), .A3(n3890), .A4(n3889), .ZN(n3894)
         );
  OAI21_X1 U4847 ( .B1(n3895), .B2(n3894), .A(n3893), .ZN(n3897) );
  NAND2_X1 U4848 ( .A1(n3987), .A2(EAX_REG_15__SCAN_IN), .ZN(n3896) );
  OAI211_X1 U4849 ( .C1(n3915), .C2(n5774), .A(n3897), .B(n3896), .ZN(n3898)
         );
  AOI21_X1 U4850 ( .B1(n3899), .B2(n4443), .A(n3898), .ZN(n5382) );
  NAND2_X1 U4851 ( .A1(n3902), .A2(n6934), .ZN(n3904) );
  INV_X1 U4852 ( .A(n3935), .ZN(n3903) );
  NAND2_X1 U4853 ( .A1(n3904), .A2(n3903), .ZN(n5769) );
  AOI22_X1 U4854 ( .A1(n3477), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3908) );
  AOI22_X1 U4855 ( .A1(n3137), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3907) );
  AOI22_X1 U4856 ( .A1(n4421), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4429), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3906) );
  AOI22_X1 U4857 ( .A1(n4610), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4422), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3905) );
  NAND4_X1 U4858 ( .A1(n3908), .A2(n3907), .A3(n3906), .A4(n3905), .ZN(n3914)
         );
  AOI22_X1 U4859 ( .A1(n3920), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3257), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4860 ( .A1(n4423), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4861 ( .A1(n4015), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3910) );
  AOI22_X1 U4862 ( .A1(n3644), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3584), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3909) );
  NAND4_X1 U4863 ( .A1(n3912), .A2(n3911), .A3(n3910), .A4(n3909), .ZN(n3913)
         );
  NOR2_X1 U4864 ( .A1(n3914), .A2(n3913), .ZN(n3918) );
  AOI21_X1 U4865 ( .B1(n3987), .B2(EAX_REG_16__SCAN_IN), .A(n3916), .ZN(n3917)
         );
  OAI21_X1 U4866 ( .B1(n4061), .B2(n3918), .A(n3917), .ZN(n3919) );
  AOI21_X1 U4867 ( .B1(n5769), .B2(n4443), .A(n3919), .ZN(n5556) );
  AOI22_X1 U4868 ( .A1(n3996), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3924) );
  AOI22_X1 U4869 ( .A1(n3920), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4421), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3923) );
  AOI22_X1 U4870 ( .A1(n4423), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4422), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3922) );
  AOI22_X1 U4871 ( .A1(n3137), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3584), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3921) );
  NAND4_X1 U4872 ( .A1(n3924), .A2(n3923), .A3(n3922), .A4(n3921), .ZN(n3930)
         );
  AOI22_X1 U4873 ( .A1(n3644), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3928) );
  AOI22_X1 U4874 ( .A1(n4429), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3257), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3927) );
  AOI22_X1 U4875 ( .A1(n4610), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3926) );
  AOI22_X1 U4876 ( .A1(n4015), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3925) );
  NAND4_X1 U4877 ( .A1(n3928), .A2(n3927), .A3(n3926), .A4(n3925), .ZN(n3929)
         );
  NOR2_X1 U4878 ( .A1(n3930), .A2(n3929), .ZN(n3934) );
  OAI21_X1 U4879 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6064), .A(n6937), 
        .ZN(n3931) );
  INV_X1 U4880 ( .A(n3931), .ZN(n3932) );
  AOI21_X1 U4881 ( .B1(n3987), .B2(EAX_REG_17__SCAN_IN), .A(n3932), .ZN(n3933)
         );
  OAI21_X1 U4882 ( .B1(n4061), .B2(n3934), .A(n3933), .ZN(n3937) );
  OAI21_X1 U4883 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n3935), .A(n3951), 
        .ZN(n6092) );
  OR2_X1 U4884 ( .A1(n3150), .A2(n6092), .ZN(n3936) );
  AOI22_X1 U4885 ( .A1(n3137), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4015), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3941) );
  AOI22_X1 U4886 ( .A1(n3975), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4610), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3940) );
  AOI22_X1 U4887 ( .A1(n3477), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3939) );
  AOI22_X1 U4888 ( .A1(n4423), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4422), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3938) );
  NAND4_X1 U4889 ( .A1(n3941), .A2(n3940), .A3(n3939), .A4(n3938), .ZN(n3947)
         );
  AOI22_X1 U4890 ( .A1(n3920), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4421), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3945) );
  AOI22_X1 U4891 ( .A1(n4429), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3257), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3944) );
  AOI22_X1 U4892 ( .A1(n3644), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U4893 ( .A1(n4431), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3584), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3942) );
  NAND4_X1 U4894 ( .A1(n3945), .A2(n3944), .A3(n3943), .A4(n3942), .ZN(n3946)
         );
  NOR2_X1 U4895 ( .A1(n3947), .A2(n3946), .ZN(n3950) );
  AOI21_X1 U4896 ( .B1(n5760), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3948) );
  AOI21_X1 U4897 ( .B1(n3987), .B2(EAX_REG_18__SCAN_IN), .A(n3948), .ZN(n3949)
         );
  OAI21_X1 U4898 ( .B1(n4061), .B2(n3950), .A(n3949), .ZN(n3953) );
  XNOR2_X1 U4899 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n3951), .ZN(n5762)
         );
  NAND2_X1 U4900 ( .A1(n4443), .A2(n5762), .ZN(n3952) );
  NAND2_X1 U4901 ( .A1(n3953), .A2(n3952), .ZN(n5538) );
  AOI22_X1 U4902 ( .A1(n3996), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3476), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3957) );
  AOI22_X1 U4903 ( .A1(n4423), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4015), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3956) );
  AOI22_X1 U4904 ( .A1(n3470), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3257), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U4905 ( .A1(n3644), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3954) );
  NAND4_X1 U4906 ( .A1(n3957), .A2(n3956), .A3(n3955), .A4(n3954), .ZN(n3963)
         );
  AOI22_X1 U4907 ( .A1(n3920), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4421), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3961) );
  AOI22_X1 U4908 ( .A1(n4610), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3960) );
  AOI22_X1 U4909 ( .A1(n3137), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4422), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3959) );
  AOI22_X1 U4910 ( .A1(n4431), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3958) );
  NAND4_X1 U4911 ( .A1(n3961), .A2(n3960), .A3(n3959), .A4(n3958), .ZN(n3962)
         );
  NOR2_X1 U4912 ( .A1(n3963), .A2(n3962), .ZN(n3967) );
  NAND2_X1 U4913 ( .A1(n6937), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3964)
         );
  NAND2_X1 U4914 ( .A1(n3150), .A2(n3964), .ZN(n3965) );
  AOI21_X1 U4915 ( .B1(n3987), .B2(EAX_REG_19__SCAN_IN), .A(n3965), .ZN(n3966)
         );
  OAI21_X1 U4916 ( .B1(n4061), .B2(n3967), .A(n3966), .ZN(n3974) );
  INV_X1 U4917 ( .A(n3990), .ZN(n3972) );
  INV_X1 U4918 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3970) );
  INV_X1 U4919 ( .A(n3968), .ZN(n3969) );
  NAND2_X1 U4920 ( .A1(n3970), .A2(n3969), .ZN(n3971) );
  NAND2_X1 U4921 ( .A1(n3972), .A2(n3971), .ZN(n5993) );
  NAND2_X1 U4922 ( .A1(n3974), .A2(n3973), .ZN(n5663) );
  AOI22_X1 U4923 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n3644), .B1(n4423), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3979) );
  AOI22_X1 U4924 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n3920), .B1(n4429), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U4925 ( .A1(n3996), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U4926 ( .A1(n3975), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4422), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3976) );
  NAND4_X1 U4927 ( .A1(n3979), .A2(n3978), .A3(n3977), .A4(n3976), .ZN(n3985)
         );
  AOI22_X1 U4928 ( .A1(n3137), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4610), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3983) );
  AOI22_X1 U4929 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n4421), .B1(n3257), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3982) );
  AOI22_X1 U4930 ( .A1(n4015), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3981) );
  AOI22_X1 U4931 ( .A1(n4431), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3980) );
  NAND4_X1 U4932 ( .A1(n3983), .A2(n3982), .A3(n3981), .A4(n3980), .ZN(n3984)
         );
  NOR2_X1 U4933 ( .A1(n3985), .A2(n3984), .ZN(n3989) );
  INV_X1 U4934 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5946) );
  OAI21_X1 U4935 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5946), .A(n3150), .ZN(
        n3986) );
  AOI21_X1 U4936 ( .B1(n3987), .B2(EAX_REG_20__SCAN_IN), .A(n3986), .ZN(n3988)
         );
  OAI21_X1 U4937 ( .B1(n4061), .B2(n3989), .A(n3988), .ZN(n3992) );
  XNOR2_X1 U4938 ( .A(n3990), .B(n5946), .ZN(n5938) );
  NAND2_X1 U4939 ( .A1(n5938), .A2(n4443), .ZN(n3991) );
  AND2_X1 U4940 ( .A1(n3994), .A2(n3993), .ZN(n3995) );
  OR2_X1 U4941 ( .A1(n3995), .A2(n4023), .ZN(n5930) );
  INV_X1 U4942 ( .A(EAX_REG_21__SCAN_IN), .ZN(n6950) );
  AOI22_X1 U4943 ( .A1(n3996), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3476), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4000) );
  AOI22_X1 U4944 ( .A1(n4423), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3999) );
  AOI22_X1 U4945 ( .A1(n4610), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4422), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U4946 ( .A1(n4431), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3997) );
  NAND4_X1 U4947 ( .A1(n4000), .A2(n3999), .A3(n3998), .A4(n3997), .ZN(n4007)
         );
  AOI22_X1 U4948 ( .A1(n3920), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4421), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4005) );
  AOI22_X1 U4949 ( .A1(n4429), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3257), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4004) );
  AOI22_X1 U4950 ( .A1(n3137), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4003) );
  AOI22_X1 U4951 ( .A1(n4015), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4002) );
  NAND4_X1 U4952 ( .A1(n4005), .A2(n4004), .A3(n4003), .A4(n4002), .ZN(n4006)
         );
  OAI21_X1 U4953 ( .B1(n4007), .B2(n4006), .A(n4440), .ZN(n4009) );
  OAI21_X1 U4954 ( .B1(PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6064), .A(n6937), 
        .ZN(n4008) );
  OAI211_X1 U4955 ( .C1(n3244), .C2(n6950), .A(n4009), .B(n4008), .ZN(n4010)
         );
  AOI22_X1 U4956 ( .A1(n3137), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4014) );
  AOI22_X1 U4957 ( .A1(n3476), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U4958 ( .A1(n4423), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4422), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4012) );
  AOI22_X1 U4959 ( .A1(n4429), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4011) );
  NAND4_X1 U4960 ( .A1(n4014), .A2(n4013), .A3(n4012), .A4(n4011), .ZN(n4021)
         );
  AOI22_X1 U4961 ( .A1(n3477), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4610), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4019) );
  AOI22_X1 U4962 ( .A1(n3920), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4018) );
  AOI22_X1 U4963 ( .A1(n4421), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3257), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U4964 ( .A1(n4015), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4016) );
  NAND4_X1 U4965 ( .A1(n4019), .A2(n4018), .A3(n4017), .A4(n4016), .ZN(n4020)
         );
  OAI21_X1 U4966 ( .B1(n4021), .B2(n4020), .A(n4440), .ZN(n4025) );
  INV_X1 U4967 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5741) );
  NOR2_X1 U4968 ( .A1(n5741), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4022) );
  AOI211_X1 U4969 ( .C1(n3987), .C2(EAX_REG_22__SCAN_IN), .A(n4443), .B(n4022), 
        .ZN(n4024) );
  XNOR2_X1 U4970 ( .A(n4023), .B(n5741), .ZN(n5920) );
  AOI22_X1 U4971 ( .A1(n4025), .A2(n4024), .B1(n4443), .B2(n5920), .ZN(n5643)
         );
  NOR2_X1 U4972 ( .A1(n4026), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4027)
         );
  OR2_X1 U4973 ( .A1(n4036), .A2(n4027), .ZN(n5918) );
  XNOR2_X1 U4974 ( .A(n4029), .B(n4028), .ZN(n4032) );
  AOI21_X1 U4975 ( .B1(PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n6937), .A(n4443), 
        .ZN(n4031) );
  NAND2_X1 U4976 ( .A1(n3987), .A2(EAX_REG_23__SCAN_IN), .ZN(n4030) );
  OAI211_X1 U4977 ( .C1(n4061), .C2(n4032), .A(n4031), .B(n4030), .ZN(n4033)
         );
  XNOR2_X1 U4978 ( .A(n4035), .B(n4034), .ZN(n4039) );
  AOI22_X1 U4979 ( .A1(n3987), .A2(EAX_REG_24__SCAN_IN), .B1(n4447), .B2(
        PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4038) );
  XNOR2_X1 U4980 ( .A(n4036), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5728)
         );
  NAND2_X1 U4981 ( .A1(n5728), .A2(n4443), .ZN(n4037) );
  OAI211_X1 U4982 ( .C1(n4039), .C2(n4061), .A(n4038), .B(n4037), .ZN(n5523)
         );
  INV_X1 U4983 ( .A(n4040), .ZN(n4041) );
  OAI21_X1 U4984 ( .B1(PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n4041), .A(n4052), 
        .ZN(n5980) );
  XNOR2_X1 U4985 ( .A(n4043), .B(n4042), .ZN(n4046) );
  AOI21_X1 U4986 ( .B1(PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6937), .A(n4443), 
        .ZN(n4045) );
  NAND2_X1 U4987 ( .A1(n3987), .A2(EAX_REG_25__SCAN_IN), .ZN(n4044) );
  OAI211_X1 U4988 ( .C1(n4046), .C2(n4061), .A(n4045), .B(n4044), .ZN(n4047)
         );
  XOR2_X1 U4989 ( .A(n4049), .B(n4048), .Z(n4050) );
  NAND2_X1 U4990 ( .A1(n4050), .A2(n4440), .ZN(n4054) );
  INV_X1 U4991 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5511) );
  NOR2_X1 U4992 ( .A1(n5511), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4051) );
  AOI211_X1 U4993 ( .C1(n3987), .C2(EAX_REG_26__SCAN_IN), .A(n4443), .B(n4051), 
        .ZN(n4053) );
  XNOR2_X1 U4994 ( .A(n4052), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5510)
         );
  AOI22_X1 U4995 ( .A1(n4054), .A2(n4053), .B1(n4443), .B2(n5510), .ZN(n5509)
         );
  NAND2_X1 U4996 ( .A1(n4055), .A2(n7097), .ZN(n4056) );
  NAND2_X1 U4997 ( .A1(n4068), .A2(n4056), .ZN(n5704) );
  XNOR2_X1 U4998 ( .A(n4058), .B(n4057), .ZN(n4062) );
  NOR2_X1 U4999 ( .A1(n7097), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4059) );
  AOI211_X1 U5000 ( .C1(n3987), .C2(EAX_REG_27__SCAN_IN), .A(n4443), .B(n4059), 
        .ZN(n4060) );
  OAI21_X1 U5001 ( .B1(n4062), .B2(n4061), .A(n4060), .ZN(n4063) );
  XOR2_X1 U5002 ( .A(n4065), .B(n4064), .Z(n4066) );
  NAND2_X1 U5003 ( .A1(n4066), .A2(n4440), .ZN(n4070) );
  NOR2_X1 U5004 ( .A1(n5488), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4067) );
  AOI211_X1 U5005 ( .C1(n3987), .C2(EAX_REG_28__SCAN_IN), .A(n4443), .B(n4067), 
        .ZN(n4069) );
  XNOR2_X1 U5006 ( .A(n4068), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5487)
         );
  AOI22_X1 U5007 ( .A1(n4070), .A2(n4069), .B1(n4443), .B2(n5487), .ZN(n5486)
         );
  INV_X1 U5008 ( .A(n5691), .ZN(n5674) );
  OR2_X1 U5009 ( .A1(n4073), .A2(n3174), .ZN(n4081) );
  OAI21_X1 U5010 ( .B1(n4076), .B2(n5400), .A(n6782), .ZN(n4075) );
  OAI21_X1 U5011 ( .B1(n4074), .B2(n4076), .A(n4075), .ZN(n4356) );
  OR2_X1 U5012 ( .A1(n4077), .A2(n4585), .ZN(n4478) );
  NAND2_X1 U5013 ( .A1(n4470), .A2(n4478), .ZN(n4078) );
  NAND2_X1 U5014 ( .A1(n4078), .A2(n4354), .ZN(n4080) );
  NAND2_X1 U5015 ( .A1(n4368), .A2(n4373), .ZN(n4079) );
  NAND2_X1 U5016 ( .A1(n4083), .A2(n4082), .ZN(n4487) );
  INV_X1 U5017 ( .A(n4085), .ZN(n4086) );
  NAND2_X1 U5018 ( .A1(n4492), .A2(n4086), .ZN(n4612) );
  OR2_X1 U5019 ( .A1(n4087), .A2(n3425), .ZN(n4088) );
  OAI211_X1 U5020 ( .C1(n4084), .C2(n3118), .A(n4612), .B(n4088), .ZN(n4089)
         );
  NOR2_X1 U5021 ( .A1(n4487), .A2(n4089), .ZN(n4384) );
  NOR2_X1 U5022 ( .A1(n6619), .A2(n4585), .ZN(n4359) );
  INV_X1 U5023 ( .A(n4090), .ZN(n4091) );
  NAND2_X1 U5024 ( .A1(n6556), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4106) );
  XNOR2_X1 U5025 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4100) );
  NAND2_X1 U5026 ( .A1(n4102), .A2(n4100), .ZN(n4093) );
  NAND2_X1 U5027 ( .A1(n7064), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4092) );
  NAND2_X1 U5028 ( .A1(n4093), .A2(n4092), .ZN(n4120) );
  XNOR2_X1 U5029 ( .A(n6925), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4118)
         );
  NAND2_X1 U5030 ( .A1(n4120), .A2(n4118), .ZN(n4095) );
  NAND2_X1 U5031 ( .A1(n6631), .A2(n6925), .ZN(n4094) );
  NAND2_X1 U5032 ( .A1(n4095), .A2(n4094), .ZN(n4128) );
  XNOR2_X1 U5033 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4126) );
  NAND2_X1 U5034 ( .A1(n4128), .A2(n4126), .ZN(n4097) );
  NAND2_X1 U5035 ( .A1(n7081), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4096) );
  NAND2_X1 U5036 ( .A1(n4097), .A2(n4096), .ZN(n4135) );
  AND2_X1 U5037 ( .A1(n6637), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4098)
         );
  NAND2_X1 U5038 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n4627), .ZN(n4134) );
  INV_X1 U5039 ( .A(n4100), .ZN(n4101) );
  XNOR2_X1 U5040 ( .A(n4102), .B(n4101), .ZN(n4361) );
  NAND2_X1 U5041 ( .A1(n4361), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4108) );
  INV_X1 U5042 ( .A(n4108), .ZN(n4113) );
  OR2_X1 U5043 ( .A1(n4138), .A2(n4585), .ZN(n4103) );
  AND2_X1 U5044 ( .A1(n4103), .A2(n3493), .ZN(n4109) );
  INV_X1 U5045 ( .A(n4109), .ZN(n4112) );
  OR2_X1 U5046 ( .A1(n5400), .A2(n3493), .ZN(n4104) );
  NAND2_X1 U5047 ( .A1(n4104), .A2(n4585), .ZN(n4121) );
  OAI21_X1 U5048 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6556), .A(n4106), 
        .ZN(n4110) );
  OAI21_X1 U5049 ( .B1(n4379), .B2(n4110), .A(n3118), .ZN(n4107) );
  AOI22_X1 U5050 ( .A1(n4109), .A2(n4108), .B1(n4121), .B2(n4107), .ZN(n4116)
         );
  NOR2_X1 U5051 ( .A1(n4138), .A2(n4110), .ZN(n4111) );
  AOI22_X1 U5052 ( .A1(n4113), .A2(n4112), .B1(n4116), .B2(n4111), .ZN(n4125)
         );
  INV_X1 U5053 ( .A(n4361), .ZN(n4117) );
  INV_X1 U5054 ( .A(n4114), .ZN(n4115) );
  OAI21_X1 U5055 ( .B1(n4117), .B2(n4116), .A(n4115), .ZN(n4124) );
  INV_X1 U5056 ( .A(n4118), .ZN(n4119) );
  XNOR2_X1 U5057 ( .A(n4120), .B(n4119), .ZN(n4362) );
  INV_X1 U5058 ( .A(n4121), .ZN(n4130) );
  NOR2_X1 U5059 ( .A1(n4362), .A2(n3555), .ZN(n4122) );
  AOI211_X1 U5060 ( .C1(n4362), .C2(n4129), .A(n4130), .B(n4122), .ZN(n4123)
         );
  AOI21_X1 U5061 ( .B1(n4125), .B2(n4124), .A(n4123), .ZN(n4133) );
  INV_X1 U5062 ( .A(n4126), .ZN(n4127) );
  XNOR2_X1 U5063 ( .A(n4128), .B(n4127), .ZN(n4363) );
  NAND3_X1 U5064 ( .A1(n4362), .A2(n4130), .A3(n4129), .ZN(n4131) );
  OAI21_X1 U5065 ( .B1(n4363), .B2(n4091), .A(n4131), .ZN(n4132) );
  INV_X1 U5066 ( .A(n4366), .ZN(n4137) );
  AOI222_X1 U5067 ( .A1(n4141), .A2(n4140), .B1(n4141), .B2(n4139), .C1(n4140), 
        .C2(n4139), .ZN(n4142) );
  INV_X1 U5068 ( .A(n4142), .ZN(n4143) );
  NAND3_X1 U5069 ( .A1(n6640), .A2(n6672), .A3(n6645), .ZN(n4154) );
  INV_X1 U5070 ( .A(n4147), .ZN(n4152) );
  INV_X1 U5071 ( .A(n3488), .ZN(n4148) );
  AND3_X1 U5072 ( .A1(n3510), .A2(n4149), .A3(n4148), .ZN(n4150) );
  NAND3_X1 U5073 ( .A1(n4152), .A2(n4151), .A3(n4150), .ZN(n4523) );
  NAND2_X2 U5074 ( .A1(n6231), .A2(n3488), .ZN(n5670) );
  INV_X1 U5075 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4541) );
  NAND2_X1 U5076 ( .A1(n4164), .A2(n4541), .ZN(n4158) );
  INV_X1 U5077 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4155) );
  NAND2_X1 U5078 ( .A1(n4230), .A2(n4155), .ZN(n4156) );
  OAI211_X1 U5079 ( .C1(n4168), .C2(EBX_REG_1__SCAN_IN), .A(n4156), .B(n3174), 
        .ZN(n4157) );
  INV_X1 U5080 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5618) );
  NAND2_X1 U5081 ( .A1(n3174), .A2(n5618), .ZN(n4160) );
  NAND2_X1 U5082 ( .A1(n4230), .A2(EBX_REG_0__SCAN_IN), .ZN(n4159) );
  NOR2_X1 U5083 ( .A1(n4539), .A2(n4168), .ZN(n4163) );
  INV_X1 U5084 ( .A(n4161), .ZN(n4162) );
  INV_X1 U5085 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4549) );
  NAND2_X1 U5086 ( .A1(n4164), .A2(n4549), .ZN(n4167) );
  NAND2_X1 U5087 ( .A1(n4238), .A2(n4168), .ZN(n4204) );
  NAND2_X1 U5088 ( .A1(n4238), .A2(EBX_REG_2__SCAN_IN), .ZN(n4166) );
  NAND2_X1 U5089 ( .A1(n4168), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4165)
         );
  NAND4_X1 U5090 ( .A1(n4167), .A2(n4204), .A3(n4166), .A4(n4165), .ZN(n4545)
         );
  NAND2_X1 U5091 ( .A1(n4546), .A2(n4545), .ZN(n4533) );
  INV_X1 U5092 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n7057) );
  INV_X1 U5093 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4169) );
  NAND2_X1 U5094 ( .A1(n4540), .A2(n4169), .ZN(n4170) );
  OAI211_X1 U5095 ( .C1(n5540), .C2(n7057), .A(n4170), .B(n4230), .ZN(n4171)
         );
  OAI21_X1 U5096 ( .B1(n4201), .B2(EBX_REG_3__SCAN_IN), .A(n4171), .ZN(n4534)
         );
  INV_X1 U5097 ( .A(n4164), .ZN(n4198) );
  INV_X1 U5098 ( .A(EBX_REG_4__SCAN_IN), .ZN(n6900) );
  NAND2_X1 U5099 ( .A1(n4540), .A2(n6900), .ZN(n4172) );
  OAI211_X1 U5100 ( .C1(n4238), .C2(INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4172), 
        .B(n3174), .ZN(n4173) );
  OAI21_X1 U5101 ( .B1(n4198), .B2(EBX_REG_4__SCAN_IN), .A(n4173), .ZN(n4559)
         );
  NAND2_X1 U5102 ( .A1(EBX_REG_5__SCAN_IN), .A2(n5540), .ZN(n4175) );
  INV_X1 U5103 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4667) );
  NAND2_X1 U5104 ( .A1(n4470), .A2(n4667), .ZN(n4174) );
  OAI211_X1 U5105 ( .C1(EBX_REG_5__SCAN_IN), .C2(n4201), .A(n4175), .B(n4174), 
        .ZN(n4553) );
  INV_X1 U5106 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6151) );
  NAND2_X1 U5107 ( .A1(n4164), .A2(n6151), .ZN(n4178) );
  INV_X1 U5108 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4302) );
  NAND2_X1 U5109 ( .A1(n4230), .A2(n4302), .ZN(n4176) );
  OAI211_X1 U5110 ( .C1(n4168), .C2(EBX_REG_6__SCAN_IN), .A(n4176), .B(n3174), 
        .ZN(n4177) );
  NAND2_X1 U5111 ( .A1(n4178), .A2(n4177), .ZN(n4680) );
  NAND2_X1 U5112 ( .A1(n5540), .A2(EBX_REG_7__SCAN_IN), .ZN(n4180) );
  INV_X1 U5113 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6395) );
  NAND2_X1 U5114 ( .A1(n4470), .A2(n6395), .ZN(n4179) );
  OAI211_X1 U5115 ( .C1(EBX_REG_7__SCAN_IN), .C2(n4201), .A(n4180), .B(n4179), 
        .ZN(n4800) );
  INV_X1 U5116 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5599) );
  NAND2_X1 U5117 ( .A1(n4164), .A2(n5599), .ZN(n4183) );
  INV_X1 U5118 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4323) );
  NAND2_X1 U5119 ( .A1(n4230), .A2(n4323), .ZN(n4181) );
  OAI211_X1 U5120 ( .C1(n4168), .C2(EBX_REG_8__SCAN_IN), .A(n4181), .B(n3174), 
        .ZN(n4182) );
  NAND2_X1 U5121 ( .A1(n4183), .A2(n4182), .ZN(n4900) );
  NOR2_X1 U5122 ( .A1(n4201), .A2(EBX_REG_9__SCAN_IN), .ZN(n4184) );
  AOI21_X1 U5123 ( .B1(EBX_REG_9__SCAN_IN), .B2(n5540), .A(n4184), .ZN(n4185)
         );
  OAI21_X1 U5124 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n5460), .A(n4185), 
        .ZN(n5178) );
  INV_X1 U5125 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5270) );
  NAND2_X1 U5126 ( .A1(n4164), .A2(n5270), .ZN(n4188) );
  NAND2_X1 U5127 ( .A1(n4238), .A2(EBX_REG_10__SCAN_IN), .ZN(n4187) );
  NAND2_X1 U5128 ( .A1(n4168), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4186) );
  NAND4_X1 U5129 ( .A1(n4188), .A2(n4204), .A3(n4187), .A4(n4186), .ZN(n5268)
         );
  INV_X1 U5130 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4330) );
  INV_X1 U5131 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5585) );
  NAND2_X1 U5132 ( .A1(n4540), .A2(n5585), .ZN(n4189) );
  OAI211_X1 U5133 ( .C1(n5540), .C2(n4330), .A(n4189), .B(n4230), .ZN(n4190)
         );
  OAI21_X1 U5134 ( .B1(n4201), .B2(EBX_REG_11__SCAN_IN), .A(n4190), .ZN(n5275)
         );
  INV_X1 U5135 ( .A(n4204), .ZN(n4195) );
  AOI21_X1 U5136 ( .B1(n4238), .B2(EBX_REG_12__SCAN_IN), .A(n4195), .ZN(n4192)
         );
  NAND2_X1 U5137 ( .A1(n4168), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4191) );
  OAI211_X1 U5138 ( .C1(EBX_REG_12__SCAN_IN), .C2(n4198), .A(n4192), .B(n4191), 
        .ZN(n5346) );
  NAND2_X1 U5139 ( .A1(n5347), .A2(n5346), .ZN(n5359) );
  INV_X1 U5140 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4389) );
  INV_X1 U5141 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6939) );
  NAND2_X1 U5142 ( .A1(n4540), .A2(n6939), .ZN(n4193) );
  OAI211_X1 U5143 ( .C1(n5540), .C2(n4389), .A(n4193), .B(n4230), .ZN(n4194)
         );
  OAI21_X1 U5144 ( .B1(n4201), .B2(EBX_REG_13__SCAN_IN), .A(n4194), .ZN(n5360)
         );
  NOR2_X2 U5145 ( .A1(n5359), .A2(n5360), .ZN(n5377) );
  AOI21_X1 U5146 ( .B1(n4238), .B2(EBX_REG_14__SCAN_IN), .A(n4195), .ZN(n4197)
         );
  NAND2_X1 U5147 ( .A1(n4168), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4196) );
  OAI211_X1 U5148 ( .C1(EBX_REG_14__SCAN_IN), .C2(n4198), .A(n4197), .B(n4196), 
        .ZN(n5378) );
  INV_X1 U5149 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n7094) );
  INV_X1 U5150 ( .A(EBX_REG_15__SCAN_IN), .ZN(n6956) );
  NAND2_X1 U5151 ( .A1(n4540), .A2(n6956), .ZN(n4199) );
  OAI211_X1 U5152 ( .C1(n5540), .C2(n7094), .A(n4199), .B(n4230), .ZN(n4200)
         );
  OAI21_X1 U5153 ( .B1(n4201), .B2(EBX_REG_15__SCAN_IN), .A(n4200), .ZN(n5396)
         );
  INV_X1 U5154 ( .A(EBX_REG_16__SCAN_IN), .ZN(n4202) );
  NAND2_X1 U5155 ( .A1(n4164), .A2(n4202), .ZN(n4206) );
  NAND2_X1 U5156 ( .A1(n4238), .A2(EBX_REG_16__SCAN_IN), .ZN(n4205) );
  NAND2_X1 U5157 ( .A1(n4168), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4203) );
  NAND4_X1 U5158 ( .A1(n4206), .A2(n4205), .A3(n4204), .A4(n4203), .ZN(n5560)
         );
  INV_X1 U5159 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6225) );
  NAND2_X1 U5160 ( .A1(n4234), .A2(n6225), .ZN(n4209) );
  NAND2_X1 U5161 ( .A1(n3174), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4207) );
  OAI211_X1 U5162 ( .C1(n4168), .C2(EBX_REG_17__SCAN_IN), .A(n4230), .B(n4207), 
        .ZN(n4208) );
  NAND2_X1 U5163 ( .A1(n4209), .A2(n4208), .ZN(n6021) );
  INV_X1 U5164 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5667) );
  NAND2_X1 U5165 ( .A1(n4164), .A2(n5667), .ZN(n4211) );
  AOI22_X1 U5166 ( .A1(n4238), .A2(EBX_REG_19__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n4168), .ZN(n4210) );
  INV_X1 U5167 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5879) );
  NAND2_X1 U5168 ( .A1(n4470), .A2(n5879), .ZN(n4213) );
  INV_X1 U5169 ( .A(EBX_REG_18__SCAN_IN), .ZN(n4212) );
  NAND2_X1 U5170 ( .A1(n4540), .A2(n4212), .ZN(n5539) );
  OAI22_X1 U5171 ( .A1(n5460), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        EBX_REG_20__SCAN_IN), .B2(n4168), .ZN(n5659) );
  NAND2_X1 U5172 ( .A1(n5656), .A2(n5659), .ZN(n4215) );
  NAND2_X1 U5173 ( .A1(n5540), .A2(EBX_REG_20__SCAN_IN), .ZN(n4214) );
  OAI211_X1 U5174 ( .C1(n5656), .C2(n5540), .A(n4215), .B(n4214), .ZN(n4216)
         );
  INV_X1 U5175 ( .A(n4216), .ZN(n4217) );
  NAND2_X1 U5176 ( .A1(n5658), .A2(n4217), .ZN(n5651) );
  INV_X1 U5177 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5653) );
  NAND2_X1 U5178 ( .A1(n4234), .A2(n5653), .ZN(n4219) );
  NAND2_X1 U5179 ( .A1(n5540), .A2(EBX_REG_21__SCAN_IN), .ZN(n4218) );
  OAI211_X1 U5180 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5460), .A(n4219), .B(n4218), .ZN(n5650) );
  OR2_X2 U5181 ( .A1(n5651), .A2(n5650), .ZN(n5648) );
  INV_X1 U5182 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5645) );
  NAND2_X1 U5183 ( .A1(n4164), .A2(n5645), .ZN(n4221) );
  AOI22_X1 U5184 ( .A1(n4238), .A2(EBX_REG_22__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n4168), .ZN(n4220) );
  INV_X1 U5185 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5639) );
  NAND2_X1 U5186 ( .A1(n4234), .A2(n5639), .ZN(n4224) );
  NAND2_X1 U5187 ( .A1(n3174), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4222) );
  OAI211_X1 U5188 ( .C1(n4168), .C2(EBX_REG_23__SCAN_IN), .A(n4230), .B(n4222), 
        .ZN(n4223) );
  AND2_X1 U5189 ( .A1(n4224), .A2(n4223), .ZN(n5636) );
  INV_X1 U5190 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5529) );
  NAND2_X1 U5191 ( .A1(n4164), .A2(n5529), .ZN(n4226) );
  AOI22_X1 U5192 ( .A1(n4238), .A2(EBX_REG_24__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n4168), .ZN(n4225) );
  NAND2_X1 U5193 ( .A1(n4226), .A2(n4225), .ZN(n5525) );
  INV_X1 U5194 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5631) );
  NAND2_X1 U5195 ( .A1(n4234), .A2(n5631), .ZN(n4228) );
  NAND2_X1 U5196 ( .A1(n5540), .A2(EBX_REG_25__SCAN_IN), .ZN(n4227) );
  OAI211_X1 U5197 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n5460), .A(n4228), .B(n4227), .ZN(n5629) );
  INV_X1 U5198 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5627) );
  NAND2_X1 U5199 ( .A1(n4164), .A2(n5627), .ZN(n4233) );
  INV_X1 U5200 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4229) );
  NAND2_X1 U5201 ( .A1(n4230), .A2(n4229), .ZN(n4231) );
  OAI211_X1 U5202 ( .C1(n4168), .C2(EBX_REG_26__SCAN_IN), .A(n4231), .B(n3174), 
        .ZN(n4232) );
  NAND2_X1 U5203 ( .A1(n4233), .A2(n4232), .ZN(n5514) );
  NAND2_X1 U5204 ( .A1(n5512), .A2(n5514), .ZN(n5513) );
  INV_X1 U5205 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5626) );
  NAND2_X1 U5206 ( .A1(n4234), .A2(n5626), .ZN(n4236) );
  NAND2_X1 U5207 ( .A1(n5540), .A2(EBX_REG_27__SCAN_IN), .ZN(n4235) );
  OAI211_X1 U5208 ( .C1(INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n5460), .A(n4236), .B(n4235), .ZN(n5498) );
  INV_X1 U5209 ( .A(n4237), .ZN(n5500) );
  INV_X1 U5210 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5624) );
  NAND2_X1 U5211 ( .A1(n4164), .A2(n5624), .ZN(n4240) );
  AOI22_X1 U5212 ( .A1(n4238), .A2(EBX_REG_28__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n4168), .ZN(n4239) );
  AND2_X1 U5213 ( .A1(n4240), .A2(n4239), .ZN(n4404) );
  OAI22_X1 U5214 ( .A1(n5460), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        EBX_REG_29__SCAN_IN), .B2(n4168), .ZN(n4242) );
  INV_X1 U5215 ( .A(EBX_REG_29__SCAN_IN), .ZN(n4245) );
  NAND2_X1 U5216 ( .A1(n4164), .A2(n4245), .ZN(n4241) );
  OAI22_X1 U5217 ( .A1(n5446), .A2(n5540), .B1(n4241), .B2(n5445), .ZN(n5462)
         );
  OAI211_X1 U5218 ( .C1(n5540), .C2(n4242), .A(n5445), .B(n4241), .ZN(n4243)
         );
  INV_X1 U5219 ( .A(n4243), .ZN(n4244) );
  INV_X1 U5220 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4347) );
  INV_X1 U5221 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n7001) );
  NAND2_X1 U5222 ( .A1(n4347), .A2(n7001), .ZN(n5417) );
  NAND2_X1 U5223 ( .A1(n4574), .A2(n4090), .ZN(n4252) );
  AND2_X1 U5224 ( .A1(n5400), .A2(n4656), .ZN(n4265) );
  INV_X1 U5225 ( .A(n4265), .ZN(n4249) );
  OAI21_X1 U5226 ( .B1(n6782), .B2(n4254), .A(n4249), .ZN(n4250) );
  INV_X1 U5227 ( .A(n4250), .ZN(n4251) );
  NAND2_X1 U5228 ( .A1(n4252), .A2(n4251), .ZN(n6362) );
  NAND2_X1 U5229 ( .A1(n4573), .A2(n4090), .ZN(n4259) );
  NAND2_X1 U5230 ( .A1(n4253), .A2(n4254), .ZN(n4263) );
  OAI21_X1 U5231 ( .B1(n4254), .B2(n4253), .A(n4263), .ZN(n4256) );
  INV_X1 U5232 ( .A(n4354), .ZN(n4255) );
  OAI211_X1 U5233 ( .C1(n4256), .C2(n6782), .A(n4255), .B(n3493), .ZN(n4257)
         );
  INV_X1 U5234 ( .A(n4257), .ZN(n4258) );
  NAND2_X1 U5235 ( .A1(n4259), .A2(n4258), .ZN(n4562) );
  NAND2_X1 U5236 ( .A1(n4563), .A2(n4562), .ZN(n4561) );
  INV_X1 U5237 ( .A(n4260), .ZN(n4261) );
  NAND2_X1 U5238 ( .A1(n4261), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4262)
         );
  AND2_X1 U5239 ( .A1(n4561), .A2(n4262), .ZN(n6355) );
  NAND2_X1 U5240 ( .A1(n4571), .A2(n4090), .ZN(n4268) );
  NAND2_X1 U5241 ( .A1(n4263), .A2(n4264), .ZN(n4273) );
  OAI21_X1 U5242 ( .B1(n4264), .B2(n4263), .A(n4273), .ZN(n4266) );
  AOI21_X1 U5243 ( .B1(n4266), .B2(n4309), .A(n4265), .ZN(n4267) );
  NAND2_X1 U5244 ( .A1(n4269), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6352)
         );
  NAND2_X1 U5245 ( .A1(n6355), .A2(n6352), .ZN(n4272) );
  NAND2_X1 U5246 ( .A1(n4271), .A2(n4270), .ZN(n6353) );
  AND2_X1 U5247 ( .A1(n4272), .A2(n6353), .ZN(n4762) );
  NAND2_X1 U5248 ( .A1(n4273), .A2(n4274), .ZN(n4290) );
  OAI211_X1 U5249 ( .C1(n4274), .C2(n4273), .A(n4290), .B(n4309), .ZN(n4275)
         );
  XNOR2_X1 U5250 ( .A(n4277), .B(n7057), .ZN(n4763) );
  NAND2_X1 U5251 ( .A1(n4762), .A2(n4763), .ZN(n4279) );
  NAND2_X1 U5252 ( .A1(n4277), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4278)
         );
  NAND2_X1 U5253 ( .A1(n4279), .A2(n4278), .ZN(n4777) );
  NAND2_X1 U5254 ( .A1(n4280), .A2(n4090), .ZN(n4284) );
  XNOR2_X1 U5255 ( .A(n4290), .B(n4281), .ZN(n4282) );
  NAND2_X1 U5256 ( .A1(n4282), .A2(n4309), .ZN(n4283) );
  NAND2_X1 U5257 ( .A1(n4284), .A2(n4283), .ZN(n4286) );
  INV_X1 U5258 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4285) );
  NAND2_X1 U5259 ( .A1(n4777), .A2(n4778), .ZN(n4288) );
  NAND2_X1 U5260 ( .A1(n4286), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4287)
         );
  NOR2_X1 U5261 ( .A1(n4290), .A2(n4289), .ZN(n4292) );
  NAND2_X1 U5262 ( .A1(n4292), .A2(n4291), .ZN(n4306) );
  OAI211_X1 U5263 ( .C1(n4292), .C2(n4291), .A(n4306), .B(n4309), .ZN(n4293)
         );
  XNOR2_X1 U5264 ( .A(n4295), .B(n4667), .ZN(n4661) );
  NAND2_X1 U5265 ( .A1(n4662), .A2(n4661), .ZN(n4297) );
  NAND2_X1 U5266 ( .A1(n4295), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4296)
         );
  NAND3_X1 U5267 ( .A1(n4316), .A2(n4298), .A3(n4090), .ZN(n4301) );
  XNOR2_X1 U5268 ( .A(n4306), .B(n4307), .ZN(n4299) );
  NAND2_X1 U5269 ( .A1(n4299), .A2(n4309), .ZN(n4300) );
  NAND2_X1 U5270 ( .A1(n4303), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4304)
         );
  NAND2_X1 U5271 ( .A1(n4305), .A2(n4090), .ZN(n4312) );
  INV_X1 U5272 ( .A(n4306), .ZN(n4308) );
  NAND2_X1 U5273 ( .A1(n4308), .A2(n4307), .ZN(n4321) );
  XNOR2_X1 U5274 ( .A(n4321), .B(n4319), .ZN(n4310) );
  NAND2_X1 U5275 ( .A1(n4310), .A2(n4309), .ZN(n4311) );
  NAND2_X1 U5276 ( .A1(n4312), .A2(n4311), .ZN(n4313) );
  XNOR2_X1 U5277 ( .A(n4313), .B(n6395), .ZN(n5262) );
  NAND2_X1 U5278 ( .A1(n4313), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4314)
         );
  NAND2_X1 U5279 ( .A1(n4315), .A2(n4314), .ZN(n5205) );
  NOR2_X1 U5280 ( .A1(n4317), .A2(n4091), .ZN(n4318) );
  NAND2_X1 U5281 ( .A1(n4309), .A2(n4319), .ZN(n4320) );
  OR2_X1 U5282 ( .A1(n4321), .A2(n4320), .ZN(n4322) );
  NAND2_X1 U5283 ( .A1(n4327), .A2(n4322), .ZN(n4324) );
  XNOR2_X1 U5284 ( .A(n4324), .B(n4323), .ZN(n5206) );
  NAND2_X1 U5285 ( .A1(n5205), .A2(n5206), .ZN(n4326) );
  NAND2_X1 U5286 ( .A1(n4324), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4325)
         );
  INV_X1 U5287 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5300) );
  NAND2_X1 U5288 ( .A1(n4327), .A2(n5300), .ZN(n4328) );
  INV_X1 U5289 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5291) );
  AND2_X1 U5290 ( .A1(n4327), .A2(n5291), .ZN(n5283) );
  NAND2_X1 U5291 ( .A1(n4327), .A2(n4330), .ZN(n5319) );
  OR2_X1 U5292 ( .A1(n4327), .A2(n4330), .ZN(n5320) );
  INV_X1 U5293 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4332) );
  NOR2_X1 U5294 ( .A1(n4327), .A2(n4332), .ZN(n5329) );
  INV_X1 U5295 ( .A(n5329), .ZN(n4331) );
  NAND2_X1 U5296 ( .A1(n4327), .A2(n4332), .ZN(n5328) );
  XNOR2_X1 U5297 ( .A(n4327), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5363)
         );
  NAND2_X1 U5298 ( .A1(n4327), .A2(n4389), .ZN(n4334) );
  INV_X1 U5299 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6047) );
  OR2_X1 U5300 ( .A1(n4327), .A2(n6047), .ZN(n4335) );
  NAND2_X1 U5301 ( .A1(n4327), .A2(n6047), .ZN(n4336) );
  XNOR2_X1 U5302 ( .A(n4327), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5773)
         );
  NAND2_X1 U5303 ( .A1(n4327), .A2(n7094), .ZN(n4338) );
  INV_X1 U5304 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5893) );
  NAND2_X1 U5305 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4393) );
  AND2_X1 U5306 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5848) );
  AND2_X1 U5307 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5863) );
  AND2_X1 U5308 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4410) );
  NAND3_X1 U5309 ( .A1(n5848), .A2(n5863), .A3(n4410), .ZN(n4340) );
  NOR2_X1 U5310 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5847) );
  NOR2_X1 U5311 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5832) );
  NOR2_X1 U5312 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5864) );
  AND3_X1 U5313 ( .A1(n5847), .A2(n5832), .A3(n5864), .ZN(n4342) );
  OR2_X1 U5314 ( .A1(n4327), .A2(n4342), .ZN(n4343) );
  INV_X1 U5315 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6010) );
  XNOR2_X1 U5316 ( .A(n4327), .B(n6010), .ZN(n5975) );
  INV_X1 U5317 ( .A(n5975), .ZN(n4344) );
  INV_X1 U5318 ( .A(n4346), .ZN(n5974) );
  NOR2_X1 U5319 ( .A1(n4327), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5709)
         );
  NAND2_X1 U5320 ( .A1(n4327), .A2(n6010), .ZN(n4345) );
  AND2_X2 U5321 ( .A1(n4346), .A2(n4345), .ZN(n5416) );
  AND2_X1 U5322 ( .A1(n4327), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5708)
         );
  INV_X1 U5323 ( .A(n4417), .ZN(n5686) );
  NAND3_X1 U5324 ( .A1(n5686), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n4347), .ZN(n4349) );
  NAND3_X1 U5325 ( .A1(n5701), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .A3(n7001), .ZN(n4348) );
  OAI211_X1 U5326 ( .C1(n5417), .C2(n5701), .A(n4349), .B(n4348), .ZN(n4351)
         );
  AND2_X1 U5327 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5805) );
  NOR2_X1 U5328 ( .A1(n4351), .A2(n4350), .ZN(n5700) );
  AND2_X1 U5329 ( .A1(n4379), .A2(n5400), .ZN(n4353) );
  INV_X1 U5330 ( .A(n6644), .ZN(n4358) );
  AOI21_X1 U5331 ( .B1(n6619), .B2(n5400), .A(n4354), .ZN(n4355) );
  AND2_X1 U5332 ( .A1(n4073), .A2(n4355), .ZN(n4380) );
  NAND2_X1 U5333 ( .A1(n4380), .A2(n4356), .ZN(n4357) );
  NAND2_X1 U5334 ( .A1(n4358), .A2(n4357), .ZN(n4481) );
  NAND2_X1 U5335 ( .A1(n6645), .A2(n4359), .ZN(n4370) );
  OR2_X1 U5336 ( .A1(n4360), .A2(STATE_REG_0__SCAN_IN), .ZN(n6689) );
  INV_X1 U5337 ( .A(n6689), .ZN(n4705) );
  NAND3_X1 U5338 ( .A1(n4363), .A2(n4362), .A3(n4361), .ZN(n4364) );
  NAND2_X1 U5339 ( .A1(n4365), .A2(n4364), .ZN(n4367) );
  NOR2_X1 U5340 ( .A1(n6643), .A2(READY_N), .ZN(n4524) );
  OAI211_X1 U5341 ( .C1(n4585), .C2(n4705), .A(n4368), .B(n4524), .ZN(n4369)
         );
  NAND3_X1 U5342 ( .A1(n4481), .A2(n4370), .A3(n4369), .ZN(n4371) );
  NAND2_X1 U5343 ( .A1(n4371), .A2(n6672), .ZN(n4377) );
  NAND2_X1 U5344 ( .A1(n4585), .A2(n6689), .ZN(n5401) );
  NAND2_X1 U5345 ( .A1(n5401), .A2(n6778), .ZN(n4374) );
  OAI211_X1 U5346 ( .C1(n4372), .C2(n4374), .A(n3118), .B(n4373), .ZN(n4375)
         );
  NAND3_X1 U5347 ( .A1(n4703), .A2(n4599), .A3(n4375), .ZN(n4376) );
  AND2_X1 U5348 ( .A1(n4380), .A2(n5606), .ZN(n4525) );
  AND2_X1 U5349 ( .A1(n4380), .A2(n4379), .ZN(n6649) );
  NOR2_X1 U5350 ( .A1(n4525), .A2(n6649), .ZN(n6642) );
  OR2_X1 U5351 ( .A1(n4372), .A2(n4168), .ZN(n4520) );
  INV_X1 U5352 ( .A(n4381), .ZN(n4400) );
  NAND2_X1 U5353 ( .A1(n4400), .A2(n3487), .ZN(n4382) );
  AND4_X1 U5354 ( .A1(n4378), .A2(n6642), .A3(n4520), .A4(n4382), .ZN(n4383)
         );
  NAND2_X1 U5355 ( .A1(n6644), .A2(n3492), .ZN(n6622) );
  OR2_X1 U5356 ( .A1(n4384), .A2(n4403), .ZN(n4387) );
  INV_X1 U5357 ( .A(n4387), .ZN(n5338) );
  INV_X1 U5358 ( .A(n4403), .ZN(n4385) );
  INV_X1 U5359 ( .A(n5370), .ZN(n4386) );
  NAND2_X1 U5360 ( .A1(n6419), .A2(n4386), .ZN(n5887) );
  AND2_X1 U5361 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4411) );
  NAND2_X1 U5362 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4399) );
  NAND2_X1 U5363 ( .A1(n4387), .A2(n6419), .ZN(n5335) );
  INV_X1 U5364 ( .A(n6419), .ZN(n5344) );
  NOR2_X1 U5365 ( .A1(n5344), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4564)
         );
  INV_X1 U5366 ( .A(n4564), .ZN(n4388) );
  NAND2_X1 U5367 ( .A1(n5335), .A2(n4388), .ZN(n4764) );
  NAND2_X1 U5368 ( .A1(n4764), .A2(n6403), .ZN(n4398) );
  NOR2_X1 U5369 ( .A1(n6395), .A2(n4323), .ZN(n5290) );
  NAND3_X1 U5370 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n5290), .ZN(n5339) );
  NAND2_X1 U5371 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5372) );
  NOR2_X1 U5372 ( .A1(n4389), .A2(n5372), .ZN(n5889) );
  NAND2_X1 U5373 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5889), .ZN(n5888) );
  NAND2_X1 U5374 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5891) );
  OR3_X1 U5375 ( .A1(n5339), .A2(n5888), .A3(n5891), .ZN(n4395) );
  NAND2_X1 U5376 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4392) );
  INV_X1 U5377 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6757) );
  OAI21_X1 U5378 ( .B1(n4155), .B2(n6757), .A(n4270), .ZN(n6399) );
  INV_X1 U5379 ( .A(n6399), .ZN(n4390) );
  NAND2_X1 U5380 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4779) );
  NOR2_X1 U5381 ( .A1(n4390), .A2(n4779), .ZN(n4790) );
  NAND2_X1 U5382 ( .A1(n4391), .A2(n4790), .ZN(n4666) );
  NOR2_X1 U5383 ( .A1(n4395), .A2(n5341), .ZN(n5866) );
  NAND2_X1 U5384 ( .A1(n4403), .A2(n6401), .ZN(n6418) );
  NAND2_X1 U5385 ( .A1(n6757), .A2(n5370), .ZN(n6411) );
  NAND2_X1 U5386 ( .A1(n6418), .A2(n6411), .ZN(n4663) );
  INV_X1 U5387 ( .A(n4663), .ZN(n4570) );
  NAND2_X1 U5388 ( .A1(n6403), .A2(n4570), .ZN(n5204) );
  INV_X1 U5389 ( .A(n5204), .ZN(n5867) );
  NOR2_X1 U5390 ( .A1(n5866), .A2(n5867), .ZN(n4394) );
  INV_X1 U5391 ( .A(n4393), .ZN(n5862) );
  NAND2_X1 U5392 ( .A1(n5862), .A2(n5863), .ZN(n4407) );
  OAI22_X1 U5393 ( .A1(n4394), .A2(n4407), .B1(n5204), .B2(n5335), .ZN(n4397)
         );
  NAND2_X1 U5394 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4765) );
  NOR2_X1 U5395 ( .A1(n4765), .A2(n4779), .ZN(n4665) );
  NAND3_X1 U5396 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n4665), .ZN(n5342) );
  NOR2_X1 U5397 ( .A1(n5342), .A2(n4395), .ZN(n4406) );
  INV_X1 U5398 ( .A(n4406), .ZN(n4396) );
  NAND2_X1 U5399 ( .A1(n5335), .A2(n4396), .ZN(n5865) );
  OAI21_X1 U5400 ( .B1(n5848), .B2(n5288), .A(n5861), .ZN(n5843) );
  AOI21_X1 U5401 ( .B1(n4399), .B2(n4398), .A(n5843), .ZN(n6011) );
  OAI21_X1 U5402 ( .B1(n5288), .B2(n4411), .A(n6011), .ZN(n5818) );
  OR2_X1 U5403 ( .A1(n4372), .A2(n6782), .ZN(n4701) );
  NAND2_X1 U5404 ( .A1(n4400), .A2(n4848), .ZN(n4401) );
  AND2_X1 U5405 ( .A1(n4701), .A2(n4401), .ZN(n4402) );
  INV_X1 U5406 ( .A(n4404), .ZN(n4405) );
  OAI21_X1 U5407 ( .B1(n4237), .B2(n4405), .A(n5445), .ZN(n5625) );
  INV_X1 U5408 ( .A(n4764), .ZN(n6397) );
  OR2_X1 U5409 ( .A1(n5866), .A2(n5868), .ZN(n6026) );
  INV_X1 U5410 ( .A(n4407), .ZN(n4408) );
  NAND2_X1 U5411 ( .A1(n6026), .A2(n4408), .ZN(n5855) );
  INV_X1 U5412 ( .A(n5848), .ZN(n4409) );
  NOR2_X1 U5413 ( .A1(n5855), .A2(n4409), .ZN(n5831) );
  NAND2_X1 U5414 ( .A1(n5831), .A2(n4410), .ZN(n5826) );
  INV_X1 U5415 ( .A(n4411), .ZN(n4412) );
  NOR2_X1 U5416 ( .A1(n5826), .A2(n4412), .ZN(n5817) );
  INV_X1 U5417 ( .A(n5805), .ZN(n5788) );
  NAND3_X1 U5418 ( .A1(n5817), .A2(n5417), .A3(n5788), .ZN(n4414) );
  AND2_X1 U5419 ( .A1(n6351), .A2(REIP_REG_28__SCAN_IN), .ZN(n5694) );
  INV_X1 U5420 ( .A(n5694), .ZN(n4413) );
  OAI211_X1 U5421 ( .C1(n6413), .C2(n5625), .A(n4414), .B(n4413), .ZN(n4415)
         );
  AOI21_X1 U5422 ( .B1(n5818), .B2(INSTADDRPOINTER_REG_28__SCAN_IN), .A(n4415), 
        .ZN(n4416) );
  INV_X1 U5423 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5790) );
  INV_X1 U5424 ( .A(n5796), .ZN(n4418) );
  NAND2_X1 U5425 ( .A1(n4418), .A2(n6367), .ZN(n4460) );
  NOR2_X1 U5426 ( .A1(n4420), .A2(n4419), .ZN(n4439) );
  AOI22_X1 U5427 ( .A1(n4421), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3257), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4427) );
  AOI22_X1 U5428 ( .A1(n4610), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4426) );
  AOI22_X1 U5429 ( .A1(n4423), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4422), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4425) );
  AOI22_X1 U5430 ( .A1(n3644), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3584), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4424) );
  NAND4_X1 U5431 ( .A1(n4427), .A2(n4426), .A3(n4425), .A4(n4424), .ZN(n4437)
         );
  AOI22_X1 U5432 ( .A1(n3477), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3476), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4435) );
  AOI22_X1 U5433 ( .A1(n3560), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4428), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4434) );
  AOI22_X1 U5434 ( .A1(n3920), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4429), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4433) );
  AOI22_X1 U5435 ( .A1(n4431), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4430), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4432) );
  NAND4_X1 U5436 ( .A1(n4435), .A2(n4434), .A3(n4433), .A4(n4432), .ZN(n4436)
         );
  NOR2_X1 U5437 ( .A1(n4437), .A2(n4436), .ZN(n4438) );
  XNOR2_X1 U5438 ( .A(n4439), .B(n4438), .ZN(n4441) );
  NAND2_X1 U5439 ( .A1(n4441), .A2(n4440), .ZN(n4446) );
  INV_X1 U5440 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n6923) );
  OAI21_X1 U5441 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6923), .A(n3150), .ZN(
        n4442) );
  AOI21_X1 U5442 ( .B1(n3987), .B2(EAX_REG_30__SCAN_IN), .A(n4442), .ZN(n4445)
         );
  XNOR2_X1 U5443 ( .A(n4454), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5449)
         );
  AOI21_X1 U5444 ( .B1(n4446), .B2(n4445), .A(n4444), .ZN(n5422) );
  AOI22_X1 U5445 ( .A1(n3987), .A2(EAX_REG_31__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n4447), .ZN(n4448) );
  XNOR2_X2 U5446 ( .A(n4449), .B(n4448), .ZN(n5466) );
  AND2_X1 U5447 ( .A1(n6872), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5385) );
  NAND2_X1 U5448 ( .A1(n5385), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6679) );
  NAND2_X1 U5449 ( .A1(n6564), .A2(n4450), .ZN(n6777) );
  NAND2_X1 U5450 ( .A1(n6777), .A2(n6872), .ZN(n4451) );
  NAND2_X1 U5451 ( .A1(n6872), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4453) );
  NAND2_X1 U5452 ( .A1(n6064), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4452) );
  AND2_X1 U5453 ( .A1(n4453), .A2(n4452), .ZN(n6364) );
  INV_X1 U5454 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n6869) );
  NAND2_X1 U5455 ( .A1(n6368), .A2(REIP_REG_31__SCAN_IN), .ZN(n5791) );
  OAI21_X1 U5456 ( .B1(n6365), .B2(n6869), .A(n5791), .ZN(n4456) );
  NAND2_X1 U5457 ( .A1(n4460), .A2(n4459), .ZN(U2955) );
  NOR2_X1 U5458 ( .A1(n6643), .A2(n6660), .ZN(n4461) );
  NAND2_X1 U5459 ( .A1(n6644), .A2(n4461), .ZN(n4465) );
  INV_X1 U5460 ( .A(n4465), .ZN(n4464) );
  INV_X1 U5461 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n4463) );
  NAND2_X1 U5462 ( .A1(n6520), .A2(n5389), .ZN(n6060) );
  INV_X1 U5463 ( .A(n6641), .ZN(n4462) );
  OAI211_X1 U5464 ( .C1(n4464), .C2(n4463), .A(n6060), .B(n6265), .ZN(U2788)
         );
  INV_X1 U5465 ( .A(n6776), .ZN(n4468) );
  AND2_X1 U5466 ( .A1(n5400), .A2(n3492), .ZN(n5605) );
  INV_X1 U5467 ( .A(n5605), .ZN(n4466) );
  NAND2_X1 U5468 ( .A1(n4466), .A2(n6782), .ZN(n6065) );
  INV_X1 U5469 ( .A(n6060), .ZN(n5397) );
  OAI21_X1 U5470 ( .B1(n5397), .B2(READREQUEST_REG_SCAN_IN), .A(n4468), .ZN(
        n4467) );
  OAI21_X1 U5471 ( .B1(n4468), .B2(n6065), .A(n4467), .ZN(U3474) );
  INV_X1 U5472 ( .A(n4469), .ZN(n4472) );
  NAND2_X1 U5473 ( .A1(n4470), .A2(n6757), .ZN(n4471) );
  NAND2_X1 U5474 ( .A1(n4472), .A2(n4471), .ZN(n6412) );
  OAI21_X1 U5475 ( .B1(n4475), .B2(n4474), .A(n4473), .ZN(n6371) );
  OAI222_X1 U5476 ( .A1(n6412), .A2(n5671), .B1(n6231), .B2(n5618), .C1(n5670), 
        .C2(n6371), .ZN(U2859) );
  NAND2_X1 U5477 ( .A1(n6622), .A2(n4372), .ZN(n4477) );
  AOI21_X1 U5478 ( .B1(n4168), .B2(n6689), .A(READY_N), .ZN(n4476) );
  INV_X1 U5479 ( .A(n6645), .ZN(n6639) );
  NAND3_X1 U5480 ( .A1(n4477), .A2(n4476), .A3(n6639), .ZN(n4483) );
  INV_X1 U5481 ( .A(n4478), .ZN(n4479) );
  AOI21_X1 U5482 ( .B1(n6639), .B2(n4525), .A(n4479), .ZN(n4482) );
  INV_X1 U5483 ( .A(n4378), .ZN(n6049) );
  NAND2_X1 U5484 ( .A1(n6049), .A2(n4524), .ZN(n4480) );
  NAND4_X1 U5485 ( .A1(n4483), .A2(n4482), .A3(n4481), .A4(n4480), .ZN(n4484)
         );
  AOI21_X1 U5486 ( .B1(n6640), .B2(n6645), .A(n4484), .ZN(n4619) );
  INV_X1 U5487 ( .A(n4619), .ZN(n6624) );
  INV_X1 U5488 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6069) );
  NAND2_X1 U5489 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .ZN(n4707) );
  INV_X1 U5490 ( .A(n4707), .ZN(n4634) );
  NAND2_X1 U5491 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4634), .ZN(n6753) );
  NOR2_X1 U5492 ( .A1(n6069), .A2(n6753), .ZN(n4485) );
  AOI21_X1 U5493 ( .B1(n6624), .B2(n6672), .A(n4485), .ZN(n6053) );
  NAND2_X1 U5494 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6872), .ZN(n6754) );
  NAND2_X1 U5495 ( .A1(n6053), .A2(n6754), .ZN(n6761) );
  INV_X1 U5496 ( .A(n6761), .ZN(n4514) );
  INV_X1 U5497 ( .A(n4487), .ZN(n4489) );
  AND4_X1 U5498 ( .A1(n4378), .A2(n4084), .A3(n4372), .A4(n4087), .ZN(n4488)
         );
  NAND2_X1 U5499 ( .A1(n4489), .A2(n4488), .ZN(n6621) );
  NAND2_X1 U5500 ( .A1(n4486), .A2(n6621), .ZN(n4494) );
  INV_X1 U5501 ( .A(n4490), .ZN(n4624) );
  INV_X1 U5502 ( .A(n4491), .ZN(n4498) );
  NAND3_X1 U5503 ( .A1(n4492), .A2(n4624), .A3(n4498), .ZN(n4493) );
  OAI211_X1 U5504 ( .C1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n6622), .A(n4494), .B(n4493), .ZN(n6625) );
  AOI22_X1 U5505 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5790), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4155), .ZN(n4510) );
  NOR2_X1 U5506 ( .A1(n5389), .A2(n6757), .ZN(n4508) );
  AOI222_X1 U5507 ( .A1(n6625), .A2(n6050), .B1(n4510), .B2(n4508), .C1(n4495), 
        .C2(n4576), .ZN(n4497) );
  INV_X1 U5508 ( .A(n4576), .ZN(n6664) );
  NOR2_X1 U5509 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6664), .ZN(n6756)
         );
  OAI21_X1 U5510 ( .B1(n4514), .B2(n6756), .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), 
        .ZN(n4496) );
  OAI21_X1 U5511 ( .B1(n4514), .B2(n4497), .A(n4496), .ZN(U3460) );
  AOI21_X1 U5512 ( .B1(n4576), .B2(n4498), .A(n4514), .ZN(n4516) );
  NAND2_X1 U5513 ( .A1(n4499), .A2(n6621), .ZN(n4507) );
  INV_X1 U5514 ( .A(n6640), .ZN(n4501) );
  INV_X1 U5515 ( .A(n4525), .ZN(n4500) );
  NAND2_X1 U5516 ( .A1(n4501), .A2(n4500), .ZN(n4616) );
  XNOR2_X1 U5517 ( .A(n4491), .B(n6925), .ZN(n4502) );
  NAND2_X1 U5518 ( .A1(n4616), .A2(n4502), .ZN(n4506) );
  XNOR2_X1 U5519 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n6925), .ZN(n4503)
         );
  OAI22_X1 U5520 ( .A1(n6622), .A2(n4503), .B1(n4612), .B2(n4502), .ZN(n4504)
         );
  INV_X1 U5521 ( .A(n4504), .ZN(n4505) );
  NAND3_X1 U5522 ( .A1(n4507), .A2(n4506), .A3(n4505), .ZN(n4620) );
  INV_X1 U5523 ( .A(n4508), .ZN(n4511) );
  NAND3_X1 U5524 ( .A1(n4491), .A2(n4576), .A3(n4515), .ZN(n4509) );
  OAI21_X1 U5525 ( .B1(n4511), .B2(n4510), .A(n4509), .ZN(n4512) );
  AOI21_X1 U5526 ( .B1(n4620), .B2(n6050), .A(n4512), .ZN(n4513) );
  OAI22_X1 U5527 ( .A1(n4516), .A2(n4515), .B1(n4514), .B2(n4513), .ZN(U3459)
         );
  NOR2_X1 U5528 ( .A1(n4517), .A2(n4519), .ZN(n6357) );
  INV_X1 U5529 ( .A(n6357), .ZN(n4548) );
  NOR2_X1 U5530 ( .A1(n4520), .A2(READY_N), .ZN(n4521) );
  OR2_X1 U5531 ( .A1(n4523), .A2(n4522), .ZN(n4528) );
  NAND3_X1 U5532 ( .A1(n6049), .A2(n6672), .A3(n4524), .ZN(n4527) );
  NAND2_X1 U5533 ( .A1(n4703), .A2(n4525), .ZN(n4526) );
  NAND2_X1 U5534 ( .A1(n3536), .A2(n3488), .ZN(n4529) );
  INV_X1 U5535 ( .A(n4529), .ZN(n4530) );
  AOI22_X1 U5536 ( .A1(n5414), .A2(DATAI_2_), .B1(n6241), .B2(
        EAX_REG_2__SCAN_IN), .ZN(n4531) );
  OAI21_X1 U5537 ( .B1(n4548), .B2(n5684), .A(n4531), .ZN(U2889) );
  OAI21_X1 U5538 ( .B1(n4517), .B2(n4532), .A(n4555), .ZN(n5137) );
  AOI21_X1 U5539 ( .B1(n4534), .B2(n4533), .A(n4558), .ZN(n6197) );
  INV_X1 U5540 ( .A(n6231), .ZN(n5412) );
  AOI22_X1 U5541 ( .A1(n6227), .A2(n6197), .B1(n5412), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4535) );
  OAI21_X1 U5542 ( .B1(n5137), .B2(n5670), .A(n4535), .ZN(U2856) );
  NOR2_X1 U5543 ( .A1(n4536), .A2(n4537), .ZN(n4538) );
  NOR2_X1 U5544 ( .A1(n3660), .A2(n4538), .ZN(n5609) );
  INV_X1 U5545 ( .A(n5670), .ZN(n6228) );
  XNOR2_X1 U5546 ( .A(n4539), .B(n4540), .ZN(n4565) );
  OAI22_X1 U5547 ( .A1(n5671), .A2(n4565), .B1(n4541), .B2(n6231), .ZN(n4542)
         );
  AOI21_X1 U5548 ( .B1(n5609), .B2(n6228), .A(n4542), .ZN(n4543) );
  INV_X1 U5549 ( .A(n4543), .ZN(U2858) );
  INV_X1 U5550 ( .A(DATAI_3_), .ZN(n6890) );
  INV_X1 U5551 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6315) );
  OAI222_X1 U5552 ( .A1(n5137), .A2(n5684), .B1(n5381), .B2(n6890), .C1(n5467), 
        .C2(n6315), .ZN(U2888) );
  INV_X1 U5553 ( .A(DATAI_0_), .ZN(n4544) );
  INV_X1 U5554 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6949) );
  OAI222_X1 U5555 ( .A1(n6371), .A2(n5684), .B1(n5381), .B2(n4544), .C1(n5467), 
        .C2(n6949), .ZN(U2891) );
  OR2_X1 U5556 ( .A1(n4546), .A2(n4545), .ZN(n4547) );
  NAND2_X1 U5557 ( .A1(n4547), .A2(n4533), .ZN(n6398) );
  OAI222_X1 U5558 ( .A1(n6398), .A2(n5671), .B1(n4549), .B2(n6231), .C1(n5670), 
        .C2(n4548), .ZN(U2857) );
  OAI21_X1 U5559 ( .B1(n4550), .B2(n4552), .A(n4551), .ZN(n6167) );
  AOI21_X1 U5560 ( .B1(n4553), .B2(n4557), .A(n3142), .ZN(n6162) );
  AOI22_X1 U5561 ( .A1(n6227), .A2(n6162), .B1(n5412), .B2(EBX_REG_5__SCAN_IN), 
        .ZN(n4554) );
  OAI21_X1 U5562 ( .B1(n6167), .B2(n5670), .A(n4554), .ZN(U2854) );
  AOI21_X1 U5563 ( .B1(n4556), .B2(n4555), .A(n4550), .ZN(n6189) );
  INV_X1 U5564 ( .A(n6189), .ZN(n4710) );
  OAI21_X1 U5565 ( .B1(n4559), .B2(n4558), .A(n4557), .ZN(n4781) );
  INV_X1 U5566 ( .A(n4781), .ZN(n6185) );
  AOI22_X1 U5567 ( .A1(n6227), .A2(n6185), .B1(n5412), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4560) );
  OAI21_X1 U5568 ( .B1(n4710), .B2(n5670), .A(n4560), .ZN(U2855) );
  OAI21_X1 U5569 ( .B1(n4563), .B2(n4562), .A(n4561), .ZN(n5136) );
  INV_X1 U5570 ( .A(n5136), .ZN(n4568) );
  NOR3_X1 U5571 ( .A1(n5288), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n4564), 
        .ZN(n4567) );
  NAND2_X1 U5572 ( .A1(n6351), .A2(REIP_REG_1__SCAN_IN), .ZN(n5131) );
  OAI21_X1 U5573 ( .B1(n6413), .B2(n4565), .A(n5131), .ZN(n4566) );
  AOI211_X1 U5574 ( .C1(n4568), .C2(n6415), .A(n4567), .B(n4566), .ZN(n4569)
         );
  OAI21_X1 U5575 ( .B1(n4570), .B2(n4155), .A(n4569), .ZN(U3017) );
  INV_X1 U5576 ( .A(n4743), .ZN(n4715) );
  INV_X1 U5577 ( .A(n5030), .ZN(n4641) );
  NAND2_X1 U5578 ( .A1(n6423), .A2(n4641), .ZN(n4827) );
  INV_X1 U5579 ( .A(DATAI_17_), .ZN(n6893) );
  NOR2_X1 U5580 ( .A1(n5989), .A2(n6893), .ZN(n6575) );
  INV_X1 U5581 ( .A(n6575), .ZN(n6797) );
  NAND3_X1 U5582 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n7081), .A3(n7064), .ZN(n4818) );
  NOR2_X1 U5583 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4818), .ZN(n4927)
         );
  INV_X1 U5584 ( .A(n4927), .ZN(n4593) );
  NOR2_X1 U5585 ( .A1(n4583), .A2(n6937), .ZN(n6430) );
  INV_X1 U5586 ( .A(n4718), .ZN(n4575) );
  OR2_X1 U5587 ( .A1(n6424), .A2(n4575), .ZN(n5225) );
  INV_X1 U5588 ( .A(n5225), .ZN(n4577) );
  NAND2_X1 U5589 ( .A1(n5389), .A2(n6937), .ZN(n6677) );
  OAI21_X1 U5590 ( .B1(n4577), .B2(n6937), .A(n4860), .ZN(n5219) );
  AOI211_X1 U5591 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4593), .A(n6430), .B(
        n5219), .ZN(n4582) );
  INV_X1 U5592 ( .A(n4572), .ZN(n5146) );
  NAND3_X1 U5593 ( .A1(n4276), .A2(n5146), .A3(n5030), .ZN(n4642) );
  AND2_X1 U5594 ( .A1(n6520), .A2(n6064), .ZN(n5032) );
  NOR2_X1 U5595 ( .A1(n5030), .A2(n6064), .ZN(n4579) );
  AOI21_X1 U5596 ( .B1(n6423), .B2(n4579), .A(n6564), .ZN(n4821) );
  INV_X1 U5597 ( .A(n4486), .ZN(n5616) );
  AND2_X1 U5598 ( .A1(n4499), .A2(n5616), .ZN(n6557) );
  INV_X1 U5599 ( .A(n4717), .ZN(n6467) );
  AND2_X1 U5600 ( .A1(n6557), .A2(n6467), .ZN(n4817) );
  INV_X1 U5601 ( .A(n4817), .ZN(n4580) );
  OAI211_X1 U5602 ( .C1(n6796), .C2(n5032), .A(n4821), .B(n4580), .ZN(n4581)
         );
  INV_X1 U5603 ( .A(n4934), .ZN(n4591) );
  NAND2_X1 U5604 ( .A1(n4591), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4589) );
  INV_X1 U5605 ( .A(DATAI_1_), .ZN(n4735) );
  OR2_X1 U5606 ( .A1(n5074), .A2(n6564), .ZN(n6428) );
  INV_X1 U5607 ( .A(n6557), .ZN(n4722) );
  AND2_X1 U5608 ( .A1(n4583), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6425) );
  INV_X1 U5609 ( .A(n6425), .ZN(n5076) );
  OAI22_X1 U5610 ( .A1(n6428), .A2(n4722), .B1(n5076), .B2(n5225), .ZN(n4928)
         );
  NOR2_X2 U5611 ( .A1(n4862), .A2(n4585), .ZN(n6574) );
  INV_X1 U5612 ( .A(n6574), .ZN(n6795) );
  INV_X1 U5613 ( .A(DATAI_25_), .ZN(n4586) );
  NOR2_X1 U5614 ( .A1(n5989), .A2(n4586), .ZN(n6573) );
  INV_X1 U5615 ( .A(n6573), .ZN(n6793) );
  OAI22_X1 U5616 ( .A1(n6795), .A2(n4593), .B1(n6793), .B2(n6796), .ZN(n4587)
         );
  AOI21_X1 U5617 ( .B1(n6437), .B2(n4928), .A(n4587), .ZN(n4588) );
  OAI211_X1 U5618 ( .C1(n4865), .C2(n6797), .A(n4589), .B(n4588), .ZN(U3053)
         );
  INV_X1 U5619 ( .A(DATAI_22_), .ZN(n4590) );
  INV_X1 U5620 ( .A(n6604), .ZN(n6457) );
  NAND2_X1 U5621 ( .A1(n4591), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4596) );
  INV_X1 U5622 ( .A(DATAI_6_), .ZN(n4700) );
  NOR2_X2 U5623 ( .A1(n4862), .A2(n3392), .ZN(n6603) );
  INV_X1 U5624 ( .A(n6603), .ZN(n5105) );
  INV_X1 U5625 ( .A(DATAI_30_), .ZN(n4592) );
  NOR2_X1 U5626 ( .A1(n6370), .A2(n4592), .ZN(n6602) );
  INV_X1 U5627 ( .A(n6602), .ZN(n6540) );
  OAI22_X1 U5628 ( .A1(n5105), .A2(n4593), .B1(n6540), .B2(n6796), .ZN(n4594)
         );
  AOI21_X1 U5629 ( .B1(n6454), .B2(n4928), .A(n4594), .ZN(n4595) );
  OAI211_X1 U5630 ( .C1(n4865), .C2(n6457), .A(n4596), .B(n4595), .ZN(U3058)
         );
  INV_X1 U5631 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4603) );
  INV_X1 U5632 ( .A(DATAI_18_), .ZN(n4597) );
  NOR2_X1 U5633 ( .A1(n5989), .A2(n4597), .ZN(n6580) );
  INV_X1 U5634 ( .A(n4865), .ZN(n4931) );
  INV_X1 U5635 ( .A(DATAI_26_), .ZN(n4598) );
  NOR2_X1 U5636 ( .A1(n6370), .A2(n4598), .ZN(n6578) );
  INV_X1 U5637 ( .A(n6578), .ZN(n6526) );
  NAND2_X1 U5638 ( .A1(DATAI_2_), .A2(n4860), .ZN(n6583) );
  NOR2_X2 U5639 ( .A1(n4862), .A2(n4599), .ZN(n6579) );
  AOI22_X1 U5640 ( .A1(n6440), .A2(n4928), .B1(n6579), .B2(n4927), .ZN(n4600)
         );
  OAI21_X1 U5641 ( .B1(n6526), .B2(n6796), .A(n4600), .ZN(n4601) );
  AOI21_X1 U5642 ( .B1(n6580), .B2(n4931), .A(n4601), .ZN(n4602) );
  OAI21_X1 U5643 ( .B1(n4934), .B2(n4603), .A(n4602), .ZN(U3054) );
  NAND2_X1 U5644 ( .A1(n5074), .A2(n6621), .ZN(n4618) );
  MUX2_X1 U5645 ( .A(n4604), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4491), 
        .Z(n4605) );
  NOR2_X1 U5646 ( .A1(n4605), .A2(n4621), .ZN(n4615) );
  NAND2_X1 U5647 ( .A1(n6925), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4607) );
  INV_X1 U5648 ( .A(n4607), .ZN(n4606) );
  MUX2_X1 U5649 ( .A(n4607), .B(n4606), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4613) );
  INV_X1 U5650 ( .A(n4608), .ZN(n4609) );
  OAI21_X1 U5651 ( .B1(n4491), .B2(n3690), .A(n4609), .ZN(n4611) );
  NOR2_X1 U5652 ( .A1(n4611), .A2(n4610), .ZN(n5900) );
  OAI22_X1 U5653 ( .A1(n6622), .A2(n4613), .B1(n5900), .B2(n4612), .ZN(n4614)
         );
  AOI21_X1 U5654 ( .B1(n4616), .B2(n4615), .A(n4614), .ZN(n4617) );
  NAND2_X1 U5655 ( .A1(n4618), .A2(n4617), .ZN(n5899) );
  MUX2_X1 U5656 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5899), .S(n6624), 
        .Z(n6633) );
  MUX2_X1 U5657 ( .A(n4620), .B(n6925), .S(n4619), .Z(n6630) );
  NAND3_X1 U5658 ( .A1(n6633), .A2(n6630), .A3(n5389), .ZN(n4623) );
  AND2_X1 U5659 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6069), .ZN(n4629) );
  NAND2_X1 U5660 ( .A1(n4621), .A2(n4629), .ZN(n4622) );
  NAND2_X1 U5661 ( .A1(n4623), .A2(n4622), .ZN(n6656) );
  NAND2_X1 U5662 ( .A1(n6656), .A2(n4624), .ZN(n4636) );
  OR2_X1 U5663 ( .A1(n4625), .A2(n6467), .ZN(n4626) );
  XNOR2_X1 U5664 ( .A(n4626), .B(n4627), .ZN(n6187) );
  OAI22_X1 U5665 ( .A1(n6187), .A2(n4378), .B1(n4627), .B2(n6624), .ZN(n4628)
         );
  NAND2_X1 U5666 ( .A1(n4628), .A2(n5389), .ZN(n4631) );
  NAND2_X1 U5667 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n4629), .ZN(n4630) );
  NAND2_X1 U5668 ( .A1(n4631), .A2(n4630), .ZN(n6654) );
  NOR2_X1 U5669 ( .A1(n6654), .A2(FLUSH_REG_SCAN_IN), .ZN(n4632) );
  AOI21_X1 U5670 ( .B1(n4636), .B2(n4632), .A(n6753), .ZN(n4633) );
  INV_X1 U5671 ( .A(n6654), .ZN(n4635) );
  NAND3_X1 U5672 ( .A1(n4636), .A2(n4635), .A3(n4634), .ZN(n6671) );
  INV_X1 U5673 ( .A(n6671), .ZN(n4639) );
  INV_X1 U5674 ( .A(n3133), .ZN(n6510) );
  NAND2_X1 U5675 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n3515), .ZN(n4814) );
  INV_X1 U5676 ( .A(n4814), .ZN(n4637) );
  OAI22_X1 U5677 ( .A1(n4578), .A2(n6564), .B1(n6510), .B2(n4637), .ZN(n4638)
         );
  OAI21_X1 U5678 ( .B1(n4639), .B2(n4638), .A(n6420), .ZN(n4640) );
  OAI21_X1 U5679 ( .B1(n6420), .B2(n6556), .A(n4640), .ZN(U3465) );
  NAND3_X1 U5680 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n7081), .A3(n6631), .ZN(n5143) );
  NOR2_X1 U5681 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5143), .ZN(n4935)
         );
  INV_X1 U5682 ( .A(n4935), .ZN(n4646) );
  NAND3_X1 U5683 ( .A1(n4276), .A2(n4641), .A3(n5146), .ZN(n5009) );
  INV_X1 U5684 ( .A(n5009), .ZN(n5005) );
  NAND2_X1 U5685 ( .A1(n5005), .A2(n4574), .ZN(n4647) );
  AOI21_X1 U5686 ( .B1(n4647), .B2(n6792), .A(n5032), .ZN(n4643) );
  INV_X1 U5687 ( .A(n5074), .ZN(n6200) );
  NOR2_X1 U5688 ( .A1(n4499), .A2(n5616), .ZN(n5034) );
  AND2_X1 U5689 ( .A1(n6200), .A2(n5034), .ZN(n5144) );
  OAI21_X1 U5690 ( .B1(n4643), .B2(n5144), .A(n3515), .ZN(n4645) );
  OAI21_X1 U5691 ( .B1(n6424), .B2(n6937), .A(n4860), .ZN(n6429) );
  NOR2_X1 U5692 ( .A1(n6425), .A2(n6429), .ZN(n5036) );
  INV_X1 U5693 ( .A(n5036), .ZN(n4644) );
  INV_X1 U5694 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4653) );
  INV_X1 U5695 ( .A(n6580), .ZN(n6443) );
  INV_X1 U5696 ( .A(n5144), .ZN(n4649) );
  NAND3_X1 U5697 ( .A1(n6430), .A2(n6424), .A3(n7081), .ZN(n4648) );
  OAI21_X1 U5698 ( .B1(n4649), .B2(n6564), .A(n4648), .ZN(n4936) );
  AOI22_X1 U5699 ( .A1(n6440), .A2(n4936), .B1(n6579), .B2(n4935), .ZN(n4650)
         );
  OAI21_X1 U5700 ( .B1(n6443), .B2(n6792), .A(n4650), .ZN(n4651) );
  AOI21_X1 U5701 ( .B1(n6578), .B2(n5201), .A(n4651), .ZN(n4652) );
  OAI21_X1 U5702 ( .B1(n4941), .B2(n4653), .A(n4652), .ZN(U3038) );
  INV_X1 U5703 ( .A(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4660) );
  INV_X1 U5704 ( .A(DATAI_27_), .ZN(n4654) );
  NOR2_X1 U5705 ( .A1(n5989), .A2(n4654), .ZN(n6584) );
  INV_X1 U5706 ( .A(DATAI_19_), .ZN(n4655) );
  NOR2_X1 U5707 ( .A1(n5989), .A2(n4655), .ZN(n6586) );
  INV_X1 U5708 ( .A(n6586), .ZN(n6530) );
  NAND2_X1 U5709 ( .A1(DATAI_3_), .A2(n4860), .ZN(n6589) );
  NOR2_X2 U5710 ( .A1(n4862), .A2(n3531), .ZN(n6585) );
  AOI22_X1 U5711 ( .A1(n6444), .A2(n4936), .B1(n6585), .B2(n4935), .ZN(n4657)
         );
  OAI21_X1 U5712 ( .B1(n6530), .B2(n6792), .A(n4657), .ZN(n4658) );
  AOI21_X1 U5713 ( .B1(n6584), .B2(n5201), .A(n4658), .ZN(n4659) );
  OAI21_X1 U5714 ( .B1(n4941), .B2(n4660), .A(n4659), .ZN(U3039) );
  XNOR2_X1 U5715 ( .A(n4661), .B(n3120), .ZN(n5185) );
  AND2_X1 U5716 ( .A1(n4790), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4664)
         );
  AOI22_X1 U5717 ( .A1(n5335), .A2(n4765), .B1(n6403), .B2(n4663), .ZN(n6408)
         );
  OAI21_X1 U5718 ( .B1(n5288), .B2(n4664), .A(n6408), .ZN(n4794) );
  INV_X1 U5719 ( .A(n4665), .ZN(n4668) );
  OAI211_X1 U5720 ( .C1(n4668), .C2(n4764), .A(n4667), .B(n4666), .ZN(n4669)
         );
  NAND2_X1 U5721 ( .A1(n4794), .A2(n4669), .ZN(n4672) );
  INV_X1 U5722 ( .A(REIP_REG_5__SCAN_IN), .ZN(n4670) );
  NOR2_X1 U5723 ( .A1(n6401), .A2(n4670), .ZN(n5180) );
  AOI21_X1 U5724 ( .B1(n6389), .B2(n6162), .A(n5180), .ZN(n4671) );
  OAI211_X1 U5725 ( .C1(n5185), .C2(n6014), .A(n4672), .B(n4671), .ZN(U3013)
         );
  INV_X1 U5726 ( .A(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4676) );
  INV_X1 U5727 ( .A(n6584), .ZN(n5163) );
  AOI22_X1 U5728 ( .A1(n6444), .A2(n4928), .B1(n6585), .B2(n4927), .ZN(n4673)
         );
  OAI21_X1 U5729 ( .B1(n5163), .B2(n6796), .A(n4673), .ZN(n4674) );
  AOI21_X1 U5730 ( .B1(n6586), .B2(n4931), .A(n4674), .ZN(n4675) );
  OAI21_X1 U5731 ( .B1(n4934), .B2(n4676), .A(n4675), .ZN(U3055) );
  NAND2_X1 U5732 ( .A1(n4551), .A2(n4678), .ZN(n4679) );
  NAND2_X1 U5733 ( .A1(n4677), .A2(n4679), .ZN(n6157) );
  OR2_X1 U5734 ( .A1(n4680), .A2(n3142), .ZN(n4681) );
  NAND2_X1 U5735 ( .A1(n4681), .A2(n4799), .ZN(n4791) );
  INV_X1 U5736 ( .A(n4791), .ZN(n6149) );
  AOI22_X1 U5737 ( .A1(n6227), .A2(n6149), .B1(n5412), .B2(EBX_REG_6__SCAN_IN), 
        .ZN(n4682) );
  OAI21_X1 U5738 ( .B1(n6157), .B2(n5670), .A(n4682), .ZN(U2853) );
  INV_X1 U5739 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4687) );
  INV_X1 U5740 ( .A(DATAI_16_), .ZN(n6968) );
  NOR2_X1 U5741 ( .A1(n5989), .A2(n6968), .ZN(n6569) );
  INV_X1 U5742 ( .A(DATAI_24_), .ZN(n4683) );
  NOR2_X1 U5743 ( .A1(n5989), .A2(n4683), .ZN(n6561) );
  INV_X1 U5744 ( .A(n6561), .ZN(n5194) );
  NAND2_X1 U5745 ( .A1(DATAI_0_), .A2(n4860), .ZN(n6572) );
  NOR2_X2 U5746 ( .A1(n4862), .A2(n5400), .ZN(n6562) );
  AOI22_X1 U5747 ( .A1(n6498), .A2(n4928), .B1(n6562), .B2(n4927), .ZN(n4684)
         );
  OAI21_X1 U5748 ( .B1(n5194), .B2(n6796), .A(n4684), .ZN(n4685) );
  AOI21_X1 U5749 ( .B1(n6569), .B2(n4931), .A(n4685), .ZN(n4686) );
  OAI21_X1 U5750 ( .B1(n4934), .B2(n4687), .A(n4686), .ZN(U3052) );
  INV_X1 U5751 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4691) );
  INV_X1 U5752 ( .A(n6569), .ZN(n6436) );
  AOI22_X1 U5753 ( .A1(n6498), .A2(n4936), .B1(n6562), .B2(n4935), .ZN(n4688)
         );
  OAI21_X1 U5754 ( .B1(n6436), .B2(n6792), .A(n4688), .ZN(n4689) );
  AOI21_X1 U5755 ( .B1(n6561), .B2(n5201), .A(n4689), .ZN(n4690) );
  OAI21_X1 U5756 ( .B1(n4941), .B2(n4691), .A(n4690), .ZN(U3036) );
  INV_X1 U5757 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4695) );
  NOR2_X1 U5758 ( .A1(n6792), .A2(n6797), .ZN(n4692) );
  AOI21_X1 U5759 ( .B1(n6574), .B2(n4935), .A(n4692), .ZN(n4694) );
  AOI22_X1 U5760 ( .A1(n6437), .A2(n4936), .B1(n6573), .B2(n5201), .ZN(n4693)
         );
  OAI211_X1 U5761 ( .C1(n4941), .C2(n4695), .A(n4694), .B(n4693), .ZN(U3037)
         );
  INV_X1 U5762 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4699) );
  NOR2_X1 U5763 ( .A1(n6792), .A2(n6457), .ZN(n4696) );
  AOI21_X1 U5764 ( .B1(n6603), .B2(n4935), .A(n4696), .ZN(n4698) );
  AOI22_X1 U5765 ( .A1(n6454), .A2(n4936), .B1(n6602), .B2(n5201), .ZN(n4697)
         );
  OAI211_X1 U5766 ( .C1(n4941), .C2(n4699), .A(n4698), .B(n4697), .ZN(U3042)
         );
  INV_X1 U5767 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6324) );
  OAI222_X1 U5768 ( .A1(n6157), .A2(n5684), .B1(n5381), .B2(n4700), .C1(n5467), 
        .C2(n6324), .ZN(U2885) );
  INV_X1 U5769 ( .A(EAX_REG_17__SCAN_IN), .ZN(n6269) );
  INV_X1 U5770 ( .A(n4703), .ZN(n4704) );
  OAI21_X1 U5771 ( .B1(n4704), .B2(n6622), .A(n6348), .ZN(n4706) );
  NOR2_X1 U5772 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4707), .ZN(n5128) );
  INV_X1 U5773 ( .A(n5128), .ZN(n6659) );
  AOI22_X1 U5774 ( .A1(DATAO_REG_17__SCAN_IN), .A2(n6260), .B1(n6779), .B2(
        UWORD_REG_1__SCAN_IN), .ZN(n4708) );
  OAI21_X1 U5775 ( .B1(n6269), .B2(n5130), .A(n4708), .ZN(U2906) );
  AOI22_X1 U5776 ( .A1(n5414), .A2(DATAI_4_), .B1(n6241), .B2(
        EAX_REG_4__SCAN_IN), .ZN(n4709) );
  OAI21_X1 U5777 ( .B1(n4710), .B2(n5684), .A(n4709), .ZN(U2887) );
  INV_X1 U5778 ( .A(EAX_REG_25__SCAN_IN), .ZN(n6288) );
  AOI22_X1 U5779 ( .A1(UWORD_REG_9__SCAN_IN), .A2(n5128), .B1(n6260), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4711) );
  OAI21_X1 U5780 ( .B1(n6288), .B2(n5130), .A(n4711), .ZN(U2898) );
  INV_X1 U5781 ( .A(EAX_REG_29__SCAN_IN), .ZN(n6300) );
  AOI22_X1 U5782 ( .A1(UWORD_REG_13__SCAN_IN), .A2(n5128), .B1(n6260), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4712) );
  OAI21_X1 U5783 ( .B1(n6300), .B2(n5130), .A(n4712), .ZN(U2894) );
  INV_X1 U5784 ( .A(EAX_REG_27__SCAN_IN), .ZN(n6294) );
  AOI22_X1 U5785 ( .A1(n6779), .A2(UWORD_REG_11__SCAN_IN), .B1(n6260), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4713) );
  OAI21_X1 U5786 ( .B1(n6294), .B2(n5130), .A(n4713), .ZN(U2896) );
  AND2_X1 U5787 ( .A1(n5030), .A2(n4574), .ZN(n5072) );
  INV_X1 U5788 ( .A(n5072), .ZN(n4714) );
  NOR2_X1 U5789 ( .A1(n5030), .A2(n4715), .ZN(n4716) );
  OAI21_X1 U5790 ( .B1(n6543), .B2(n6612), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4721) );
  AOI21_X1 U5791 ( .B1(n6557), .B2(n4717), .A(n6564), .ZN(n4720) );
  NOR3_X1 U5792 ( .A1(n6631), .A2(n7081), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n6560) );
  INV_X1 U5793 ( .A(n6560), .ZN(n6563) );
  NOR2_X1 U5794 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6563), .ZN(n4942)
         );
  OR2_X1 U5795 ( .A1(n6424), .A2(n4718), .ZN(n5080) );
  AOI21_X1 U5796 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5080), .A(n4819), .ZN(
        n5071) );
  INV_X1 U5797 ( .A(n6430), .ZN(n5226) );
  OAI211_X1 U5798 ( .C1(n4942), .C2(n3515), .A(n5071), .B(n5226), .ZN(n4719)
         );
  INV_X1 U5799 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n7032) );
  INV_X1 U5800 ( .A(n6612), .ZN(n4945) );
  NOR2_X1 U5801 ( .A1(n6200), .A2(n6564), .ZN(n5083) );
  INV_X1 U5802 ( .A(n5083), .ZN(n4723) );
  OAI22_X1 U5803 ( .A1(n4723), .A2(n4722), .B1(n5080), .B2(n5076), .ZN(n4943)
         );
  AOI22_X1 U5804 ( .A1(n6498), .A2(n4943), .B1(n6562), .B2(n4942), .ZN(n4724)
         );
  OAI21_X1 U5805 ( .B1(n6436), .B2(n4945), .A(n4724), .ZN(n4725) );
  AOI21_X1 U5806 ( .B1(n6561), .B2(n6543), .A(n4725), .ZN(n4726) );
  OAI21_X1 U5807 ( .B1(n4949), .B2(n7032), .A(n4726), .ZN(U3116) );
  INV_X1 U5808 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4730) );
  AOI22_X1 U5809 ( .A1(n6440), .A2(n4943), .B1(n6579), .B2(n4942), .ZN(n4727)
         );
  OAI21_X1 U5810 ( .B1(n6443), .B2(n4945), .A(n4727), .ZN(n4728) );
  AOI21_X1 U5811 ( .B1(n6578), .B2(n6543), .A(n4728), .ZN(n4729) );
  OAI21_X1 U5812 ( .B1(n4949), .B2(n4730), .A(n4729), .ZN(U3118) );
  INV_X1 U5813 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4734) );
  AOI22_X1 U5814 ( .A1(n6444), .A2(n4943), .B1(n6585), .B2(n4942), .ZN(n4731)
         );
  OAI21_X1 U5815 ( .B1(n6530), .B2(n4945), .A(n4731), .ZN(n4732) );
  AOI21_X1 U5816 ( .B1(n6584), .B2(n6543), .A(n4732), .ZN(n4733) );
  OAI21_X1 U5817 ( .B1(n4949), .B2(n4734), .A(n4733), .ZN(U3119) );
  INV_X1 U5818 ( .A(n5609), .ZN(n4736) );
  INV_X1 U5819 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6309) );
  OAI222_X1 U5820 ( .A1(n4736), .A2(n5684), .B1(n5381), .B2(n4735), .C1(n5467), 
        .C2(n6309), .ZN(U2890) );
  INV_X1 U5821 ( .A(DATAI_5_), .ZN(n7016) );
  INV_X1 U5822 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6321) );
  OAI222_X1 U5823 ( .A1(n6167), .A2(n5684), .B1(n5381), .B2(n7016), .C1(n5467), 
        .C2(n6321), .ZN(U2886) );
  INV_X1 U5824 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4739) );
  AOI22_X1 U5825 ( .A1(n6437), .A2(n4943), .B1(n6573), .B2(n6543), .ZN(n4738)
         );
  AOI22_X1 U5826 ( .A1(n6574), .A2(n4942), .B1(n6575), .B2(n6612), .ZN(n4737)
         );
  OAI211_X1 U5827 ( .C1(n4949), .C2(n4739), .A(n4738), .B(n4737), .ZN(U3117)
         );
  INV_X1 U5828 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4742) );
  AOI22_X1 U5829 ( .A1(n6454), .A2(n4943), .B1(n6602), .B2(n6543), .ZN(n4741)
         );
  AOI22_X1 U5830 ( .A1(n6603), .A2(n4942), .B1(n6604), .B2(n6612), .ZN(n4740)
         );
  OAI211_X1 U5831 ( .C1(n4949), .C2(n4742), .A(n4741), .B(n4740), .ZN(U3122)
         );
  NAND3_X1 U5832 ( .A1(n4572), .A2(n4743), .A3(n5030), .ZN(n4953) );
  INV_X1 U5833 ( .A(n4953), .ZN(n4950) );
  OR2_X1 U5834 ( .A1(n6430), .A2(n6429), .ZN(n4749) );
  AND2_X1 U5835 ( .A1(n4499), .A2(n4486), .ZN(n6468) );
  NOR2_X1 U5836 ( .A1(n6468), .A2(n6564), .ZN(n6432) );
  INV_X1 U5837 ( .A(n6432), .ZN(n4745) );
  INV_X1 U5838 ( .A(n6608), .ZN(n4758) );
  AOI21_X1 U5839 ( .B1(n4758), .B2(n5003), .A(n6064), .ZN(n4744) );
  AOI21_X1 U5840 ( .B1(n6428), .B2(n4745), .A(n4744), .ZN(n4748) );
  INV_X1 U5841 ( .A(n4955), .ZN(n4746) );
  NOR2_X1 U5842 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4746), .ZN(n4771)
         );
  NAND2_X1 U5843 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n7081), .ZN(n5035) );
  OAI21_X1 U5844 ( .B1(n3515), .B2(n4771), .A(n5035), .ZN(n4747) );
  NAND2_X1 U5845 ( .A1(n4972), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4753)
         );
  NOR2_X1 U5846 ( .A1(n5076), .A2(n7081), .ZN(n4750) );
  AOI22_X1 U5847 ( .A1(n5083), .A2(n6468), .B1(n6424), .B2(n4750), .ZN(n4974)
         );
  INV_X1 U5848 ( .A(n6579), .ZN(n5089) );
  INV_X1 U5849 ( .A(n4771), .ZN(n4973) );
  OAI22_X1 U5850 ( .A1(n6583), .A2(n4974), .B1(n5089), .B2(n4973), .ZN(n4751)
         );
  AOI21_X1 U5851 ( .B1(n6578), .B2(n6608), .A(n4751), .ZN(n4752) );
  OAI211_X1 U5852 ( .C1(n5003), .C2(n6443), .A(n4753), .B(n4752), .ZN(U3134)
         );
  NAND2_X1 U5853 ( .A1(n4972), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4756)
         );
  INV_X1 U5854 ( .A(n6562), .ZN(n5096) );
  OAI22_X1 U5855 ( .A1(n6572), .A2(n4974), .B1(n5096), .B2(n4973), .ZN(n4754)
         );
  AOI21_X1 U5856 ( .B1(n6561), .B2(n6608), .A(n4754), .ZN(n4755) );
  OAI211_X1 U5857 ( .C1(n5003), .C2(n6436), .A(n4756), .B(n4755), .ZN(U3132)
         );
  INV_X1 U5858 ( .A(n4972), .ZN(n4776) );
  INV_X1 U5859 ( .A(n5003), .ZN(n4986) );
  INV_X1 U5860 ( .A(n4974), .ZN(n4772) );
  AOI22_X1 U5861 ( .A1(n6444), .A2(n4772), .B1(n6585), .B2(n4771), .ZN(n4757)
         );
  OAI21_X1 U5862 ( .B1(n5163), .B2(n4758), .A(n4757), .ZN(n4759) );
  AOI21_X1 U5863 ( .B1(n6586), .B2(n4986), .A(n4759), .ZN(n4760) );
  OAI21_X1 U5864 ( .B1(n4776), .B2(n4761), .A(n4760), .ZN(U3135) );
  XNOR2_X1 U5865 ( .A(n4762), .B(n4763), .ZN(n5142) );
  OAI21_X1 U5866 ( .B1(n6403), .B2(n6399), .A(n6408), .ZN(n4784) );
  OAI21_X1 U5867 ( .B1(n4765), .B2(n4764), .A(n6403), .ZN(n4789) );
  AND2_X1 U5868 ( .A1(n6399), .A2(n4789), .ZN(n4780) );
  AOI22_X1 U5869 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n4784), .B1(n4780), 
        .B2(n7057), .ZN(n4767) );
  INV_X1 U5870 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6204) );
  NOR2_X1 U5871 ( .A1(n6401), .A2(n6204), .ZN(n5138) );
  AOI21_X1 U5872 ( .B1(n6389), .B2(n6197), .A(n5138), .ZN(n4766) );
  OAI211_X1 U5873 ( .C1(n5142), .C2(n6014), .A(n4767), .B(n4766), .ZN(U3015)
         );
  INV_X1 U5874 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4770) );
  AOI22_X1 U5875 ( .A1(n6574), .A2(n4771), .B1(n6573), .B2(n6608), .ZN(n4769)
         );
  AOI22_X1 U5876 ( .A1(n6437), .A2(n4772), .B1(n6575), .B2(n4986), .ZN(n4768)
         );
  OAI211_X1 U5877 ( .C1(n4776), .C2(n4770), .A(n4769), .B(n4768), .ZN(U3133)
         );
  INV_X1 U5878 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4775) );
  AOI22_X1 U5879 ( .A1(n6603), .A2(n4771), .B1(n6602), .B2(n6608), .ZN(n4774)
         );
  AOI22_X1 U5880 ( .A1(n6454), .A2(n4772), .B1(n6604), .B2(n4986), .ZN(n4773)
         );
  OAI211_X1 U5881 ( .C1(n4776), .C2(n4775), .A(n4774), .B(n4773), .ZN(U3138)
         );
  XNOR2_X1 U5882 ( .A(n4777), .B(n4778), .ZN(n5298) );
  OAI211_X1 U5883 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4780), .B(n4779), .ZN(n4786) );
  INV_X1 U5884 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6706) );
  NOR2_X1 U5885 ( .A1(n6401), .A2(n6706), .ZN(n4783) );
  NOR2_X1 U5886 ( .A1(n6413), .A2(n4781), .ZN(n4782) );
  AOI211_X1 U5887 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n4784), .A(n4783), 
        .B(n4782), .ZN(n4785) );
  OAI211_X1 U5888 ( .C1(n6014), .C2(n5298), .A(n4786), .B(n4785), .ZN(U3014)
         );
  XNOR2_X1 U5889 ( .A(n4788), .B(n4787), .ZN(n5282) );
  NAND3_X1 U5890 ( .A1(n4790), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n4789), 
        .ZN(n5207) );
  NOR2_X1 U5891 ( .A1(n5207), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4793)
         );
  NAND2_X1 U5892 ( .A1(n6368), .A2(REIP_REG_6__SCAN_IN), .ZN(n5277) );
  OAI21_X1 U5893 ( .B1(n6413), .B2(n4791), .A(n5277), .ZN(n4792) );
  AOI211_X1 U5894 ( .C1(n4794), .C2(INSTADDRPOINTER_REG_6__SCAN_IN), .A(n4793), 
        .B(n4792), .ZN(n4795) );
  OAI21_X1 U5895 ( .B1(n6014), .B2(n5282), .A(n4795), .ZN(U3012) );
  OAI21_X1 U5896 ( .B1(n3767), .B2(n4798), .A(n4797), .ZN(n6141) );
  AOI21_X1 U5897 ( .B1(n4800), .B2(n4799), .A(n4899), .ZN(n6388) );
  AOI22_X1 U5898 ( .A1(n6227), .A2(n6388), .B1(n5412), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n4801) );
  OAI21_X1 U5899 ( .B1(n6141), .B2(n5670), .A(n4801), .ZN(U2852) );
  INV_X1 U5900 ( .A(n6420), .ZN(n4811) );
  NOR2_X1 U5901 ( .A1(n4811), .A2(n6564), .ZN(n4813) );
  INV_X1 U5902 ( .A(n6508), .ZN(n4812) );
  XNOR2_X1 U5903 ( .A(n4572), .B(n4812), .ZN(n4802) );
  NAND2_X1 U5904 ( .A1(n4813), .A2(n4802), .ZN(n4804) );
  NAND3_X1 U5905 ( .A1(n6420), .A2(n4814), .A3(n4499), .ZN(n4803) );
  OAI211_X1 U5906 ( .C1(n6420), .C2(n6631), .A(n4804), .B(n4803), .ZN(U3463)
         );
  INV_X1 U5907 ( .A(n6423), .ZN(n4805) );
  NOR2_X1 U5908 ( .A1(n4805), .A2(n4812), .ZN(n6466) );
  INV_X1 U5909 ( .A(n4276), .ZN(n4806) );
  AOI222_X1 U5910 ( .A1(n5074), .A2(n4814), .B1(n6520), .B2(n6466), .C1(n5032), 
        .C2(n4806), .ZN(n4810) );
  INV_X1 U5911 ( .A(n5031), .ZN(n6509) );
  NOR2_X1 U5912 ( .A1(n6509), .A2(n6555), .ZN(n5147) );
  INV_X1 U5913 ( .A(n5147), .ZN(n4808) );
  AOI22_X1 U5914 ( .A1(n4813), .A2(n4808), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n4811), .ZN(n4809) );
  OAI21_X1 U5915 ( .B1(n4811), .B2(n4810), .A(n4809), .ZN(U3462) );
  OAI211_X1 U5916 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n5030), .A(n4813), .B(
        n4812), .ZN(n4816) );
  NAND3_X1 U5917 ( .A1(n6420), .A2(n4486), .A3(n4814), .ZN(n4815) );
  OAI211_X1 U5918 ( .C1(n6420), .C2(n7064), .A(n4816), .B(n4815), .ZN(U3464)
         );
  INV_X1 U5919 ( .A(DATAI_7_), .ZN(n6991) );
  OAI222_X1 U5920 ( .A1(n6141), .A2(n5684), .B1(n5381), .B2(n6991), .C1(n5467), 
        .C2(n3763), .ZN(U2884) );
  NOR2_X1 U5921 ( .A1(n6556), .A2(n4818), .ZN(n4863) );
  AOI21_X1 U5922 ( .B1(n4817), .B2(n3133), .A(n4863), .ZN(n4822) );
  INV_X1 U5923 ( .A(n4818), .ZN(n4824) );
  OAI21_X1 U5924 ( .B1(n6520), .B2(n4824), .A(n6568), .ZN(n4820) );
  INV_X1 U5925 ( .A(n4821), .ZN(n4823) );
  OR2_X1 U5926 ( .A1(n4823), .A2(n4822), .ZN(n4826) );
  NAND2_X1 U5927 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n4824), .ZN(n4825) );
  NAND2_X1 U5928 ( .A1(n4826), .A2(n4825), .ZN(n4867) );
  NOR2_X2 U5929 ( .A1(n4827), .A2(n4578), .ZN(n6461) );
  AOI22_X1 U5930 ( .A1(n6574), .A2(n4863), .B1(n6575), .B2(n6461), .ZN(n4828)
         );
  OAI21_X1 U5931 ( .B1(n6793), .B2(n4865), .A(n4828), .ZN(n4829) );
  AOI21_X1 U5932 ( .B1(n6437), .B2(n4867), .A(n4829), .ZN(n4830) );
  OAI21_X1 U5933 ( .B1(n4870), .B2(n6859), .A(n4830), .ZN(U3061) );
  INV_X1 U5934 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4834) );
  AOI22_X1 U5935 ( .A1(n6603), .A2(n4863), .B1(n6604), .B2(n6461), .ZN(n4831)
         );
  OAI21_X1 U5936 ( .B1(n6540), .B2(n4865), .A(n4831), .ZN(n4832) );
  AOI21_X1 U5937 ( .B1(n6454), .B2(n4867), .A(n4832), .ZN(n4833) );
  OAI21_X1 U5938 ( .B1(n4870), .B2(n4834), .A(n4833), .ZN(U3066) );
  INV_X1 U5939 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4838) );
  AOI22_X1 U5940 ( .A1(n6562), .A2(n4863), .B1(n6461), .B2(n6569), .ZN(n4835)
         );
  OAI21_X1 U5941 ( .B1(n5194), .B2(n4865), .A(n4835), .ZN(n4836) );
  AOI21_X1 U5942 ( .B1(n6498), .B2(n4867), .A(n4836), .ZN(n4837) );
  OAI21_X1 U5943 ( .B1(n4870), .B2(n4838), .A(n4837), .ZN(U3060) );
  INV_X1 U5944 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4842) );
  AOI22_X1 U5945 ( .A1(n6579), .A2(n4863), .B1(n6580), .B2(n6461), .ZN(n4839)
         );
  OAI21_X1 U5946 ( .B1(n6526), .B2(n4865), .A(n4839), .ZN(n4840) );
  AOI21_X1 U5947 ( .B1(n6440), .B2(n4867), .A(n4840), .ZN(n4841) );
  OAI21_X1 U5948 ( .B1(n4870), .B2(n4842), .A(n4841), .ZN(U3062) );
  INV_X1 U5949 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4846) );
  AOI22_X1 U5950 ( .A1(n6585), .A2(n4863), .B1(n6586), .B2(n6461), .ZN(n4843)
         );
  OAI21_X1 U5951 ( .B1(n5163), .B2(n4865), .A(n4843), .ZN(n4844) );
  AOI21_X1 U5952 ( .B1(n6444), .B2(n4867), .A(n4844), .ZN(n4845) );
  OAI21_X1 U5953 ( .B1(n4870), .B2(n4846), .A(n4845), .ZN(U3063) );
  INV_X1 U5954 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4853) );
  NAND2_X1 U5955 ( .A1(DATAI_4_), .A2(n4860), .ZN(n6595) );
  INV_X1 U5956 ( .A(DATAI_28_), .ZN(n4847) );
  NOR2_X1 U5957 ( .A1(n5989), .A2(n4847), .ZN(n6592) );
  INV_X1 U5958 ( .A(n6592), .ZN(n6534) );
  NOR2_X2 U5959 ( .A1(n4862), .A2(n4848), .ZN(n6591) );
  INV_X1 U5960 ( .A(DATAI_20_), .ZN(n4849) );
  NOR2_X1 U5961 ( .A1(n5989), .A2(n4849), .ZN(n6590) );
  AOI22_X1 U5962 ( .A1(n6591), .A2(n4863), .B1(n6590), .B2(n6461), .ZN(n4850)
         );
  OAI21_X1 U5963 ( .B1(n6534), .B2(n4865), .A(n4850), .ZN(n4851) );
  AOI21_X1 U5964 ( .B1(n6447), .B2(n4867), .A(n4851), .ZN(n4852) );
  OAI21_X1 U5965 ( .B1(n4870), .B2(n4853), .A(n4852), .ZN(U3064) );
  INV_X1 U5966 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4859) );
  NAND2_X1 U5967 ( .A1(DATAI_7_), .A2(n4860), .ZN(n6617) );
  INV_X1 U5968 ( .A(DATAI_31_), .ZN(n4854) );
  NOR2_X1 U5969 ( .A1(n6370), .A2(n4854), .ZN(n6613) );
  INV_X1 U5970 ( .A(n6613), .ZN(n5170) );
  NOR2_X2 U5971 ( .A1(n4862), .A2(n4148), .ZN(n6611) );
  INV_X1 U5972 ( .A(DATAI_23_), .ZN(n4855) );
  NOR2_X1 U5973 ( .A1(n6370), .A2(n4855), .ZN(n6609) );
  AOI22_X1 U5974 ( .A1(n6611), .A2(n4863), .B1(n6609), .B2(n6461), .ZN(n4856)
         );
  OAI21_X1 U5975 ( .B1(n5170), .B2(n4865), .A(n4856), .ZN(n4857) );
  AOI21_X1 U5976 ( .B1(n6460), .B2(n4867), .A(n4857), .ZN(n4858) );
  OAI21_X1 U5977 ( .B1(n4870), .B2(n4859), .A(n4858), .ZN(U3067) );
  INV_X1 U5978 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4869) );
  NAND2_X1 U5979 ( .A1(DATAI_5_), .A2(n4860), .ZN(n6601) );
  INV_X1 U5980 ( .A(DATAI_29_), .ZN(n4861) );
  NOR2_X1 U5981 ( .A1(n6370), .A2(n4861), .ZN(n6596) );
  INV_X1 U5982 ( .A(n6596), .ZN(n5187) );
  NOR2_X2 U5983 ( .A1(n4862), .A2(n5455), .ZN(n6597) );
  NAND2_X1 U5984 ( .A1(n6356), .A2(DATAI_21_), .ZN(n6453) );
  INV_X1 U5985 ( .A(n6453), .ZN(n6598) );
  AOI22_X1 U5986 ( .A1(n6597), .A2(n4863), .B1(n6461), .B2(n6598), .ZN(n4864)
         );
  OAI21_X1 U5987 ( .B1(n5187), .B2(n4865), .A(n4864), .ZN(n4866) );
  AOI21_X1 U5988 ( .B1(n6503), .B2(n4867), .A(n4866), .ZN(n4868) );
  OAI21_X1 U5989 ( .B1(n4870), .B2(n4869), .A(n4868), .ZN(U3065) );
  INV_X1 U5990 ( .A(n4876), .ZN(n4871) );
  OAI21_X1 U5991 ( .B1(n4871), .B2(n6064), .A(n6520), .ZN(n4875) );
  AND2_X1 U5992 ( .A1(n5074), .A2(n3133), .ZN(n6558) );
  OR2_X1 U5993 ( .A1(n4499), .A2(n4486), .ZN(n5227) );
  NAND3_X1 U5994 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6631), .A3(n7064), .ZN(n5075) );
  NOR2_X1 U5995 ( .A1(n6556), .A2(n5075), .ZN(n4893) );
  AOI21_X1 U5996 ( .B1(n6558), .B2(n5082), .A(n4893), .ZN(n4874) );
  INV_X1 U5997 ( .A(n4874), .ZN(n4873) );
  NAND2_X1 U5998 ( .A1(n6564), .A2(n5075), .ZN(n4872) );
  OAI211_X1 U5999 ( .C1(n4875), .C2(n4873), .A(n6568), .B(n4872), .ZN(n4892)
         );
  OAI22_X1 U6000 ( .A1(n4875), .A2(n4874), .B1(n6937), .B2(n5075), .ZN(n4891)
         );
  AOI22_X1 U6001 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4892), .B1(n6444), 
        .B2(n4891), .ZN(n4878) );
  NAND2_X1 U6002 ( .A1(n4876), .A2(n4574), .ZN(n5063) );
  AOI22_X1 U6003 ( .A1(n6502), .A2(n6586), .B1(n6585), .B2(n4893), .ZN(n4877)
         );
  OAI211_X1 U6004 ( .C1(n5163), .C2(n5121), .A(n4878), .B(n4877), .ZN(U3095)
         );
  AOI22_X1 U6005 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4892), .B1(n6503), 
        .B2(n4891), .ZN(n4880) );
  AOI22_X1 U6006 ( .A1(n6502), .A2(n6598), .B1(n6597), .B2(n4893), .ZN(n4879)
         );
  OAI211_X1 U6007 ( .C1(n5187), .C2(n5121), .A(n4880), .B(n4879), .ZN(U3097)
         );
  AOI22_X1 U6008 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4892), .B1(n6498), 
        .B2(n4891), .ZN(n4882) );
  AOI22_X1 U6009 ( .A1(n6502), .A2(n6569), .B1(n6562), .B2(n4893), .ZN(n4881)
         );
  OAI211_X1 U6010 ( .C1(n5194), .C2(n5121), .A(n4882), .B(n4881), .ZN(U3092)
         );
  AOI22_X1 U6011 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4892), .B1(n6440), 
        .B2(n4891), .ZN(n4884) );
  AOI22_X1 U6012 ( .A1(n6502), .A2(n6580), .B1(n6579), .B2(n4893), .ZN(n4883)
         );
  OAI211_X1 U6013 ( .C1(n6526), .C2(n5121), .A(n4884), .B(n4883), .ZN(U3094)
         );
  AOI22_X1 U6014 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4892), .B1(n6437), 
        .B2(n4891), .ZN(n4886) );
  AOI22_X1 U6015 ( .A1(n6502), .A2(n6575), .B1(n6574), .B2(n4893), .ZN(n4885)
         );
  OAI211_X1 U6016 ( .C1(n6793), .C2(n5121), .A(n4886), .B(n4885), .ZN(U3093)
         );
  AOI22_X1 U6017 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4892), .B1(n6454), 
        .B2(n4891), .ZN(n4888) );
  AOI22_X1 U6018 ( .A1(n6502), .A2(n6604), .B1(n6603), .B2(n4893), .ZN(n4887)
         );
  OAI211_X1 U6019 ( .C1(n6540), .C2(n5121), .A(n4888), .B(n4887), .ZN(U3098)
         );
  AOI22_X1 U6020 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4892), .B1(n6447), 
        .B2(n4891), .ZN(n4890) );
  AOI22_X1 U6021 ( .A1(n6502), .A2(n6590), .B1(n6591), .B2(n4893), .ZN(n4889)
         );
  OAI211_X1 U6022 ( .C1(n6534), .C2(n5121), .A(n4890), .B(n4889), .ZN(U3096)
         );
  AOI22_X1 U6023 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4892), .B1(n6460), 
        .B2(n4891), .ZN(n4895) );
  AOI22_X1 U6024 ( .A1(n6502), .A2(n6609), .B1(n6611), .B2(n4893), .ZN(n4894)
         );
  OAI211_X1 U6025 ( .C1(n5170), .C2(n5121), .A(n4895), .B(n4894), .ZN(U3099)
         );
  AOI21_X1 U6026 ( .B1(n4897), .B2(n4797), .A(n4896), .ZN(n4898) );
  INV_X1 U6027 ( .A(n4898), .ZN(n5604) );
  OR2_X1 U6028 ( .A1(n4900), .A2(n4899), .ZN(n4901) );
  NAND2_X1 U6029 ( .A1(n4901), .A2(n5177), .ZN(n5209) );
  INV_X1 U6030 ( .A(n5209), .ZN(n5602) );
  AOI22_X1 U6031 ( .A1(n6227), .A2(n5602), .B1(n5412), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n4902) );
  OAI21_X1 U6032 ( .B1(n5604), .B2(n5670), .A(n4902), .ZN(U2851) );
  AOI22_X1 U6033 ( .A1(n5414), .A2(DATAI_8_), .B1(n6241), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n4903) );
  OAI21_X1 U6034 ( .B1(n5604), .B2(n5684), .A(n4903), .ZN(U2883) );
  INV_X1 U6035 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4907) );
  AOI22_X1 U6036 ( .A1(n6503), .A2(n4928), .B1(n6597), .B2(n4927), .ZN(n4904)
         );
  OAI21_X1 U6037 ( .B1(n5187), .B2(n6796), .A(n4904), .ZN(n4905) );
  AOI21_X1 U6038 ( .B1(n6598), .B2(n4931), .A(n4905), .ZN(n4906) );
  OAI21_X1 U6039 ( .B1(n4934), .B2(n4907), .A(n4906), .ZN(U3057) );
  INV_X1 U6040 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n7029) );
  INV_X1 U6041 ( .A(n6590), .ZN(n6450) );
  AOI22_X1 U6042 ( .A1(n6447), .A2(n4943), .B1(n6591), .B2(n4942), .ZN(n4908)
         );
  OAI21_X1 U6043 ( .B1(n6450), .B2(n4945), .A(n4908), .ZN(n4909) );
  AOI21_X1 U6044 ( .B1(n6592), .B2(n6543), .A(n4909), .ZN(n4910) );
  OAI21_X1 U6045 ( .B1(n4949), .B2(n7029), .A(n4910), .ZN(U3120) );
  INV_X1 U6046 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4914) );
  AOI22_X1 U6047 ( .A1(n6447), .A2(n4936), .B1(n6591), .B2(n4935), .ZN(n4911)
         );
  OAI21_X1 U6048 ( .B1(n6450), .B2(n6792), .A(n4911), .ZN(n4912) );
  AOI21_X1 U6049 ( .B1(n6592), .B2(n5201), .A(n4912), .ZN(n4913) );
  OAI21_X1 U6050 ( .B1(n4941), .B2(n4914), .A(n4913), .ZN(U3040) );
  INV_X1 U6051 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4918) );
  INV_X1 U6052 ( .A(n6609), .ZN(n6546) );
  AOI22_X1 U6053 ( .A1(n6460), .A2(n4936), .B1(n6611), .B2(n4935), .ZN(n4915)
         );
  OAI21_X1 U6054 ( .B1(n6546), .B2(n6792), .A(n4915), .ZN(n4916) );
  AOI21_X1 U6055 ( .B1(n6613), .B2(n5201), .A(n4916), .ZN(n4917) );
  OAI21_X1 U6056 ( .B1(n4941), .B2(n4918), .A(n4917), .ZN(U3043) );
  INV_X1 U6057 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4922) );
  AOI22_X1 U6058 ( .A1(n6460), .A2(n4943), .B1(n6611), .B2(n4942), .ZN(n4919)
         );
  OAI21_X1 U6059 ( .B1(n6546), .B2(n4945), .A(n4919), .ZN(n4920) );
  AOI21_X1 U6060 ( .B1(n6613), .B2(n6543), .A(n4920), .ZN(n4921) );
  OAI21_X1 U6061 ( .B1(n4949), .B2(n4922), .A(n4921), .ZN(U3123) );
  INV_X1 U6062 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4926) );
  AOI22_X1 U6063 ( .A1(n6460), .A2(n4928), .B1(n6611), .B2(n4927), .ZN(n4923)
         );
  OAI21_X1 U6064 ( .B1(n5170), .B2(n6796), .A(n4923), .ZN(n4924) );
  AOI21_X1 U6065 ( .B1(n6609), .B2(n4931), .A(n4924), .ZN(n4925) );
  OAI21_X1 U6066 ( .B1(n4934), .B2(n4926), .A(n4925), .ZN(U3059) );
  INV_X1 U6067 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4933) );
  AOI22_X1 U6068 ( .A1(n6447), .A2(n4928), .B1(n6591), .B2(n4927), .ZN(n4929)
         );
  OAI21_X1 U6069 ( .B1(n6534), .B2(n6796), .A(n4929), .ZN(n4930) );
  AOI21_X1 U6070 ( .B1(n6590), .B2(n4931), .A(n4930), .ZN(n4932) );
  OAI21_X1 U6071 ( .B1(n4934), .B2(n4933), .A(n4932), .ZN(U3056) );
  INV_X1 U6072 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4940) );
  AOI22_X1 U6073 ( .A1(n6503), .A2(n4936), .B1(n6597), .B2(n4935), .ZN(n4937)
         );
  OAI21_X1 U6074 ( .B1(n6453), .B2(n6792), .A(n4937), .ZN(n4938) );
  AOI21_X1 U6075 ( .B1(n6596), .B2(n5201), .A(n4938), .ZN(n4939) );
  OAI21_X1 U6076 ( .B1(n4941), .B2(n4940), .A(n4939), .ZN(U3041) );
  INV_X1 U6077 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4948) );
  AOI22_X1 U6078 ( .A1(n6503), .A2(n4943), .B1(n6597), .B2(n4942), .ZN(n4944)
         );
  OAI21_X1 U6079 ( .B1(n6453), .B2(n4945), .A(n4944), .ZN(n4946) );
  AOI21_X1 U6080 ( .B1(n6596), .B2(n6543), .A(n4946), .ZN(n4947) );
  OAI21_X1 U6081 ( .B1(n4949), .B2(n4948), .A(n4947), .ZN(U3121) );
  NOR2_X1 U6082 ( .A1(n4950), .A2(n6370), .ZN(n4951) );
  INV_X1 U6083 ( .A(n4998), .ZN(n4985) );
  AOI21_X1 U6084 ( .B1(n6558), .B2(n6468), .A(n4985), .ZN(n4954) );
  OAI21_X1 U6085 ( .B1(n4951), .B2(n5032), .A(n4954), .ZN(n4952) );
  OAI211_X1 U6086 ( .C1(n4955), .C2(n6520), .A(n6568), .B(n4952), .ZN(n4997)
         );
  NAND2_X1 U6087 ( .A1(n4997), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4959)
         );
  NOR2_X2 U6088 ( .A1(n4953), .A2(n4578), .ZN(n5256) );
  INV_X1 U6089 ( .A(n4954), .ZN(n4956) );
  AOI22_X1 U6090 ( .A1(n4956), .A2(n6520), .B1(n4955), .B2(
        STATE2_REG_2__SCAN_IN), .ZN(n4999) );
  OAI22_X1 U6091 ( .A1(n6583), .A2(n4999), .B1(n4998), .B2(n5089), .ZN(n4957)
         );
  AOI21_X1 U6092 ( .B1(n6580), .B2(n5256), .A(n4957), .ZN(n4958) );
  OAI211_X1 U6093 ( .C1(n5003), .C2(n6526), .A(n4959), .B(n4958), .ZN(U3142)
         );
  NAND2_X1 U6094 ( .A1(n4997), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4962)
         );
  INV_X1 U6095 ( .A(n6585), .ZN(n5110) );
  OAI22_X1 U6096 ( .A1(n6589), .A2(n4999), .B1(n4998), .B2(n5110), .ZN(n4960)
         );
  AOI21_X1 U6097 ( .B1(n6586), .B2(n5256), .A(n4960), .ZN(n4961) );
  OAI211_X1 U6098 ( .C1(n5003), .C2(n5163), .A(n4962), .B(n4961), .ZN(U3143)
         );
  NAND2_X1 U6099 ( .A1(n4997), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4965)
         );
  OAI22_X1 U6100 ( .A1(n6572), .A2(n4999), .B1(n4998), .B2(n5096), .ZN(n4963)
         );
  AOI21_X1 U6101 ( .B1(n6569), .B2(n5256), .A(n4963), .ZN(n4964) );
  OAI211_X1 U6102 ( .C1(n5003), .C2(n5194), .A(n4965), .B(n4964), .ZN(U3140)
         );
  NAND2_X1 U6103 ( .A1(n4972), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4968)
         );
  INV_X1 U6104 ( .A(n6591), .ZN(n5116) );
  OAI22_X1 U6105 ( .A1(n6595), .A2(n4974), .B1(n5116), .B2(n4973), .ZN(n4966)
         );
  AOI21_X1 U6106 ( .B1(n6592), .B2(n6608), .A(n4966), .ZN(n4967) );
  OAI211_X1 U6107 ( .C1(n5003), .C2(n6450), .A(n4968), .B(n4967), .ZN(U3136)
         );
  NAND2_X1 U6108 ( .A1(n4972), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4971)
         );
  INV_X1 U6109 ( .A(n6611), .ZN(n5100) );
  OAI22_X1 U6110 ( .A1(n6617), .A2(n4974), .B1(n5100), .B2(n4973), .ZN(n4969)
         );
  AOI21_X1 U6111 ( .B1(n6613), .B2(n6608), .A(n4969), .ZN(n4970) );
  OAI211_X1 U6112 ( .C1(n5003), .C2(n6546), .A(n4971), .B(n4970), .ZN(U3139)
         );
  NAND2_X1 U6113 ( .A1(n4972), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4977)
         );
  INV_X1 U6114 ( .A(n6597), .ZN(n5085) );
  OAI22_X1 U6115 ( .A1(n6601), .A2(n4974), .B1(n5085), .B2(n4973), .ZN(n4975)
         );
  AOI21_X1 U6116 ( .B1(n6596), .B2(n6608), .A(n4975), .ZN(n4976) );
  OAI211_X1 U6117 ( .C1(n5003), .C2(n6453), .A(n4977), .B(n4976), .ZN(U3137)
         );
  NOR2_X1 U6118 ( .A1(n4896), .A2(n4979), .ZN(n4980) );
  OR2_X1 U6119 ( .A1(n4978), .A2(n4980), .ZN(n6131) );
  AOI22_X1 U6120 ( .A1(n5414), .A2(DATAI_9_), .B1(n6241), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n4981) );
  OAI21_X1 U6121 ( .B1(n6131), .B2(n5684), .A(n4981), .ZN(U2882) );
  INV_X1 U6122 ( .A(n4997), .ZN(n4990) );
  INV_X1 U6123 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4984) );
  AOI22_X1 U6124 ( .A1(n6603), .A2(n4985), .B1(n6604), .B2(n5256), .ZN(n4983)
         );
  INV_X1 U6125 ( .A(n4999), .ZN(n4987) );
  AOI22_X1 U6126 ( .A1(n6454), .A2(n4987), .B1(n6602), .B2(n4986), .ZN(n4982)
         );
  OAI211_X1 U6127 ( .C1(n4990), .C2(n4984), .A(n4983), .B(n4982), .ZN(U3146)
         );
  AOI22_X1 U6128 ( .A1(n6574), .A2(n4985), .B1(n6575), .B2(n5256), .ZN(n4989)
         );
  AOI22_X1 U6129 ( .A1(n6437), .A2(n4987), .B1(n6573), .B2(n4986), .ZN(n4988)
         );
  OAI211_X1 U6130 ( .C1(n4990), .C2(n6959), .A(n4989), .B(n4988), .ZN(U3141)
         );
  NAND2_X1 U6131 ( .A1(n4997), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4993)
         );
  OAI22_X1 U6132 ( .A1(n6617), .A2(n4999), .B1(n4998), .B2(n5100), .ZN(n4991)
         );
  AOI21_X1 U6133 ( .B1(n6609), .B2(n5256), .A(n4991), .ZN(n4992) );
  OAI211_X1 U6134 ( .C1(n5003), .C2(n5170), .A(n4993), .B(n4992), .ZN(U3147)
         );
  NAND2_X1 U6135 ( .A1(n4997), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4996)
         );
  OAI22_X1 U6136 ( .A1(n6595), .A2(n4999), .B1(n4998), .B2(n5116), .ZN(n4994)
         );
  AOI21_X1 U6137 ( .B1(n6590), .B2(n5256), .A(n4994), .ZN(n4995) );
  OAI211_X1 U6138 ( .C1(n5003), .C2(n6534), .A(n4996), .B(n4995), .ZN(U3144)
         );
  NAND2_X1 U6139 ( .A1(n4997), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n5002)
         );
  OAI22_X1 U6140 ( .A1(n6601), .A2(n4999), .B1(n4998), .B2(n5085), .ZN(n5000)
         );
  AOI21_X1 U6141 ( .B1(n6598), .B2(n5256), .A(n5000), .ZN(n5001) );
  OAI211_X1 U6142 ( .C1(n5003), .C2(n5187), .A(n5002), .B(n5001), .ZN(U3145)
         );
  INV_X1 U6143 ( .A(n5032), .ZN(n5004) );
  OAI21_X1 U6144 ( .B1(n5005), .B2(n6564), .A(n5004), .ZN(n5011) );
  NAND2_X1 U6145 ( .A1(n6200), .A2(n5082), .ZN(n5221) );
  OR2_X1 U6146 ( .A1(n5221), .A2(n6510), .ZN(n5007) );
  NAND3_X1 U6147 ( .A1(n7081), .A2(n6631), .A3(n7064), .ZN(n5218) );
  NOR2_X1 U6148 ( .A1(n6556), .A2(n5218), .ZN(n5198) );
  INV_X1 U6149 ( .A(n5198), .ZN(n5006) );
  NAND2_X1 U6150 ( .A1(n5007), .A2(n5006), .ZN(n5010) );
  INV_X1 U6151 ( .A(n5218), .ZN(n5008) );
  AOI22_X1 U6152 ( .A1(n5011), .A2(n5010), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5008), .ZN(n5203) );
  INV_X1 U6153 ( .A(n5010), .ZN(n5012) );
  AOI22_X1 U6154 ( .A1(n5012), .A2(n5011), .B1(n5218), .B2(n6564), .ZN(n5013)
         );
  NAND2_X1 U6155 ( .A1(n6568), .A2(n5013), .ZN(n5197) );
  AOI22_X1 U6156 ( .A1(n6579), .A2(n5198), .B1(INSTQUEUE_REG_1__2__SCAN_IN), 
        .B2(n5197), .ZN(n5015) );
  NAND2_X1 U6157 ( .A1(n5201), .A2(n6580), .ZN(n5014) );
  OAI211_X1 U6158 ( .C1(n5248), .C2(n6526), .A(n5015), .B(n5014), .ZN(n5016)
         );
  INV_X1 U6159 ( .A(n5016), .ZN(n5017) );
  OAI21_X1 U6160 ( .B1(n5203), .B2(n6583), .A(n5017), .ZN(U3030) );
  AOI22_X1 U6161 ( .A1(n6585), .A2(n5198), .B1(INSTQUEUE_REG_1__3__SCAN_IN), 
        .B2(n5197), .ZN(n5019) );
  NAND2_X1 U6162 ( .A1(n5201), .A2(n6586), .ZN(n5018) );
  OAI211_X1 U6163 ( .C1(n5248), .C2(n5163), .A(n5019), .B(n5018), .ZN(n5020)
         );
  INV_X1 U6164 ( .A(n5020), .ZN(n5021) );
  OAI21_X1 U6165 ( .B1(n5203), .B2(n6589), .A(n5021), .ZN(U3031) );
  AOI22_X1 U6166 ( .A1(n6611), .A2(n5198), .B1(INSTQUEUE_REG_1__7__SCAN_IN), 
        .B2(n5197), .ZN(n5023) );
  NAND2_X1 U6167 ( .A1(n5201), .A2(n6609), .ZN(n5022) );
  OAI211_X1 U6168 ( .C1(n5248), .C2(n5170), .A(n5023), .B(n5022), .ZN(n5024)
         );
  INV_X1 U6169 ( .A(n5024), .ZN(n5025) );
  OAI21_X1 U6170 ( .B1(n5203), .B2(n6617), .A(n5025), .ZN(U3035) );
  AOI22_X1 U6171 ( .A1(n6591), .A2(n5198), .B1(INSTQUEUE_REG_1__4__SCAN_IN), 
        .B2(n5197), .ZN(n5027) );
  NAND2_X1 U6172 ( .A1(n5201), .A2(n6590), .ZN(n5026) );
  OAI211_X1 U6173 ( .C1(n5248), .C2(n6534), .A(n5027), .B(n5026), .ZN(n5028)
         );
  INV_X1 U6174 ( .A(n5028), .ZN(n5029) );
  OAI21_X1 U6175 ( .B1(n5203), .B2(n6595), .A(n5029), .ZN(U3032) );
  NOR3_X1 U6176 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n7081), .A3(n7064), 
        .ZN(n6519) );
  NAND2_X1 U6177 ( .A1(n6519), .A2(n6556), .ZN(n5041) );
  NAND2_X1 U6178 ( .A1(n5030), .A2(n4578), .ZN(n6421) );
  NOR2_X1 U6179 ( .A1(n6550), .A2(n6564), .ZN(n5033) );
  AOI21_X1 U6180 ( .B1(n5033), .B2(n5063), .A(n5032), .ZN(n5040) );
  NAND2_X1 U6181 ( .A1(n5034), .A2(n5074), .ZN(n6511) );
  INV_X1 U6182 ( .A(n6511), .ZN(n5037) );
  OAI211_X1 U6183 ( .C1(n5040), .C2(n5037), .A(n5036), .B(n5035), .ZN(n5038)
         );
  INV_X1 U6184 ( .A(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5045) );
  NAND3_X1 U6185 ( .A1(n6430), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6424), .ZN(n5039) );
  OAI21_X1 U6186 ( .B1(n5040), .B2(n6511), .A(n5039), .ZN(n6504) );
  INV_X1 U6187 ( .A(n5041), .ZN(n6501) );
  AOI22_X1 U6188 ( .A1(n6603), .A2(n6501), .B1(n6550), .B2(n6604), .ZN(n5042)
         );
  OAI21_X1 U6189 ( .B1(n5063), .B2(n6540), .A(n5042), .ZN(n5043) );
  AOI21_X1 U6190 ( .B1(n6504), .B2(n6454), .A(n5043), .ZN(n5044) );
  OAI21_X1 U6191 ( .B1(n6507), .B2(n5045), .A(n5044), .ZN(U3106) );
  AOI22_X1 U6192 ( .A1(n6585), .A2(n6501), .B1(n6550), .B2(n6586), .ZN(n5046)
         );
  OAI21_X1 U6193 ( .B1(n5063), .B2(n5163), .A(n5046), .ZN(n5047) );
  AOI21_X1 U6194 ( .B1(n6504), .B2(n6444), .A(n5047), .ZN(n5048) );
  OAI21_X1 U6195 ( .B1(n6507), .B2(n5049), .A(n5048), .ZN(U3103) );
  INV_X1 U6196 ( .A(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5053) );
  AOI22_X1 U6197 ( .A1(n6579), .A2(n6501), .B1(n6550), .B2(n6580), .ZN(n5050)
         );
  OAI21_X1 U6198 ( .B1(n5063), .B2(n6526), .A(n5050), .ZN(n5051) );
  AOI21_X1 U6199 ( .B1(n6504), .B2(n6440), .A(n5051), .ZN(n5052) );
  OAI21_X1 U6200 ( .B1(n6507), .B2(n5053), .A(n5052), .ZN(U3102) );
  INV_X1 U6201 ( .A(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5057) );
  AOI22_X1 U6202 ( .A1(n6574), .A2(n6501), .B1(n6550), .B2(n6575), .ZN(n5054)
         );
  OAI21_X1 U6203 ( .B1(n5063), .B2(n6793), .A(n5054), .ZN(n5055) );
  AOI21_X1 U6204 ( .B1(n6504), .B2(n6437), .A(n5055), .ZN(n5056) );
  OAI21_X1 U6205 ( .B1(n6507), .B2(n5057), .A(n5056), .ZN(U3101) );
  INV_X1 U6206 ( .A(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5061) );
  AOI22_X1 U6207 ( .A1(n6591), .A2(n6501), .B1(n6550), .B2(n6590), .ZN(n5058)
         );
  OAI21_X1 U6208 ( .B1(n5063), .B2(n6534), .A(n5058), .ZN(n5059) );
  AOI21_X1 U6209 ( .B1(n6504), .B2(n6447), .A(n5059), .ZN(n5060) );
  OAI21_X1 U6210 ( .B1(n6507), .B2(n5061), .A(n5060), .ZN(U3104) );
  INV_X1 U6211 ( .A(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5066) );
  AOI22_X1 U6212 ( .A1(n6611), .A2(n6501), .B1(n6550), .B2(n6609), .ZN(n5062)
         );
  OAI21_X1 U6213 ( .B1(n5063), .B2(n5170), .A(n5062), .ZN(n5064) );
  AOI21_X1 U6214 ( .B1(n6504), .B2(n6460), .A(n5064), .ZN(n5065) );
  OAI21_X1 U6215 ( .B1(n6507), .B2(n5066), .A(n5065), .ZN(U3107) );
  INV_X1 U6216 ( .A(EAX_REG_24__SCAN_IN), .ZN(n6285) );
  AOI22_X1 U6217 ( .A1(UWORD_REG_8__SCAN_IN), .A2(n5128), .B1(n6262), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n5067) );
  OAI21_X1 U6218 ( .B1(n6285), .B2(n5130), .A(n5067), .ZN(U2899) );
  INV_X1 U6219 ( .A(EAX_REG_19__SCAN_IN), .ZN(n6274) );
  AOI22_X1 U6220 ( .A1(UWORD_REG_3__SCAN_IN), .A2(n5128), .B1(n6262), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n5068) );
  OAI21_X1 U6221 ( .B1(n6274), .B2(n5130), .A(n5068), .ZN(U2904) );
  INV_X1 U6222 ( .A(EAX_REG_16__SCAN_IN), .ZN(n7031) );
  AOI22_X1 U6223 ( .A1(UWORD_REG_0__SCAN_IN), .A2(n5128), .B1(n6262), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n5069) );
  OAI21_X1 U6224 ( .B1(n7031), .B2(n5130), .A(n5069), .ZN(U2907) );
  INV_X1 U6225 ( .A(EAX_REG_28__SCAN_IN), .ZN(n6297) );
  AOI22_X1 U6226 ( .A1(UWORD_REG_12__SCAN_IN), .A2(n5128), .B1(n6262), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n5070) );
  OAI21_X1 U6227 ( .B1(n6297), .B2(n5130), .A(n5070), .ZN(U2895) );
  INV_X1 U6228 ( .A(n5071), .ZN(n5079) );
  INV_X1 U6229 ( .A(n6493), .ZN(n5104) );
  AOI21_X1 U6230 ( .B1(n5121), .B2(n5104), .A(n6064), .ZN(n5073) );
  AOI211_X1 U6231 ( .C1(n5082), .C2(n5074), .A(n6564), .B(n5073), .ZN(n5078)
         );
  NOR2_X1 U6232 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5075), .ZN(n5084)
         );
  OAI21_X1 U6233 ( .B1(n3515), .B2(n5084), .A(n5076), .ZN(n5077) );
  NAND2_X1 U6234 ( .A1(n5114), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5088) );
  INV_X1 U6235 ( .A(n5080), .ZN(n5081) );
  AOI22_X1 U6236 ( .A1(n5083), .A2(n5082), .B1(n6430), .B2(n5081), .ZN(n5117)
         );
  INV_X1 U6237 ( .A(n5084), .ZN(n5115) );
  OAI22_X1 U6238 ( .A1(n6601), .A2(n5117), .B1(n5085), .B2(n5115), .ZN(n5086)
         );
  AOI21_X1 U6239 ( .B1(n6596), .B2(n6493), .A(n5086), .ZN(n5087) );
  OAI211_X1 U6240 ( .C1(n6453), .C2(n5121), .A(n5088), .B(n5087), .ZN(U3089)
         );
  NAND2_X1 U6241 ( .A1(n5114), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5092) );
  OAI22_X1 U6242 ( .A1(n6583), .A2(n5117), .B1(n5089), .B2(n5115), .ZN(n5090)
         );
  AOI21_X1 U6243 ( .B1(n6578), .B2(n6493), .A(n5090), .ZN(n5091) );
  OAI211_X1 U6244 ( .C1(n5121), .C2(n6443), .A(n5092), .B(n5091), .ZN(U3086)
         );
  NAND2_X1 U6245 ( .A1(n5114), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5095) );
  INV_X1 U6246 ( .A(n5117), .ZN(n5107) );
  OAI22_X1 U6247 ( .A1(n6795), .A2(n5115), .B1(n6793), .B2(n5104), .ZN(n5093)
         );
  AOI21_X1 U6248 ( .B1(n6437), .B2(n5107), .A(n5093), .ZN(n5094) );
  OAI211_X1 U6249 ( .C1(n5121), .C2(n6797), .A(n5095), .B(n5094), .ZN(U3085)
         );
  NAND2_X1 U6250 ( .A1(n5114), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5099) );
  OAI22_X1 U6251 ( .A1(n6572), .A2(n5117), .B1(n5096), .B2(n5115), .ZN(n5097)
         );
  AOI21_X1 U6252 ( .B1(n6561), .B2(n6493), .A(n5097), .ZN(n5098) );
  OAI211_X1 U6253 ( .C1(n6436), .C2(n5121), .A(n5099), .B(n5098), .ZN(U3084)
         );
  NAND2_X1 U6254 ( .A1(n5114), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5103) );
  OAI22_X1 U6255 ( .A1(n6617), .A2(n5117), .B1(n5100), .B2(n5115), .ZN(n5101)
         );
  AOI21_X1 U6256 ( .B1(n6613), .B2(n6493), .A(n5101), .ZN(n5102) );
  OAI211_X1 U6257 ( .C1(n5121), .C2(n6546), .A(n5103), .B(n5102), .ZN(U3091)
         );
  NAND2_X1 U6258 ( .A1(n5114), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5109) );
  OAI22_X1 U6259 ( .A1(n5105), .A2(n5115), .B1(n6540), .B2(n5104), .ZN(n5106)
         );
  AOI21_X1 U6260 ( .B1(n6454), .B2(n5107), .A(n5106), .ZN(n5108) );
  OAI211_X1 U6261 ( .C1(n5121), .C2(n6457), .A(n5109), .B(n5108), .ZN(U3090)
         );
  NAND2_X1 U6262 ( .A1(n5114), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5113) );
  OAI22_X1 U6263 ( .A1(n6589), .A2(n5117), .B1(n5110), .B2(n5115), .ZN(n5111)
         );
  AOI21_X1 U6264 ( .B1(n6584), .B2(n6493), .A(n5111), .ZN(n5112) );
  OAI211_X1 U6265 ( .C1(n5121), .C2(n6530), .A(n5113), .B(n5112), .ZN(U3087)
         );
  NAND2_X1 U6266 ( .A1(n5114), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5120) );
  OAI22_X1 U6267 ( .A1(n6595), .A2(n5117), .B1(n5116), .B2(n5115), .ZN(n5118)
         );
  AOI21_X1 U6268 ( .B1(n6592), .B2(n6493), .A(n5118), .ZN(n5119) );
  OAI211_X1 U6269 ( .C1(n5121), .C2(n6450), .A(n5120), .B(n5119), .ZN(U3088)
         );
  INV_X1 U6270 ( .A(EAX_REG_26__SCAN_IN), .ZN(n6291) );
  AOI22_X1 U6271 ( .A1(n6779), .A2(UWORD_REG_10__SCAN_IN), .B1(n6262), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n5122) );
  OAI21_X1 U6272 ( .B1(n6291), .B2(n5130), .A(n5122), .ZN(U2897) );
  INV_X1 U6273 ( .A(EAX_REG_22__SCAN_IN), .ZN(n6279) );
  AOI22_X1 U6274 ( .A1(n6779), .A2(UWORD_REG_6__SCAN_IN), .B1(n6262), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n5123) );
  OAI21_X1 U6275 ( .B1(n6279), .B2(n5130), .A(n5123), .ZN(U2901) );
  INV_X1 U6276 ( .A(EAX_REG_23__SCAN_IN), .ZN(n6281) );
  AOI22_X1 U6277 ( .A1(n6779), .A2(UWORD_REG_7__SCAN_IN), .B1(n6262), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n5124) );
  OAI21_X1 U6278 ( .B1(n6281), .B2(n5130), .A(n5124), .ZN(U2900) );
  INV_X1 U6279 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6304) );
  AOI22_X1 U6280 ( .A1(n5128), .A2(UWORD_REG_14__SCAN_IN), .B1(n6262), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n5125) );
  OAI21_X1 U6281 ( .B1(n6304), .B2(n5130), .A(n5125), .ZN(U2893) );
  INV_X1 U6282 ( .A(EAX_REG_20__SCAN_IN), .ZN(n7100) );
  AOI22_X1 U6283 ( .A1(n5128), .A2(UWORD_REG_4__SCAN_IN), .B1(n6262), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n5126) );
  OAI21_X1 U6284 ( .B1(n7100), .B2(n5130), .A(n5126), .ZN(U2903) );
  AOI22_X1 U6285 ( .A1(n5128), .A2(UWORD_REG_5__SCAN_IN), .B1(n6262), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n5127) );
  OAI21_X1 U6286 ( .B1(n6950), .B2(n5130), .A(n5127), .ZN(U2902) );
  INV_X1 U6287 ( .A(EAX_REG_18__SCAN_IN), .ZN(n6272) );
  AOI22_X1 U6288 ( .A1(n5128), .A2(UWORD_REG_2__SCAN_IN), .B1(n6262), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n5129) );
  OAI21_X1 U6289 ( .B1(n6272), .B2(n5130), .A(n5129), .ZN(U2905) );
  INV_X1 U6290 ( .A(n5131), .ZN(n5132) );
  AOI21_X1 U6291 ( .B1(n6350), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n5132), 
        .ZN(n5133) );
  OAI21_X1 U6292 ( .B1(n6361), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n5133), 
        .ZN(n5134) );
  AOI21_X1 U6293 ( .B1(n5609), .B2(n6356), .A(n5134), .ZN(n5135) );
  OAI21_X1 U6294 ( .B1(n6068), .B2(n5136), .A(n5135), .ZN(U2985) );
  INV_X1 U6295 ( .A(n5137), .ZN(n6202) );
  AOI21_X1 U6296 ( .B1(n6350), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n5138), 
        .ZN(n5139) );
  OAI21_X1 U6297 ( .B1(n6361), .B2(n6194), .A(n5139), .ZN(n5140) );
  AOI21_X1 U6298 ( .B1(n6202), .B2(n6356), .A(n5140), .ZN(n5141) );
  OAI21_X1 U6299 ( .B1(n5142), .B2(n6068), .A(n5141), .ZN(U2983) );
  INV_X1 U6300 ( .A(n5143), .ZN(n5151) );
  NOR2_X1 U6301 ( .A1(n6512), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6791)
         );
  AOI21_X1 U6302 ( .B1(n5144), .B2(n3133), .A(n6791), .ZN(n5149) );
  NOR2_X1 U6303 ( .A1(n5149), .A2(n6564), .ZN(n5145) );
  AOI21_X1 U6304 ( .B1(n5151), .B2(STATE2_REG_2__SCAN_IN), .A(n5145), .ZN(
        n6799) );
  NAND3_X1 U6305 ( .A1(n5147), .A2(n6508), .A3(n5146), .ZN(n5148) );
  NAND2_X1 U6306 ( .A1(n5149), .A2(n5148), .ZN(n5150) );
  MUX2_X1 U6307 ( .A(n5151), .B(n5150), .S(n6520), .Z(n5152) );
  NAND2_X1 U6308 ( .A1(n6568), .A2(n5152), .ZN(n6802) );
  AOI22_X1 U6309 ( .A1(n6562), .A2(n6791), .B1(INSTQUEUE_REG_3__0__SCAN_IN), 
        .B2(n6802), .ZN(n5153) );
  OAI21_X1 U6310 ( .B1(n5194), .B2(n6792), .A(n5153), .ZN(n5154) );
  AOI21_X1 U6311 ( .B1(n6569), .B2(n5175), .A(n5154), .ZN(n5155) );
  OAI21_X1 U6312 ( .B1(n6799), .B2(n6572), .A(n5155), .ZN(U3044) );
  AOI22_X1 U6313 ( .A1(n6597), .A2(n6791), .B1(INSTQUEUE_REG_3__5__SCAN_IN), 
        .B2(n6802), .ZN(n5156) );
  OAI21_X1 U6314 ( .B1(n5187), .B2(n6792), .A(n5156), .ZN(n5157) );
  AOI21_X1 U6315 ( .B1(n6598), .B2(n5175), .A(n5157), .ZN(n5158) );
  OAI21_X1 U6316 ( .B1(n6799), .B2(n6601), .A(n5158), .ZN(U3049) );
  AOI22_X1 U6317 ( .A1(n6579), .A2(n6791), .B1(INSTQUEUE_REG_3__2__SCAN_IN), 
        .B2(n6802), .ZN(n5159) );
  OAI21_X1 U6318 ( .B1(n6526), .B2(n6792), .A(n5159), .ZN(n5160) );
  AOI21_X1 U6319 ( .B1(n6580), .B2(n5175), .A(n5160), .ZN(n5161) );
  OAI21_X1 U6320 ( .B1(n6799), .B2(n6583), .A(n5161), .ZN(U3046) );
  AOI22_X1 U6321 ( .A1(n6585), .A2(n6791), .B1(INSTQUEUE_REG_3__3__SCAN_IN), 
        .B2(n6802), .ZN(n5162) );
  OAI21_X1 U6322 ( .B1(n5163), .B2(n6792), .A(n5162), .ZN(n5164) );
  AOI21_X1 U6323 ( .B1(n6586), .B2(n5175), .A(n5164), .ZN(n5165) );
  OAI21_X1 U6324 ( .B1(n6799), .B2(n6589), .A(n5165), .ZN(U3047) );
  INV_X1 U6325 ( .A(n6454), .ZN(n6607) );
  AOI22_X1 U6326 ( .A1(n6603), .A2(n6791), .B1(INSTQUEUE_REG_3__6__SCAN_IN), 
        .B2(n6802), .ZN(n5166) );
  OAI21_X1 U6327 ( .B1(n6540), .B2(n6792), .A(n5166), .ZN(n5167) );
  AOI21_X1 U6328 ( .B1(n6604), .B2(n5175), .A(n5167), .ZN(n5168) );
  OAI21_X1 U6329 ( .B1(n6607), .B2(n6799), .A(n5168), .ZN(U3050) );
  AOI22_X1 U6330 ( .A1(n6611), .A2(n6791), .B1(INSTQUEUE_REG_3__7__SCAN_IN), 
        .B2(n6802), .ZN(n5169) );
  OAI21_X1 U6331 ( .B1(n5170), .B2(n6792), .A(n5169), .ZN(n5171) );
  AOI21_X1 U6332 ( .B1(n6609), .B2(n5175), .A(n5171), .ZN(n5172) );
  OAI21_X1 U6333 ( .B1(n6799), .B2(n6617), .A(n5172), .ZN(U3051) );
  AOI22_X1 U6334 ( .A1(n6591), .A2(n6791), .B1(INSTQUEUE_REG_3__4__SCAN_IN), 
        .B2(n6802), .ZN(n5173) );
  OAI21_X1 U6335 ( .B1(n6534), .B2(n6792), .A(n5173), .ZN(n5174) );
  AOI21_X1 U6336 ( .B1(n6590), .B2(n5175), .A(n5174), .ZN(n5176) );
  OAI21_X1 U6337 ( .B1(n6799), .B2(n6595), .A(n5176), .ZN(U3048) );
  AOI21_X1 U6338 ( .B1(n5178), .B2(n5177), .A(n5267), .ZN(n6381) );
  INV_X1 U6339 ( .A(n6381), .ZN(n5179) );
  INV_X1 U6340 ( .A(EBX_REG_9__SCAN_IN), .ZN(n6137) );
  OAI222_X1 U6341 ( .A1(n5179), .A2(n5671), .B1(n6231), .B2(n6137), .C1(n5670), 
        .C2(n6131), .ZN(U2850) );
  INV_X1 U6342 ( .A(n6167), .ZN(n5183) );
  AOI21_X1 U6343 ( .B1(n6350), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n5180), 
        .ZN(n5181) );
  OAI21_X1 U6344 ( .B1(n6361), .B2(n6176), .A(n5181), .ZN(n5182) );
  AOI21_X1 U6345 ( .B1(n5183), .B2(n6356), .A(n5182), .ZN(n5184) );
  OAI21_X1 U6346 ( .B1(n6068), .B2(n5185), .A(n5184), .ZN(U2981) );
  AOI22_X1 U6347 ( .A1(n6597), .A2(n5198), .B1(INSTQUEUE_REG_1__5__SCAN_IN), 
        .B2(n5197), .ZN(n5186) );
  OAI21_X1 U6348 ( .B1(n5187), .B2(n5248), .A(n5186), .ZN(n5188) );
  AOI21_X1 U6349 ( .B1(n6598), .B2(n5201), .A(n5188), .ZN(n5189) );
  OAI21_X1 U6350 ( .B1(n5203), .B2(n6601), .A(n5189), .ZN(U3033) );
  INV_X1 U6351 ( .A(n6437), .ZN(n6798) );
  AOI22_X1 U6352 ( .A1(n6574), .A2(n5198), .B1(INSTQUEUE_REG_1__1__SCAN_IN), 
        .B2(n5197), .ZN(n5190) );
  OAI21_X1 U6353 ( .B1(n6793), .B2(n5248), .A(n5190), .ZN(n5191) );
  AOI21_X1 U6354 ( .B1(n6575), .B2(n5201), .A(n5191), .ZN(n5192) );
  OAI21_X1 U6355 ( .B1(n6798), .B2(n5203), .A(n5192), .ZN(U3029) );
  AOI22_X1 U6356 ( .A1(n6562), .A2(n5198), .B1(INSTQUEUE_REG_1__0__SCAN_IN), 
        .B2(n5197), .ZN(n5193) );
  OAI21_X1 U6357 ( .B1(n5194), .B2(n5248), .A(n5193), .ZN(n5195) );
  AOI21_X1 U6358 ( .B1(n6569), .B2(n5201), .A(n5195), .ZN(n5196) );
  OAI21_X1 U6359 ( .B1(n5203), .B2(n6572), .A(n5196), .ZN(U3028) );
  AOI22_X1 U6360 ( .A1(n6603), .A2(n5198), .B1(INSTQUEUE_REG_1__6__SCAN_IN), 
        .B2(n5197), .ZN(n5199) );
  OAI21_X1 U6361 ( .B1(n6540), .B2(n5248), .A(n5199), .ZN(n5200) );
  AOI21_X1 U6362 ( .B1(n6604), .B2(n5201), .A(n5200), .ZN(n5202) );
  OAI21_X1 U6363 ( .B1(n6607), .B2(n5203), .A(n5202), .ZN(U3034) );
  AOI22_X1 U6364 ( .A1(n5341), .A2(n5204), .B1(n5342), .B2(n5335), .ZN(n6396)
         );
  XOR2_X1 U6365 ( .A(n5205), .B(n5206), .Z(n5305) );
  NAND2_X1 U6366 ( .A1(n5305), .A2(n6415), .ZN(n5213) );
  AOI21_X1 U6367 ( .B1(n6395), .B2(n4323), .A(n5290), .ZN(n5211) );
  INV_X1 U6368 ( .A(n5207), .ZN(n5208) );
  NAND2_X1 U6369 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n5208), .ZN(n6391)
         );
  INV_X1 U6370 ( .A(n6391), .ZN(n5289) );
  AND2_X1 U6371 ( .A1(n6368), .A2(REIP_REG_8__SCAN_IN), .ZN(n5307) );
  NOR2_X1 U6372 ( .A1(n6413), .A2(n5209), .ZN(n5210) );
  AOI211_X1 U6373 ( .C1(n5211), .C2(n5289), .A(n5307), .B(n5210), .ZN(n5212)
         );
  OAI211_X1 U6374 ( .C1(n6396), .C2(n4323), .A(n5213), .B(n5212), .ZN(U3010)
         );
  NOR2_X1 U6375 ( .A1(n4978), .A2(n5215), .ZN(n5216) );
  OR2_X1 U6376 ( .A1(n5214), .A2(n5216), .ZN(n6119) );
  AOI22_X1 U6377 ( .A1(n5414), .A2(DATAI_10_), .B1(n6241), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n5217) );
  OAI21_X1 U6378 ( .B1(n6119), .B2(n5684), .A(n5217), .ZN(U2881) );
  NOR2_X1 U6379 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5218), .ZN(n5255)
         );
  INV_X1 U6380 ( .A(n5255), .ZN(n5220) );
  AOI211_X1 U6381 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5220), .A(n6425), .B(
        n5219), .ZN(n5224) );
  INV_X1 U6382 ( .A(n5248), .ZN(n5254) );
  OAI21_X1 U6383 ( .B1(n5254), .B2(n5256), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5222) );
  NAND3_X1 U6384 ( .A1(n5222), .A2(n6520), .A3(n5221), .ZN(n5223) );
  OAI22_X1 U6385 ( .A1(n6428), .A2(n5227), .B1(n5226), .B2(n5225), .ZN(n5257)
         );
  AOI22_X1 U6386 ( .A1(n6503), .A2(n5257), .B1(n6597), .B2(n5255), .ZN(n5228)
         );
  OAI21_X1 U6387 ( .B1(n6453), .B2(n5248), .A(n5228), .ZN(n5229) );
  AOI21_X1 U6388 ( .B1(n6596), .B2(n5256), .A(n5229), .ZN(n5230) );
  OAI21_X1 U6389 ( .B1(n5261), .B2(n5231), .A(n5230), .ZN(U3025) );
  AOI22_X1 U6390 ( .A1(n6460), .A2(n5257), .B1(n6611), .B2(n5255), .ZN(n5232)
         );
  OAI21_X1 U6391 ( .B1(n6546), .B2(n5248), .A(n5232), .ZN(n5233) );
  AOI21_X1 U6392 ( .B1(n6613), .B2(n5256), .A(n5233), .ZN(n5234) );
  OAI21_X1 U6393 ( .B1(n5261), .B2(n5235), .A(n5234), .ZN(U3027) );
  AOI22_X1 U6394 ( .A1(n6498), .A2(n5257), .B1(n6562), .B2(n5255), .ZN(n5236)
         );
  OAI21_X1 U6395 ( .B1(n6436), .B2(n5248), .A(n5236), .ZN(n5237) );
  AOI21_X1 U6396 ( .B1(n6561), .B2(n5256), .A(n5237), .ZN(n5238) );
  OAI21_X1 U6397 ( .B1(n5261), .B2(n6902), .A(n5238), .ZN(U3020) );
  AOI22_X1 U6398 ( .A1(n6440), .A2(n5257), .B1(n6579), .B2(n5255), .ZN(n5239)
         );
  OAI21_X1 U6399 ( .B1(n6443), .B2(n5248), .A(n5239), .ZN(n5240) );
  AOI21_X1 U6400 ( .B1(n6578), .B2(n5256), .A(n5240), .ZN(n5241) );
  OAI21_X1 U6401 ( .B1(n5261), .B2(n5242), .A(n5241), .ZN(U3022) );
  AOI22_X1 U6402 ( .A1(n6447), .A2(n5257), .B1(n6591), .B2(n5255), .ZN(n5243)
         );
  OAI21_X1 U6403 ( .B1(n6450), .B2(n5248), .A(n5243), .ZN(n5244) );
  AOI21_X1 U6404 ( .B1(n6592), .B2(n5256), .A(n5244), .ZN(n5245) );
  OAI21_X1 U6405 ( .B1(n5261), .B2(n5246), .A(n5245), .ZN(U3024) );
  AOI22_X1 U6406 ( .A1(n6444), .A2(n5257), .B1(n6585), .B2(n5255), .ZN(n5247)
         );
  OAI21_X1 U6407 ( .B1(n6530), .B2(n5248), .A(n5247), .ZN(n5249) );
  AOI21_X1 U6408 ( .B1(n6584), .B2(n5256), .A(n5249), .ZN(n5250) );
  OAI21_X1 U6409 ( .B1(n5261), .B2(n3679), .A(n5250), .ZN(U3023) );
  AOI22_X1 U6410 ( .A1(n6603), .A2(n5255), .B1(n6604), .B2(n5254), .ZN(n5252)
         );
  AOI22_X1 U6411 ( .A1(n6454), .A2(n5257), .B1(n6602), .B2(n5256), .ZN(n5251)
         );
  OAI211_X1 U6412 ( .C1(n5261), .C2(n5253), .A(n5252), .B(n5251), .ZN(U3026)
         );
  AOI22_X1 U6413 ( .A1(n6574), .A2(n5255), .B1(n6575), .B2(n5254), .ZN(n5259)
         );
  AOI22_X1 U6414 ( .A1(n6437), .A2(n5257), .B1(n6573), .B2(n5256), .ZN(n5258)
         );
  OAI211_X1 U6415 ( .C1(n5261), .C2(n5260), .A(n5259), .B(n5258), .ZN(U3021)
         );
  XOR2_X1 U6416 ( .A(n5262), .B(n5263), .Z(n6393) );
  INV_X1 U6417 ( .A(n6068), .ZN(n6367) );
  NAND2_X1 U6418 ( .A1(n6393), .A2(n6367), .ZN(n5266) );
  INV_X1 U6419 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6905) );
  NOR2_X1 U6420 ( .A1(n6401), .A2(n6905), .ZN(n6387) );
  NOR2_X1 U6421 ( .A1(n6361), .A2(n6140), .ZN(n5264) );
  AOI211_X1 U6422 ( .C1(n6350), .C2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n6387), 
        .B(n5264), .ZN(n5265) );
  OAI211_X1 U6423 ( .C1(n5989), .C2(n6141), .A(n5266), .B(n5265), .ZN(U2979)
         );
  OR2_X1 U6424 ( .A1(n5268), .A2(n5267), .ZN(n5269) );
  NAND2_X1 U6425 ( .A1(n5269), .A2(n5274), .ZN(n6114) );
  OAI222_X1 U6426 ( .A1(n6114), .A2(n5671), .B1(n5270), .B2(n6231), .C1(n6119), 
        .C2(n5670), .ZN(U2849) );
  OAI21_X1 U6427 ( .B1(n5214), .B2(n5272), .A(n5271), .ZN(n5591) );
  AOI22_X1 U6428 ( .A1(n5414), .A2(DATAI_11_), .B1(n6241), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n5273) );
  OAI21_X1 U6429 ( .B1(n5591), .B2(n5684), .A(n5273), .ZN(U2880) );
  AOI21_X1 U6430 ( .B1(n5275), .B2(n5274), .A(n5347), .ZN(n6373) );
  AOI22_X1 U6431 ( .A1(n6227), .A2(n6373), .B1(n5412), .B2(EBX_REG_11__SCAN_IN), .ZN(n5276) );
  OAI21_X1 U6432 ( .B1(n5591), .B2(n5670), .A(n5276), .ZN(U2848) );
  OAI21_X1 U6433 ( .B1(n6365), .B2(n5278), .A(n5277), .ZN(n5280) );
  NOR2_X1 U6434 ( .A1(n6157), .A2(n6370), .ZN(n5279) );
  AOI211_X1 U6435 ( .C1(n5776), .C2(n6154), .A(n5280), .B(n5279), .ZN(n5281)
         );
  OAI21_X1 U6436 ( .B1(n6068), .B2(n5282), .A(n5281), .ZN(U2980) );
  INV_X1 U6437 ( .A(n5283), .ZN(n5285) );
  NAND2_X1 U6438 ( .A1(n5285), .A2(n5284), .ZN(n5286) );
  XNOR2_X1 U6439 ( .A(n5287), .B(n5286), .ZN(n5315) );
  OAI21_X1 U6440 ( .B1(n5288), .B2(n5290), .A(n6396), .ZN(n6382) );
  INV_X1 U6441 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6713) );
  OAI22_X1 U6442 ( .A1(n6413), .A2(n6114), .B1(n6713), .B2(n6401), .ZN(n5293)
         );
  NAND2_X1 U6443 ( .A1(n5290), .A2(n5289), .ZN(n6386) );
  AOI221_X1 U6444 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .C1(n5300), .C2(n5291), .A(n6386), 
        .ZN(n5292) );
  AOI211_X1 U6445 ( .C1(INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n6382), .A(n5293), .B(n5292), .ZN(n5294) );
  OAI21_X1 U6446 ( .B1(n6014), .B2(n5315), .A(n5294), .ZN(U3008) );
  NAND2_X1 U6447 ( .A1(n6189), .A2(n6356), .ZN(n5297) );
  OAI22_X1 U6448 ( .A1(n6365), .A2(n6180), .B1(n6401), .B2(n6706), .ZN(n5295)
         );
  AOI21_X1 U6449 ( .B1(n6177), .B2(n5776), .A(n5295), .ZN(n5296) );
  OAI211_X1 U6450 ( .C1(n5298), .C2(n6068), .A(n5297), .B(n5296), .ZN(U2982)
         );
  XNOR2_X1 U6451 ( .A(n4327), .B(n5300), .ZN(n5301) );
  XNOR2_X1 U6452 ( .A(n5299), .B(n5301), .ZN(n6383) );
  NAND2_X1 U6453 ( .A1(n6383), .A2(n6367), .ZN(n5304) );
  NAND2_X1 U6454 ( .A1(n6368), .A2(REIP_REG_9__SCAN_IN), .ZN(n6379) );
  OAI21_X1 U6455 ( .B1(n6365), .B2(n6128), .A(n6379), .ZN(n5302) );
  AOI21_X1 U6456 ( .B1(n6134), .B2(n5776), .A(n5302), .ZN(n5303) );
  OAI211_X1 U6457 ( .C1(n5989), .C2(n6131), .A(n5304), .B(n5303), .ZN(U2977)
         );
  NAND2_X1 U6458 ( .A1(n5305), .A2(n6367), .ZN(n5309) );
  AND2_X1 U6459 ( .A1(n6350), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5306)
         );
  AOI211_X1 U6460 ( .C1(n5776), .C2(n5592), .A(n5307), .B(n5306), .ZN(n5308)
         );
  OAI211_X1 U6461 ( .C1(n6370), .C2(n5604), .A(n5309), .B(n5308), .ZN(U2978)
         );
  INV_X1 U6462 ( .A(n6119), .ZN(n5313) );
  INV_X1 U6463 ( .A(n5310), .ZN(n6118) );
  AOI22_X1 U6464 ( .A1(n6350), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6368), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5311) );
  OAI21_X1 U6465 ( .B1(n6361), .B2(n6118), .A(n5311), .ZN(n5312) );
  AOI21_X1 U6466 ( .B1(n5313), .B2(n6356), .A(n5312), .ZN(n5314) );
  OAI21_X1 U6467 ( .B1(n5315), .B2(n6068), .A(n5314), .ZN(U2976) );
  AOI21_X1 U6468 ( .B1(n5316), .B2(n5271), .A(n3129), .ZN(n6229) );
  INV_X1 U6469 ( .A(n6229), .ZN(n5318) );
  INV_X1 U6470 ( .A(DATAI_12_), .ZN(n6295) );
  OAI222_X1 U6471 ( .A1(n5318), .A2(n5684), .B1(n5467), .B2(n5317), .C1(n6295), 
        .C2(n5381), .ZN(U2879) );
  NAND2_X1 U6472 ( .A1(n5320), .A2(n5319), .ZN(n5321) );
  XNOR2_X1 U6473 ( .A(n5322), .B(n5321), .ZN(n6375) );
  NAND2_X1 U6474 ( .A1(n6375), .A2(n6367), .ZN(n5326) );
  INV_X1 U6475 ( .A(REIP_REG_11__SCAN_IN), .ZN(n5323) );
  NOR2_X1 U6476 ( .A1(n6401), .A2(n5323), .ZN(n6372) );
  NOR2_X1 U6477 ( .A1(n6361), .A2(n5582), .ZN(n5324) );
  AOI211_X1 U6478 ( .C1(n6350), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6372), 
        .B(n5324), .ZN(n5325) );
  OAI211_X1 U6479 ( .C1(n5989), .C2(n5591), .A(n5326), .B(n5325), .ZN(U2975)
         );
  NOR2_X1 U6480 ( .A1(n5329), .A2(n3225), .ZN(n5330) );
  XNOR2_X1 U6481 ( .A(n5327), .B(n5330), .ZN(n5351) );
  INV_X1 U6482 ( .A(n6109), .ZN(n5332) );
  AND2_X1 U6483 ( .A1(n6351), .A2(REIP_REG_12__SCAN_IN), .ZN(n5348) );
  AOI21_X1 U6484 ( .B1(n6350), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n5348), 
        .ZN(n5331) );
  OAI21_X1 U6485 ( .B1(n6361), .B2(n5332), .A(n5331), .ZN(n5333) );
  AOI21_X1 U6486 ( .B1(n6229), .B2(n6356), .A(n5333), .ZN(n5334) );
  OAI21_X1 U6487 ( .B1(n5351), .B2(n6068), .A(n5334), .ZN(U2974) );
  NOR2_X1 U6488 ( .A1(n5339), .A2(n5341), .ZN(n5337) );
  INV_X1 U6489 ( .A(n5335), .ZN(n5336) );
  NOR2_X1 U6490 ( .A1(n5342), .A2(n5339), .ZN(n5343) );
  OAI22_X1 U6491 ( .A1(n5337), .A2(n5867), .B1(n5336), .B2(n5343), .ZN(n6374)
         );
  NAND2_X1 U6492 ( .A1(n5338), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5340)
         );
  AOI221_X1 U6493 ( .B1(n5342), .B2(n5341), .C1(n5340), .C2(n5341), .A(n5339), 
        .ZN(n6039) );
  AOI21_X1 U6494 ( .B1(n5344), .B2(n5343), .A(n6039), .ZN(n6378) );
  INV_X1 U6495 ( .A(n6378), .ZN(n5890) );
  XOR2_X1 U6496 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .B(
        INSTADDRPOINTER_REG_11__SCAN_IN), .Z(n5345) );
  AOI22_X1 U6497 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n6374), .B1(n5890), .B2(n5345), .ZN(n5350) );
  XOR2_X1 U6498 ( .A(n5347), .B(n5346), .Z(n6226) );
  AOI21_X1 U6499 ( .B1(n6389), .B2(n6226), .A(n5348), .ZN(n5349) );
  OAI211_X1 U6500 ( .C1(n5351), .C2(n6014), .A(n5350), .B(n5349), .ZN(U3006)
         );
  OAI21_X1 U6501 ( .B1(n3123), .B2(n5355), .A(n5354), .ZN(n5787) );
  AOI22_X1 U6502 ( .A1(n5414), .A2(DATAI_14_), .B1(n6241), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5356) );
  OAI21_X1 U6503 ( .B1(n5787), .B2(n5684), .A(n5356), .ZN(U2877) );
  XOR2_X1 U6504 ( .A(n5358), .B(n5357), .Z(n6099) );
  INV_X1 U6505 ( .A(n6099), .ZN(n5380) );
  AOI21_X1 U6506 ( .B1(n5360), .B2(n5359), .A(n5377), .ZN(n6093) );
  AOI22_X1 U6507 ( .A1(n6227), .A2(n6093), .B1(n5412), .B2(EBX_REG_13__SCAN_IN), .ZN(n5361) );
  OAI21_X1 U6508 ( .B1(n5380), .B2(n5670), .A(n5361), .ZN(U2846) );
  OAI21_X1 U6509 ( .B1(n5364), .B2(n5363), .A(n5362), .ZN(n5365) );
  INV_X1 U6510 ( .A(n5365), .ZN(n5376) );
  INV_X1 U6511 ( .A(REIP_REG_13__SCAN_IN), .ZN(n5366) );
  NOR2_X1 U6512 ( .A1(n6401), .A2(n5366), .ZN(n5373) );
  AOI21_X1 U6513 ( .B1(n6350), .B2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5373), 
        .ZN(n5367) );
  OAI21_X1 U6514 ( .B1(n6361), .B2(n6097), .A(n5367), .ZN(n5368) );
  AOI21_X1 U6515 ( .B1(n6099), .B2(n6356), .A(n5368), .ZN(n5369) );
  OAI21_X1 U6516 ( .B1(n5376), .B2(n6068), .A(n5369), .ZN(U2973) );
  AOI21_X1 U6517 ( .B1(n5372), .B2(n5370), .A(n6374), .ZN(n5371) );
  OAI21_X1 U6518 ( .B1(n5889), .B2(n6419), .A(n5371), .ZN(n6038) );
  NOR2_X1 U6519 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5372), .ZN(n6040)
         );
  AOI22_X1 U6520 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n6038), .B1(n6040), .B2(n5890), .ZN(n5375) );
  AOI21_X1 U6521 ( .B1(n6389), .B2(n6093), .A(n5373), .ZN(n5374) );
  OAI211_X1 U6522 ( .C1(n5376), .C2(n6014), .A(n5375), .B(n5374), .ZN(U3005)
         );
  XNOR2_X1 U6523 ( .A(n5378), .B(n5377), .ZN(n5571) );
  INV_X1 U6524 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5379) );
  OAI222_X1 U6525 ( .A1(n5787), .A2(n5670), .B1(n5671), .B2(n5571), .C1(n6231), 
        .C2(n5379), .ZN(U2845) );
  INV_X1 U6526 ( .A(DATAI_13_), .ZN(n6298) );
  INV_X1 U6527 ( .A(EAX_REG_13__SCAN_IN), .ZN(n7003) );
  OAI222_X1 U6528 ( .A1(n5381), .A2(n6298), .B1(n5684), .B2(n5380), .C1(n7003), 
        .C2(n5467), .ZN(U2878) );
  INV_X1 U6529 ( .A(n5354), .ZN(n5384) );
  OAI21_X1 U6530 ( .B1(n5384), .B2(n3900), .A(n5557), .ZN(n5780) );
  NAND2_X1 U6531 ( .A1(n5385), .A2(n4443), .ZN(n6675) );
  INV_X1 U6532 ( .A(n6677), .ZN(n6783) );
  NAND3_X1 U6533 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), 
        .A3(n6783), .ZN(n6669) );
  NAND2_X1 U6534 ( .A1(n6675), .A2(n6669), .ZN(n5386) );
  NOR2_X1 U6535 ( .A1(n5390), .A2(n5389), .ZN(n5391) );
  NOR2_X1 U6536 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5399) );
  OR2_X1 U6537 ( .A1(n5400), .A2(n5399), .ZN(n5406) );
  NAND2_X1 U6538 ( .A1(n3492), .A2(EBX_REG_31__SCAN_IN), .ZN(n5392) );
  NOR2_X1 U6539 ( .A1(n5406), .A2(n5392), .ZN(n5393) );
  AOI21_X1 U6540 ( .B1(n5396), .B2(n5395), .A(n5394), .ZN(n6031) );
  NAND2_X1 U6541 ( .A1(n6214), .A2(n6031), .ZN(n5398) );
  NAND2_X1 U6542 ( .A1(n6193), .A2(n5397), .ZN(n6163) );
  OAI211_X1 U6543 ( .C1(n6212), .C2(n5774), .A(n5398), .B(n6163), .ZN(n5410)
         );
  INV_X1 U6544 ( .A(n5399), .ZN(n5405) );
  NOR2_X1 U6545 ( .A1(n5400), .A2(n5405), .ZN(n5402) );
  AND2_X1 U6546 ( .A1(n5402), .A2(n5401), .ZN(n5403) );
  NAND2_X2 U6547 ( .A1(n5607), .A2(n5403), .ZN(n6206) );
  INV_X1 U6548 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6719) );
  INV_X1 U6549 ( .A(REIP_REG_12__SCAN_IN), .ZN(n5404) );
  INV_X1 U6550 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6711) );
  INV_X1 U6551 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6999) );
  NAND3_X1 U6552 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .A3(
        REIP_REG_3__SCAN_IN), .ZN(n6183) );
  NOR2_X1 U6553 ( .A1(n6706), .A2(n6183), .ZN(n6170) );
  NAND2_X1 U6554 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6170), .ZN(n6139) );
  NOR2_X1 U6555 ( .A1(n6999), .A2(n6139), .ZN(n6143) );
  NAND2_X1 U6556 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6143), .ZN(n5593) );
  NOR2_X1 U6557 ( .A1(n6711), .A2(n5593), .ZN(n5597) );
  NAND2_X1 U6558 ( .A1(REIP_REG_9__SCAN_IN), .A2(n5597), .ZN(n6116) );
  NOR2_X1 U6559 ( .A1(n6713), .A2(n6116), .ZN(n5588) );
  NAND2_X1 U6560 ( .A1(REIP_REG_11__SCAN_IN), .A2(n5588), .ZN(n6100) );
  NOR2_X1 U6561 ( .A1(n5404), .A2(n6100), .ZN(n6101) );
  NAND2_X1 U6562 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6101), .ZN(n5577) );
  NOR2_X1 U6563 ( .A1(n6719), .A2(n5577), .ZN(n5430) );
  NAND2_X1 U6564 ( .A1(n6171), .A2(n5430), .ZN(n5566) );
  NOR2_X1 U6565 ( .A1(n6689), .A2(n5405), .ZN(n5470) );
  OAI22_X1 U6566 ( .A1(n5470), .A2(n6782), .B1(n5406), .B2(EBX_REG_31__SCAN_IN), .ZN(n5407) );
  OAI21_X1 U6567 ( .B1(n6206), .B2(n5430), .A(n6193), .ZN(n5574) );
  AOI22_X1 U6568 ( .A1(EBX_REG_15__SCAN_IN), .A2(n6209), .B1(
        REIP_REG_15__SCAN_IN), .B2(n5574), .ZN(n5408) );
  OAI21_X1 U6569 ( .B1(REIP_REG_15__SCAN_IN), .B2(n5566), .A(n5408), .ZN(n5409) );
  AOI211_X1 U6570 ( .C1(n5777), .C2(n6133), .A(n5410), .B(n5409), .ZN(n5411)
         );
  OAI21_X1 U6571 ( .B1(n5780), .B2(n6156), .A(n5411), .ZN(U2812) );
  AOI22_X1 U6572 ( .A1(n6227), .A2(n6031), .B1(n5412), .B2(EBX_REG_15__SCAN_IN), .ZN(n5413) );
  OAI21_X1 U6573 ( .B1(n5780), .B2(n5670), .A(n5413), .ZN(U2844) );
  AOI22_X1 U6574 ( .A1(n5414), .A2(DATAI_15_), .B1(n6241), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5415) );
  OAI21_X1 U6575 ( .B1(n5780), .B2(n5684), .A(n5415), .ZN(U2876) );
  INV_X1 U6576 ( .A(n5417), .ZN(n5418) );
  NAND2_X1 U6577 ( .A1(n5709), .A2(n5418), .ZN(n5419) );
  NOR2_X1 U6578 ( .A1(n5416), .A2(n5419), .ZN(n5685) );
  INV_X1 U6579 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n7006) );
  AOI21_X1 U6580 ( .B1(n5685), .B2(n7006), .A(n5420), .ZN(n5421) );
  XOR2_X1 U6581 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .B(n5421), .Z(n5803) );
  NOR2_X1 U6582 ( .A1(n5429), .A2(n6370), .ZN(n5427) );
  INV_X1 U6583 ( .A(n5449), .ZN(n5424) );
  NOR2_X1 U6584 ( .A1(n5424), .A2(n6361), .ZN(n5426) );
  NAND2_X1 U6585 ( .A1(n6368), .A2(REIP_REG_30__SCAN_IN), .ZN(n5797) );
  OAI21_X1 U6586 ( .B1(n6365), .B2(n6923), .A(n5797), .ZN(n5425) );
  OAI21_X1 U6587 ( .B1(n5803), .B2(n6068), .A(n5428), .ZN(U2956) );
  INV_X1 U6588 ( .A(REIP_REG_18__SCAN_IN), .ZN(n5878) );
  NAND2_X1 U6589 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n5563) );
  NAND2_X1 U6590 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6085), .ZN(n5947) );
  NAND3_X1 U6591 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        n5950), .ZN(n5924) );
  NAND3_X1 U6592 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n5432) );
  NAND2_X1 U6593 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n5905) );
  INV_X1 U6594 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6734) );
  NOR2_X1 U6595 ( .A1(n5905), .A2(n6734), .ZN(n5434) );
  NAND2_X1 U6596 ( .A1(n5906), .A2(n5434), .ZN(n5507) );
  INV_X1 U6597 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6737) );
  INV_X1 U6598 ( .A(REIP_REG_28__SCAN_IN), .ZN(n5437) );
  AND2_X1 U6599 ( .A1(REIP_REG_30__SCAN_IN), .A2(REIP_REG_29__SCAN_IN), .ZN(
        n5473) );
  INV_X1 U6600 ( .A(n6193), .ZN(n6179) );
  INV_X1 U6601 ( .A(REIP_REG_17__SCAN_IN), .ZN(n7037) );
  INV_X1 U6602 ( .A(n5430), .ZN(n5573) );
  NOR4_X1 U6603 ( .A1(n6179), .A2(n7037), .A3(n5573), .A4(n5563), .ZN(n5550)
         );
  NAND4_X1 U6604 ( .A1(REIP_REG_18__SCAN_IN), .A2(n5550), .A3(
        REIP_REG_20__SCAN_IN), .A4(REIP_REG_19__SCAN_IN), .ZN(n5431) );
  NAND2_X1 U6605 ( .A1(n6206), .A2(n6193), .ZN(n6178) );
  NAND2_X1 U6606 ( .A1(n5431), .A2(n6178), .ZN(n5941) );
  NAND2_X1 U6607 ( .A1(n6171), .A2(n5432), .ZN(n5433) );
  NAND2_X1 U6608 ( .A1(n5941), .A2(n5433), .ZN(n5911) );
  INV_X1 U6609 ( .A(n5434), .ZN(n5435) );
  AND2_X1 U6610 ( .A1(n6178), .A2(n5435), .ZN(n5436) );
  NOR2_X1 U6611 ( .A1(n5437), .A2(n6737), .ZN(n5438) );
  NOR2_X1 U6612 ( .A1(n6206), .A2(n5438), .ZN(n5439) );
  NOR2_X1 U6613 ( .A1(n5517), .A2(n5439), .ZN(n5477) );
  OAI21_X1 U6614 ( .B1(n5484), .B2(n5473), .A(n5477), .ZN(n5476) );
  INV_X1 U6615 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6742) );
  INV_X1 U6616 ( .A(REIP_REG_30__SCAN_IN), .ZN(n5440) );
  OAI21_X1 U6617 ( .B1(n5484), .B2(n6742), .A(n5440), .ZN(n5453) );
  NOR2_X1 U6618 ( .A1(n5444), .A2(n5540), .ZN(n5461) );
  NAND2_X1 U6619 ( .A1(n5460), .A2(EBX_REG_30__SCAN_IN), .ZN(n5442) );
  NAND2_X1 U6620 ( .A1(n4168), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5441) );
  AND2_X1 U6621 ( .A1(n5442), .A2(n5441), .ZN(n5463) );
  INV_X1 U6622 ( .A(n5463), .ZN(n5443) );
  OAI21_X1 U6623 ( .B1(n5444), .B2(n5445), .A(n5443), .ZN(n5448) );
  OAI211_X1 U6624 ( .C1(n3173), .C2(n3174), .A(n5446), .B(n5463), .ZN(n5447)
         );
  OAI21_X1 U6625 ( .B1(n5461), .B2(n5448), .A(n5447), .ZN(n5799) );
  AOI22_X1 U6626 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n6148), .B1(n6133), 
        .B2(n5449), .ZN(n5451) );
  NAND2_X1 U6627 ( .A1(n6209), .A2(EBX_REG_30__SCAN_IN), .ZN(n5450) );
  OAI211_X1 U6628 ( .C1(n5799), .C2(n6095), .A(n5451), .B(n5450), .ZN(n5452)
         );
  AOI21_X1 U6629 ( .B1(n5476), .B2(n5453), .A(n5452), .ZN(n5454) );
  OAI21_X1 U6630 ( .B1(n5429), .B2(n6156), .A(n5454), .ZN(U2797) );
  AOI22_X1 U6631 ( .A1(n6238), .A2(DATAI_30_), .B1(n6241), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5458) );
  AND2_X1 U6632 ( .A1(n5455), .A2(n3488), .ZN(n5456) );
  NAND2_X1 U6633 ( .A1(n6242), .A2(DATAI_14_), .ZN(n5457) );
  OAI211_X1 U6634 ( .C1(n5429), .C2(n5684), .A(n5458), .B(n5457), .ZN(U2861)
         );
  INV_X1 U6635 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5459) );
  OAI22_X1 U6636 ( .A1(n5460), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4168), .ZN(n5465) );
  AOI21_X1 U6637 ( .B1(n5463), .B2(n5462), .A(n5461), .ZN(n5464) );
  INV_X1 U6638 ( .A(EBX_REG_31__SCAN_IN), .ZN(n7103) );
  OAI22_X1 U6639 ( .A1(n5793), .A2(n5671), .B1(n7103), .B2(n6231), .ZN(U2828)
         );
  NAND2_X1 U6640 ( .A1(n5467), .A2(n4148), .ZN(n5469) );
  AOI22_X1 U6641 ( .A1(n6238), .A2(DATAI_31_), .B1(n6241), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n5468) );
  OAI21_X1 U6642 ( .B1(n5466), .B2(n5469), .A(n5468), .ZN(U2860) );
  NAND2_X1 U6643 ( .A1(n6148), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5472)
         );
  INV_X1 U6644 ( .A(n5470), .ZN(n6661) );
  NAND4_X1 U6645 ( .A1(n5607), .A2(n4309), .A3(EBX_REG_31__SCAN_IN), .A4(n6661), .ZN(n5471) );
  INV_X1 U6646 ( .A(n5473), .ZN(n5474) );
  NOR3_X1 U6647 ( .A1(n5484), .A2(REIP_REG_31__SCAN_IN), .A3(n5474), .ZN(n5475) );
  NAND2_X1 U6648 ( .A1(n5691), .A2(n6110), .ZN(n5483) );
  INV_X1 U6649 ( .A(n5477), .ZN(n5493) );
  INV_X1 U6650 ( .A(n5689), .ZN(n5478) );
  AOI22_X1 U6651 ( .A1(PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n6148), .B1(n6133), 
        .B2(n5478), .ZN(n5480) );
  NAND2_X1 U6652 ( .A1(n6209), .A2(EBX_REG_29__SCAN_IN), .ZN(n5479) );
  OAI211_X1 U6653 ( .C1(n5809), .C2(n6095), .A(n5480), .B(n5479), .ZN(n5481)
         );
  AOI21_X1 U6654 ( .B1(n5493), .B2(REIP_REG_29__SCAN_IN), .A(n5481), .ZN(n5482) );
  OAI211_X1 U6655 ( .C1(REIP_REG_29__SCAN_IN), .C2(n5484), .A(n5483), .B(n5482), .ZN(U2798) );
  OAI21_X1 U6656 ( .B1(n5485), .B2(n5486), .A(n4071), .ZN(n5693) );
  INV_X1 U6657 ( .A(n5487), .ZN(n5696) );
  OAI22_X1 U6658 ( .A1(n5488), .A2(n6212), .B1(n6222), .B2(n5696), .ZN(n5489)
         );
  AOI21_X1 U6659 ( .B1(n6209), .B2(EBX_REG_28__SCAN_IN), .A(n5489), .ZN(n5490)
         );
  OAI21_X1 U6660 ( .B1(n5625), .B2(n6095), .A(n5490), .ZN(n5492) );
  NOR3_X1 U6661 ( .A1(n5507), .A2(REIP_REG_28__SCAN_IN), .A3(n6737), .ZN(n5491) );
  AOI211_X1 U6662 ( .C1(REIP_REG_28__SCAN_IN), .C2(n5493), .A(n5492), .B(n5491), .ZN(n5494) );
  OAI21_X1 U6663 ( .B1(n5693), .B2(n6156), .A(n5494), .ZN(U2799) );
  NAND2_X1 U6664 ( .A1(n5706), .A2(n6110), .ZN(n5506) );
  NAND2_X1 U6665 ( .A1(n5513), .A2(n5498), .ZN(n5499) );
  NAND2_X1 U6666 ( .A1(n5500), .A2(n5499), .ZN(n5814) );
  INV_X1 U6667 ( .A(n5704), .ZN(n5501) );
  AOI22_X1 U6668 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n6148), .B1(n6133), 
        .B2(n5501), .ZN(n5503) );
  NAND2_X1 U6669 ( .A1(n6209), .A2(EBX_REG_27__SCAN_IN), .ZN(n5502) );
  OAI211_X1 U6670 ( .C1(n5814), .C2(n6095), .A(n5503), .B(n5502), .ZN(n5504)
         );
  AOI21_X1 U6671 ( .B1(n5517), .B2(REIP_REG_27__SCAN_IN), .A(n5504), .ZN(n5505) );
  OAI211_X1 U6672 ( .C1(REIP_REG_27__SCAN_IN), .C2(n5507), .A(n5506), .B(n5505), .ZN(U2800) );
  OAI21_X1 U6673 ( .B1(n5508), .B2(n5509), .A(n5496), .ZN(n5711) );
  INV_X1 U6674 ( .A(n5510), .ZN(n5713) );
  OAI22_X1 U6675 ( .A1(n5511), .A2(n6212), .B1(n6222), .B2(n5713), .ZN(n5516)
         );
  OAI21_X1 U6676 ( .B1(n5512), .B2(n5514), .A(n5513), .ZN(n5822) );
  NOR2_X1 U6677 ( .A1(n5822), .A2(n6095), .ZN(n5515) );
  AOI211_X1 U6678 ( .C1(EBX_REG_26__SCAN_IN), .C2(n6209), .A(n5516), .B(n5515), 
        .ZN(n5520) );
  INV_X1 U6679 ( .A(n5906), .ZN(n5530) );
  NOR2_X1 U6680 ( .A1(n5530), .A2(n5905), .ZN(n5518) );
  OAI21_X1 U6681 ( .B1(n5518), .B2(REIP_REG_26__SCAN_IN), .A(n5517), .ZN(n5519) );
  OAI211_X1 U6682 ( .C1(n5711), .C2(n6156), .A(n5520), .B(n5519), .ZN(U2801)
         );
  OAI21_X1 U6683 ( .B1(n5521), .B2(n5523), .A(n5522), .ZN(n5726) );
  OAI21_X1 U6684 ( .B1(n5524), .B2(n5525), .A(n3141), .ZN(n5633) );
  INV_X1 U6685 ( .A(n5633), .ZN(n5836) );
  INV_X1 U6686 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5526) );
  OAI22_X1 U6687 ( .A1(n5526), .A2(n6212), .B1(n6222), .B2(n5728), .ZN(n5527)
         );
  AOI21_X1 U6688 ( .B1(n5836), .B2(n6214), .A(n5527), .ZN(n5528) );
  OAI21_X1 U6689 ( .B1(n5529), .B2(n6150), .A(n5528), .ZN(n5532) );
  NOR2_X1 U6690 ( .A1(n5530), .A2(REIP_REG_24__SCAN_IN), .ZN(n5531) );
  AOI211_X1 U6691 ( .C1(REIP_REG_24__SCAN_IN), .C2(n5911), .A(n5532), .B(n5531), .ZN(n5533) );
  OAI21_X1 U6692 ( .B1(n5726), .B2(n6156), .A(n5533), .ZN(U2803) );
  INV_X1 U6693 ( .A(n5536), .ZN(n5537) );
  AOI21_X1 U6694 ( .B1(n5538), .B2(n5534), .A(n5537), .ZN(n6232) );
  INV_X1 U6695 ( .A(n6232), .ZN(n5668) );
  INV_X1 U6696 ( .A(n5762), .ZN(n5549) );
  NAND2_X1 U6697 ( .A1(n5656), .A2(n3174), .ZN(n5543) );
  INV_X1 U6698 ( .A(n5539), .ZN(n5541) );
  NAND2_X1 U6699 ( .A1(n5541), .A2(n5540), .ZN(n5542) );
  NAND2_X1 U6700 ( .A1(n5543), .A2(n5542), .ZN(n5546) );
  INV_X1 U6701 ( .A(n5546), .ZN(n5545) );
  NAND2_X1 U6702 ( .A1(n5545), .A2(n5544), .ZN(n5548) );
  INV_X1 U6703 ( .A(n5544), .ZN(n5547) );
  NAND2_X1 U6704 ( .A1(n5547), .A2(n5546), .ZN(n5666) );
  AND2_X1 U6705 ( .A1(n5548), .A2(n5666), .ZN(n5883) );
  INV_X1 U6706 ( .A(n5883), .ZN(n5669) );
  OAI22_X1 U6707 ( .A1(n5549), .A2(n6222), .B1(n6095), .B2(n5669), .ZN(n5554)
         );
  INV_X1 U6708 ( .A(n5550), .ZN(n5551) );
  NAND2_X1 U6709 ( .A1(n6178), .A2(n5551), .ZN(n6087) );
  AOI21_X1 U6710 ( .B1(n6148), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6182), 
        .ZN(n5552) );
  OAI221_X1 U6711 ( .B1(REIP_REG_18__SCAN_IN), .B2(n5947), .C1(n5878), .C2(
        n6087), .A(n5552), .ZN(n5553) );
  AOI211_X1 U6712 ( .C1(n6209), .C2(EBX_REG_18__SCAN_IN), .A(n5554), .B(n5553), 
        .ZN(n5555) );
  OAI21_X1 U6713 ( .B1(n5668), .B2(n6156), .A(n5555), .ZN(U2809) );
  AND2_X1 U6714 ( .A1(n5557), .A2(n5556), .ZN(n5559) );
  OR2_X1 U6715 ( .A1(n5559), .A2(n5558), .ZN(n5767) );
  INV_X1 U6716 ( .A(n5769), .ZN(n5569) );
  OR2_X1 U6717 ( .A1(n5560), .A2(n5394), .ZN(n5561) );
  NAND2_X1 U6718 ( .A1(n5561), .A2(n6020), .ZN(n5886) );
  AOI21_X1 U6719 ( .B1(n6148), .B2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6182), 
        .ZN(n5562) );
  OAI21_X1 U6720 ( .B1(n6095), .B2(n5886), .A(n5562), .ZN(n5568) );
  OAI21_X1 U6721 ( .B1(REIP_REG_16__SCAN_IN), .B2(REIP_REG_15__SCAN_IN), .A(
        n5563), .ZN(n5565) );
  AOI22_X1 U6722 ( .A1(EBX_REG_16__SCAN_IN), .A2(n6209), .B1(
        REIP_REG_16__SCAN_IN), .B2(n5574), .ZN(n5564) );
  OAI21_X1 U6723 ( .B1(n5566), .B2(n5565), .A(n5564), .ZN(n5567) );
  AOI211_X1 U6724 ( .C1(n6133), .C2(n5569), .A(n5568), .B(n5567), .ZN(n5570)
         );
  OAI21_X1 U6725 ( .B1(n5767), .B2(n6156), .A(n5570), .ZN(U2811) );
  INV_X1 U6726 ( .A(n5571), .ZN(n6042) );
  AOI21_X1 U6727 ( .B1(n6148), .B2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n6182), 
        .ZN(n5572) );
  OAI21_X1 U6728 ( .B1(n5783), .B2(n6222), .A(n5572), .ZN(n5579) );
  NAND2_X1 U6729 ( .A1(n6171), .A2(n5573), .ZN(n5576) );
  AOI22_X1 U6730 ( .A1(EBX_REG_14__SCAN_IN), .A2(n6209), .B1(
        REIP_REG_14__SCAN_IN), .B2(n5574), .ZN(n5575) );
  OAI21_X1 U6731 ( .B1(n5577), .B2(n5576), .A(n5575), .ZN(n5578) );
  AOI211_X1 U6732 ( .C1(n6214), .C2(n6042), .A(n5579), .B(n5578), .ZN(n5580)
         );
  OAI21_X1 U6733 ( .B1(n5787), .B2(n6156), .A(n5580), .ZN(U2813) );
  NAND2_X1 U6734 ( .A1(n6171), .A2(n6100), .ZN(n5583) );
  INV_X1 U6735 ( .A(n5583), .ZN(n5589) );
  INV_X1 U6736 ( .A(n6373), .ZN(n5581) );
  OAI22_X1 U6737 ( .A1(n5582), .A2(n6222), .B1(n6095), .B2(n5581), .ZN(n5587)
         );
  NAND2_X1 U6738 ( .A1(n6193), .A2(n5583), .ZN(n6108) );
  AOI22_X1 U6739 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n6148), .B1(
        REIP_REG_11__SCAN_IN), .B2(n6108), .ZN(n5584) );
  OAI211_X1 U6740 ( .C1(n6150), .C2(n5585), .A(n5584), .B(n6163), .ZN(n5586)
         );
  AOI211_X1 U6741 ( .C1(n5589), .C2(n5588), .A(n5587), .B(n5586), .ZN(n5590)
         );
  OAI21_X1 U6742 ( .B1(n6156), .B2(n5591), .A(n5590), .ZN(U2816) );
  INV_X1 U6743 ( .A(n5592), .ZN(n5596) );
  INV_X1 U6744 ( .A(n5597), .ZN(n6121) );
  INV_X1 U6745 ( .A(n5593), .ZN(n5594) );
  NAND3_X1 U6746 ( .A1(n6171), .A2(n6121), .A3(n5594), .ZN(n5595) );
  OAI21_X1 U6747 ( .B1(n5596), .B2(n6222), .A(n5595), .ZN(n5601) );
  OAI21_X1 U6748 ( .B1(n6206), .B2(n5597), .A(n6193), .ZN(n6127) );
  AOI22_X1 U6749 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n6148), .B1(
        REIP_REG_8__SCAN_IN), .B2(n6127), .ZN(n5598) );
  OAI211_X1 U6750 ( .C1(n6150), .C2(n5599), .A(n5598), .B(n6163), .ZN(n5600)
         );
  AOI211_X1 U6751 ( .C1(n5602), .C2(n6214), .A(n5601), .B(n5600), .ZN(n5603)
         );
  OAI21_X1 U6752 ( .B1(n6156), .B2(n5604), .A(n5603), .ZN(U2819) );
  NAND2_X1 U6753 ( .A1(n5607), .A2(n5605), .ZN(n6217) );
  NAND2_X1 U6754 ( .A1(n5607), .A2(n5606), .ZN(n5608) );
  NAND2_X1 U6755 ( .A1(n5609), .A2(n6220), .ZN(n5615) );
  NAND2_X1 U6756 ( .A1(n6209), .A2(EBX_REG_1__SCAN_IN), .ZN(n5611) );
  AOI22_X1 U6757 ( .A1(n6148), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6179), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n5610) );
  OAI211_X1 U6758 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n6222), .A(n5611), 
        .B(n5610), .ZN(n5613) );
  OAI22_X1 U6759 ( .A1(n4539), .A2(n6095), .B1(n6206), .B2(REIP_REG_1__SCAN_IN), .ZN(n5612) );
  NOR2_X1 U6760 ( .A1(n5613), .A2(n5612), .ZN(n5614) );
  OAI211_X1 U6761 ( .C1(n6217), .C2(n5616), .A(n5615), .B(n5614), .ZN(U2826)
         );
  OAI21_X1 U6762 ( .B1(n6148), .B2(n6133), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5617) );
  OAI21_X1 U6763 ( .B1(n6412), .B2(n6095), .A(n5617), .ZN(n5620) );
  NOR2_X1 U6764 ( .A1(n6150), .A2(n5618), .ZN(n5619) );
  AOI211_X1 U6765 ( .C1(REIP_REG_0__SCAN_IN), .C2(n6178), .A(n5620), .B(n5619), 
        .ZN(n5623) );
  INV_X1 U6766 ( .A(n6217), .ZN(n5621) );
  NAND2_X1 U6767 ( .A1(n5621), .A2(n3133), .ZN(n5622) );
  OAI211_X1 U6768 ( .C1(n6371), .C2(n6166), .A(n5623), .B(n5622), .ZN(U2827)
         );
  OAI222_X1 U6769 ( .A1(n5625), .A2(n5671), .B1(n5624), .B2(n6231), .C1(n5693), 
        .C2(n5670), .ZN(U2831) );
  INV_X1 U6770 ( .A(n5706), .ZN(n5679) );
  OAI222_X1 U6771 ( .A1(n5626), .A2(n6231), .B1(n5671), .B2(n5814), .C1(n5679), 
        .C2(n5670), .ZN(U2832) );
  OAI222_X1 U6772 ( .A1(n5627), .A2(n6231), .B1(n5671), .B2(n5822), .C1(n5711), 
        .C2(n5670), .ZN(U2833) );
  AOI21_X1 U6773 ( .B1(n5628), .B2(n5522), .A(n5508), .ZN(n5977) );
  INV_X1 U6774 ( .A(n5977), .ZN(n5632) );
  AND2_X1 U6775 ( .A1(n3141), .A2(n5629), .ZN(n5630) );
  OR2_X1 U6776 ( .A1(n5512), .A2(n5630), .ZN(n5904) );
  OAI222_X1 U6777 ( .A1(n5632), .A2(n5670), .B1(n6231), .B2(n5631), .C1(n5904), 
        .C2(n5671), .ZN(U2834) );
  OAI222_X1 U6778 ( .A1(n5670), .A2(n5726), .B1(n6231), .B2(n5529), .C1(n5633), 
        .C2(n5671), .ZN(U2835) );
  AOI21_X1 U6779 ( .B1(n5635), .B2(n5634), .A(n5521), .ZN(n5958) );
  NOR2_X1 U6780 ( .A1(n5637), .A2(n5636), .ZN(n5638) );
  OR2_X1 U6781 ( .A1(n5524), .A2(n5638), .ZN(n5912) );
  OAI22_X1 U6782 ( .A1(n5671), .A2(n5912), .B1(n5639), .B2(n6231), .ZN(n5640)
         );
  AOI21_X1 U6783 ( .B1(n5958), .B2(n6228), .A(n5640), .ZN(n5641) );
  INV_X1 U6784 ( .A(n5641), .ZN(U2836) );
  OAI21_X1 U6785 ( .B1(n5642), .B2(n5643), .A(n5634), .ZN(n5921) );
  XNOR2_X1 U6786 ( .A(n5648), .B(n5644), .ZN(n5922) );
  OAI222_X1 U6787 ( .A1(n5670), .A2(n5921), .B1(n5671), .B2(n5922), .C1(n5645), 
        .C2(n6231), .ZN(U2837) );
  AOI21_X1 U6788 ( .B1(n5647), .B2(n5646), .A(n5642), .ZN(n5964) );
  INV_X1 U6789 ( .A(n5964), .ZN(n5752) );
  INV_X1 U6790 ( .A(n5648), .ZN(n5649) );
  AOI21_X1 U6791 ( .B1(n5651), .B2(n5650), .A(n5649), .ZN(n5932) );
  INV_X1 U6792 ( .A(n5932), .ZN(n5652) );
  OAI222_X1 U6793 ( .A1(n5752), .A2(n5670), .B1(n6231), .B2(n5653), .C1(n5652), 
        .C2(n5671), .ZN(U2838) );
  OAI21_X1 U6794 ( .B1(n5654), .B2(n5655), .A(n5646), .ZN(n5939) );
  NAND2_X1 U6795 ( .A1(n5658), .A2(n5656), .ZN(n5657) );
  OAI21_X1 U6796 ( .B1(n5658), .B2(n3174), .A(n5657), .ZN(n5661) );
  INV_X1 U6797 ( .A(n5659), .ZN(n5660) );
  XNOR2_X1 U6798 ( .A(n5661), .B(n5660), .ZN(n5940) );
  INV_X1 U6799 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5662) );
  OAI222_X1 U6800 ( .A1(n5939), .A2(n5670), .B1(n5671), .B2(n5940), .C1(n6231), 
        .C2(n5662), .ZN(U2839) );
  AND2_X1 U6801 ( .A1(n5536), .A2(n5663), .ZN(n5664) );
  OR2_X1 U6802 ( .A1(n5654), .A2(n5664), .ZN(n5988) );
  XNOR2_X1 U6803 ( .A(n5666), .B(n5665), .ZN(n6013) );
  OAI222_X1 U6804 ( .A1(n5988), .A2(n5670), .B1(n5671), .B2(n6013), .C1(n5667), 
        .C2(n6231), .ZN(U2840) );
  OAI222_X1 U6805 ( .A1(n5669), .A2(n5671), .B1(n6231), .B2(n4212), .C1(n5670), 
        .C2(n5668), .ZN(U2841) );
  OAI222_X1 U6806 ( .A1(n5886), .A2(n5671), .B1(n6231), .B2(n4202), .C1(n5670), 
        .C2(n5767), .ZN(U2843) );
  AOI22_X1 U6807 ( .A1(n6238), .A2(DATAI_29_), .B1(n6241), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5673) );
  NAND2_X1 U6808 ( .A1(n6242), .A2(DATAI_13_), .ZN(n5672) );
  OAI211_X1 U6809 ( .C1(n5674), .C2(n5684), .A(n5673), .B(n5672), .ZN(U2862)
         );
  AOI22_X1 U6810 ( .A1(n6238), .A2(DATAI_28_), .B1(n6241), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5676) );
  NAND2_X1 U6811 ( .A1(n6242), .A2(DATAI_12_), .ZN(n5675) );
  OAI211_X1 U6812 ( .C1(n5693), .C2(n5684), .A(n5676), .B(n5675), .ZN(U2863)
         );
  AOI22_X1 U6813 ( .A1(n6238), .A2(DATAI_27_), .B1(n6241), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5678) );
  NAND2_X1 U6814 ( .A1(n6242), .A2(DATAI_11_), .ZN(n5677) );
  OAI211_X1 U6815 ( .C1(n5679), .C2(n5684), .A(n5678), .B(n5677), .ZN(U2864)
         );
  AOI22_X1 U6816 ( .A1(n6238), .A2(DATAI_26_), .B1(n6241), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5681) );
  NAND2_X1 U6817 ( .A1(n6242), .A2(DATAI_10_), .ZN(n5680) );
  OAI211_X1 U6818 ( .C1(n5711), .C2(n5684), .A(n5681), .B(n5680), .ZN(U2865)
         );
  AOI22_X1 U6819 ( .A1(n6238), .A2(DATAI_24_), .B1(n6241), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5683) );
  NAND2_X1 U6820 ( .A1(n6242), .A2(DATAI_8_), .ZN(n5682) );
  OAI211_X1 U6821 ( .C1(n5726), .C2(n5684), .A(n5683), .B(n5682), .ZN(U2867)
         );
  AOI21_X1 U6822 ( .B1(n5805), .B2(n5686), .A(n5685), .ZN(n5687) );
  XNOR2_X1 U6823 ( .A(n5687), .B(n7006), .ZN(n5813) );
  AND2_X1 U6824 ( .A1(n6351), .A2(REIP_REG_29__SCAN_IN), .ZN(n5806) );
  AOI21_X1 U6825 ( .B1(n6350), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5806), 
        .ZN(n5688) );
  OAI21_X1 U6826 ( .B1(n6361), .B2(n5689), .A(n5688), .ZN(n5690) );
  AOI21_X1 U6827 ( .B1(n5691), .B2(n6356), .A(n5690), .ZN(n5692) );
  OAI21_X1 U6828 ( .B1(n5813), .B2(n6068), .A(n5692), .ZN(U2957) );
  INV_X1 U6829 ( .A(n5693), .ZN(n5698) );
  AOI21_X1 U6830 ( .B1(n6350), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5694), 
        .ZN(n5695) );
  OAI21_X1 U6831 ( .B1(n6361), .B2(n5696), .A(n5695), .ZN(n5697) );
  AOI21_X1 U6832 ( .B1(n5698), .B2(n6356), .A(n5697), .ZN(n5699) );
  OAI21_X1 U6833 ( .B1(n5700), .B2(n6068), .A(n5699), .ZN(U2958) );
  NAND2_X1 U6834 ( .A1(n4417), .A2(n5701), .ZN(n5702) );
  XNOR2_X1 U6835 ( .A(n5702), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5821)
         );
  AND2_X1 U6836 ( .A1(n6351), .A2(REIP_REG_27__SCAN_IN), .ZN(n5815) );
  AOI21_X1 U6837 ( .B1(n6350), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5815), 
        .ZN(n5703) );
  OAI21_X1 U6838 ( .B1(n6361), .B2(n5704), .A(n5703), .ZN(n5705) );
  AOI21_X1 U6839 ( .B1(n5706), .B2(n6356), .A(n5705), .ZN(n5707) );
  OAI21_X1 U6840 ( .B1(n5821), .B2(n6068), .A(n5707), .ZN(U2959) );
  NOR2_X1 U6841 ( .A1(n5709), .A2(n5708), .ZN(n5710) );
  XOR2_X1 U6842 ( .A(n5710), .B(n5416), .Z(n5830) );
  INV_X1 U6843 ( .A(n5711), .ZN(n5715) );
  AND2_X1 U6844 ( .A1(n6351), .A2(REIP_REG_26__SCAN_IN), .ZN(n5824) );
  AOI21_X1 U6845 ( .B1(n6350), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5824), 
        .ZN(n5712) );
  OAI21_X1 U6846 ( .B1(n6361), .B2(n5713), .A(n5712), .ZN(n5714) );
  AOI21_X1 U6847 ( .B1(n5715), .B2(n6356), .A(n5714), .ZN(n5716) );
  OAI21_X1 U6848 ( .B1(n5830), .B2(n6068), .A(n5716), .ZN(U2960) );
  INV_X1 U6849 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n7085) );
  NAND2_X1 U6850 ( .A1(n4327), .A2(n7085), .ZN(n5718) );
  OR2_X1 U6851 ( .A1(n4327), .A2(n7085), .ZN(n5981) );
  INV_X1 U6852 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5719) );
  NAND2_X1 U6853 ( .A1(n4327), .A2(n5719), .ZN(n5721) );
  NOR2_X1 U6854 ( .A1(n4327), .A2(n5719), .ZN(n5720) );
  XNOR2_X1 U6855 ( .A(n4327), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5748)
         );
  NOR2_X1 U6856 ( .A1(n4327), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5738)
         );
  INV_X1 U6857 ( .A(n5732), .ZN(n5723) );
  INV_X1 U6858 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5722) );
  INV_X1 U6859 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5860) );
  INV_X1 U6860 ( .A(n5726), .ZN(n5730) );
  INV_X1 U6861 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6732) );
  NOR2_X1 U6862 ( .A1(n6401), .A2(n6732), .ZN(n5835) );
  AOI21_X1 U6863 ( .B1(n6350), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5835), 
        .ZN(n5727) );
  OAI21_X1 U6864 ( .B1(n6361), .B2(n5728), .A(n5727), .ZN(n5729) );
  AOI21_X1 U6865 ( .B1(n5730), .B2(n6356), .A(n5729), .ZN(n5731) );
  OAI21_X1 U6866 ( .B1(n5838), .B2(n6068), .A(n5731), .ZN(U2962) );
  INV_X1 U6867 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6909) );
  OR3_X1 U6868 ( .A1(n3246), .A2(n5994), .A3(n6909), .ZN(n5997) );
  NAND3_X1 U6869 ( .A1(n5848), .A2(n5863), .A3(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5733) );
  OAI21_X1 U6870 ( .B1(n5997), .B2(n5733), .A(n5732), .ZN(n5734) );
  XNOR2_X1 U6871 ( .A(n5734), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5845)
         );
  NAND2_X1 U6872 ( .A1(n6368), .A2(REIP_REG_23__SCAN_IN), .ZN(n5839) );
  NAND2_X1 U6873 ( .A1(n6350), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5735)
         );
  OAI211_X1 U6874 ( .C1(n6361), .C2(n5918), .A(n5839), .B(n5735), .ZN(n5736)
         );
  AOI21_X1 U6875 ( .B1(n5958), .B2(n6356), .A(n5736), .ZN(n5737) );
  OAI21_X1 U6876 ( .B1(n5845), .B2(n6068), .A(n5737), .ZN(U2963) );
  AOI21_X1 U6877 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n4327), .A(n5738), 
        .ZN(n5740) );
  XOR2_X1 U6878 ( .A(n5740), .B(n5739), .Z(n5853) );
  NAND2_X1 U6879 ( .A1(n6368), .A2(REIP_REG_22__SCAN_IN), .ZN(n5846) );
  OAI21_X1 U6880 ( .B1(n6365), .B2(n5741), .A(n5846), .ZN(n5743) );
  NOR2_X1 U6881 ( .A1(n5921), .A2(n6370), .ZN(n5742) );
  AOI211_X1 U6882 ( .C1(n5776), .C2(n5920), .A(n5743), .B(n5742), .ZN(n5744)
         );
  OAI21_X1 U6883 ( .B1(n5853), .B2(n6068), .A(n5744), .ZN(U2964) );
  INV_X1 U6884 ( .A(n5745), .ZN(n5746) );
  OAI21_X1 U6885 ( .B1(n5748), .B2(n5747), .A(n5746), .ZN(n5854) );
  NAND2_X1 U6886 ( .A1(n5854), .A2(n6367), .ZN(n5751) );
  AND2_X1 U6887 ( .A1(n6351), .A2(REIP_REG_21__SCAN_IN), .ZN(n5857) );
  NOR2_X1 U6888 ( .A1(n6361), .A2(n5930), .ZN(n5749) );
  AOI211_X1 U6889 ( .C1(n6350), .C2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n5857), 
        .B(n5749), .ZN(n5750) );
  OAI211_X1 U6890 ( .C1(n5989), .C2(n5752), .A(n5751), .B(n5750), .ZN(U2965)
         );
  XNOR2_X1 U6891 ( .A(n4327), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5753)
         );
  XNOR2_X1 U6892 ( .A(n5754), .B(n5753), .ZN(n5876) );
  NAND2_X1 U6893 ( .A1(n6368), .A2(REIP_REG_20__SCAN_IN), .ZN(n5870) );
  OAI21_X1 U6894 ( .B1(n6365), .B2(n5946), .A(n5870), .ZN(n5756) );
  NOR2_X1 U6895 ( .A1(n5939), .A2(n6370), .ZN(n5755) );
  AOI211_X1 U6896 ( .C1(n5776), .C2(n5938), .A(n5756), .B(n5755), .ZN(n5757)
         );
  OAI21_X1 U6897 ( .B1(n5876), .B2(n6068), .A(n5757), .ZN(U2966) );
  OR4_X1 U6898 ( .A1(n5758), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A4(n4327), .ZN(n5998) );
  NAND2_X1 U6899 ( .A1(n5997), .A2(n5998), .ZN(n5759) );
  XNOR2_X1 U6900 ( .A(n5759), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5885)
         );
  OAI22_X1 U6901 ( .A1(n6365), .A2(n5760), .B1(n6401), .B2(n5878), .ZN(n5761)
         );
  AOI21_X1 U6902 ( .B1(n5776), .B2(n5762), .A(n5761), .ZN(n5764) );
  NAND2_X1 U6903 ( .A1(n6232), .A2(n6356), .ZN(n5763) );
  OAI211_X1 U6904 ( .C1(n5885), .C2(n6068), .A(n5764), .B(n5763), .ZN(U2968)
         );
  XNOR2_X1 U6905 ( .A(n4327), .B(n5893), .ZN(n5766) );
  XNOR2_X1 U6906 ( .A(n5765), .B(n5766), .ZN(n5898) );
  INV_X1 U6907 ( .A(n5767), .ZN(n6240) );
  AND2_X1 U6908 ( .A1(n6351), .A2(REIP_REG_16__SCAN_IN), .ZN(n5895) );
  AOI21_X1 U6909 ( .B1(n6350), .B2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n5895), 
        .ZN(n5768) );
  OAI21_X1 U6910 ( .B1(n5769), .B2(n6361), .A(n5768), .ZN(n5770) );
  AOI21_X1 U6911 ( .B1(n6240), .B2(n6356), .A(n5770), .ZN(n5771) );
  OAI21_X1 U6912 ( .B1(n5898), .B2(n6068), .A(n5771), .ZN(U2970) );
  XNOR2_X1 U6913 ( .A(n5772), .B(n5773), .ZN(n6034) );
  NAND2_X1 U6914 ( .A1(n6034), .A2(n6367), .ZN(n5779) );
  NAND2_X1 U6915 ( .A1(n6368), .A2(REIP_REG_15__SCAN_IN), .ZN(n6029) );
  OAI21_X1 U6916 ( .B1(n6365), .B2(n5774), .A(n6029), .ZN(n5775) );
  AOI21_X1 U6917 ( .B1(n5777), .B2(n5776), .A(n5775), .ZN(n5778) );
  OAI211_X1 U6918 ( .C1(n6370), .C2(n5780), .A(n5779), .B(n5778), .ZN(U2971)
         );
  XNOR2_X1 U6919 ( .A(n4327), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5781)
         );
  XNOR2_X1 U6920 ( .A(n5782), .B(n5781), .ZN(n6044) );
  NAND2_X1 U6921 ( .A1(n6044), .A2(n6367), .ZN(n5786) );
  NOR2_X1 U6922 ( .A1(n6401), .A2(n6719), .ZN(n6041) );
  NOR2_X1 U6923 ( .A1(n6361), .A2(n5783), .ZN(n5784) );
  AOI211_X1 U6924 ( .C1(n6350), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n6041), 
        .B(n5784), .ZN(n5785) );
  OAI211_X1 U6925 ( .C1(n5989), .C2(n5787), .A(n5786), .B(n5785), .ZN(U2972)
         );
  AOI21_X1 U6926 ( .B1(n5788), .B2(n5887), .A(n5818), .ZN(n5804) );
  OAI21_X1 U6927 ( .B1(n7006), .B2(n3222), .A(n5887), .ZN(n5789) );
  NAND2_X1 U6928 ( .A1(n5804), .A2(n5789), .ZN(n5801) );
  NAND4_X1 U6929 ( .A1(n5817), .A2(n3156), .A3(INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n5790), .ZN(n5792) );
  OAI211_X1 U6930 ( .C1(n5793), .C2(n6413), .A(n5792), .B(n5791), .ZN(n5794)
         );
  AOI21_X1 U6931 ( .B1(n5801), .B2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n5794), 
        .ZN(n5795) );
  OAI21_X1 U6932 ( .B1(n5796), .B2(n6014), .A(n5795), .ZN(U2987) );
  NAND3_X1 U6933 ( .A1(n5817), .A2(n3156), .A3(n3222), .ZN(n5798) );
  OAI211_X1 U6934 ( .C1(n6413), .C2(n5799), .A(n5798), .B(n5797), .ZN(n5800)
         );
  AOI21_X1 U6935 ( .B1(n5801), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5800), 
        .ZN(n5802) );
  OAI21_X1 U6936 ( .B1(n5803), .B2(n6014), .A(n5802), .ZN(U2988) );
  INV_X1 U6937 ( .A(n5804), .ZN(n5811) );
  NAND3_X1 U6938 ( .A1(n5817), .A2(n5805), .A3(n7006), .ZN(n5808) );
  INV_X1 U6939 ( .A(n5806), .ZN(n5807) );
  OAI211_X1 U6940 ( .C1(n6413), .C2(n5809), .A(n5808), .B(n5807), .ZN(n5810)
         );
  AOI21_X1 U6941 ( .B1(n5811), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5810), 
        .ZN(n5812) );
  OAI21_X1 U6942 ( .B1(n5813), .B2(n6014), .A(n5812), .ZN(U2989) );
  NOR2_X1 U6943 ( .A1(n5814), .A2(n6413), .ZN(n5816) );
  AOI211_X1 U6944 ( .C1(n5817), .C2(n7001), .A(n5816), .B(n5815), .ZN(n5820)
         );
  NAND2_X1 U6945 ( .A1(n5818), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5819) );
  OAI211_X1 U6946 ( .C1(n5821), .C2(n6014), .A(n5820), .B(n5819), .ZN(U2991)
         );
  INV_X1 U6947 ( .A(n5822), .ZN(n5825) );
  NOR3_X1 U6948 ( .A1(n5826), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .A3(n6010), 
        .ZN(n5823) );
  AOI211_X1 U6949 ( .C1(n6389), .C2(n5825), .A(n5824), .B(n5823), .ZN(n5829)
         );
  INV_X1 U6950 ( .A(n6011), .ZN(n5827) );
  NOR2_X1 U6951 ( .A1(n5826), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6005)
         );
  OAI21_X1 U6952 ( .B1(n5827), .B2(n6005), .A(INSTADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n5828) );
  OAI211_X1 U6953 ( .C1(n5830), .C2(n6014), .A(n5829), .B(n5828), .ZN(U2992)
         );
  INV_X1 U6954 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5833) );
  INV_X1 U6955 ( .A(n5831), .ZN(n5840) );
  AOI211_X1 U6956 ( .C1(n5833), .C2(n5840), .A(n5832), .B(n6011), .ZN(n5834)
         );
  AOI211_X1 U6957 ( .C1(n6389), .C2(n5836), .A(n5835), .B(n5834), .ZN(n5837)
         );
  OAI21_X1 U6958 ( .B1(n5838), .B2(n6014), .A(n5837), .ZN(U2994) );
  OAI21_X1 U6959 ( .B1(n5912), .B2(n6413), .A(n5839), .ZN(n5842) );
  NOR2_X1 U6960 ( .A1(n5840), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5841)
         );
  AOI211_X1 U6961 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n5843), .A(n5842), .B(n5841), .ZN(n5844) );
  OAI21_X1 U6962 ( .B1(n5845), .B2(n6014), .A(n5844), .ZN(U2995) );
  INV_X1 U6963 ( .A(n5861), .ZN(n5851) );
  OAI21_X1 U6964 ( .B1(n6413), .B2(n5922), .A(n5846), .ZN(n5850) );
  NOR3_X1 U6965 ( .A1(n5855), .A2(n5848), .A3(n5847), .ZN(n5849) );
  AOI211_X1 U6966 ( .C1(n5851), .C2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n5850), .B(n5849), .ZN(n5852) );
  OAI21_X1 U6967 ( .B1(n5853), .B2(n6014), .A(n5852), .ZN(U2996) );
  NAND2_X1 U6968 ( .A1(n5854), .A2(n6415), .ZN(n5859) );
  NOR2_X1 U6969 ( .A1(n5855), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5856)
         );
  AOI211_X1 U6970 ( .C1(n6389), .C2(n5932), .A(n5857), .B(n5856), .ZN(n5858)
         );
  OAI211_X1 U6971 ( .C1(n5861), .C2(n5860), .A(n5859), .B(n5858), .ZN(U2997)
         );
  NAND2_X1 U6972 ( .A1(n6026), .A2(n5862), .ZN(n6019) );
  INV_X1 U6973 ( .A(n6019), .ZN(n5874) );
  NOR2_X1 U6974 ( .A1(n5864), .A2(n5863), .ZN(n5873) );
  OAI221_X1 U6975 ( .B1(n5867), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .C1(
        n5867), .C2(n5866), .A(n5865), .ZN(n6025) );
  AOI21_X1 U6976 ( .B1(n5868), .B2(n6909), .A(n6025), .ZN(n5880) );
  NAND2_X1 U6977 ( .A1(n5887), .A2(n5879), .ZN(n5869) );
  NAND2_X1 U6978 ( .A1(n5880), .A2(n5869), .ZN(n6012) );
  NAND2_X1 U6979 ( .A1(n6012), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5871) );
  OAI211_X1 U6980 ( .C1(n5940), .C2(n6413), .A(n5871), .B(n5870), .ZN(n5872)
         );
  AOI21_X1 U6981 ( .B1(n5874), .B2(n5873), .A(n5872), .ZN(n5875) );
  OAI21_X1 U6982 ( .B1(n5876), .B2(n6014), .A(n5875), .ZN(U2998) );
  NAND3_X1 U6983 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n6026), .A3(n5879), .ZN(n5877) );
  OAI21_X1 U6984 ( .B1(n6401), .B2(n5878), .A(n5877), .ZN(n5882) );
  NOR2_X1 U6985 ( .A1(n5880), .A2(n5879), .ZN(n5881) );
  AOI211_X1 U6986 ( .C1(n6389), .C2(n5883), .A(n5882), .B(n5881), .ZN(n5884)
         );
  OAI21_X1 U6987 ( .B1(n5885), .B2(n6014), .A(n5884), .ZN(U3000) );
  INV_X1 U6988 ( .A(n5886), .ZN(n5896) );
  AOI21_X1 U6989 ( .B1(n5888), .B2(n5887), .A(n6374), .ZN(n6037) );
  NAND2_X1 U6990 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6043), .ZN(n6032) );
  OAI21_X1 U6991 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A(n5891), .ZN(n5892) );
  OAI22_X1 U6992 ( .A1(n6037), .A2(n5893), .B1(n6032), .B2(n5892), .ZN(n5894)
         );
  AOI211_X1 U6993 ( .C1(n6389), .C2(n5896), .A(n5895), .B(n5894), .ZN(n5897)
         );
  OAI21_X1 U6994 ( .B1(n5898), .B2(n6014), .A(n5897), .ZN(U3002) );
  INV_X1 U6995 ( .A(n5899), .ZN(n5901) );
  OAI22_X1 U6996 ( .A1(n5901), .A2(n6763), .B1(n5900), .B2(n6664), .ZN(n5902)
         );
  MUX2_X1 U6997 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5902), .S(n6761), 
        .Z(U3456) );
  AND2_X1 U6998 ( .A1(n6262), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI22_X1 U6999 ( .A1(EBX_REG_25__SCAN_IN), .A2(n6209), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6148), .ZN(n5910) );
  INV_X1 U7000 ( .A(n5980), .ZN(n5903) );
  AOI22_X1 U7001 ( .A1(n5903), .A2(n6133), .B1(REIP_REG_25__SCAN_IN), .B2(
        n5911), .ZN(n5909) );
  INV_X1 U7002 ( .A(n5904), .ZN(n6006) );
  AOI22_X1 U7003 ( .A1(n5977), .A2(n6110), .B1(n6214), .B2(n6006), .ZN(n5908)
         );
  OAI211_X1 U7004 ( .C1(REIP_REG_24__SCAN_IN), .C2(REIP_REG_25__SCAN_IN), .A(
        n5906), .B(n5905), .ZN(n5907) );
  NAND4_X1 U7005 ( .A1(n5910), .A2(n5909), .A3(n5908), .A4(n5907), .ZN(U2802)
         );
  AOI22_X1 U7006 ( .A1(EBX_REG_23__SCAN_IN), .A2(n6209), .B1(
        PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n6148), .ZN(n5917) );
  INV_X1 U7007 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6726) );
  NOR2_X1 U7008 ( .A1(n6726), .A2(n5924), .ZN(n5919) );
  AOI21_X1 U7009 ( .B1(REIP_REG_22__SCAN_IN), .B2(n5919), .A(
        REIP_REG_23__SCAN_IN), .ZN(n5914) );
  INV_X1 U7010 ( .A(n5911), .ZN(n5913) );
  OAI22_X1 U7011 ( .A1(n5914), .A2(n5913), .B1(n5912), .B2(n6095), .ZN(n5915)
         );
  AOI21_X1 U7012 ( .B1(n5958), .B2(n6110), .A(n5915), .ZN(n5916) );
  OAI211_X1 U7013 ( .C1(n5918), .C2(n6222), .A(n5917), .B(n5916), .ZN(U2804)
         );
  AOI22_X1 U7014 ( .A1(EBX_REG_22__SCAN_IN), .A2(n6209), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6148), .ZN(n5929) );
  INV_X1 U7015 ( .A(REIP_REG_22__SCAN_IN), .ZN(n7063) );
  AOI22_X1 U7016 ( .A1(n5920), .A2(n6133), .B1(n5919), .B2(n7063), .ZN(n5928)
         );
  INV_X1 U7017 ( .A(n5921), .ZN(n5961) );
  INV_X1 U7018 ( .A(n5922), .ZN(n5923) );
  AOI22_X1 U7019 ( .A1(n5961), .A2(n6110), .B1(n6214), .B2(n5923), .ZN(n5927)
         );
  INV_X1 U7020 ( .A(n5941), .ZN(n5925) );
  NOR2_X1 U7021 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5924), .ZN(n5933) );
  OAI21_X1 U7022 ( .B1(n5925), .B2(n5933), .A(REIP_REG_22__SCAN_IN), .ZN(n5926) );
  NAND4_X1 U7023 ( .A1(n5929), .A2(n5928), .A3(n5927), .A4(n5926), .ZN(U2805)
         );
  AOI22_X1 U7024 ( .A1(EBX_REG_21__SCAN_IN), .A2(n6209), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6148), .ZN(n5937) );
  OAI22_X1 U7025 ( .A1(n5930), .A2(n6222), .B1(n6726), .B2(n5941), .ZN(n5931)
         );
  INV_X1 U7026 ( .A(n5931), .ZN(n5936) );
  AOI22_X1 U7027 ( .A1(n5964), .A2(n6110), .B1(n6214), .B2(n5932), .ZN(n5935)
         );
  INV_X1 U7028 ( .A(n5933), .ZN(n5934) );
  NAND4_X1 U7029 ( .A1(n5937), .A2(n5936), .A3(n5935), .A4(n5934), .ZN(U2806)
         );
  AOI22_X1 U7030 ( .A1(EBX_REG_20__SCAN_IN), .A2(n6209), .B1(n5938), .B2(n6133), .ZN(n5945) );
  INV_X1 U7031 ( .A(n5939), .ZN(n5967) );
  AOI21_X1 U7032 ( .B1(REIP_REG_19__SCAN_IN), .B2(n5950), .A(
        REIP_REG_20__SCAN_IN), .ZN(n5942) );
  OAI22_X1 U7033 ( .A1(n5942), .A2(n5941), .B1(n5940), .B2(n6095), .ZN(n5943)
         );
  AOI21_X1 U7034 ( .B1(n5967), .B2(n6110), .A(n5943), .ZN(n5944) );
  OAI211_X1 U7035 ( .C1(n5946), .C2(n6212), .A(n5945), .B(n5944), .ZN(U2807)
         );
  INV_X1 U7036 ( .A(n5993), .ZN(n5949) );
  OAI21_X1 U7037 ( .B1(REIP_REG_18__SCAN_IN), .B2(n5947), .A(n6087), .ZN(n5948) );
  AOI22_X1 U7038 ( .A1(n5949), .A2(n6133), .B1(REIP_REG_19__SCAN_IN), .B2(
        n5948), .ZN(n5955) );
  AOI22_X1 U7039 ( .A1(EBX_REG_19__SCAN_IN), .A2(n6209), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6148), .ZN(n5954) );
  INV_X1 U7040 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6973) );
  AOI21_X1 U7041 ( .B1(n5950), .B2(n6973), .A(n6182), .ZN(n5953) );
  OAI22_X1 U7042 ( .A1(n5988), .A2(n6156), .B1(n6013), .B2(n6095), .ZN(n5951)
         );
  INV_X1 U7043 ( .A(n5951), .ZN(n5952) );
  NAND4_X1 U7044 ( .A1(n5955), .A2(n5954), .A3(n5953), .A4(n5952), .ZN(U2808)
         );
  AOI22_X1 U7045 ( .A1(n5977), .A2(n6239), .B1(n6238), .B2(DATAI_25_), .ZN(
        n5957) );
  AOI22_X1 U7046 ( .A1(n6242), .A2(DATAI_9_), .B1(n6241), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5956) );
  NAND2_X1 U7047 ( .A1(n5957), .A2(n5956), .ZN(U2866) );
  AOI22_X1 U7048 ( .A1(n5958), .A2(n6239), .B1(n6238), .B2(DATAI_23_), .ZN(
        n5960) );
  AOI22_X1 U7049 ( .A1(n6242), .A2(DATAI_7_), .B1(n6241), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5959) );
  NAND2_X1 U7050 ( .A1(n5960), .A2(n5959), .ZN(U2868) );
  AOI22_X1 U7051 ( .A1(n5961), .A2(n6239), .B1(n6238), .B2(DATAI_22_), .ZN(
        n5963) );
  AOI22_X1 U7052 ( .A1(n6242), .A2(DATAI_6_), .B1(n6241), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5962) );
  NAND2_X1 U7053 ( .A1(n5963), .A2(n5962), .ZN(U2869) );
  AOI22_X1 U7054 ( .A1(n5964), .A2(n6239), .B1(n6238), .B2(DATAI_21_), .ZN(
        n5966) );
  AOI22_X1 U7055 ( .A1(n6242), .A2(DATAI_5_), .B1(n6241), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5965) );
  NAND2_X1 U7056 ( .A1(n5966), .A2(n5965), .ZN(U2870) );
  AOI22_X1 U7057 ( .A1(n5967), .A2(n6239), .B1(n6238), .B2(DATAI_20_), .ZN(
        n5969) );
  AOI22_X1 U7058 ( .A1(n6242), .A2(DATAI_4_), .B1(n6241), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5968) );
  NAND2_X1 U7059 ( .A1(n5969), .A2(n5968), .ZN(U2871) );
  INV_X1 U7060 ( .A(n5988), .ZN(n5970) );
  AOI22_X1 U7061 ( .A1(n5970), .A2(n6239), .B1(n6238), .B2(DATAI_19_), .ZN(
        n5972) );
  AOI22_X1 U7062 ( .A1(n6242), .A2(DATAI_3_), .B1(n6241), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5971) );
  NAND2_X1 U7063 ( .A1(n5972), .A2(n5971), .ZN(U2872) );
  AOI22_X1 U7064 ( .A1(n6351), .A2(REIP_REG_25__SCAN_IN), .B1(n6350), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5979) );
  AOI21_X1 U7065 ( .B1(n5975), .B2(n5973), .A(n5974), .ZN(n5976) );
  INV_X1 U7066 ( .A(n5976), .ZN(n6007) );
  AOI22_X1 U7067 ( .A1(n5977), .A2(n6356), .B1(n6367), .B2(n6007), .ZN(n5978)
         );
  OAI211_X1 U7068 ( .C1(n6361), .C2(n5980), .A(n5979), .B(n5978), .ZN(U2961)
         );
  AOI22_X1 U7069 ( .A1(n6351), .A2(REIP_REG_19__SCAN_IN), .B1(n6350), .B2(
        PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5992) );
  INV_X1 U7070 ( .A(n5981), .ZN(n5982) );
  OR2_X1 U7071 ( .A1(n5983), .A2(n5982), .ZN(n5987) );
  INV_X1 U7072 ( .A(n5717), .ZN(n5985) );
  XNOR2_X1 U7073 ( .A(n4327), .B(n7085), .ZN(n5984) );
  NAND2_X1 U7074 ( .A1(n5985), .A2(n5984), .ZN(n5986) );
  NAND2_X1 U7075 ( .A1(n5987), .A2(n5986), .ZN(n6015) );
  OAI22_X1 U7076 ( .A1(n6015), .A2(n6068), .B1(n5989), .B2(n5988), .ZN(n5990)
         );
  INV_X1 U7077 ( .A(n5990), .ZN(n5991) );
  OAI211_X1 U7078 ( .C1(n6361), .C2(n5993), .A(n5992), .B(n5991), .ZN(U2967)
         );
  AOI22_X1 U7079 ( .A1(n6351), .A2(REIP_REG_17__SCAN_IN), .B1(n6350), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6004) );
  AOI21_X1 U7080 ( .B1(n3246), .B2(n6909), .A(n5994), .ZN(n5995) );
  AOI21_X1 U7081 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5996), .A(n5995), 
        .ZN(n6000) );
  INV_X1 U7082 ( .A(n5997), .ZN(n5999) );
  OAI21_X1 U7083 ( .B1(n6000), .B2(n5999), .A(n5998), .ZN(n6023) );
  OR2_X1 U7084 ( .A1(n5558), .A2(n6001), .ZN(n6002) );
  AND2_X1 U7085 ( .A1(n5534), .A2(n6002), .ZN(n6235) );
  AOI22_X1 U7086 ( .A1(n6023), .A2(n6367), .B1(n6356), .B2(n6235), .ZN(n6003)
         );
  OAI211_X1 U7087 ( .C1(n6361), .C2(n6092), .A(n6004), .B(n6003), .ZN(U2969)
         );
  AOI21_X1 U7088 ( .B1(n6351), .B2(REIP_REG_25__SCAN_IN), .A(n6005), .ZN(n6009) );
  AOI22_X1 U7089 ( .A1(n6007), .A2(n6415), .B1(n6389), .B2(n6006), .ZN(n6008)
         );
  OAI211_X1 U7090 ( .C1(n6011), .C2(n6010), .A(n6009), .B(n6008), .ZN(U2993)
         );
  AOI22_X1 U7091 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n6012), .B1(n6351), .B2(REIP_REG_19__SCAN_IN), .ZN(n6018) );
  OAI22_X1 U7092 ( .A1(n6015), .A2(n6014), .B1(n6013), .B2(n6413), .ZN(n6016)
         );
  INV_X1 U7093 ( .A(n6016), .ZN(n6017) );
  OAI211_X1 U7094 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n6019), .A(n6018), .B(n6017), .ZN(U2999) );
  NAND2_X1 U7095 ( .A1(n6021), .A2(n6020), .ZN(n6022) );
  AND2_X1 U7096 ( .A1(n5544), .A2(n6022), .ZN(n6223) );
  AOI22_X1 U7097 ( .A1(n6023), .A2(n6415), .B1(n6389), .B2(n6223), .ZN(n6028)
         );
  NOR2_X1 U7098 ( .A1(n6401), .A2(n7037), .ZN(n6024) );
  AOI221_X1 U7099 ( .B1(n6026), .B2(n6909), .C1(n6025), .C2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A(n6024), .ZN(n6027) );
  NAND2_X1 U7100 ( .A1(n6028), .A2(n6027), .ZN(U3001) );
  INV_X1 U7101 ( .A(n6029), .ZN(n6030) );
  AOI21_X1 U7102 ( .B1(n6389), .B2(n6031), .A(n6030), .ZN(n6036) );
  INV_X1 U7103 ( .A(n6032), .ZN(n6033) );
  AOI22_X1 U7104 ( .A1(n6034), .A2(n6415), .B1(n6033), .B2(n7094), .ZN(n6035)
         );
  OAI211_X1 U7105 ( .C1(n6037), .C2(n7094), .A(n6036), .B(n6035), .ZN(U3003)
         );
  AOI21_X1 U7106 ( .B1(n6040), .B2(n6039), .A(n6038), .ZN(n6048) );
  AOI21_X1 U7107 ( .B1(n6389), .B2(n6042), .A(n6041), .ZN(n6046) );
  AOI22_X1 U7108 ( .A1(n6044), .A2(n6415), .B1(n6043), .B2(n6047), .ZN(n6045)
         );
  OAI211_X1 U7109 ( .C1(n6048), .C2(n6047), .A(n6046), .B(n6045), .ZN(U3004)
         );
  INV_X1 U7110 ( .A(n6187), .ZN(n6051) );
  NAND3_X1 U7111 ( .A1(n6051), .A2(n6050), .A3(n6049), .ZN(n6052) );
  OAI22_X1 U7112 ( .A1(n6053), .A2(n6052), .B1(n4627), .B2(n6761), .ZN(U3455)
         );
  INV_X1 U7113 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6701) );
  INV_X1 U7114 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6683) );
  AOI21_X1 U7115 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6701), .A(n6683), .ZN(n6062) );
  INV_X1 U7116 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6054) );
  AOI21_X1 U7117 ( .B1(n6062), .B2(n6054), .A(n6788), .ZN(U2789) );
  INV_X1 U7118 ( .A(n6643), .ZN(n6055) );
  NAND2_X1 U7119 ( .A1(n6644), .A2(n6055), .ZN(n6057) );
  AND2_X1 U7120 ( .A1(n6645), .A2(n4522), .ZN(n6056) );
  AOI21_X1 U7121 ( .B1(n6057), .B2(n6641), .A(n6056), .ZN(n6067) );
  INV_X1 U7122 ( .A(n6067), .ZN(n6058) );
  OAI21_X1 U7123 ( .B1(n6058), .B2(n6660), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6059) );
  OAI21_X1 U7124 ( .B1(n6060), .B2(n6872), .A(n6059), .ZN(U2790) );
  INV_X2 U7125 ( .A(n6788), .ZN(n6789) );
  NOR2_X1 U7126 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n6063) );
  OAI21_X1 U7127 ( .B1(D_C_N_REG_SCAN_IN), .B2(n6063), .A(n6789), .ZN(n6061)
         );
  OAI21_X1 U7128 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6789), .A(n6061), .ZN(
        U2791) );
  NOR2_X1 U7129 ( .A1(n6788), .A2(n6062), .ZN(n6751) );
  OAI21_X1 U7130 ( .B1(BS16_N), .B2(n6063), .A(n6751), .ZN(n6749) );
  OAI21_X1 U7131 ( .B1(n6751), .B2(n6064), .A(n6749), .ZN(U2792) );
  NAND2_X1 U7132 ( .A1(n6065), .A2(n6689), .ZN(n6066) );
  NAND2_X1 U7133 ( .A1(n6066), .A2(n6778), .ZN(n6780) );
  AND2_X1 U7134 ( .A1(n6067), .A2(n6780), .ZN(n6650) );
  NOR2_X1 U7135 ( .A1(n6650), .A2(n6660), .ZN(n6775) );
  OAI21_X1 U7136 ( .B1(n6775), .B2(n6069), .A(n6068), .ZN(U2793) );
  NOR4_X1 U7137 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_21__SCAN_IN), .A4(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n6073) );
  NOR4_X1 U7138 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(
        DATAWIDTH_REG_15__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(
        DATAWIDTH_REG_17__SCAN_IN), .ZN(n6072) );
  NOR4_X1 U7139 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6071) );
  NOR4_X1 U7140 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n6070) );
  NAND4_X1 U7141 ( .A1(n6073), .A2(n6072), .A3(n6071), .A4(n6070), .ZN(n6079)
         );
  NOR4_X1 U7142 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(DATAWIDTH_REG_24__SCAN_IN), .A3(DATAWIDTH_REG_14__SCAN_IN), .A4(DATAWIDTH_REG_4__SCAN_IN), .ZN(n6077) );
  AOI211_X1 U7143 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_9__SCAN_IN), .B(
        DATAWIDTH_REG_13__SCAN_IN), .ZN(n6076) );
  NOR4_X1 U7144 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), 
        .A3(DATAWIDTH_REG_10__SCAN_IN), .A4(DATAWIDTH_REG_11__SCAN_IN), .ZN(
        n6075) );
  NOR4_X1 U7145 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(DATAWIDTH_REG_7__SCAN_IN), .A3(DATAWIDTH_REG_2__SCAN_IN), .A4(DATAWIDTH_REG_3__SCAN_IN), .ZN(n6074) );
  NAND4_X1 U7146 ( .A1(n6077), .A2(n6076), .A3(n6075), .A4(n6074), .ZN(n6078)
         );
  NOR2_X1 U7147 ( .A1(n6079), .A2(n6078), .ZN(n6770) );
  INV_X1 U7148 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6081) );
  NOR3_X1 U7149 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), 
        .A3(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6082) );
  OAI21_X1 U7150 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6082), .A(n6770), .ZN(n6080)
         );
  OAI21_X1 U7151 ( .B1(n6770), .B2(n6081), .A(n6080), .ZN(U2794) );
  INV_X1 U7152 ( .A(REIP_REG_1__SCAN_IN), .ZN(n7072) );
  INV_X1 U7153 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6750) );
  AOI21_X1 U7154 ( .B1(n7072), .B2(n6750), .A(n6082), .ZN(n6084) );
  INV_X1 U7155 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6083) );
  INV_X1 U7156 ( .A(n6770), .ZN(n6766) );
  AOI22_X1 U7157 ( .A1(n6770), .A2(n6084), .B1(n6083), .B2(n6766), .ZN(U2795)
         );
  NOR2_X1 U7158 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6085), .ZN(n6088) );
  INV_X1 U7159 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6086) );
  OAI22_X1 U7160 ( .A1(n6088), .A2(n6087), .B1(n6086), .B2(n6212), .ZN(n6089)
         );
  AOI211_X1 U7161 ( .C1(n6209), .C2(EBX_REG_17__SCAN_IN), .A(n6182), .B(n6089), 
        .ZN(n6091) );
  AOI22_X1 U7162 ( .A1(n6235), .A2(n6110), .B1(n6214), .B2(n6223), .ZN(n6090)
         );
  OAI211_X1 U7163 ( .C1(n6092), .C2(n6222), .A(n6091), .B(n6090), .ZN(U2810)
         );
  INV_X1 U7164 ( .A(n6093), .ZN(n6094) );
  OAI22_X1 U7165 ( .A1(n6150), .A2(n6939), .B1(n6095), .B2(n6094), .ZN(n6096)
         );
  AOI211_X1 U7166 ( .C1(n6148), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6182), 
        .B(n6096), .ZN(n6105) );
  INV_X1 U7167 ( .A(n6097), .ZN(n6098) );
  AOI22_X1 U7168 ( .A1(n6099), .A2(n6110), .B1(n6098), .B2(n6133), .ZN(n6104)
         );
  NOR3_X1 U7169 ( .A1(n6206), .A2(REIP_REG_12__SCAN_IN), .A3(n6100), .ZN(n6107) );
  OAI21_X1 U7170 ( .B1(n6107), .B2(n6108), .A(REIP_REG_13__SCAN_IN), .ZN(n6103) );
  NAND3_X1 U7171 ( .A1(n6171), .A2(n5366), .A3(n6101), .ZN(n6102) );
  NAND4_X1 U7172 ( .A1(n6105), .A2(n6104), .A3(n6103), .A4(n6102), .ZN(U2814)
         );
  AOI22_X1 U7173 ( .A1(n6214), .A2(n6226), .B1(n6148), .B2(
        PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n6113) );
  INV_X1 U7174 ( .A(EBX_REG_12__SCAN_IN), .ZN(n7051) );
  NOR2_X1 U7175 ( .A1(n7051), .A2(n6150), .ZN(n6106) );
  AOI211_X1 U7176 ( .C1(REIP_REG_12__SCAN_IN), .C2(n6108), .A(n6107), .B(n6106), .ZN(n6112) );
  AOI22_X1 U7177 ( .A1(n6229), .A2(n6110), .B1(n6109), .B2(n6133), .ZN(n6111)
         );
  NAND4_X1 U7178 ( .A1(n6113), .A2(n6112), .A3(n6111), .A4(n6163), .ZN(U2815)
         );
  INV_X1 U7179 ( .A(n6114), .ZN(n6115) );
  AOI22_X1 U7180 ( .A1(n6214), .A2(n6115), .B1(n6209), .B2(EBX_REG_10__SCAN_IN), .ZN(n6125) );
  NOR3_X1 U7181 ( .A1(n6206), .A2(REIP_REG_10__SCAN_IN), .A3(n6116), .ZN(n6117) );
  AOI211_X1 U7182 ( .C1(n6148), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6182), 
        .B(n6117), .ZN(n6124) );
  OAI22_X1 U7183 ( .A1(n6119), .A2(n6156), .B1(n6222), .B2(n6118), .ZN(n6120)
         );
  INV_X1 U7184 ( .A(n6120), .ZN(n6123) );
  NOR3_X1 U7185 ( .A1(n6206), .A2(REIP_REG_9__SCAN_IN), .A3(n6121), .ZN(n6126)
         );
  OAI21_X1 U7186 ( .B1(n6126), .B2(n6127), .A(REIP_REG_10__SCAN_IN), .ZN(n6122) );
  NAND4_X1 U7187 ( .A1(n6125), .A2(n6124), .A3(n6123), .A4(n6122), .ZN(U2817)
         );
  AOI21_X1 U7188 ( .B1(REIP_REG_9__SCAN_IN), .B2(n6127), .A(n6126), .ZN(n6136)
         );
  OAI21_X1 U7189 ( .B1(n6212), .B2(n6128), .A(n6163), .ZN(n6129) );
  AOI21_X1 U7190 ( .B1(n6214), .B2(n6381), .A(n6129), .ZN(n6130) );
  OAI21_X1 U7191 ( .B1(n6131), .B2(n6156), .A(n6130), .ZN(n6132) );
  AOI21_X1 U7192 ( .B1(n6134), .B2(n6133), .A(n6132), .ZN(n6135) );
  OAI211_X1 U7193 ( .C1(n6137), .C2(n6150), .A(n6136), .B(n6135), .ZN(U2818)
         );
  AOI21_X1 U7194 ( .B1(n6148), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n6182), 
        .ZN(n6147) );
  AOI22_X1 U7195 ( .A1(n6214), .A2(n6388), .B1(n6209), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n6146) );
  INV_X1 U7196 ( .A(n6139), .ZN(n6138) );
  OAI21_X1 U7197 ( .B1(n6206), .B2(n6138), .A(n6193), .ZN(n6172) );
  NOR3_X1 U7198 ( .A1(n6206), .A2(REIP_REG_6__SCAN_IN), .A3(n6139), .ZN(n6153)
         );
  OAI22_X1 U7199 ( .A1(n6141), .A2(n6156), .B1(n6140), .B2(n6222), .ZN(n6142)
         );
  AOI221_X1 U7200 ( .B1(n6172), .B2(REIP_REG_7__SCAN_IN), .C1(n6153), .C2(
        REIP_REG_7__SCAN_IN), .A(n6142), .ZN(n6145) );
  NAND3_X1 U7201 ( .A1(n6171), .A2(n6905), .A3(n6143), .ZN(n6144) );
  NAND4_X1 U7202 ( .A1(n6147), .A2(n6146), .A3(n6145), .A4(n6144), .ZN(U2820)
         );
  AOI22_X1 U7203 ( .A1(n6214), .A2(n6149), .B1(n6148), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6161) );
  NOR2_X1 U7204 ( .A1(n6151), .A2(n6150), .ZN(n6152) );
  AOI211_X1 U7205 ( .C1(n6172), .C2(REIP_REG_6__SCAN_IN), .A(n6153), .B(n6152), 
        .ZN(n6160) );
  INV_X1 U7206 ( .A(n6154), .ZN(n6155) );
  OAI22_X1 U7207 ( .A1(n6157), .A2(n6156), .B1(n6155), .B2(n6222), .ZN(n6158)
         );
  INV_X1 U7208 ( .A(n6158), .ZN(n6159) );
  NAND4_X1 U7209 ( .A1(n6161), .A2(n6160), .A3(n6159), .A4(n6163), .ZN(U2821)
         );
  INV_X1 U7210 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6165) );
  NAND2_X1 U7211 ( .A1(n6214), .A2(n6162), .ZN(n6164) );
  OAI211_X1 U7212 ( .C1(n6165), .C2(n6212), .A(n6164), .B(n6163), .ZN(n6169)
         );
  NOR2_X1 U7213 ( .A1(n6167), .A2(n6166), .ZN(n6168) );
  AOI211_X1 U7214 ( .C1(n6209), .C2(EBX_REG_5__SCAN_IN), .A(n6169), .B(n6168), 
        .ZN(n6175) );
  AND2_X1 U7215 ( .A1(n6171), .A2(n6170), .ZN(n6173) );
  OAI21_X1 U7216 ( .B1(n6173), .B2(REIP_REG_5__SCAN_IN), .A(n6172), .ZN(n6174)
         );
  OAI211_X1 U7217 ( .C1(n6222), .C2(n6176), .A(n6175), .B(n6174), .ZN(U2822)
         );
  INV_X1 U7218 ( .A(n6177), .ZN(n6192) );
  OAI21_X1 U7219 ( .B1(n6179), .B2(n6183), .A(n6178), .ZN(n6205) );
  OAI22_X1 U7220 ( .A1(n6180), .A2(n6212), .B1(n6706), .B2(n6205), .ZN(n6181)
         );
  AOI211_X1 U7221 ( .C1(n6209), .C2(EBX_REG_4__SCAN_IN), .A(n6182), .B(n6181), 
        .ZN(n6191) );
  NOR3_X1 U7222 ( .A1(n6206), .A2(REIP_REG_4__SCAN_IN), .A3(n6183), .ZN(n6184)
         );
  AOI21_X1 U7223 ( .B1(n6185), .B2(n6214), .A(n6184), .ZN(n6186) );
  OAI21_X1 U7224 ( .B1(n6187), .B2(n6217), .A(n6186), .ZN(n6188) );
  AOI21_X1 U7225 ( .B1(n6189), .B2(n6220), .A(n6188), .ZN(n6190) );
  OAI211_X1 U7226 ( .C1(n6192), .C2(n6222), .A(n6191), .B(n6190), .ZN(U2823)
         );
  OAI211_X1 U7227 ( .C1(n6206), .C2(REIP_REG_1__SCAN_IN), .A(
        REIP_REG_2__SCAN_IN), .B(n6193), .ZN(n6208) );
  INV_X1 U7228 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6195) );
  OAI22_X1 U7229 ( .A1(n6195), .A2(n6212), .B1(n6222), .B2(n6194), .ZN(n6196)
         );
  AOI21_X1 U7230 ( .B1(n6214), .B2(n6197), .A(n6196), .ZN(n6199) );
  NAND2_X1 U7231 ( .A1(n6209), .A2(EBX_REG_3__SCAN_IN), .ZN(n6198) );
  OAI211_X1 U7232 ( .C1(n6200), .C2(n6217), .A(n6199), .B(n6198), .ZN(n6201)
         );
  AOI21_X1 U7233 ( .B1(n6202), .B2(n6220), .A(n6201), .ZN(n6203) );
  OAI221_X1 U7234 ( .B1(n6205), .B2(n6204), .C1(n6205), .C2(n6208), .A(n6203), 
        .ZN(U2824) );
  INV_X1 U7235 ( .A(n4499), .ZN(n6218) );
  INV_X1 U7236 ( .A(n6398), .ZN(n6215) );
  INV_X1 U7237 ( .A(REIP_REG_2__SCAN_IN), .ZN(n7102) );
  OAI21_X1 U7238 ( .B1(n7072), .B2(n6206), .A(n7102), .ZN(n6207) );
  AOI22_X1 U7239 ( .A1(EBX_REG_2__SCAN_IN), .A2(n6209), .B1(n6208), .B2(n6207), 
        .ZN(n6210) );
  OAI21_X1 U7240 ( .B1(n6212), .B2(n6211), .A(n6210), .ZN(n6213) );
  AOI21_X1 U7241 ( .B1(n6215), .B2(n6214), .A(n6213), .ZN(n6216) );
  OAI21_X1 U7242 ( .B1(n6218), .B2(n6217), .A(n6216), .ZN(n6219) );
  AOI21_X1 U7243 ( .B1(n6357), .B2(n6220), .A(n6219), .ZN(n6221) );
  OAI21_X1 U7244 ( .B1(n6360), .B2(n6222), .A(n6221), .ZN(U2825) );
  AOI22_X1 U7245 ( .A1(n6235), .A2(n6228), .B1(n6227), .B2(n6223), .ZN(n6224)
         );
  OAI21_X1 U7246 ( .B1(n6225), .B2(n6231), .A(n6224), .ZN(U2842) );
  AOI22_X1 U7247 ( .A1(n6229), .A2(n6228), .B1(n6227), .B2(n6226), .ZN(n6230)
         );
  OAI21_X1 U7248 ( .B1(n7051), .B2(n6231), .A(n6230), .ZN(U2847) );
  AOI22_X1 U7249 ( .A1(n6232), .A2(n6239), .B1(n6238), .B2(DATAI_18_), .ZN(
        n6234) );
  AOI22_X1 U7250 ( .A1(n6242), .A2(DATAI_2_), .B1(n6241), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6233) );
  NAND2_X1 U7251 ( .A1(n6234), .A2(n6233), .ZN(U2873) );
  AOI22_X1 U7252 ( .A1(n6235), .A2(n6239), .B1(n6238), .B2(DATAI_17_), .ZN(
        n6237) );
  AOI22_X1 U7253 ( .A1(n6242), .A2(DATAI_1_), .B1(n6241), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U7254 ( .A1(n6237), .A2(n6236), .ZN(U2874) );
  AOI22_X1 U7255 ( .A1(n6240), .A2(n6239), .B1(n6238), .B2(DATAI_16_), .ZN(
        n6244) );
  AOI22_X1 U7256 ( .A1(n6242), .A2(DATAI_0_), .B1(n6241), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6243) );
  NAND2_X1 U7257 ( .A1(n6244), .A2(n6243), .ZN(U2875) );
  INV_X1 U7258 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6349) );
  AOI22_X1 U7259 ( .A1(n6779), .A2(LWORD_REG_15__SCAN_IN), .B1(n6262), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6246) );
  OAI21_X1 U7260 ( .B1(n6349), .B2(n6264), .A(n6246), .ZN(U2908) );
  INV_X1 U7261 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6344) );
  AOI22_X1 U7262 ( .A1(n6779), .A2(LWORD_REG_14__SCAN_IN), .B1(n6262), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6247) );
  OAI21_X1 U7263 ( .B1(n6344), .B2(n6264), .A(n6247), .ZN(U2909) );
  AOI22_X1 U7264 ( .A1(DATAO_REG_13__SCAN_IN), .A2(n6262), .B1(n6779), .B2(
        LWORD_REG_13__SCAN_IN), .ZN(n6248) );
  OAI21_X1 U7265 ( .B1(n7003), .B2(n6264), .A(n6248), .ZN(U2910) );
  AOI22_X1 U7266 ( .A1(LWORD_REG_12__SCAN_IN), .A2(n6779), .B1(n6262), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6249) );
  OAI21_X1 U7267 ( .B1(n5317), .B2(n6264), .A(n6249), .ZN(U2911) );
  INV_X1 U7268 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6875) );
  AOI22_X1 U7269 ( .A1(LWORD_REG_11__SCAN_IN), .A2(n6779), .B1(n6262), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6250) );
  OAI21_X1 U7270 ( .B1(n6875), .B2(n6264), .A(n6250), .ZN(U2912) );
  INV_X1 U7271 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6335) );
  AOI22_X1 U7272 ( .A1(n6779), .A2(LWORD_REG_10__SCAN_IN), .B1(n6260), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6251) );
  OAI21_X1 U7273 ( .B1(n6335), .B2(n6264), .A(n6251), .ZN(U2913) );
  INV_X1 U7274 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6332) );
  AOI22_X1 U7275 ( .A1(LWORD_REG_9__SCAN_IN), .A2(n6779), .B1(n6260), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6252) );
  OAI21_X1 U7276 ( .B1(n6332), .B2(n6264), .A(n6252), .ZN(U2914) );
  INV_X1 U7277 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6329) );
  AOI22_X1 U7278 ( .A1(n6779), .A2(LWORD_REG_8__SCAN_IN), .B1(n6260), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6253) );
  OAI21_X1 U7279 ( .B1(n6329), .B2(n6264), .A(n6253), .ZN(U2915) );
  AOI22_X1 U7280 ( .A1(n6779), .A2(LWORD_REG_7__SCAN_IN), .B1(n6260), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6254) );
  OAI21_X1 U7281 ( .B1(n3763), .B2(n6264), .A(n6254), .ZN(U2916) );
  AOI22_X1 U7282 ( .A1(LWORD_REG_6__SCAN_IN), .A2(n6779), .B1(
        DATAO_REG_6__SCAN_IN), .B2(n6260), .ZN(n6255) );
  OAI21_X1 U7283 ( .B1(n6324), .B2(n6264), .A(n6255), .ZN(U2917) );
  AOI22_X1 U7284 ( .A1(DATAO_REG_5__SCAN_IN), .A2(n6262), .B1(
        LWORD_REG_5__SCAN_IN), .B2(n6779), .ZN(n6256) );
  OAI21_X1 U7285 ( .B1(n6321), .B2(n6264), .A(n6256), .ZN(U2918) );
  INV_X1 U7286 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6318) );
  AOI22_X1 U7287 ( .A1(LWORD_REG_4__SCAN_IN), .A2(n6779), .B1(n6262), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6257) );
  OAI21_X1 U7288 ( .B1(n6318), .B2(n6264), .A(n6257), .ZN(U2919) );
  AOI22_X1 U7289 ( .A1(n6779), .A2(LWORD_REG_3__SCAN_IN), .B1(n6260), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6258) );
  OAI21_X1 U7290 ( .B1(n6315), .B2(n6264), .A(n6258), .ZN(U2920) );
  INV_X1 U7291 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6312) );
  AOI22_X1 U7292 ( .A1(LWORD_REG_2__SCAN_IN), .A2(n6779), .B1(n6262), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6259) );
  OAI21_X1 U7293 ( .B1(n6312), .B2(n6264), .A(n6259), .ZN(U2921) );
  AOI22_X1 U7294 ( .A1(LWORD_REG_1__SCAN_IN), .A2(n6779), .B1(
        DATAO_REG_1__SCAN_IN), .B2(n6260), .ZN(n6261) );
  OAI21_X1 U7295 ( .B1(n6309), .B2(n6264), .A(n6261), .ZN(U2922) );
  AOI22_X1 U7296 ( .A1(n6779), .A2(LWORD_REG_0__SCAN_IN), .B1(n6262), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6263) );
  OAI21_X1 U7297 ( .B1(n6949), .B2(n6264), .A(n6263), .ZN(U2923) );
  INV_X1 U7298 ( .A(READY_N), .ZN(n6778) );
  INV_X1 U7299 ( .A(n6265), .ZN(n6266) );
  INV_X1 U7300 ( .A(n6302), .ZN(n6345) );
  AND2_X1 U7301 ( .A1(n6345), .A2(DATAI_0_), .ZN(n6305) );
  AOI21_X1 U7302 ( .B1(UWORD_REG_0__SCAN_IN), .B2(n6346), .A(n6305), .ZN(n6267) );
  OAI21_X1 U7303 ( .B1(n7031), .B2(n6348), .A(n6267), .ZN(U2924) );
  AND2_X1 U7304 ( .A1(n6345), .A2(DATAI_1_), .ZN(n6307) );
  AOI21_X1 U7305 ( .B1(UWORD_REG_1__SCAN_IN), .B2(n6346), .A(n6307), .ZN(n6268) );
  OAI21_X1 U7306 ( .B1(n6269), .B2(n6348), .A(n6268), .ZN(U2925) );
  INV_X1 U7307 ( .A(DATAI_2_), .ZN(n6270) );
  NOR2_X1 U7308 ( .A1(n6302), .A2(n6270), .ZN(n6310) );
  AOI21_X1 U7309 ( .B1(UWORD_REG_2__SCAN_IN), .B2(n6283), .A(n6310), .ZN(n6271) );
  OAI21_X1 U7310 ( .B1(n6272), .B2(n6348), .A(n6271), .ZN(U2926) );
  AND2_X1 U7311 ( .A1(n6345), .A2(DATAI_3_), .ZN(n6313) );
  AOI21_X1 U7312 ( .B1(UWORD_REG_3__SCAN_IN), .B2(n6283), .A(n6313), .ZN(n6273) );
  OAI21_X1 U7313 ( .B1(n6274), .B2(n6348), .A(n6273), .ZN(U2927) );
  INV_X1 U7314 ( .A(DATAI_4_), .ZN(n6275) );
  NOR2_X1 U7315 ( .A1(n6302), .A2(n6275), .ZN(n6316) );
  AOI21_X1 U7316 ( .B1(UWORD_REG_4__SCAN_IN), .B2(n6283), .A(n6316), .ZN(n6276) );
  OAI21_X1 U7317 ( .B1(n7100), .B2(n6348), .A(n6276), .ZN(U2928) );
  AND2_X1 U7318 ( .A1(n6345), .A2(DATAI_5_), .ZN(n6319) );
  AOI21_X1 U7319 ( .B1(UWORD_REG_5__SCAN_IN), .B2(n6283), .A(n6319), .ZN(n6277) );
  OAI21_X1 U7320 ( .B1(n6950), .B2(n6348), .A(n6277), .ZN(U2929) );
  AND2_X1 U7321 ( .A1(n6345), .A2(DATAI_6_), .ZN(n6322) );
  AOI21_X1 U7322 ( .B1(UWORD_REG_6__SCAN_IN), .B2(n6283), .A(n6322), .ZN(n6278) );
  OAI21_X1 U7323 ( .B1(n6279), .B2(n6348), .A(n6278), .ZN(U2930) );
  AND2_X1 U7324 ( .A1(n6345), .A2(DATAI_7_), .ZN(n6325) );
  AOI21_X1 U7325 ( .B1(UWORD_REG_7__SCAN_IN), .B2(n6346), .A(n6325), .ZN(n6280) );
  OAI21_X1 U7326 ( .B1(n6281), .B2(n6348), .A(n6280), .ZN(U2931) );
  INV_X1 U7327 ( .A(DATAI_8_), .ZN(n6282) );
  NOR2_X1 U7328 ( .A1(n6302), .A2(n6282), .ZN(n6327) );
  AOI21_X1 U7329 ( .B1(UWORD_REG_8__SCAN_IN), .B2(n6283), .A(n6327), .ZN(n6284) );
  OAI21_X1 U7330 ( .B1(n6285), .B2(n6348), .A(n6284), .ZN(U2932) );
  INV_X1 U7331 ( .A(DATAI_9_), .ZN(n6286) );
  NOR2_X1 U7332 ( .A1(n6302), .A2(n6286), .ZN(n6330) );
  AOI21_X1 U7333 ( .B1(UWORD_REG_9__SCAN_IN), .B2(n6346), .A(n6330), .ZN(n6287) );
  OAI21_X1 U7334 ( .B1(n6288), .B2(n6348), .A(n6287), .ZN(U2933) );
  INV_X1 U7335 ( .A(DATAI_10_), .ZN(n6289) );
  NOR2_X1 U7336 ( .A1(n6302), .A2(n6289), .ZN(n6333) );
  AOI21_X1 U7337 ( .B1(UWORD_REG_10__SCAN_IN), .B2(n6346), .A(n6333), .ZN(
        n6290) );
  OAI21_X1 U7338 ( .B1(n6291), .B2(n6348), .A(n6290), .ZN(U2934) );
  INV_X1 U7339 ( .A(DATAI_11_), .ZN(n6292) );
  NOR2_X1 U7340 ( .A1(n6302), .A2(n6292), .ZN(n6336) );
  AOI21_X1 U7341 ( .B1(UWORD_REG_11__SCAN_IN), .B2(n6346), .A(n6336), .ZN(
        n6293) );
  OAI21_X1 U7342 ( .B1(n6294), .B2(n6348), .A(n6293), .ZN(U2935) );
  NOR2_X1 U7343 ( .A1(n6302), .A2(n6295), .ZN(n6338) );
  AOI21_X1 U7344 ( .B1(UWORD_REG_12__SCAN_IN), .B2(n6346), .A(n6338), .ZN(
        n6296) );
  OAI21_X1 U7345 ( .B1(n6297), .B2(n6348), .A(n6296), .ZN(U2936) );
  NOR2_X1 U7346 ( .A1(n6302), .A2(n6298), .ZN(n6340) );
  AOI21_X1 U7347 ( .B1(UWORD_REG_13__SCAN_IN), .B2(n6346), .A(n6340), .ZN(
        n6299) );
  OAI21_X1 U7348 ( .B1(n6300), .B2(n6348), .A(n6299), .ZN(U2937) );
  INV_X1 U7349 ( .A(DATAI_14_), .ZN(n6301) );
  NOR2_X1 U7350 ( .A1(n6302), .A2(n6301), .ZN(n6342) );
  AOI21_X1 U7351 ( .B1(UWORD_REG_14__SCAN_IN), .B2(n6346), .A(n6342), .ZN(
        n6303) );
  OAI21_X1 U7352 ( .B1(n6304), .B2(n6348), .A(n6303), .ZN(U2938) );
  AOI21_X1 U7353 ( .B1(LWORD_REG_0__SCAN_IN), .B2(n6346), .A(n6305), .ZN(n6306) );
  OAI21_X1 U7354 ( .B1(n6949), .B2(n6348), .A(n6306), .ZN(U2939) );
  AOI21_X1 U7355 ( .B1(LWORD_REG_1__SCAN_IN), .B2(n6346), .A(n6307), .ZN(n6308) );
  OAI21_X1 U7356 ( .B1(n6309), .B2(n6348), .A(n6308), .ZN(U2940) );
  AOI21_X1 U7357 ( .B1(LWORD_REG_2__SCAN_IN), .B2(n6346), .A(n6310), .ZN(n6311) );
  OAI21_X1 U7358 ( .B1(n6312), .B2(n6348), .A(n6311), .ZN(U2941) );
  AOI21_X1 U7359 ( .B1(LWORD_REG_3__SCAN_IN), .B2(n6346), .A(n6313), .ZN(n6314) );
  OAI21_X1 U7360 ( .B1(n6315), .B2(n6348), .A(n6314), .ZN(U2942) );
  AOI21_X1 U7361 ( .B1(LWORD_REG_4__SCAN_IN), .B2(n6346), .A(n6316), .ZN(n6317) );
  OAI21_X1 U7362 ( .B1(n6318), .B2(n6348), .A(n6317), .ZN(U2943) );
  AOI21_X1 U7363 ( .B1(LWORD_REG_5__SCAN_IN), .B2(n6346), .A(n6319), .ZN(n6320) );
  OAI21_X1 U7364 ( .B1(n6321), .B2(n6348), .A(n6320), .ZN(U2944) );
  AOI21_X1 U7365 ( .B1(LWORD_REG_6__SCAN_IN), .B2(n6346), .A(n6322), .ZN(n6323) );
  OAI21_X1 U7366 ( .B1(n6324), .B2(n6348), .A(n6323), .ZN(U2945) );
  AOI21_X1 U7367 ( .B1(LWORD_REG_7__SCAN_IN), .B2(n6346), .A(n6325), .ZN(n6326) );
  OAI21_X1 U7368 ( .B1(n3763), .B2(n6348), .A(n6326), .ZN(U2946) );
  AOI21_X1 U7369 ( .B1(LWORD_REG_8__SCAN_IN), .B2(n6346), .A(n6327), .ZN(n6328) );
  OAI21_X1 U7370 ( .B1(n6329), .B2(n6348), .A(n6328), .ZN(U2947) );
  AOI21_X1 U7371 ( .B1(LWORD_REG_9__SCAN_IN), .B2(n6346), .A(n6330), .ZN(n6331) );
  OAI21_X1 U7372 ( .B1(n6332), .B2(n6348), .A(n6331), .ZN(U2948) );
  AOI21_X1 U7373 ( .B1(LWORD_REG_10__SCAN_IN), .B2(n6346), .A(n6333), .ZN(
        n6334) );
  OAI21_X1 U7374 ( .B1(n6335), .B2(n6348), .A(n6334), .ZN(U2949) );
  AOI21_X1 U7375 ( .B1(LWORD_REG_11__SCAN_IN), .B2(n6346), .A(n6336), .ZN(
        n6337) );
  OAI21_X1 U7376 ( .B1(n6875), .B2(n6348), .A(n6337), .ZN(U2950) );
  AOI21_X1 U7377 ( .B1(LWORD_REG_12__SCAN_IN), .B2(n6346), .A(n6338), .ZN(
        n6339) );
  OAI21_X1 U7378 ( .B1(n5317), .B2(n6348), .A(n6339), .ZN(U2951) );
  AOI21_X1 U7379 ( .B1(LWORD_REG_13__SCAN_IN), .B2(n6346), .A(n6340), .ZN(
        n6341) );
  OAI21_X1 U7380 ( .B1(n7003), .B2(n6348), .A(n6341), .ZN(U2952) );
  AOI21_X1 U7381 ( .B1(LWORD_REG_14__SCAN_IN), .B2(n6346), .A(n6342), .ZN(
        n6343) );
  OAI21_X1 U7382 ( .B1(n6344), .B2(n6348), .A(n6343), .ZN(U2953) );
  AOI22_X1 U7383 ( .A1(n6346), .A2(LWORD_REG_15__SCAN_IN), .B1(n6345), .B2(
        DATAI_15_), .ZN(n6347) );
  OAI21_X1 U7384 ( .B1(n6349), .B2(n6348), .A(n6347), .ZN(U2954) );
  AOI22_X1 U7385 ( .A1(n6351), .A2(REIP_REG_2__SCAN_IN), .B1(n6350), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6359) );
  NAND2_X1 U7386 ( .A1(n6353), .A2(n6352), .ZN(n6354) );
  XOR2_X1 U7387 ( .A(n6355), .B(n6354), .Z(n6406) );
  AOI22_X1 U7388 ( .A1(n6406), .A2(n6367), .B1(n6357), .B2(n6356), .ZN(n6358)
         );
  OAI211_X1 U7389 ( .C1(n6361), .C2(n6360), .A(n6359), .B(n6358), .ZN(U2984)
         );
  OAI21_X1 U7390 ( .B1(n6362), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4260), 
        .ZN(n6363) );
  INV_X1 U7391 ( .A(n6363), .ZN(n6416) );
  NAND2_X1 U7392 ( .A1(n6365), .A2(n6364), .ZN(n6366) );
  AOI22_X1 U7393 ( .A1(n6416), .A2(n6367), .B1(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n6366), .ZN(n6369) );
  NAND2_X1 U7394 ( .A1(n6368), .A2(REIP_REG_0__SCAN_IN), .ZN(n6410) );
  OAI211_X1 U7395 ( .C1(n6371), .C2(n6370), .A(n6369), .B(n6410), .ZN(U2986)
         );
  AOI21_X1 U7396 ( .B1(n6389), .B2(n6373), .A(n6372), .ZN(n6377) );
  AOI22_X1 U7397 ( .A1(n6375), .A2(n6415), .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6374), .ZN(n6376) );
  OAI211_X1 U7398 ( .C1(INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n6378), .A(n6377), .B(n6376), .ZN(U3007) );
  INV_X1 U7399 ( .A(n6379), .ZN(n6380) );
  AOI21_X1 U7400 ( .B1(n6389), .B2(n6381), .A(n6380), .ZN(n6385) );
  AOI22_X1 U7401 ( .A1(n6383), .A2(n6415), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6382), .ZN(n6384) );
  OAI211_X1 U7402 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6386), .A(n6385), 
        .B(n6384), .ZN(U3009) );
  AOI21_X1 U7403 ( .B1(n6389), .B2(n6388), .A(n6387), .ZN(n6390) );
  OAI21_X1 U7404 ( .B1(n6391), .B2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n6390), 
        .ZN(n6392) );
  AOI21_X1 U7405 ( .B1(n6393), .B2(n6415), .A(n6392), .ZN(n6394) );
  OAI21_X1 U7406 ( .B1(n6396), .B2(n6395), .A(n6394), .ZN(U3011) );
  NAND2_X1 U7407 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6397), .ZN(n6409)
         );
  NOR2_X1 U7408 ( .A1(n6398), .A2(n6413), .ZN(n6405) );
  NAND3_X1 U7409 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A3(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6400) );
  AND2_X1 U7410 ( .A1(n6400), .A2(n6399), .ZN(n6402) );
  OAI22_X1 U7411 ( .A1(n6403), .A2(n6402), .B1(n7102), .B2(n6401), .ZN(n6404)
         );
  AOI211_X1 U7412 ( .C1(n6406), .C2(n6415), .A(n6405), .B(n6404), .ZN(n6407)
         );
  OAI221_X1 U7413 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6409), .C1(n4270), .C2(n6408), .A(n6407), .ZN(U3016) );
  OAI211_X1 U7414 ( .C1(n6413), .C2(n6412), .A(n6411), .B(n6410), .ZN(n6414)
         );
  AOI21_X1 U7415 ( .B1(n6416), .B2(n6415), .A(n6414), .ZN(n6417) );
  OAI221_X1 U7416 ( .B1(n6757), .B2(n6419), .C1(n6757), .C2(n6418), .A(n6417), 
        .ZN(U3018) );
  NOR2_X1 U7417 ( .A1(n6637), .A2(n6420), .ZN(U3019) );
  INV_X1 U7418 ( .A(n6421), .ZN(n6422) );
  INV_X1 U7419 ( .A(n6468), .ZN(n6427) );
  NAND3_X1 U7420 ( .A1(n6425), .A2(n6424), .A3(n7081), .ZN(n6426) );
  OAI21_X1 U7421 ( .B1(n6428), .B2(n6427), .A(n6426), .ZN(n6459) );
  NOR2_X1 U7422 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6473), .ZN(n6458)
         );
  AOI22_X1 U7423 ( .A1(n6498), .A2(n6459), .B1(n6562), .B2(n6458), .ZN(n6435)
         );
  OAI21_X1 U7424 ( .B1(n6461), .B2(n6491), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6431) );
  AOI211_X1 U7425 ( .C1(n6432), .C2(n6431), .A(n6430), .B(n6429), .ZN(n6433)
         );
  AOI22_X1 U7426 ( .A1(n6462), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6561), 
        .B2(n6461), .ZN(n6434) );
  OAI211_X1 U7427 ( .C1(n6436), .C2(n6465), .A(n6435), .B(n6434), .ZN(U3068)
         );
  AOI22_X1 U7428 ( .A1(n6437), .A2(n6459), .B1(n6574), .B2(n6458), .ZN(n6439)
         );
  AOI22_X1 U7429 ( .A1(n6462), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6573), 
        .B2(n6461), .ZN(n6438) );
  OAI211_X1 U7430 ( .C1(n6797), .C2(n6465), .A(n6439), .B(n6438), .ZN(U3069)
         );
  AOI22_X1 U7431 ( .A1(n6440), .A2(n6459), .B1(n6579), .B2(n6458), .ZN(n6442)
         );
  AOI22_X1 U7432 ( .A1(n6462), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6578), 
        .B2(n6461), .ZN(n6441) );
  OAI211_X1 U7433 ( .C1(n6443), .C2(n6465), .A(n6442), .B(n6441), .ZN(U3070)
         );
  AOI22_X1 U7434 ( .A1(n6444), .A2(n6459), .B1(n6585), .B2(n6458), .ZN(n6446)
         );
  AOI22_X1 U7435 ( .A1(n6462), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6584), 
        .B2(n6461), .ZN(n6445) );
  OAI211_X1 U7436 ( .C1(n6530), .C2(n6465), .A(n6446), .B(n6445), .ZN(U3071)
         );
  AOI22_X1 U7437 ( .A1(n6447), .A2(n6459), .B1(n6591), .B2(n6458), .ZN(n6449)
         );
  AOI22_X1 U7438 ( .A1(n6462), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6592), 
        .B2(n6461), .ZN(n6448) );
  OAI211_X1 U7439 ( .C1(n6450), .C2(n6465), .A(n6449), .B(n6448), .ZN(U3072)
         );
  AOI22_X1 U7440 ( .A1(n6503), .A2(n6459), .B1(n6597), .B2(n6458), .ZN(n6452)
         );
  AOI22_X1 U7441 ( .A1(n6462), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6461), 
        .B2(n6596), .ZN(n6451) );
  OAI211_X1 U7442 ( .C1(n6453), .C2(n6465), .A(n6452), .B(n6451), .ZN(U3073)
         );
  AOI22_X1 U7443 ( .A1(n6454), .A2(n6459), .B1(n6603), .B2(n6458), .ZN(n6456)
         );
  AOI22_X1 U7444 ( .A1(n6462), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6602), 
        .B2(n6461), .ZN(n6455) );
  OAI211_X1 U7445 ( .C1(n6457), .C2(n6465), .A(n6456), .B(n6455), .ZN(U3074)
         );
  AOI22_X1 U7446 ( .A1(n6460), .A2(n6459), .B1(n6611), .B2(n6458), .ZN(n6464)
         );
  AOI22_X1 U7447 ( .A1(n6462), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6613), 
        .B2(n6461), .ZN(n6463) );
  OAI211_X1 U7448 ( .C1(n6546), .C2(n6465), .A(n6464), .B(n6463), .ZN(U3075)
         );
  NOR2_X1 U7449 ( .A1(n6466), .A2(n6564), .ZN(n6475) );
  NAND3_X1 U7450 ( .A1(n6468), .A2(n6467), .A3(n3133), .ZN(n6469) );
  AND2_X1 U7451 ( .A1(n6469), .A2(n6472), .ZN(n6474) );
  INV_X1 U7452 ( .A(n6474), .ZN(n6470) );
  AOI22_X1 U7453 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6471), .B1(n6475), .B2(
        n6470), .ZN(n6497) );
  INV_X1 U7454 ( .A(n6472), .ZN(n6492) );
  AOI22_X1 U7455 ( .A1(n6562), .A2(n6492), .B1(n6561), .B2(n6491), .ZN(n6478)
         );
  AOI22_X1 U7456 ( .A1(n6475), .A2(n6474), .B1(n6473), .B2(n6564), .ZN(n6476)
         );
  NAND2_X1 U7457 ( .A1(n6568), .A2(n6476), .ZN(n6494) );
  AOI22_X1 U7458 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6494), .B1(n6569), 
        .B2(n6493), .ZN(n6477) );
  OAI211_X1 U7459 ( .C1(n6497), .C2(n6572), .A(n6478), .B(n6477), .ZN(U3076)
         );
  AOI22_X1 U7460 ( .A1(n6574), .A2(n6492), .B1(n6573), .B2(n6491), .ZN(n6480)
         );
  AOI22_X1 U7461 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6494), .B1(n6575), 
        .B2(n6493), .ZN(n6479) );
  OAI211_X1 U7462 ( .C1(n6497), .C2(n6798), .A(n6480), .B(n6479), .ZN(U3077)
         );
  AOI22_X1 U7463 ( .A1(n6579), .A2(n6492), .B1(n6580), .B2(n6493), .ZN(n6482)
         );
  AOI22_X1 U7464 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6494), .B1(n6578), 
        .B2(n6491), .ZN(n6481) );
  OAI211_X1 U7465 ( .C1(n6497), .C2(n6583), .A(n6482), .B(n6481), .ZN(U3078)
         );
  AOI22_X1 U7466 ( .A1(n6585), .A2(n6492), .B1(n6584), .B2(n6491), .ZN(n6484)
         );
  AOI22_X1 U7467 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6494), .B1(n6586), 
        .B2(n6493), .ZN(n6483) );
  OAI211_X1 U7468 ( .C1(n6497), .C2(n6589), .A(n6484), .B(n6483), .ZN(U3079)
         );
  AOI22_X1 U7469 ( .A1(n6591), .A2(n6492), .B1(n6590), .B2(n6493), .ZN(n6486)
         );
  AOI22_X1 U7470 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6494), .B1(n6592), 
        .B2(n6491), .ZN(n6485) );
  OAI211_X1 U7471 ( .C1(n6497), .C2(n6595), .A(n6486), .B(n6485), .ZN(U3080)
         );
  AOI22_X1 U7472 ( .A1(n6597), .A2(n6492), .B1(n6598), .B2(n6493), .ZN(n6488)
         );
  AOI22_X1 U7473 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6494), .B1(n6596), 
        .B2(n6491), .ZN(n6487) );
  OAI211_X1 U7474 ( .C1(n6497), .C2(n6601), .A(n6488), .B(n6487), .ZN(U3081)
         );
  AOI22_X1 U7475 ( .A1(n6603), .A2(n6492), .B1(n6604), .B2(n6493), .ZN(n6490)
         );
  AOI22_X1 U7476 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6494), .B1(n6602), 
        .B2(n6491), .ZN(n6489) );
  OAI211_X1 U7477 ( .C1(n6497), .C2(n6607), .A(n6490), .B(n6489), .ZN(U3082)
         );
  AOI22_X1 U7478 ( .A1(n6611), .A2(n6492), .B1(n6613), .B2(n6491), .ZN(n6496)
         );
  AOI22_X1 U7479 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6494), .B1(n6609), 
        .B2(n6493), .ZN(n6495) );
  OAI211_X1 U7480 ( .C1(n6497), .C2(n6617), .A(n6496), .B(n6495), .ZN(U3083)
         );
  INV_X1 U7481 ( .A(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n6884) );
  AOI22_X1 U7482 ( .A1(n6562), .A2(n6501), .B1(n6550), .B2(n6569), .ZN(n6500)
         );
  AOI22_X1 U7483 ( .A1(n6504), .A2(n6498), .B1(n6502), .B2(n6561), .ZN(n6499)
         );
  OAI211_X1 U7484 ( .C1(n6507), .C2(n6884), .A(n6500), .B(n6499), .ZN(U3100)
         );
  INV_X1 U7485 ( .A(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n7022) );
  AOI22_X1 U7486 ( .A1(n6597), .A2(n6501), .B1(n6550), .B2(n6598), .ZN(n6506)
         );
  AOI22_X1 U7487 ( .A1(n6504), .A2(n6503), .B1(n6502), .B2(n6596), .ZN(n6505)
         );
  OAI211_X1 U7488 ( .C1(n6507), .C2(n7022), .A(n6506), .B(n6505), .ZN(U3105)
         );
  AOI21_X1 U7489 ( .B1(n6509), .B2(n6508), .A(n6564), .ZN(n6517) );
  OR2_X1 U7490 ( .A1(n6511), .A2(n6510), .ZN(n6514) );
  NOR2_X1 U7491 ( .A1(n6512), .A2(n7081), .ZN(n6549) );
  INV_X1 U7492 ( .A(n6549), .ZN(n6513) );
  NAND2_X1 U7493 ( .A1(n6514), .A2(n6513), .ZN(n6515) );
  AOI22_X1 U7494 ( .A1(n6517), .A2(n6515), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6519), .ZN(n6554) );
  AOI22_X1 U7495 ( .A1(n6562), .A2(n6549), .B1(n6550), .B2(n6561), .ZN(n6522)
         );
  INV_X1 U7496 ( .A(n6515), .ZN(n6516) );
  NAND2_X1 U7497 ( .A1(n6517), .A2(n6516), .ZN(n6518) );
  OAI211_X1 U7498 ( .C1(n6520), .C2(n6519), .A(n6568), .B(n6518), .ZN(n6551)
         );
  AOI22_X1 U7499 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6551), .B1(n6569), 
        .B2(n6543), .ZN(n6521) );
  OAI211_X1 U7500 ( .C1(n6554), .C2(n6572), .A(n6522), .B(n6521), .ZN(U3108)
         );
  NOR2_X1 U7501 ( .A1(n6547), .A2(n6797), .ZN(n6523) );
  AOI21_X1 U7502 ( .B1(n6574), .B2(n6549), .A(n6523), .ZN(n6525) );
  AOI22_X1 U7503 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6551), .B1(n6573), 
        .B2(n6550), .ZN(n6524) );
  OAI211_X1 U7504 ( .C1(n6554), .C2(n6798), .A(n6525), .B(n6524), .ZN(U3109)
         );
  NOR2_X1 U7505 ( .A1(n6541), .A2(n6526), .ZN(n6527) );
  AOI21_X1 U7506 ( .B1(n6579), .B2(n6549), .A(n6527), .ZN(n6529) );
  AOI22_X1 U7507 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6551), .B1(n6580), 
        .B2(n6543), .ZN(n6528) );
  OAI211_X1 U7508 ( .C1(n6554), .C2(n6583), .A(n6529), .B(n6528), .ZN(U3110)
         );
  NOR2_X1 U7509 ( .A1(n6547), .A2(n6530), .ZN(n6531) );
  AOI21_X1 U7510 ( .B1(n6585), .B2(n6549), .A(n6531), .ZN(n6533) );
  AOI22_X1 U7511 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6551), .B1(n6584), 
        .B2(n6550), .ZN(n6532) );
  OAI211_X1 U7512 ( .C1(n6554), .C2(n6589), .A(n6533), .B(n6532), .ZN(U3111)
         );
  NOR2_X1 U7513 ( .A1(n6541), .A2(n6534), .ZN(n6535) );
  AOI21_X1 U7514 ( .B1(n6591), .B2(n6549), .A(n6535), .ZN(n6537) );
  AOI22_X1 U7515 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6551), .B1(n6590), 
        .B2(n6543), .ZN(n6536) );
  OAI211_X1 U7516 ( .C1(n6554), .C2(n6595), .A(n6537), .B(n6536), .ZN(U3112)
         );
  AOI22_X1 U7517 ( .A1(n6597), .A2(n6549), .B1(n6598), .B2(n6543), .ZN(n6539)
         );
  AOI22_X1 U7518 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6551), .B1(n6596), 
        .B2(n6550), .ZN(n6538) );
  OAI211_X1 U7519 ( .C1(n6554), .C2(n6601), .A(n6539), .B(n6538), .ZN(U3113)
         );
  NOR2_X1 U7520 ( .A1(n6541), .A2(n6540), .ZN(n6542) );
  AOI21_X1 U7521 ( .B1(n6603), .B2(n6549), .A(n6542), .ZN(n6545) );
  AOI22_X1 U7522 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6551), .B1(n6604), 
        .B2(n6543), .ZN(n6544) );
  OAI211_X1 U7523 ( .C1(n6554), .C2(n6607), .A(n6545), .B(n6544), .ZN(U3114)
         );
  NOR2_X1 U7524 ( .A1(n6547), .A2(n6546), .ZN(n6548) );
  AOI21_X1 U7525 ( .B1(n6611), .B2(n6549), .A(n6548), .ZN(n6553) );
  AOI22_X1 U7526 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6551), .B1(n6613), 
        .B2(n6550), .ZN(n6552) );
  OAI211_X1 U7527 ( .C1(n6554), .C2(n6617), .A(n6553), .B(n6552), .ZN(U3115)
         );
  NOR2_X1 U7528 ( .A1(n6555), .A2(n6564), .ZN(n6566) );
  NOR2_X1 U7529 ( .A1(n6556), .A2(n6563), .ZN(n6610) );
  AOI21_X1 U7530 ( .B1(n6558), .B2(n6557), .A(n6610), .ZN(n6565) );
  INV_X1 U7531 ( .A(n6565), .ZN(n6559) );
  AOI22_X1 U7532 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6560), .B1(n6566), .B2(
        n6559), .ZN(n6618) );
  AOI22_X1 U7533 ( .A1(n6562), .A2(n6610), .B1(n6561), .B2(n6612), .ZN(n6571)
         );
  AOI22_X1 U7534 ( .A1(n6566), .A2(n6565), .B1(n6564), .B2(n6563), .ZN(n6567)
         );
  NAND2_X1 U7535 ( .A1(n6568), .A2(n6567), .ZN(n6614) );
  AOI22_X1 U7536 ( .A1(n6614), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n6569), 
        .B2(n6608), .ZN(n6570) );
  OAI211_X1 U7537 ( .C1(n6618), .C2(n6572), .A(n6571), .B(n6570), .ZN(U3124)
         );
  AOI22_X1 U7538 ( .A1(n6574), .A2(n6610), .B1(n6573), .B2(n6612), .ZN(n6577)
         );
  AOI22_X1 U7539 ( .A1(n6614), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n6575), 
        .B2(n6608), .ZN(n6576) );
  OAI211_X1 U7540 ( .C1(n6618), .C2(n6798), .A(n6577), .B(n6576), .ZN(U3125)
         );
  AOI22_X1 U7541 ( .A1(n6579), .A2(n6610), .B1(n6578), .B2(n6612), .ZN(n6582)
         );
  AOI22_X1 U7542 ( .A1(n6614), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n6580), 
        .B2(n6608), .ZN(n6581) );
  OAI211_X1 U7543 ( .C1(n6618), .C2(n6583), .A(n6582), .B(n6581), .ZN(U3126)
         );
  AOI22_X1 U7544 ( .A1(n6585), .A2(n6610), .B1(n6584), .B2(n6612), .ZN(n6588)
         );
  AOI22_X1 U7545 ( .A1(n6614), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n6586), 
        .B2(n6608), .ZN(n6587) );
  OAI211_X1 U7546 ( .C1(n6618), .C2(n6589), .A(n6588), .B(n6587), .ZN(U3127)
         );
  AOI22_X1 U7547 ( .A1(n6591), .A2(n6610), .B1(n6590), .B2(n6608), .ZN(n6594)
         );
  AOI22_X1 U7548 ( .A1(n6614), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n6592), 
        .B2(n6612), .ZN(n6593) );
  OAI211_X1 U7549 ( .C1(n6618), .C2(n6595), .A(n6594), .B(n6593), .ZN(U3128)
         );
  AOI22_X1 U7550 ( .A1(n6597), .A2(n6610), .B1(n6596), .B2(n6612), .ZN(n6600)
         );
  AOI22_X1 U7551 ( .A1(n6614), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n6598), 
        .B2(n6608), .ZN(n6599) );
  OAI211_X1 U7552 ( .C1(n6618), .C2(n6601), .A(n6600), .B(n6599), .ZN(U3129)
         );
  AOI22_X1 U7553 ( .A1(n6603), .A2(n6610), .B1(n6602), .B2(n6612), .ZN(n6606)
         );
  AOI22_X1 U7554 ( .A1(n6614), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n6604), 
        .B2(n6608), .ZN(n6605) );
  OAI211_X1 U7555 ( .C1(n6618), .C2(n6607), .A(n6606), .B(n6605), .ZN(U3130)
         );
  AOI22_X1 U7556 ( .A1(n6611), .A2(n6610), .B1(n6609), .B2(n6608), .ZN(n6616)
         );
  AOI22_X1 U7557 ( .A1(n6614), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n6613), 
        .B2(n6612), .ZN(n6615) );
  OAI211_X1 U7558 ( .C1(n6618), .C2(n6617), .A(n6616), .B(n6615), .ZN(U3131)
         );
  INV_X1 U7559 ( .A(n6633), .ZN(n6636) );
  NOR2_X1 U7560 ( .A1(n6619), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6620)
         );
  AOI21_X1 U7561 ( .B1(n3133), .B2(n6621), .A(n6620), .ZN(n6759) );
  INV_X1 U7562 ( .A(n6622), .ZN(n6623) );
  NAND2_X1 U7563 ( .A1(n6623), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6764) );
  NAND3_X1 U7564 ( .A1(n6759), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6764), .ZN(n6626) );
  INV_X1 U7565 ( .A(n6626), .ZN(n6628) );
  OAI211_X1 U7566 ( .C1(n7064), .C2(n6626), .A(n6625), .B(n6624), .ZN(n6627)
         );
  OAI21_X1 U7567 ( .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n6628), .A(n6627), 
        .ZN(n6629) );
  AOI222_X1 U7568 ( .A1(n6631), .A2(n6630), .B1(n6631), .B2(n6629), .C1(n6630), 
        .C2(n6629), .ZN(n6635) );
  INV_X1 U7569 ( .A(n6635), .ZN(n6632) );
  OAI21_X1 U7570 ( .B1(n6633), .B2(n6632), .A(n7081), .ZN(n6634) );
  OAI21_X1 U7571 ( .B1(n6636), .B2(n6635), .A(n6634), .ZN(n6638) );
  NAND2_X1 U7572 ( .A1(n6638), .A2(n6637), .ZN(n6658) );
  NAND2_X1 U7573 ( .A1(n6640), .A2(n6639), .ZN(n6648) );
  NAND2_X1 U7574 ( .A1(n6642), .A2(n6641), .ZN(n6646) );
  AOI22_X1 U7575 ( .A1(n6646), .A2(n6645), .B1(n6644), .B2(n6643), .ZN(n6647)
         );
  AND2_X1 U7576 ( .A1(n6648), .A2(n6647), .ZN(n6774) );
  INV_X1 U7577 ( .A(n6649), .ZN(n6652) );
  OAI21_X1 U7578 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6650), 
        .ZN(n6651) );
  NAND3_X1 U7579 ( .A1(n6774), .A2(n6652), .A3(n6651), .ZN(n6653) );
  OR2_X1 U7580 ( .A1(n6654), .A2(n6653), .ZN(n6655) );
  NOR2_X1 U7581 ( .A1(n6656), .A2(n6655), .ZN(n6657) );
  NAND2_X1 U7582 ( .A1(n6658), .A2(n6657), .ZN(n6668) );
  NOR2_X1 U7583 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6778), .ZN(n6681) );
  OAI22_X1 U7584 ( .A1(n6668), .A2(n6660), .B1(n6778), .B2(n6659), .ZN(n6663)
         );
  OR3_X1 U7585 ( .A1(n4372), .A2(n6782), .A3(n6661), .ZN(n6662) );
  NOR2_X1 U7586 ( .A1(n6681), .A2(n6752), .ZN(n6666) );
  OAI21_X1 U7587 ( .B1(n6677), .B2(n6664), .A(n6872), .ZN(n6665) );
  OAI22_X1 U7588 ( .A1(n6872), .A2(n6666), .B1(n6752), .B2(n6665), .ZN(n6667)
         );
  AOI21_X1 U7589 ( .B1(n6672), .B2(n6668), .A(n6667), .ZN(n6670) );
  OAI211_X1 U7590 ( .C1(n6872), .C2(n6671), .A(n6670), .B(n6669), .ZN(U3148)
         );
  NOR2_X1 U7591 ( .A1(n6872), .A2(n6763), .ZN(n6673) );
  AOI21_X1 U7592 ( .B1(n6673), .B2(n6778), .A(n6672), .ZN(n6676) );
  NAND2_X1 U7593 ( .A1(n6872), .A2(n6937), .ZN(n6678) );
  OAI211_X1 U7594 ( .C1(n6752), .C2(n6681), .A(STATE2_REG_1__SCAN_IN), .B(
        n6678), .ZN(n6674) );
  OAI211_X1 U7595 ( .C1(n6752), .C2(n6676), .A(n6675), .B(n6674), .ZN(U3149)
         );
  NAND3_X1 U7596 ( .A1(n6678), .A2(n6677), .A3(n6753), .ZN(n6680) );
  OAI21_X1 U7597 ( .B1(n6681), .B2(n6680), .A(n6679), .ZN(U3150) );
  INV_X1 U7598 ( .A(n6751), .ZN(n6682) );
  AND2_X1 U7599 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6682), .ZN(U3151) );
  AND2_X1 U7600 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6682), .ZN(U3152) );
  AND2_X1 U7601 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6682), .ZN(U3153) );
  AND2_X1 U7602 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6682), .ZN(U3154) );
  AND2_X1 U7603 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6682), .ZN(U3155) );
  AND2_X1 U7604 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6682), .ZN(U3156) );
  AND2_X1 U7605 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6682), .ZN(U3157) );
  INV_X1 U7606 ( .A(DATAWIDTH_REG_24__SCAN_IN), .ZN(n6953) );
  NOR2_X1 U7607 ( .A1(n6751), .A2(n6953), .ZN(U3158) );
  AND2_X1 U7608 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6682), .ZN(U3159) );
  AND2_X1 U7609 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6682), .ZN(U3160) );
  AND2_X1 U7610 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6682), .ZN(U3161) );
  AND2_X1 U7611 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6682), .ZN(U3162) );
  AND2_X1 U7612 ( .A1(n6682), .A2(DATAWIDTH_REG_19__SCAN_IN), .ZN(U3163) );
  AND2_X1 U7613 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6682), .ZN(U3164) );
  AND2_X1 U7614 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6682), .ZN(U3165) );
  AND2_X1 U7615 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6682), .ZN(U3166) );
  AND2_X1 U7616 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6682), .ZN(U3167) );
  INV_X1 U7617 ( .A(DATAWIDTH_REG_14__SCAN_IN), .ZN(n6989) );
  NOR2_X1 U7618 ( .A1(n6751), .A2(n6989), .ZN(U3168) );
  AND2_X1 U7619 ( .A1(n6682), .A2(DATAWIDTH_REG_13__SCAN_IN), .ZN(U3169) );
  AND2_X1 U7620 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6682), .ZN(U3170) );
  AND2_X1 U7621 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6682), .ZN(U3171) );
  AND2_X1 U7622 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6682), .ZN(U3172) );
  AND2_X1 U7623 ( .A1(n6682), .A2(DATAWIDTH_REG_9__SCAN_IN), .ZN(U3173) );
  AND2_X1 U7624 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6682), .ZN(U3174) );
  INV_X1 U7625 ( .A(DATAWIDTH_REG_7__SCAN_IN), .ZN(n6965) );
  NOR2_X1 U7626 ( .A1(n6751), .A2(n6965), .ZN(U3175) );
  INV_X1 U7627 ( .A(DATAWIDTH_REG_6__SCAN_IN), .ZN(n6952) );
  NOR2_X1 U7628 ( .A1(n6751), .A2(n6952), .ZN(U3176) );
  AND2_X1 U7629 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6682), .ZN(U3177) );
  INV_X1 U7630 ( .A(DATAWIDTH_REG_4__SCAN_IN), .ZN(n7013) );
  NOR2_X1 U7631 ( .A1(n6751), .A2(n7013), .ZN(U3178) );
  AND2_X1 U7632 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6682), .ZN(U3179) );
  AND2_X1 U7633 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6682), .ZN(U3180) );
  NAND2_X1 U7634 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6687) );
  NAND2_X1 U7635 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6692) );
  INV_X1 U7636 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6903) );
  NOR2_X1 U7637 ( .A1(n6778), .A2(n6903), .ZN(n6697) );
  INV_X1 U7638 ( .A(n6697), .ZN(n6693) );
  NAND2_X1 U7639 ( .A1(n6692), .A2(n6693), .ZN(n6685) );
  OAI211_X1 U7640 ( .C1(n6701), .C2(NA_N), .A(n6683), .B(n6694), .ZN(n6684) );
  INV_X1 U7641 ( .A(n6684), .ZN(n6700) );
  AOI21_X1 U7642 ( .B1(n6694), .B2(n6685), .A(n6700), .ZN(n6686) );
  OAI221_X1 U7643 ( .B1(n6788), .B2(REQUESTPENDING_REG_SCAN_IN), .C1(n6788), 
        .C2(n6687), .A(n6686), .ZN(U3181) );
  INV_X1 U7644 ( .A(n6692), .ZN(n6691) );
  INV_X1 U7645 ( .A(n6687), .ZN(n6688) );
  AOI21_X1 U7646 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(STATE_REG_0__SCAN_IN), 
        .A(n6688), .ZN(n6690) );
  OAI211_X1 U7647 ( .C1(n6691), .C2(n6690), .A(n6689), .B(n6693), .ZN(U3182)
         );
  AOI221_X1 U7648 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6778), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6696) );
  OAI211_X1 U7649 ( .C1(n6694), .C2(n6693), .A(STATE_REG_0__SCAN_IN), .B(n6692), .ZN(n6695) );
  AOI21_X1 U7650 ( .B1(HOLD), .B2(n6696), .A(n6695), .ZN(n6699) );
  NAND3_X1 U7651 ( .A1(STATE_REG_0__SCAN_IN), .A2(REQUESTPENDING_REG_SCAN_IN), 
        .A3(n6697), .ZN(n6698) );
  OAI22_X1 U7652 ( .A1(n6700), .A2(n6699), .B1(NA_N), .B2(n6698), .ZN(U3183)
         );
  NOR2_X1 U7653 ( .A1(n6789), .A2(STATE_REG_2__SCAN_IN), .ZN(n6730) );
  NOR2_X2 U7654 ( .A1(n6701), .A2(n6789), .ZN(n6743) );
  AOI222_X1 U7655 ( .A1(n6730), .A2(REIP_REG_2__SCAN_IN), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6789), .C1(REIP_REG_1__SCAN_IN), .C2(
        n6743), .ZN(n6702) );
  INV_X1 U7656 ( .A(n6702), .ZN(U3184) );
  INV_X1 U7657 ( .A(n6743), .ZN(n6741) );
  CLKBUF_X1 U7658 ( .A(n6730), .Z(n6739) );
  AOI22_X1 U7659 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6739), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6789), .ZN(n6703) );
  OAI21_X1 U7660 ( .B1(n7102), .B2(n6741), .A(n6703), .ZN(U3185) );
  AOI222_X1 U7661 ( .A1(n6743), .A2(REIP_REG_3__SCAN_IN), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6789), .C1(REIP_REG_4__SCAN_IN), .C2(
        n6730), .ZN(n6704) );
  INV_X1 U7662 ( .A(n6704), .ZN(U3186) );
  AOI22_X1 U7663 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6730), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6789), .ZN(n6705) );
  OAI21_X1 U7664 ( .B1(n6706), .B2(n6741), .A(n6705), .ZN(U3187) );
  AOI22_X1 U7665 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6730), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6789), .ZN(n6707) );
  OAI21_X1 U7666 ( .B1(n4670), .B2(n6741), .A(n6707), .ZN(U3188) );
  AOI22_X1 U7667 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6739), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6789), .ZN(n6708) );
  OAI21_X1 U7668 ( .B1(n6999), .B2(n6741), .A(n6708), .ZN(U3189) );
  AOI22_X1 U7669 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6739), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6789), .ZN(n6709) );
  OAI21_X1 U7670 ( .B1(n6905), .B2(n6741), .A(n6709), .ZN(U3190) );
  AOI22_X1 U7671 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6730), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6789), .ZN(n6710) );
  OAI21_X1 U7672 ( .B1(n6711), .B2(n6741), .A(n6710), .ZN(U3191) );
  INV_X1 U7673 ( .A(n6730), .ZN(n6745) );
  AOI22_X1 U7674 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6743), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6789), .ZN(n6712) );
  OAI21_X1 U7675 ( .B1(n6713), .B2(n6745), .A(n6712), .ZN(U3192) );
  AOI22_X1 U7676 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6743), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6789), .ZN(n6714) );
  OAI21_X1 U7677 ( .B1(n5323), .B2(n6745), .A(n6714), .ZN(U3193) );
  AOI222_X1 U7678 ( .A1(n6743), .A2(REIP_REG_11__SCAN_IN), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6789), .C1(REIP_REG_12__SCAN_IN), .C2(
        n6739), .ZN(n6715) );
  INV_X1 U7679 ( .A(n6715), .ZN(U3194) );
  AOI222_X1 U7680 ( .A1(n6743), .A2(REIP_REG_12__SCAN_IN), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6789), .C1(REIP_REG_13__SCAN_IN), .C2(
        n6739), .ZN(n6716) );
  INV_X1 U7681 ( .A(n6716), .ZN(U3195) );
  AOI22_X1 U7682 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6730), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6789), .ZN(n6717) );
  OAI21_X1 U7683 ( .B1(n5366), .B2(n6741), .A(n6717), .ZN(U3196) );
  AOI22_X1 U7684 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6739), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6789), .ZN(n6718) );
  OAI21_X1 U7685 ( .B1(n6719), .B2(n6741), .A(n6718), .ZN(U3197) );
  INV_X1 U7686 ( .A(REIP_REG_16__SCAN_IN), .ZN(n7084) );
  AOI22_X1 U7687 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6743), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6789), .ZN(n6720) );
  OAI21_X1 U7688 ( .B1(n7084), .B2(n6745), .A(n6720), .ZN(U3198) );
  AOI222_X1 U7689 ( .A1(n6743), .A2(REIP_REG_16__SCAN_IN), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6789), .C1(REIP_REG_17__SCAN_IN), .C2(
        n6739), .ZN(n6721) );
  INV_X1 U7690 ( .A(n6721), .ZN(U3199) );
  AOI22_X1 U7691 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6739), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6789), .ZN(n6722) );
  OAI21_X1 U7692 ( .B1(n7037), .B2(n6741), .A(n6722), .ZN(U3200) );
  AOI222_X1 U7693 ( .A1(n6739), .A2(REIP_REG_19__SCAN_IN), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6789), .C1(REIP_REG_18__SCAN_IN), .C2(
        n6743), .ZN(n6723) );
  INV_X1 U7694 ( .A(n6723), .ZN(U3201) );
  AOI222_X1 U7695 ( .A1(n6743), .A2(REIP_REG_19__SCAN_IN), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6789), .C1(REIP_REG_20__SCAN_IN), .C2(
        n6739), .ZN(n6724) );
  INV_X1 U7696 ( .A(n6724), .ZN(U3202) );
  AOI22_X1 U7697 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6743), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6789), .ZN(n6725) );
  OAI21_X1 U7698 ( .B1(n6726), .B2(n6745), .A(n6725), .ZN(U3203) );
  AOI22_X1 U7699 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6743), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6789), .ZN(n6727) );
  OAI21_X1 U7700 ( .B1(n7063), .B2(n6745), .A(n6727), .ZN(U3204) );
  AOI22_X1 U7701 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6730), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6789), .ZN(n6728) );
  OAI21_X1 U7702 ( .B1(n7063), .B2(n6741), .A(n6728), .ZN(U3205) );
  AOI22_X1 U7703 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6743), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6789), .ZN(n6729) );
  OAI21_X1 U7704 ( .B1(n6732), .B2(n6745), .A(n6729), .ZN(U3206) );
  AOI22_X1 U7705 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6730), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6789), .ZN(n6731) );
  OAI21_X1 U7706 ( .B1(n6732), .B2(n6741), .A(n6731), .ZN(U3207) );
  AOI22_X1 U7707 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6743), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6789), .ZN(n6733) );
  OAI21_X1 U7708 ( .B1(n6734), .B2(n6745), .A(n6733), .ZN(U3208) );
  AOI22_X1 U7709 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6743), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6789), .ZN(n6735) );
  OAI21_X1 U7710 ( .B1(n6737), .B2(n6745), .A(n6735), .ZN(U3209) );
  AOI22_X1 U7711 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6739), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6789), .ZN(n6736) );
  OAI21_X1 U7712 ( .B1(n6737), .B2(n6741), .A(n6736), .ZN(U3210) );
  AOI22_X1 U7713 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6743), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6789), .ZN(n6738) );
  OAI21_X1 U7714 ( .B1(n6742), .B2(n6745), .A(n6738), .ZN(U3211) );
  AOI22_X1 U7715 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6739), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6789), .ZN(n6740) );
  OAI21_X1 U7716 ( .B1(n6742), .B2(n6741), .A(n6740), .ZN(U3212) );
  INV_X1 U7717 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6746) );
  AOI22_X1 U7718 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6743), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6789), .ZN(n6744) );
  OAI21_X1 U7719 ( .B1(n6746), .B2(n6745), .A(n6744), .ZN(U3213) );
  OAI22_X1 U7720 ( .A1(n6789), .A2(BYTEENABLE_REG_3__SCAN_IN), .B1(
        BE_N_REG_3__SCAN_IN), .B2(n6788), .ZN(n6747) );
  INV_X1 U7721 ( .A(n6747), .ZN(U3445) );
  MUX2_X1 U7722 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6789), .Z(U3446) );
  MUX2_X1 U7723 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6789), .Z(U3447) );
  MUX2_X1 U7724 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6789), .Z(U3448) );
  OAI21_X1 U7725 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6751), .A(n6749), .ZN(
        n6748) );
  INV_X1 U7726 ( .A(n6748), .ZN(U3451) );
  OAI21_X1 U7727 ( .B1(n6751), .B2(n6750), .A(n6749), .ZN(U3452) );
  INV_X1 U7728 ( .A(n6752), .ZN(n6755) );
  OAI211_X1 U7729 ( .C1(n3515), .C2(n6755), .A(n6754), .B(n6753), .ZN(U3453)
         );
  AOI21_X1 U7730 ( .B1(STATE2_REG_1__SCAN_IN), .B2(n6757), .A(n6756), .ZN(
        n6758) );
  OAI211_X1 U7731 ( .C1(n6759), .C2(n6763), .A(n6761), .B(n6758), .ZN(n6760)
         );
  OAI21_X1 U7732 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6761), .A(n6760), 
        .ZN(n6762) );
  OAI21_X1 U7733 ( .B1(n6764), .B2(n6763), .A(n6762), .ZN(U3461) );
  AOI21_X1 U7734 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6765) );
  AOI22_X1 U7735 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6765), .B2(n7072), .ZN(n6768) );
  INV_X1 U7736 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6767) );
  AOI22_X1 U7737 ( .A1(n6770), .A2(n6768), .B1(n6767), .B2(n6766), .ZN(U3468)
         );
  INV_X1 U7738 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n7067) );
  OAI21_X1 U7739 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6770), .ZN(n6769) );
  OAI21_X1 U7740 ( .B1(n6770), .B2(n7067), .A(n6769), .ZN(U3469) );
  NAND2_X1 U7741 ( .A1(n6789), .A2(W_R_N_REG_SCAN_IN), .ZN(n6771) );
  OAI21_X1 U7742 ( .B1(n6789), .B2(READREQUEST_REG_SCAN_IN), .A(n6771), .ZN(
        U3470) );
  INV_X1 U7743 ( .A(MORE_REG_SCAN_IN), .ZN(n6773) );
  INV_X1 U7744 ( .A(n6775), .ZN(n6772) );
  AOI22_X1 U7745 ( .A1(n6775), .A2(n6774), .B1(n6773), .B2(n6772), .ZN(U3471)
         );
  AOI211_X1 U7746 ( .C1(n6779), .C2(n6778), .A(n6777), .B(n6776), .ZN(n6787)
         );
  INV_X1 U7747 ( .A(n6780), .ZN(n6781) );
  OAI211_X1 U7748 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6782), .A(n6781), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6784) );
  AOI21_X1 U7749 ( .B1(n6784), .B2(STATE2_REG_0__SCAN_IN), .A(n6783), .ZN(
        n6786) );
  NAND2_X1 U7750 ( .A1(n6787), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6785) );
  OAI21_X1 U7751 ( .B1(n6787), .B2(n6786), .A(n6785), .ZN(U3472) );
  OAI22_X1 U7752 ( .A1(n6789), .A2(MEMORYFETCH_REG_SCAN_IN), .B1(
        M_IO_N_REG_SCAN_IN), .B2(n6788), .ZN(n6790) );
  INV_X1 U7753 ( .A(n6790), .ZN(U3473) );
  INV_X1 U7754 ( .A(n6791), .ZN(n6794) );
  OAI22_X1 U7755 ( .A1(n6795), .A2(n6794), .B1(n6793), .B2(n6792), .ZN(n6801)
         );
  OAI22_X1 U7756 ( .A1(n6799), .A2(n6798), .B1(n6797), .B2(n6796), .ZN(n6800)
         );
  AOI211_X1 U7757 ( .C1(INSTQUEUE_REG_3__1__SCAN_IN), .C2(n6802), .A(n6801), 
        .B(n6800), .ZN(n7120) );
  INV_X1 U7758 ( .A(keyinput60), .ZN(n6805) );
  NOR2_X1 U7759 ( .A1(keyinput20), .A2(keyinput80), .ZN(n6803) );
  NAND3_X1 U7760 ( .A1(keyinput8), .A2(keyinput111), .A3(n6803), .ZN(n6804) );
  NOR3_X1 U7761 ( .A1(keyinput104), .A2(n6805), .A3(n6804), .ZN(n6816) );
  NOR4_X1 U7762 ( .A1(keyinput55), .A2(keyinput24), .A3(keyinput127), .A4(
        keyinput115), .ZN(n6806) );
  NAND3_X1 U7763 ( .A1(keyinput105), .A2(keyinput53), .A3(n6806), .ZN(n6814)
         );
  NOR4_X1 U7764 ( .A1(keyinput84), .A2(keyinput74), .A3(keyinput90), .A4(
        keyinput109), .ZN(n6812) );
  NAND2_X1 U7765 ( .A1(keyinput33), .A2(keyinput26), .ZN(n6807) );
  NOR3_X1 U7766 ( .A1(keyinput97), .A2(keyinput43), .A3(n6807), .ZN(n6811) );
  NOR4_X1 U7767 ( .A1(keyinput16), .A2(keyinput85), .A3(keyinput99), .A4(
        keyinput44), .ZN(n6810) );
  NAND2_X1 U7768 ( .A1(keyinput92), .A2(keyinput124), .ZN(n6808) );
  NOR3_X1 U7769 ( .A1(keyinput36), .A2(keyinput114), .A3(n6808), .ZN(n6809) );
  NAND4_X1 U7770 ( .A1(n6812), .A2(n6811), .A3(n6810), .A4(n6809), .ZN(n6813)
         );
  NOR4_X1 U7771 ( .A1(keyinput76), .A2(keyinput32), .A3(n6814), .A4(n6813), 
        .ZN(n6815) );
  NAND4_X1 U7772 ( .A1(keyinput78), .A2(keyinput48), .A3(n6816), .A4(n6815), 
        .ZN(n6854) );
  NOR4_X1 U7773 ( .A1(keyinput102), .A2(keyinput37), .A3(keyinput41), .A4(
        keyinput56), .ZN(n6820) );
  NOR4_X1 U7774 ( .A1(keyinput66), .A2(keyinput119), .A3(keyinput126), .A4(
        keyinput98), .ZN(n6819) );
  NOR4_X1 U7775 ( .A1(keyinput17), .A2(keyinput100), .A3(keyinput108), .A4(
        keyinput120), .ZN(n6818) );
  NOR4_X1 U7776 ( .A1(keyinput61), .A2(keyinput64), .A3(keyinput4), .A4(
        keyinput13), .ZN(n6817) );
  NAND4_X1 U7777 ( .A1(n6820), .A2(n6819), .A3(n6818), .A4(n6817), .ZN(n6853)
         );
  NOR4_X1 U7778 ( .A1(keyinput22), .A2(keyinput30), .A3(keyinput58), .A4(
        keyinput7), .ZN(n6824) );
  NOR4_X1 U7779 ( .A1(keyinput0), .A2(keyinput39), .A3(keyinput46), .A4(
        keyinput19), .ZN(n6823) );
  NOR4_X1 U7780 ( .A1(keyinput83), .A2(keyinput87), .A3(keyinput94), .A4(
        keyinput71), .ZN(n6822) );
  NOR4_X1 U7781 ( .A1(keyinput6), .A2(keyinput11), .A3(keyinput10), .A4(
        keyinput14), .ZN(n6821) );
  NAND4_X1 U7782 ( .A1(n6824), .A2(n6823), .A3(n6822), .A4(n6821), .ZN(n6852)
         );
  NAND4_X1 U7783 ( .A1(keyinput91), .A2(keyinput59), .A3(keyinput1), .A4(
        keyinput9), .ZN(n6830) );
  NOR2_X1 U7784 ( .A1(keyinput77), .A2(keyinput21), .ZN(n6825) );
  NAND3_X1 U7785 ( .A1(keyinput117), .A2(keyinput79), .A3(n6825), .ZN(n6829)
         );
  NOR2_X1 U7786 ( .A1(keyinput63), .A2(keyinput50), .ZN(n6826) );
  NAND3_X1 U7787 ( .A1(keyinput81), .A2(keyinput45), .A3(n6826), .ZN(n6828) );
  OR4_X1 U7788 ( .A1(keyinput116), .A2(keyinput67), .A3(keyinput101), .A4(
        keyinput51), .ZN(n6827) );
  NOR4_X1 U7789 ( .A1(n6830), .A2(n6829), .A3(n6828), .A4(n6827), .ZN(n6850)
         );
  NOR2_X1 U7790 ( .A1(keyinput47), .A2(keyinput69), .ZN(n6831) );
  NAND3_X1 U7791 ( .A1(keyinput29), .A2(keyinput107), .A3(n6831), .ZN(n6837)
         );
  INV_X1 U7792 ( .A(keyinput103), .ZN(n6832) );
  NAND4_X1 U7793 ( .A1(keyinput57), .A2(keyinput40), .A3(keyinput25), .A4(
        n6832), .ZN(n6836) );
  NOR2_X1 U7794 ( .A1(keyinput110), .A2(keyinput95), .ZN(n6833) );
  NAND3_X1 U7795 ( .A1(keyinput106), .A2(keyinput75), .A3(n6833), .ZN(n6835)
         );
  NAND4_X1 U7796 ( .A1(keyinput18), .A2(keyinput122), .A3(keyinput118), .A4(
        keyinput112), .ZN(n6834) );
  NOR4_X1 U7797 ( .A1(n6837), .A2(n6836), .A3(n6835), .A4(n6834), .ZN(n6849)
         );
  NAND4_X1 U7798 ( .A1(keyinput121), .A2(keyinput113), .A3(keyinput89), .A4(
        keyinput96), .ZN(n6841) );
  NAND4_X1 U7799 ( .A1(keyinput88), .A2(keyinput73), .A3(keyinput68), .A4(
        keyinput65), .ZN(n6840) );
  NAND4_X1 U7800 ( .A1(keyinput52), .A2(keyinput86), .A3(keyinput82), .A4(
        keyinput123), .ZN(n6839) );
  NAND4_X1 U7801 ( .A1(keyinput28), .A2(keyinput12), .A3(keyinput5), .A4(
        keyinput49), .ZN(n6838) );
  NOR4_X1 U7802 ( .A1(n6841), .A2(n6840), .A3(n6839), .A4(n6838), .ZN(n6848)
         );
  NAND4_X1 U7803 ( .A1(keyinput70), .A2(keyinput35), .A3(keyinput42), .A4(
        keyinput34), .ZN(n6846) );
  NOR3_X1 U7804 ( .A1(keyinput125), .A2(keyinput93), .A3(keyinput72), .ZN(
        n6842) );
  NAND2_X1 U7805 ( .A1(keyinput38), .A2(n6842), .ZN(n6845) );
  NAND4_X1 U7806 ( .A1(keyinput54), .A2(keyinput15), .A3(keyinput3), .A4(
        keyinput2), .ZN(n6844) );
  NAND4_X1 U7807 ( .A1(keyinput27), .A2(keyinput23), .A3(keyinput31), .A4(
        keyinput62), .ZN(n6843) );
  NOR4_X1 U7808 ( .A1(n6846), .A2(n6845), .A3(n6844), .A4(n6843), .ZN(n6847)
         );
  NAND4_X1 U7809 ( .A1(n6850), .A2(n6849), .A3(n6848), .A4(n6847), .ZN(n6851)
         );
  NOR4_X1 U7810 ( .A1(n6854), .A2(n6853), .A3(n6852), .A4(n6851), .ZN(n7118)
         );
  INV_X1 U7811 ( .A(keyinput86), .ZN(n6856) );
  AOI22_X1 U7812 ( .A1(n4834), .A2(keyinput66), .B1(UWORD_REG_13__SCAN_IN), 
        .B2(n6856), .ZN(n6855) );
  OAI221_X1 U7813 ( .B1(n4834), .B2(keyinput66), .C1(n6856), .C2(
        UWORD_REG_13__SCAN_IN), .A(n6855), .ZN(n6866) );
  INV_X1 U7814 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n6859) );
  INV_X1 U7815 ( .A(keyinput6), .ZN(n6858) );
  AOI22_X1 U7816 ( .A1(n6859), .A2(keyinput71), .B1(DATAO_REG_5__SCAN_IN), 
        .B2(n6858), .ZN(n6857) );
  OAI221_X1 U7817 ( .B1(n6859), .B2(keyinput71), .C1(n6858), .C2(
        DATAO_REG_5__SCAN_IN), .A(n6857), .ZN(n6865) );
  XOR2_X1 U7818 ( .A(n4846), .B(keyinput4), .Z(n6863) );
  XNOR2_X1 U7819 ( .A(INSTQUEUE_REG_9__6__SCAN_IN), .B(keyinput7), .ZN(n6862)
         );
  XNOR2_X1 U7820 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .B(keyinput61), .ZN(
        n6861) );
  XNOR2_X1 U7821 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(keyinput27), .ZN(
        n6860) );
  NAND4_X1 U7822 ( .A1(n6863), .A2(n6862), .A3(n6861), .A4(n6860), .ZN(n6864)
         );
  NOR3_X1 U7823 ( .A1(n6866), .A2(n6865), .A3(n6864), .ZN(n6917) );
  INV_X1 U7824 ( .A(keyinput12), .ZN(n6868) );
  AOI22_X1 U7825 ( .A1(n6869), .A2(keyinput108), .B1(BYTEENABLE_REG_2__SCAN_IN), .B2(n6868), .ZN(n6867) );
  OAI221_X1 U7826 ( .B1(n6869), .B2(keyinput108), .C1(n6868), .C2(
        BYTEENABLE_REG_2__SCAN_IN), .A(n6867), .ZN(n6881) );
  INV_X1 U7827 ( .A(keyinput89), .ZN(n6871) );
  AOI22_X1 U7828 ( .A1(n6872), .A2(keyinput38), .B1(LWORD_REG_12__SCAN_IN), 
        .B2(n6871), .ZN(n6870) );
  OAI221_X1 U7829 ( .B1(n6872), .B2(keyinput38), .C1(n6871), .C2(
        LWORD_REG_12__SCAN_IN), .A(n6870), .ZN(n6880) );
  INV_X1 U7830 ( .A(keyinput87), .ZN(n6874) );
  AOI22_X1 U7831 ( .A1(n5323), .A2(keyinput93), .B1(ADDRESS_REG_10__SCAN_IN), 
        .B2(n6874), .ZN(n6873) );
  OAI221_X1 U7832 ( .B1(n5323), .B2(keyinput93), .C1(n6874), .C2(
        ADDRESS_REG_10__SCAN_IN), .A(n6873), .ZN(n6879) );
  XOR2_X1 U7833 ( .A(n6875), .B(keyinput35), .Z(n6877) );
  XNOR2_X1 U7834 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .B(keyinput64), .ZN(n6876)
         );
  NAND2_X1 U7835 ( .A1(n6877), .A2(n6876), .ZN(n6878) );
  NOR4_X1 U7836 ( .A1(n6881), .A2(n6880), .A3(n6879), .A4(n6878), .ZN(n6916)
         );
  INV_X1 U7837 ( .A(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n6883) );
  AOI22_X1 U7838 ( .A1(n6884), .A2(keyinput34), .B1(keyinput5), .B2(n6883), 
        .ZN(n6882) );
  OAI221_X1 U7839 ( .B1(n6884), .B2(keyinput34), .C1(n6883), .C2(keyinput5), 
        .A(n6882), .ZN(n6897) );
  INV_X1 U7840 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n6887) );
  INV_X1 U7841 ( .A(keyinput15), .ZN(n6886) );
  AOI22_X1 U7842 ( .A1(n6887), .A2(keyinput22), .B1(LWORD_REG_6__SCAN_IN), 
        .B2(n6886), .ZN(n6885) );
  OAI221_X1 U7843 ( .B1(n6887), .B2(keyinput22), .C1(n6886), .C2(
        LWORD_REG_6__SCAN_IN), .A(n6885), .ZN(n6896) );
  AOI22_X1 U7844 ( .A1(n6890), .A2(keyinput14), .B1(n6889), .B2(keyinput121), 
        .ZN(n6888) );
  OAI221_X1 U7845 ( .B1(n6890), .B2(keyinput14), .C1(n6889), .C2(keyinput121), 
        .A(n6888), .ZN(n6895) );
  INV_X1 U7846 ( .A(keyinput39), .ZN(n6892) );
  AOI22_X1 U7847 ( .A1(n6893), .A2(keyinput28), .B1(LWORD_REG_5__SCAN_IN), 
        .B2(n6892), .ZN(n6891) );
  OAI221_X1 U7848 ( .B1(n6893), .B2(keyinput28), .C1(n6892), .C2(
        LWORD_REG_5__SCAN_IN), .A(n6891), .ZN(n6894) );
  NOR4_X1 U7849 ( .A1(n6897), .A2(n6896), .A3(n6895), .A4(n6894), .ZN(n6915)
         );
  INV_X1 U7850 ( .A(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n6899) );
  AOI22_X1 U7851 ( .A1(n6900), .A2(keyinput125), .B1(n6899), .B2(keyinput123), 
        .ZN(n6898) );
  OAI221_X1 U7852 ( .B1(n6900), .B2(keyinput125), .C1(n6899), .C2(keyinput123), 
        .A(n6898), .ZN(n6913) );
  AOI22_X1 U7853 ( .A1(n6903), .A2(keyinput62), .B1(n6902), .B2(keyinput52), 
        .ZN(n6901) );
  OAI221_X1 U7854 ( .B1(n6903), .B2(keyinput62), .C1(n6902), .C2(keyinput52), 
        .A(n6901), .ZN(n6912) );
  AOI22_X1 U7855 ( .A1(n6906), .A2(keyinput120), .B1(keyinput72), .B2(n6905), 
        .ZN(n6904) );
  OAI221_X1 U7856 ( .B1(n6906), .B2(keyinput120), .C1(n6905), .C2(keyinput72), 
        .A(n6904), .ZN(n6911) );
  INV_X1 U7857 ( .A(keyinput11), .ZN(n6908) );
  AOI22_X1 U7858 ( .A1(n6909), .A2(keyinput3), .B1(UWORD_REG_8__SCAN_IN), .B2(
        n6908), .ZN(n6907) );
  OAI221_X1 U7859 ( .B1(n6909), .B2(keyinput3), .C1(n6908), .C2(
        UWORD_REG_8__SCAN_IN), .A(n6907), .ZN(n6910) );
  NOR4_X1 U7860 ( .A1(n6913), .A2(n6912), .A3(n6911), .A4(n6910), .ZN(n6914)
         );
  NAND4_X1 U7861 ( .A1(n6917), .A2(n6916), .A3(n6915), .A4(n6914), .ZN(n7117)
         );
  INV_X1 U7862 ( .A(keyinput88), .ZN(n6919) );
  AOI22_X1 U7863 ( .A1(n4691), .A2(keyinput68), .B1(LWORD_REG_1__SCAN_IN), 
        .B2(n6919), .ZN(n6918) );
  OAI221_X1 U7864 ( .B1(n4691), .B2(keyinput68), .C1(n6919), .C2(
        LWORD_REG_1__SCAN_IN), .A(n6918), .ZN(n6931) );
  INV_X1 U7865 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n6921) );
  AOI22_X1 U7866 ( .A1(n6921), .A2(keyinput10), .B1(keyinput102), .B2(n4598), 
        .ZN(n6920) );
  OAI221_X1 U7867 ( .B1(n6921), .B2(keyinput10), .C1(n4598), .C2(keyinput102), 
        .A(n6920), .ZN(n6930) );
  AOI22_X1 U7868 ( .A1(n6924), .A2(keyinput41), .B1(keyinput23), .B2(n6923), 
        .ZN(n6922) );
  OAI221_X1 U7869 ( .B1(n6924), .B2(keyinput41), .C1(n6923), .C2(keyinput23), 
        .A(n6922), .ZN(n6929) );
  XOR2_X1 U7870 ( .A(n3434), .B(keyinput73), .Z(n6927) );
  XNOR2_X1 U7871 ( .A(n6925), .B(keyinput37), .ZN(n6926) );
  NAND2_X1 U7872 ( .A1(n6927), .A2(n6926), .ZN(n6928) );
  NOR4_X1 U7873 ( .A1(n6931), .A2(n6930), .A3(n6929), .A4(n6928), .ZN(n7115)
         );
  INV_X1 U7874 ( .A(keyinput70), .ZN(n6933) );
  INV_X1 U7875 ( .A(keyinput56), .ZN(n6936) );
  OAI22_X1 U7876 ( .A1(n6937), .A2(keyinput100), .B1(n6936), .B2(
        DATAWIDTH_REG_0__SCAN_IN), .ZN(n6935) );
  AOI221_X1 U7877 ( .B1(n6937), .B2(keyinput100), .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(n6936), .A(n6935), .ZN(n6946) );
  INV_X1 U7878 ( .A(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n6940) );
  OAI22_X1 U7879 ( .A1(n6940), .A2(keyinput30), .B1(n6939), .B2(keyinput49), 
        .ZN(n6938) );
  AOI221_X1 U7880 ( .B1(n6940), .B2(keyinput30), .C1(keyinput49), .C2(n6939), 
        .A(n6938), .ZN(n6945) );
  INV_X1 U7881 ( .A(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n6943) );
  INV_X1 U7882 ( .A(keyinput0), .ZN(n6942) );
  OAI22_X1 U7883 ( .A1(n6943), .A2(keyinput113), .B1(n6942), .B2(
        ADDRESS_REG_18__SCAN_IN), .ZN(n6941) );
  AOI221_X1 U7884 ( .B1(n6943), .B2(keyinput113), .C1(ADDRESS_REG_18__SCAN_IN), 
        .C2(n6942), .A(n6941), .ZN(n6944) );
  NAND4_X1 U7885 ( .A1(n6947), .A2(n6946), .A3(n6945), .A4(n6944), .ZN(n6982)
         );
  AOI22_X1 U7886 ( .A1(n6950), .A2(keyinput19), .B1(n6949), .B2(keyinput98), 
        .ZN(n6948) );
  OAI221_X1 U7887 ( .B1(n6950), .B2(keyinput19), .C1(n6949), .C2(keyinput98), 
        .A(n6948), .ZN(n6981) );
  OAI22_X1 U7888 ( .A1(keyinput94), .A2(n6953), .B1(n6952), .B2(keyinput31), 
        .ZN(n6951) );
  AOI221_X1 U7889 ( .B1(n6953), .B2(keyinput94), .C1(n6952), .C2(keyinput31), 
        .A(n6951), .ZN(n6962) );
  INV_X1 U7890 ( .A(keyinput13), .ZN(n6955) );
  OAI22_X1 U7891 ( .A1(n6956), .A2(keyinput54), .B1(n6955), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6954) );
  AOI221_X1 U7892 ( .B1(n6956), .B2(keyinput54), .C1(DATAO_REG_6__SCAN_IN), 
        .C2(n6955), .A(n6954), .ZN(n6961) );
  INV_X1 U7893 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n6959) );
  INV_X1 U7894 ( .A(keyinput83), .ZN(n6958) );
  OAI22_X1 U7895 ( .A1(n6959), .A2(keyinput42), .B1(n6958), .B2(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n6957) );
  AOI221_X1 U7896 ( .B1(n6959), .B2(keyinput42), .C1(DATAWIDTH_REG_19__SCAN_IN), .C2(n6958), .A(n6957), .ZN(n6960) );
  NAND3_X1 U7897 ( .A1(n6962), .A2(n6961), .A3(n6960), .ZN(n6980) );
  INV_X1 U7898 ( .A(keyinput126), .ZN(n6964) );
  OAI22_X1 U7899 ( .A1(keyinput58), .A2(n6965), .B1(n6964), .B2(
        M_IO_N_REG_SCAN_IN), .ZN(n6963) );
  AOI221_X1 U7900 ( .B1(n6965), .B2(keyinput58), .C1(n6964), .C2(
        M_IO_N_REG_SCAN_IN), .A(n6963), .ZN(n6978) );
  INV_X1 U7901 ( .A(keyinput82), .ZN(n6967) );
  OAI22_X1 U7902 ( .A1(n6968), .A2(keyinput17), .B1(n6967), .B2(HOLD), .ZN(
        n6966) );
  AOI221_X1 U7903 ( .B1(n6968), .B2(keyinput17), .C1(HOLD), .C2(n6967), .A(
        n6966), .ZN(n6977) );
  INV_X1 U7904 ( .A(keyinput46), .ZN(n6971) );
  INV_X1 U7905 ( .A(keyinput65), .ZN(n6970) );
  OAI22_X1 U7906 ( .A1(n6971), .A2(ADDRESS_REG_23__SCAN_IN), .B1(n6970), .B2(
        READREQUEST_REG_SCAN_IN), .ZN(n6969) );
  AOI221_X1 U7907 ( .B1(n6971), .B2(ADDRESS_REG_23__SCAN_IN), .C1(
        READREQUEST_REG_SCAN_IN), .C2(n6970), .A(n6969), .ZN(n6976) );
  INV_X1 U7908 ( .A(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n6974) );
  OAI22_X1 U7909 ( .A1(n6974), .A2(keyinput2), .B1(n6973), .B2(keyinput96), 
        .ZN(n6972) );
  AOI221_X1 U7910 ( .B1(n6974), .B2(keyinput2), .C1(keyinput96), .C2(n6973), 
        .A(n6972), .ZN(n6975) );
  NAND4_X1 U7911 ( .A1(n6978), .A2(n6977), .A3(n6976), .A4(n6975), .ZN(n6979)
         );
  NOR4_X1 U7912 ( .A1(n6982), .A2(n6981), .A3(n6980), .A4(n6979), .ZN(n7114)
         );
  INV_X1 U7913 ( .A(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n6984) );
  OAI22_X1 U7914 ( .A1(n3435), .A2(keyinput106), .B1(n6984), .B2(keyinput95), 
        .ZN(n6983) );
  AOI221_X1 U7915 ( .B1(n3435), .B2(keyinput106), .C1(keyinput95), .C2(n6984), 
        .A(n6983), .ZN(n6996) );
  INV_X1 U7916 ( .A(keyinput122), .ZN(n6986) );
  OAI22_X1 U7917 ( .A1(n4907), .A2(keyinput18), .B1(n6986), .B2(
        ADDRESS_REG_15__SCAN_IN), .ZN(n6985) );
  AOI221_X1 U7918 ( .B1(n4907), .B2(keyinput18), .C1(ADDRESS_REG_15__SCAN_IN), 
        .C2(n6986), .A(n6985), .ZN(n6995) );
  INV_X1 U7919 ( .A(keyinput112), .ZN(n6988) );
  OAI22_X1 U7920 ( .A1(keyinput75), .A2(n6989), .B1(n6988), .B2(
        ADDRESS_REG_14__SCAN_IN), .ZN(n6987) );
  AOI221_X1 U7921 ( .B1(n6989), .B2(keyinput75), .C1(n6988), .C2(
        ADDRESS_REG_14__SCAN_IN), .A(n6987), .ZN(n6994) );
  INV_X1 U7922 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n6992) );
  OAI22_X1 U7923 ( .A1(n6992), .A2(keyinput110), .B1(n6991), .B2(keyinput118), 
        .ZN(n6990) );
  AOI221_X1 U7924 ( .B1(n6992), .B2(keyinput110), .C1(keyinput118), .C2(n6991), 
        .A(n6990), .ZN(n6993) );
  NAND4_X1 U7925 ( .A1(n6996), .A2(n6995), .A3(n6994), .A4(n6993), .ZN(n7045)
         );
  INV_X1 U7926 ( .A(keyinput40), .ZN(n6998) );
  OAI22_X1 U7927 ( .A1(n6999), .A2(keyinput25), .B1(n6998), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n6997) );
  AOI221_X1 U7928 ( .B1(n6999), .B2(keyinput25), .C1(LWORD_REG_9__SCAN_IN), 
        .C2(n6998), .A(n6997), .ZN(n7010) );
  OAI22_X1 U7929 ( .A1(n4842), .A2(keyinput103), .B1(n7001), .B2(keyinput57), 
        .ZN(n7000) );
  AOI221_X1 U7930 ( .B1(n4842), .B2(keyinput103), .C1(keyinput57), .C2(n7001), 
        .A(n7000), .ZN(n7009) );
  OAI22_X1 U7931 ( .A1(n4695), .A2(keyinput107), .B1(n7003), .B2(keyinput69), 
        .ZN(n7002) );
  AOI221_X1 U7932 ( .B1(n4695), .B2(keyinput107), .C1(keyinput69), .C2(n7003), 
        .A(n7002), .ZN(n7008) );
  INV_X1 U7933 ( .A(keyinput47), .ZN(n7005) );
  OAI22_X1 U7934 ( .A1(n7006), .A2(keyinput29), .B1(n7005), .B2(
        DATAWIDTH_REG_9__SCAN_IN), .ZN(n7004) );
  AOI221_X1 U7935 ( .B1(n7006), .B2(keyinput29), .C1(DATAWIDTH_REG_9__SCAN_IN), 
        .C2(n7005), .A(n7004), .ZN(n7007) );
  NAND4_X1 U7936 ( .A1(n7010), .A2(n7009), .A3(n7008), .A4(n7007), .ZN(n7044)
         );
  INV_X1 U7937 ( .A(keyinput51), .ZN(n7012) );
  OAI22_X1 U7938 ( .A1(keyinput101), .A2(n7013), .B1(n7012), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n7011) );
  AOI221_X1 U7939 ( .B1(n7013), .B2(keyinput101), .C1(n7012), .C2(
        LWORD_REG_11__SCAN_IN), .A(n7011), .ZN(n7026) );
  INV_X1 U7940 ( .A(keyinput67), .ZN(n7015) );
  OAI22_X1 U7941 ( .A1(n7016), .A2(keyinput116), .B1(n7015), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n7014) );
  AOI221_X1 U7942 ( .B1(n7016), .B2(keyinput116), .C1(UWORD_REG_9__SCAN_IN), 
        .C2(n7015), .A(n7014), .ZN(n7025) );
  INV_X1 U7943 ( .A(LWORD_REG_4__SCAN_IN), .ZN(n7019) );
  INV_X1 U7944 ( .A(keyinput50), .ZN(n7018) );
  OAI22_X1 U7945 ( .A1(keyinput45), .A2(n7019), .B1(n7018), .B2(BS16_N), .ZN(
        n7017) );
  AOI221_X1 U7946 ( .B1(n7019), .B2(keyinput45), .C1(n7018), .C2(BS16_N), .A(
        n7017), .ZN(n7024) );
  OAI22_X1 U7947 ( .A1(n7022), .A2(keyinput81), .B1(n7021), .B2(keyinput63), 
        .ZN(n7020) );
  AOI221_X1 U7948 ( .B1(n7022), .B2(keyinput81), .C1(keyinput63), .C2(n7021), 
        .A(n7020), .ZN(n7023) );
  NAND4_X1 U7949 ( .A1(n7026), .A2(n7025), .A3(n7024), .A4(n7023), .ZN(n7043)
         );
  INV_X1 U7950 ( .A(keyinput21), .ZN(n7028) );
  OAI22_X1 U7951 ( .A1(n7029), .A2(keyinput59), .B1(n7028), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n7027) );
  AOI221_X1 U7952 ( .B1(n7029), .B2(keyinput59), .C1(DATAO_REG_1__SCAN_IN), 
        .C2(n7028), .A(n7027), .ZN(n7041) );
  OAI22_X1 U7953 ( .A1(n7032), .A2(keyinput117), .B1(n7031), .B2(keyinput91), 
        .ZN(n7030) );
  AOI221_X1 U7954 ( .B1(n7032), .B2(keyinput117), .C1(keyinput91), .C2(n7031), 
        .A(n7030), .ZN(n7040) );
  INV_X1 U7955 ( .A(REIP_REG_20__SCAN_IN), .ZN(n7035) );
  INV_X1 U7956 ( .A(keyinput9), .ZN(n7034) );
  OAI22_X1 U7957 ( .A1(n7035), .A2(keyinput1), .B1(n7034), .B2(
        UWORD_REG_3__SCAN_IN), .ZN(n7033) );
  AOI221_X1 U7958 ( .B1(n7035), .B2(keyinput1), .C1(UWORD_REG_3__SCAN_IN), 
        .C2(n7034), .A(n7033), .ZN(n7039) );
  OAI22_X1 U7959 ( .A1(n5667), .A2(keyinput77), .B1(n7037), .B2(keyinput79), 
        .ZN(n7036) );
  AOI221_X1 U7960 ( .B1(n5667), .B2(keyinput77), .C1(keyinput79), .C2(n7037), 
        .A(n7036), .ZN(n7038) );
  NAND4_X1 U7961 ( .A1(n7041), .A2(n7040), .A3(n7039), .A4(n7038), .ZN(n7042)
         );
  NOR4_X1 U7962 ( .A1(n7045), .A2(n7044), .A3(n7043), .A4(n7042), .ZN(n7113)
         );
  INV_X1 U7963 ( .A(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n7048) );
  INV_X1 U7964 ( .A(keyinput85), .ZN(n7047) );
  OAI22_X1 U7965 ( .A1(n7048), .A2(keyinput16), .B1(n7047), .B2(
        ADDRESS_REG_0__SCAN_IN), .ZN(n7046) );
  AOI221_X1 U7966 ( .B1(n7048), .B2(keyinput16), .C1(ADDRESS_REG_0__SCAN_IN), 
        .C2(n7047), .A(n7046), .ZN(n7061) );
  INV_X1 U7967 ( .A(keyinput124), .ZN(n7050) );
  OAI22_X1 U7968 ( .A1(n7051), .A2(keyinput36), .B1(n7050), .B2(
        UWORD_REG_0__SCAN_IN), .ZN(n7049) );
  AOI221_X1 U7969 ( .B1(n7051), .B2(keyinput36), .C1(UWORD_REG_0__SCAN_IN), 
        .C2(n7050), .A(n7049), .ZN(n7060) );
  INV_X1 U7970 ( .A(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n7054) );
  INV_X1 U7971 ( .A(keyinput92), .ZN(n7053) );
  OAI22_X1 U7972 ( .A1(n7054), .A2(keyinput44), .B1(n7053), .B2(
        ADDRESS_REG_2__SCAN_IN), .ZN(n7052) );
  AOI221_X1 U7973 ( .B1(n7054), .B2(keyinput44), .C1(ADDRESS_REG_2__SCAN_IN), 
        .C2(n7053), .A(n7052), .ZN(n7059) );
  INV_X1 U7974 ( .A(keyinput114), .ZN(n7056) );
  OAI22_X1 U7975 ( .A1(n7057), .A2(keyinput99), .B1(n7056), .B2(
        FLUSH_REG_SCAN_IN), .ZN(n7055) );
  AOI221_X1 U7976 ( .B1(n7057), .B2(keyinput99), .C1(FLUSH_REG_SCAN_IN), .C2(
        n7056), .A(n7055), .ZN(n7058) );
  NAND4_X1 U7977 ( .A1(n7061), .A2(n7060), .A3(n7059), .A4(n7058), .ZN(n7111)
         );
  OAI22_X1 U7978 ( .A1(n7064), .A2(keyinput43), .B1(n7063), .B2(keyinput74), 
        .ZN(n7062) );
  AOI221_X1 U7979 ( .B1(n7064), .B2(keyinput43), .C1(keyinput74), .C2(n7063), 
        .A(n7062), .ZN(n7076) );
  INV_X1 U7980 ( .A(keyinput84), .ZN(n7066) );
  OAI22_X1 U7981 ( .A1(keyinput26), .A2(n7067), .B1(n7066), .B2(
        LWORD_REG_2__SCAN_IN), .ZN(n7065) );
  AOI221_X1 U7982 ( .B1(n7067), .B2(keyinput26), .C1(n7066), .C2(
        LWORD_REG_2__SCAN_IN), .A(n7065), .ZN(n7075) );
  INV_X1 U7983 ( .A(keyinput33), .ZN(n7069) );
  OAI22_X1 U7984 ( .A1(n5626), .A2(keyinput109), .B1(n7069), .B2(
        ADDRESS_REG_17__SCAN_IN), .ZN(n7068) );
  AOI221_X1 U7985 ( .B1(n5626), .B2(keyinput109), .C1(ADDRESS_REG_17__SCAN_IN), 
        .C2(n7069), .A(n7068), .ZN(n7074) );
  INV_X1 U7986 ( .A(keyinput97), .ZN(n7071) );
  OAI22_X1 U7987 ( .A1(n7072), .A2(keyinput90), .B1(n7071), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n7070) );
  AOI221_X1 U7988 ( .B1(n7072), .B2(keyinput90), .C1(DATAO_REG_13__SCAN_IN), 
        .C2(n7071), .A(n7070), .ZN(n7073) );
  NAND4_X1 U7989 ( .A1(n7076), .A2(n7075), .A3(n7074), .A4(n7073), .ZN(n7110)
         );
  OAI22_X1 U7990 ( .A1(n4770), .A2(keyinput20), .B1(n7078), .B2(keyinput8), 
        .ZN(n7077) );
  AOI221_X1 U7991 ( .B1(n4770), .B2(keyinput20), .C1(keyinput8), .C2(n7078), 
        .A(n7077), .ZN(n7091) );
  INV_X1 U7992 ( .A(keyinput111), .ZN(n7080) );
  OAI22_X1 U7993 ( .A1(n7081), .A2(keyinput80), .B1(n7080), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n7079) );
  AOI221_X1 U7994 ( .B1(n7081), .B2(keyinput80), .C1(DATAO_REG_17__SCAN_IN), 
        .C2(n7080), .A(n7079), .ZN(n7090) );
  INV_X1 U7995 ( .A(keyinput78), .ZN(n7083) );
  OAI22_X1 U7996 ( .A1(n7084), .A2(keyinput48), .B1(n7083), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n7082) );
  AOI221_X1 U7997 ( .B1(n7084), .B2(keyinput48), .C1(UWORD_REG_12__SCAN_IN), 
        .C2(n7083), .A(n7082), .ZN(n7089) );
  XNOR2_X1 U7998 ( .A(n7085), .B(keyinput60), .ZN(n7087) );
  XNOR2_X1 U7999 ( .A(n3166), .B(keyinput104), .ZN(n7086) );
  NOR2_X1 U8000 ( .A1(n7087), .A2(n7086), .ZN(n7088) );
  NAND4_X1 U8001 ( .A1(n7091), .A2(n7090), .A3(n7089), .A4(n7088), .ZN(n7109)
         );
  INV_X1 U8002 ( .A(keyinput53), .ZN(n7093) );
  OAI22_X1 U8003 ( .A1(n7094), .A2(keyinput32), .B1(n7093), .B2(NA_N), .ZN(
        n7092) );
  AOI221_X1 U8004 ( .B1(n7094), .B2(keyinput32), .C1(NA_N), .C2(n7093), .A(
        n7092), .ZN(n7107) );
  INV_X1 U8005 ( .A(keyinput105), .ZN(n7096) );
  OAI22_X1 U8006 ( .A1(n7097), .A2(keyinput76), .B1(n7096), .B2(
        DATAWIDTH_REG_13__SCAN_IN), .ZN(n7095) );
  AOI221_X1 U8007 ( .B1(n7097), .B2(keyinput76), .C1(DATAWIDTH_REG_13__SCAN_IN), .C2(n7096), .A(n7095), .ZN(n7106) );
  INV_X1 U8008 ( .A(keyinput115), .ZN(n7099) );
  OAI22_X1 U8009 ( .A1(n7100), .A2(keyinput127), .B1(n7099), .B2(
        BE_N_REG_3__SCAN_IN), .ZN(n7098) );
  AOI221_X1 U8010 ( .B1(n7100), .B2(keyinput127), .C1(BE_N_REG_3__SCAN_IN), 
        .C2(n7099), .A(n7098), .ZN(n7105) );
  OAI22_X1 U8011 ( .A1(n7103), .A2(keyinput55), .B1(n7102), .B2(keyinput24), 
        .ZN(n7101) );
  AOI221_X1 U8012 ( .B1(n7103), .B2(keyinput55), .C1(keyinput24), .C2(n7102), 
        .A(n7101), .ZN(n7104) );
  NAND4_X1 U8013 ( .A1(n7107), .A2(n7106), .A3(n7105), .A4(n7104), .ZN(n7108)
         );
  NOR4_X1 U8014 ( .A1(n7111), .A2(n7110), .A3(n7109), .A4(n7108), .ZN(n7112)
         );
  NAND4_X1 U8015 ( .A1(n7115), .A2(n7114), .A3(n7113), .A4(n7112), .ZN(n7116)
         );
  NOR3_X1 U8016 ( .A1(n7118), .A2(n7117), .A3(n7116), .ZN(n7119) );
  XNOR2_X1 U8017 ( .A(n7120), .B(n7119), .ZN(U3045) );
  CLKBUF_X1 U3608 ( .A(n6260), .Z(n6262) );
  AND2_X1 U3635 ( .A1(n3654), .A2(n3915), .ZN(n7121) );
endmodule

