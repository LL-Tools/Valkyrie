

module b17_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_,
         DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
         DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
         DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
         DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
         DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1,
         READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
         n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
         n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
         n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
         n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
         n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
         n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
         n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588,
         n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
         n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,
         n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
         n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620,
         n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,
         n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636,
         n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,
         n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
         n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660,
         n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
         n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676,
         n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684,
         n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,
         n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700,
         n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708,
         n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,
         n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
         n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732,
         n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,
         n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748,
         n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756,
         n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764,
         n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772,
         n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780,
         n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788,
         n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796,
         n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804,
         n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812,
         n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820,
         n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828,
         n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836,
         n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844,
         n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852,
         n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860,
         n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868,
         n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876,
         n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884,
         n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892,
         n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900,
         n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908,
         n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916,
         n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924,
         n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932,
         n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940,
         n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948,
         n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956,
         n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964,
         n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972,
         n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980,
         n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988,
         n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996,
         n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004,
         n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012,
         n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020,
         n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028,
         n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036,
         n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044,
         n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052,
         n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060,
         n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068,
         n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076,
         n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084,
         n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092,
         n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100,
         n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108,
         n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116,
         n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124,
         n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132,
         n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140,
         n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148,
         n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156,
         n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164,
         n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172,
         n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180,
         n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188,
         n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196,
         n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204,
         n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212,
         n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220,
         n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228,
         n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236,
         n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244,
         n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252,
         n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260,
         n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268,
         n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276,
         n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284,
         n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,
         n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300,
         n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308,
         n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316,
         n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324,
         n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332,
         n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340,
         n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348,
         n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356,
         n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364,
         n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372,
         n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380,
         n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388,
         n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396,
         n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404,
         n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412,
         n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420,
         n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428,
         n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436,
         n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444,
         n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452,
         n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460,
         n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468,
         n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476,
         n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484,
         n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492,
         n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500,
         n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508,
         n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516,
         n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524,
         n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532,
         n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540,
         n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548,
         n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556,
         n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564,
         n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572,
         n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580,
         n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588,
         n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596,
         n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604,
         n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612,
         n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620,
         n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628,
         n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636,
         n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644,
         n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652,
         n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660,
         n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668,
         n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676,
         n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684,
         n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692,
         n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700,
         n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708,
         n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716,
         n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724,
         n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732,
         n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740,
         n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748,
         n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756,
         n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764,
         n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772,
         n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780,
         n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788,
         n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796,
         n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804,
         n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812,
         n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820,
         n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828,
         n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836,
         n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844,
         n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852,
         n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860,
         n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868,
         n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876,
         n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884,
         n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892,
         n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900,
         n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908,
         n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916,
         n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924,
         n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932,
         n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940,
         n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948,
         n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956,
         n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964,
         n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972,
         n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980,
         n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988,
         n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996,
         n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004,
         n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012,
         n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020,
         n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028,
         n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036,
         n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044,
         n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052,
         n17053, n17055, n17056, n17057, n17058, n17059, n17060, n17061,
         n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069,
         n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077,
         n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085,
         n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093,
         n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101,
         n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109,
         n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117,
         n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125,
         n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133,
         n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141,
         n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149,
         n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157,
         n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165,
         n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173,
         n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181,
         n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189,
         n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197,
         n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205,
         n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213,
         n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221,
         n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229,
         n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237,
         n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245,
         n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253,
         n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261,
         n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269,
         n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277,
         n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285,
         n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293,
         n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301,
         n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309,
         n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317,
         n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325,
         n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333,
         n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341,
         n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349,
         n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357,
         n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365,
         n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373,
         n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381,
         n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389,
         n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397,
         n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405,
         n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413,
         n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421,
         n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429,
         n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437,
         n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445,
         n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453,
         n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461,
         n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469,
         n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
         n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485,
         n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493,
         n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501,
         n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509,
         n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517,
         n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525,
         n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533,
         n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541,
         n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549,
         n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557,
         n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565,
         n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573,
         n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581,
         n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589,
         n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597,
         n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605,
         n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613,
         n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
         n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629,
         n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637,
         n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645,
         n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653,
         n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661,
         n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669,
         n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677,
         n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685,
         n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693,
         n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701,
         n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709,
         n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717,
         n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725,
         n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733,
         n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741,
         n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749,
         n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757,
         n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765,
         n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773,
         n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781,
         n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789,
         n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797,
         n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805,
         n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813,
         n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821,
         n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829,
         n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837,
         n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845,
         n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853,
         n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861,
         n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869,
         n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877,
         n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885,
         n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893,
         n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901,
         n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909,
         n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917,
         n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925,
         n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933,
         n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941,
         n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949,
         n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957,
         n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965,
         n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973,
         n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981,
         n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989,
         n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997,
         n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005,
         n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013,
         n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021,
         n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029,
         n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037,
         n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045,
         n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053,
         n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061,
         n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069,
         n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077,
         n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085,
         n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093,
         n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101,
         n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109,
         n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117,
         n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125,
         n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133,
         n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141,
         n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149,
         n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157,
         n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165,
         n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173,
         n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181,
         n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189,
         n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197,
         n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205,
         n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213,
         n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221,
         n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229,
         n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237,
         n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245,
         n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253,
         n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261,
         n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269,
         n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277,
         n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285,
         n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293,
         n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301,
         n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309,
         n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317,
         n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325,
         n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333,
         n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341,
         n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349,
         n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357,
         n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365,
         n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373,
         n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381,
         n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389,
         n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397,
         n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405,
         n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413,
         n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421,
         n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429,
         n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437,
         n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445,
         n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453,
         n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461,
         n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469,
         n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477,
         n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485,
         n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493,
         n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501,
         n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509,
         n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517,
         n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525,
         n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533,
         n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541,
         n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549,
         n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557,
         n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565,
         n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573,
         n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581,
         n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589,
         n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597,
         n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605,
         n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613,
         n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621,
         n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629,
         n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637,
         n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645,
         n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653,
         n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661,
         n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669,
         n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677,
         n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685,
         n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693,
         n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701,
         n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709,
         n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717,
         n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725,
         n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733,
         n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741,
         n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749,
         n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757,
         n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765,
         n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773,
         n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781,
         n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789,
         n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797,
         n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805,
         n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813,
         n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821,
         n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829,
         n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837,
         n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845,
         n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853,
         n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861,
         n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869,
         n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877,
         n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885,
         n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893,
         n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901,
         n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909,
         n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917,
         n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925,
         n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933,
         n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941,
         n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949,
         n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957,
         n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965,
         n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973,
         n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981,
         n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989,
         n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997,
         n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005,
         n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013,
         n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021,
         n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029,
         n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037,
         n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045,
         n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053,
         n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061,
         n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069,
         n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077,
         n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085,
         n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093,
         n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101,
         n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109,
         n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117,
         n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125,
         n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133,
         n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141,
         n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149,
         n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157,
         n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165,
         n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173,
         n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181,
         n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189,
         n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197,
         n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205,
         n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213,
         n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221,
         n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229,
         n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237,
         n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245,
         n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253,
         n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261,
         n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269,
         n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277,
         n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285,
         n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293,
         n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301,
         n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309,
         n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317,
         n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325,
         n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333,
         n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341,
         n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349,
         n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357,
         n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365,
         n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373,
         n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381,
         n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389,
         n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397,
         n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405,
         n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413,
         n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421,
         n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429,
         n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437,
         n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445,
         n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453,
         n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461,
         n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469,
         n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477,
         n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485,
         n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493,
         n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501,
         n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509,
         n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517,
         n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525,
         n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533,
         n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541,
         n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549,
         n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557,
         n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565,
         n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573,
         n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581,
         n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589,
         n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597,
         n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605,
         n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613,
         n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621,
         n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629,
         n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19638,
         n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646,
         n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654,
         n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662,
         n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670,
         n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678,
         n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686,
         n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694,
         n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702,
         n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710,
         n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718,
         n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726,
         n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734,
         n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742,
         n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750,
         n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758,
         n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766,
         n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774,
         n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782,
         n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790,
         n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798,
         n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806,
         n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814,
         n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822,
         n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830,
         n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838,
         n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846,
         n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854,
         n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862,
         n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870,
         n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878,
         n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886,
         n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894,
         n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902,
         n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910,
         n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918,
         n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926,
         n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934,
         n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942,
         n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950,
         n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958,
         n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966,
         n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974,
         n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982,
         n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990,
         n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998,
         n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006,
         n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014,
         n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022,
         n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030,
         n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038,
         n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046,
         n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054,
         n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062,
         n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070,
         n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078,
         n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086,
         n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094,
         n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102,
         n20103, n20104, n20105, n20107, n20108, n20109, n20110, n20111,
         n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119,
         n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127,
         n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135,
         n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143,
         n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151,
         n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159,
         n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167,
         n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175,
         n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183,
         n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191,
         n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199,
         n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207,
         n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215,
         n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223,
         n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231,
         n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239,
         n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247,
         n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255,
         n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263,
         n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271,
         n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279,
         n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287,
         n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295,
         n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303,
         n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311,
         n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319,
         n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327,
         n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335,
         n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343,
         n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351,
         n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359,
         n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367,
         n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375,
         n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383,
         n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391,
         n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399,
         n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407,
         n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415,
         n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423,
         n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431,
         n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439,
         n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447,
         n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455,
         n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463,
         n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471,
         n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479,
         n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487,
         n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495,
         n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503,
         n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511,
         n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519,
         n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527,
         n20528, n20529, n20530, n20531, n20532, n20533, n20534, n20535,
         n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543,
         n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551,
         n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559,
         n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567,
         n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575,
         n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583,
         n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591,
         n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599,
         n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607,
         n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615,
         n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623,
         n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631,
         n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639,
         n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647,
         n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655,
         n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663,
         n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671,
         n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679,
         n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687,
         n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695,
         n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703,
         n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711,
         n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719,
         n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727,
         n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735,
         n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743,
         n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751,
         n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759,
         n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767,
         n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775,
         n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783,
         n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791,
         n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799,
         n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807,
         n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815,
         n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823,
         n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831,
         n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839,
         n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847,
         n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855,
         n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863,
         n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871,
         n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879,
         n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887,
         n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895,
         n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903,
         n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911,
         n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919,
         n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927,
         n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935,
         n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943,
         n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951,
         n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959,
         n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967,
         n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975,
         n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983,
         n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991,
         n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999,
         n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007,
         n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015,
         n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023,
         n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031,
         n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039,
         n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047,
         n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055,
         n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063,
         n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071,
         n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079,
         n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087,
         n21088, n21089, n21090, n21091, n21092, n21093, n21094, n21095,
         n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103,
         n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111,
         n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119,
         n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127,
         n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135,
         n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143,
         n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151,
         n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159,
         n21160, n21161, n21162, n21163, n21164, n21165, n21166, n21167,
         n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175,
         n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183,
         n21184, n21185, n21186, n21187, n21188, n21189, n21190, n21191,
         n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199,
         n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207,
         n21208, n21209, n21210, n21211, n21212, n21213, n21214, n21215,
         n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223,
         n21224, n21225, n21226, n21227, n21228, n21229, n21230, n21231,
         n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239,
         n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247,
         n21248, n21249, n21250, n21251, n21252, n21253, n21254, n21255,
         n21256, n21257, n21258, n21259, n21260, n21261, n21262, n21263,
         n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271,
         n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279,
         n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21287,
         n21288, n21289, n21290, n21291, n21292, n21293, n21294, n21295,
         n21296, n21297, n21298, n21299, n21300, n21301, n21302, n21303,
         n21304, n21305, n21306, n21307, n21308, n21309, n21310, n21311,
         n21312, n21313, n21314, n21315, n21316, n21317, n21318, n21319,
         n21320, n21321, n21322, n21323, n21324, n21325, n21326, n21327,
         n21328, n21329, n21330, n21331, n21332, n21333, n21334, n21335,
         n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343,
         n21344, n21345, n21346, n21347, n21348, n21349, n21350, n21351,
         n21352, n21353, n21354, n21355, n21356, n21357, n21358, n21359,
         n21360, n21361, n21362, n21363, n21364, n21365, n21366, n21367,
         n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375,
         n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21383,
         n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391,
         n21392, n21393, n21394, n21395, n21396, n21397, n21398, n21399,
         n21400, n21401, n21402, n21403, n21404, n21405, n21406, n21407,
         n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415,
         n21416, n21417, n21418, n21419, n21420, n21421, n21422, n21423,
         n21424, n21425, n21426, n21427, n21428, n21429, n21430, n21431,
         n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439,
         n21440, n21441, n21442, n21443, n21444, n21445, n21446, n21447,
         n21448, n21449, n21450, n21451, n21452, n21453, n21454, n21455,
         n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463,
         n21464, n21465, n21466, n21467, n21468, n21469, n21470, n21471,
         n21472, n21473, n21474, n21475, n21476, n21477, n21478, n21479,
         n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487,
         n21488, n21489, n21490, n21491, n21492, n21493, n21494, n21495,
         n21496, n21497, n21498, n21499, n21500, n21501, n21502, n21503,
         n21504, n21505, n21506, n21507, n21508, n21509, n21510, n21511,
         n21512, n21513, n21514, n21515, n21516, n21517, n21518, n21519,
         n21520, n21521, n21522, n21523, n21524, n21525, n21526, n21527,
         n21528, n21529, n21530, n21531, n21532, n21533, n21534, n21535,
         n21536, n21537, n21538, n21539, n21540, n21541, n21542, n21543,
         n21544, n21545, n21546, n21547, n21548, n21549, n21550, n21551,
         n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559,
         n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567,
         n21568, n21569, n21570, n21571, n21572, n21573, n21574, n21575,
         n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583,
         n21584, n21585, n21586, n21587, n21588, n21589, n21590, n21591,
         n21592, n21593, n21594, n21595, n21596, n21597, n21598, n21599,
         n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607,
         n21608, n21609, n21610, n21611, n21612, n21613, n21614, n21615,
         n21616, n21617, n21618, n21619, n21620, n21621, n21622, n21623,
         n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631,
         n21632, n21633, n21634, n21635, n21636, n21637, n21638, n21639,
         n21640, n21641, n21642, n21643, n21644, n21645, n21646, n21647,
         n21648, n21649, n21650, n21651, n21652, n21653, n21654, n21655,
         n21656, n21657, n21658, n21659, n21660, n21661, n21662, n21663,
         n21664, n21665, n21666, n21667, n21668, n21669, n21670, n21671,
         n21672, n21673, n21674, n21675, n21676, n21677, n21678, n21679,
         n21680, n21681, n21682, n21683, n21684, n21685, n21686, n21687,
         n21688, n21689, n21690, n21691, n21692, n21693, n21694, n21695,
         n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703,
         n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711,
         n21712, n21713, n21714, n21715, n21716, n21717, n21718, n21719,
         n21720, n21721, n21722, n21723, n21724, n21725, n21726, n21727,
         n21728, n21729, n21730, n21731, n21732, n21733, n21734, n21735,
         n21736, n21737, n21738, n21739, n21740, n21741, n21742, n21743,
         n21744, n21745, n21746, n21747, n21748, n21749, n21750, n21751,
         n21752, n21753, n21754, n21755, n21756, n21757, n21758, n21759,
         n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767,
         n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775,
         n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783,
         n21784, n21785, n21786, n21787, n21788, n21789, n21790, n21791,
         n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799,
         n21800, n21801, n21802, n21803, n21804, n21805, n21806, n21807,
         n21808, n21809, n21810, n21811, n21812, n21813, n21814, n21815,
         n21816, n21817, n21818, n21819, n21820, n21821, n21822, n21823,
         n21824, n21825, n21826, n21827, n21828, n21829, n21830, n21831,
         n21832, n21833, n21834, n21835, n21836, n21837, n21838, n21839,
         n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847,
         n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855,
         n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21863,
         n21864, n21865, n21866, n21867, n21868, n21869, n21870, n21871,
         n21872, n21873, n21874, n21875, n21876, n21877, n21878, n21879,
         n21880, n21881, n21882, n21883, n21884, n21885, n21886, n21887,
         n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895,
         n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903,
         n21904, n21905, n21906, n21907, n21908, n21909, n21910, n21911,
         n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919,
         n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927,
         n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935,
         n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943,
         n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951,
         n21952, n21953, n21954, n21955, n21956, n21957, n21958, n21959,
         n21960, n21961, n21962, n21963, n21964, n21965, n21966, n21967,
         n21968, n21969, n21970, n21971, n21972, n21973, n21974, n21975,
         n21976, n21977, n21978, n21979, n21980, n21981, n21982, n21983,
         n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991,
         n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999,
         n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007,
         n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015,
         n22016, n22017, n22018, n22019, n22020, n22021, n22022, n22023,
         n22024, n22025, n22026, n22027, n22028, n22029, n22030, n22031,
         n22032, n22033, n22034, n22035, n22036, n22037, n22038, n22039,
         n22040, n22041, n22042, n22043, n22044, n22045, n22046, n22047,
         n22048, n22049, n22050, n22051, n22052, n22053, n22054, n22055,
         n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22063,
         n22064, n22065, n22066, n22067, n22068, n22069, n22070, n22071,
         n22072, n22073, n22074, n22075, n22076, n22077, n22078, n22079,
         n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087,
         n22088, n22089, n22090, n22091, n22092, n22093, n22094, n22095,
         n22096, n22097, n22098, n22099, n22100, n22101, n22102, n22103,
         n22104, n22105, n22106, n22107, n22108, n22109, n22110, n22111,
         n22112, n22113, n22114, n22115, n22116, n22117, n22118, n22119,
         n22120, n22121, n22122, n22123, n22124, n22125, n22126, n22127,
         n22128, n22129, n22130, n22131, n22132, n22133, n22134, n22135,
         n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143,
         n22144, n22145, n22146, n22147, n22148, n22149, n22150, n22151,
         n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159,
         n22160, n22161, n22162, n22163, n22164, n22165, n22166, n22167,
         n22168, n22169, n22170, n22171, n22172, n22173, n22174, n22175,
         n22176, n22177, n22178, n22179, n22180, n22181, n22182, n22183,
         n22184, n22185, n22186, n22187, n22188, n22189, n22190, n22191,
         n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199,
         n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207,
         n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215,
         n22216, n22217, n22218, n22219, n22220, n22221, n22222, n22223,
         n22224, n22225, n22226, n22227, n22228, n22229, n22230, n22231,
         n22232, n22233, n22234, n22235, n22236, n22237, n22238, n22239,
         n22240, n22241, n22242, n22243, n22244, n22245, n22246, n22247,
         n22248, n22249, n22250, n22251, n22252, n22253, n22254, n22255,
         n22256, n22257, n22258, n22259, n22260, n22261, n22262, n22263,
         n22264, n22265, n22266, n22267, n22268, n22269, n22270, n22271,
         n22272, n22273, n22274, n22275, n22276, n22277, n22278, n22279,
         n22280, n22281, n22282, n22283, n22284, n22285, n22286, n22287,
         n22288, n22289, n22290, n22291, n22292, n22293, n22294, n22295,
         n22296, n22297, n22298, n22299, n22300, n22301, n22302, n22303,
         n22304, n22305, n22306, n22307, n22308, n22309, n22310, n22311,
         n22312, n22313, n22314, n22315, n22316, n22317, n22318, n22319,
         n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327,
         n22328, n22329, n22330, n22331, n22332, n22333, n22334, n22335,
         n22336, n22337, n22338, n22339, n22340, n22341, n22342, n22343,
         n22344, n22345, n22346, n22347, n22348, n22349, n22350, n22351,
         n22352, n22353, n22354, n22355, n22356, n22357, n22358, n22359,
         n22360, n22361, n22362, n22363, n22364, n22365, n22366, n22367,
         n22368, n22369, n22370, n22371, n22372, n22373, n22374, n22375,
         n22376, n22377, n22378, n22379, n22380, n22381, n22382, n22383,
         n22384, n22385, n22386, n22387, n22388, n22389, n22390, n22391,
         n22392, n22393, n22394, n22395, n22396, n22397, n22398, n22399,
         n22400, n22401, n22402, n22403, n22404, n22405, n22406, n22407,
         n22408, n22409, n22410, n22411, n22412, n22413, n22414, n22415,
         n22416, n22417, n22418, n22419, n22420, n22421, n22422, n22423,
         n22424, n22425, n22426, n22427, n22428, n22429, n22430, n22431,
         n22432, n22433, n22434, n22435, n22436, n22437, n22438, n22439,
         n22440, n22441, n22442, n22443, n22444, n22445, n22446, n22447,
         n22448, n22449, n22450, n22451, n22452, n22453, n22454, n22455,
         n22456, n22457, n22458, n22459, n22460, n22461, n22462, n22463,
         n22464, n22465, n22466, n22467, n22468, n22469, n22470, n22471,
         n22472, n22473, n22474, n22475, n22476, n22477, n22478, n22479,
         n22480, n22481, n22482, n22483, n22484, n22485, n22486, n22487,
         n22488, n22489, n22490, n22491, n22492, n22493, n22494, n22495,
         n22496, n22497, n22498, n22499, n22500, n22501, n22502, n22503,
         n22504, n22505, n22506, n22507, n22508, n22509, n22510, n22511,
         n22512, n22513, n22514, n22515, n22516, n22517, n22518, n22519,
         n22520, n22521, n22522, n22523, n22524, n22525, n22526, n22527,
         n22528, n22529, n22530, n22531, n22532, n22533, n22534, n22535,
         n22536, n22537, n22538, n22539, n22540, n22541, n22542, n22543,
         n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551,
         n22552, n22553, n22554, n22555, n22556, n22557, n22558, n22559,
         n22560, n22561, n22562, n22563, n22564, n22565, n22566, n22567,
         n22568, n22569, n22570, n22571, n22572, n22573, n22574, n22575,
         n22576, n22577, n22578, n22579, n22580, n22581, n22582, n22583,
         n22584, n22585, n22586, n22587, n22588, n22589, n22590, n22591,
         n22592, n22593, n22594, n22595, n22596, n22597, n22598, n22599,
         n22600, n22601, n22602, n22603, n22604, n22605, n22606, n22607,
         n22608, n22609, n22610, n22611, n22612, n22613, n22614, n22615,
         n22616, n22617, n22618, n22619, n22620, n22621, n22622, n22623,
         n22624, n22625, n22626, n22627, n22628, n22629, n22630, n22631,
         n22632, n22633, n22634, n22635, n22636, n22637, n22638, n22639,
         n22640, n22641, n22642, n22643, n22644, n22645, n22646, n22647,
         n22648, n22649, n22650, n22651, n22652, n22653, n22654, n22655,
         n22656, n22657, n22658, n22659, n22660, n22661, n22662, n22663,
         n22664, n22665, n22666, n22667, n22668, n22669, n22670, n22671,
         n22672, n22673, n22674, n22675, n22676, n22677, n22678, n22679,
         n22680, n22681, n22682, n22683, n22684, n22685;

  NAND2_X1 U11244 ( .A1(n11577), .A2(n11576), .ZN(n17307) );
  CLKBUF_X2 U11247 ( .A(n12989), .Z(n14002) );
  OR2_X1 U11248 ( .A1(n11872), .A2(n11874), .ZN(n11977) );
  BUF_X2 U11249 ( .A(n14341), .Z(n18342) );
  BUF_X2 U11250 ( .A(n14342), .Z(n18347) );
  CLKBUF_X2 U11251 ( .A(n14447), .Z(n18165) );
  INV_X1 U11252 ( .A(n21337), .ZN(n14577) );
  CLKBUF_X2 U11253 ( .A(n13185), .Z(n13804) );
  CLKBUF_X2 U11254 ( .A(n13082), .Z(n13801) );
  INV_X1 U11255 ( .A(n11209), .ZN(n18313) );
  BUF_X2 U11256 ( .A(n14372), .Z(n18288) );
  CLKBUF_X1 U11257 ( .A(n14447), .Z(n18331) );
  CLKBUF_X1 U11258 ( .A(n14389), .Z(n18341) );
  CLKBUF_X2 U11259 ( .A(n11786), .Z(n20020) );
  INV_X2 U11260 ( .A(n11209), .ZN(n18349) );
  CLKBUF_X1 U11261 ( .A(n11784), .Z(n19970) );
  AND2_X2 U11262 ( .A1(n14139), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11909) );
  NAND2_X1 U11264 ( .A1(n11760), .A2(n14235), .ZN(n13906) );
  AND2_X1 U11265 ( .A1(n11883), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12556) );
  AND2_X1 U11266 ( .A1(n11183), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14072) );
  INV_X2 U11267 ( .A(n11760), .ZN(n11785) );
  AND2_X1 U11268 ( .A1(n14137), .A2(n11891), .ZN(n11906) );
  BUF_X1 U11269 ( .A(n12963), .Z(n15229) );
  INV_X2 U11270 ( .A(n12966), .ZN(n14899) );
  INV_X4 U11271 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11716) );
  AND2_X1 U11272 ( .A1(n12846), .A2(n12847), .ZN(n12899) );
  BUF_X2 U11273 ( .A(n11660), .Z(n11188) );
  CLKBUF_X3 U11274 ( .A(n11660), .Z(n11186) );
  CLKBUF_X1 U11275 ( .A(n13032), .Z(n11179) );
  AND2_X1 U11276 ( .A1(n14961), .A2(n12849), .ZN(n12997) );
  AND2_X1 U11277 ( .A1(n12848), .A2(n12849), .ZN(n13377) );
  BUF_X1 U11278 ( .A(n13032), .Z(n11177) );
  AND2_X1 U11279 ( .A1(n12838), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n16603) );
  INV_X1 U11281 ( .A(n22684), .ZN(n11138) );
  AND2_X1 U11282 ( .A1(n11187), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14071) );
  NAND2_X1 U11283 ( .A1(n12378), .A2(n12377), .ZN(n12387) );
  AND2_X1 U11284 ( .A1(n11170), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11942) );
  INV_X2 U11285 ( .A(n20020), .ZN(n12493) );
  INV_X1 U11286 ( .A(n13918), .ZN(n15972) );
  AND2_X1 U11289 ( .A1(n12762), .A2(n17058), .ZN(n16849) );
  NAND2_X1 U11290 ( .A1(n16907), .A2(n12414), .ZN(n16894) );
  INV_X1 U11291 ( .A(n12007), .ZN(n17363) );
  BUF_X1 U11293 ( .A(n20933), .Z(n21128) );
  INV_X2 U11294 ( .A(n21576), .ZN(n21790) );
  INV_X1 U11295 ( .A(n14555), .ZN(n19470) );
  NOR2_X1 U11296 ( .A1(n15875), .A2(n15911), .ZN(n15910) );
  INV_X1 U11297 ( .A(n18571), .ZN(n18593) );
  INV_X1 U11298 ( .A(n22260), .ZN(n22251) );
  NOR2_X1 U11299 ( .A1(n14401), .A2(n14400), .ZN(n21350) );
  INV_X1 U11300 ( .A(n18661), .ZN(n18675) );
  INV_X2 U11301 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n21382) );
  AND3_X1 U11302 ( .A1(n11956), .A2(n11957), .A3(n12030), .ZN(n11139) );
  NAND2_X1 U11303 ( .A1(n14872), .A2(n12849), .ZN(n16605) );
  XNOR2_X2 U11305 ( .A(n13054), .B(n14893), .ZN(n15070) );
  NOR2_X4 U11306 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11891) );
  AOI21_X2 U11307 ( .B1(n12709), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n11775), 
        .ZN(n11776) );
  NOR2_X2 U11309 ( .A1(n16860), .A2(n17079), .ZN(n12761) );
  XNOR2_X2 U11311 ( .A(n12155), .B(n12148), .ZN(n19024) );
  AND2_X2 U11312 ( .A1(n11299), .A2(n12054), .ZN(n11660) );
  AOI21_X2 U11313 ( .B1(n18586), .B2(n21641), .A(n14429), .ZN(n18569) );
  NOR2_X1 U11314 ( .A1(n12962), .A2(n12966), .ZN(n12974) );
  OR2_X1 U11315 ( .A1(n11213), .A2(n12807), .ZN(n11365) );
  AND2_X1 U11316 ( .A1(n11300), .A2(n11234), .ZN(n12200) );
  NAND2_X1 U11317 ( .A1(n13477), .A2(n13476), .ZN(n15934) );
  AND2_X1 U11318 ( .A1(n11293), .A2(n11291), .ZN(n11294) );
  OR2_X1 U11319 ( .A1(n16387), .A2(n13234), .ZN(n16377) );
  OR2_X1 U11320 ( .A1(n16726), .A2(n11258), .ZN(n11515) );
  INV_X4 U11321 ( .A(n16352), .ZN(n11452) );
  CLKBUF_X1 U11322 ( .A(n12386), .Z(n12396) );
  OR2_X1 U11323 ( .A1(n12813), .A2(n12814), .ZN(n12331) );
  AND2_X1 U11324 ( .A1(n21668), .A2(n18521), .ZN(n18511) );
  AND2_X1 U11325 ( .A1(n15040), .A2(n11264), .ZN(n15563) );
  AND2_X1 U11326 ( .A1(n15706), .A2(n15714), .ZN(n15713) );
  OAI21_X1 U11327 ( .B1(n18589), .B2(n21509), .A(n11316), .ZN(n18645) );
  OR2_X1 U11328 ( .A1(n14034), .A2(n11485), .ZN(n11482) );
  OAI21_X1 U11329 ( .B1(n14999), .B2(n13215), .A(n13103), .ZN(n15209) );
  AOI211_X1 U11330 ( .C1(n19825), .C2(n19933), .A(n19932), .B(n20287), .ZN(
        n19822) );
  NAND2_X1 U11331 ( .A1(n18425), .A2(n14418), .ZN(n18639) );
  NAND2_X1 U11332 ( .A1(n14994), .A2(n14995), .ZN(n14993) );
  NOR2_X4 U11333 ( .A1(n21776), .A2(n21625), .ZN(n21756) );
  INV_X2 U11334 ( .A(n21795), .ZN(n21776) );
  NAND2_X1 U11335 ( .A1(n13069), .A2(n15454), .ZN(n14968) );
  NAND2_X1 U11336 ( .A1(n17804), .A2(n15063), .ZN(n22268) );
  NAND2_X1 U11337 ( .A1(n13045), .A2(n13044), .ZN(n13065) );
  NOR2_X1 U11338 ( .A1(n21373), .A2(n14560), .ZN(n15964) );
  NOR2_X1 U11339 ( .A1(n21816), .A2(n20671), .ZN(n15963) );
  OAI211_X1 U11340 ( .C1(n11174), .C2(n18862), .A(n11803), .B(n11802), .ZN(
        n11804) );
  CLKBUF_X3 U11341 ( .A(n11824), .Z(n12700) );
  INV_X1 U11342 ( .A(n11780), .ZN(n12482) );
  NAND2_X2 U11343 ( .A1(n13009), .A2(n16023), .ZN(n12971) );
  CLKBUF_X1 U11344 ( .A(n12964), .Z(n15146) );
  INV_X1 U11345 ( .A(n13906), .ZN(n12451) );
  INV_X2 U11346 ( .A(n13009), .ZN(n16022) );
  INV_X1 U11347 ( .A(n12717), .ZN(n11770) );
  INV_X1 U11348 ( .A(n11769), .ZN(n12442) );
  OR2_X2 U11349 ( .A1(n12893), .A2(n12892), .ZN(n12966) );
  OR2_X1 U11350 ( .A1(n12883), .A2(n12882), .ZN(n13915) );
  NAND2_X1 U11351 ( .A1(n11216), .A2(n11329), .ZN(n11328) );
  NAND2_X1 U11352 ( .A1(n11215), .A2(n11327), .ZN(n11326) );
  BUF_X2 U11354 ( .A(n13032), .Z(n11146) );
  BUF_X1 U11355 ( .A(n13136), .Z(n13784) );
  CLKBUF_X2 U11356 ( .A(n13012), .Z(n13563) );
  CLKBUF_X2 U11357 ( .A(n13377), .Z(n13799) );
  CLKBUF_X2 U11358 ( .A(n13018), .Z(n13810) );
  BUF_X2 U11360 ( .A(n12894), .Z(n13779) );
  BUF_X2 U11361 ( .A(n13083), .Z(n13778) );
  CLKBUF_X2 U11362 ( .A(n11886), .Z(n14277) );
  CLKBUF_X2 U11363 ( .A(n12899), .Z(n13800) );
  CLKBUF_X2 U11364 ( .A(n20425), .Z(n21877) );
  AND2_X2 U11365 ( .A1(n12848), .A2(n12846), .ZN(n13136) );
  CLKBUF_X1 U11366 ( .A(n11668), .Z(n11184) );
  CLKBUF_X2 U11367 ( .A(n13444), .Z(n13803) );
  AND2_X2 U11368 ( .A1(n12848), .A2(n12841), .ZN(n13032) );
  CLKBUF_X1 U11369 ( .A(n11668), .Z(n11183) );
  BUF_X2 U11370 ( .A(n12997), .Z(n13432) );
  CLKBUF_X1 U11371 ( .A(n11884), .Z(n11140) );
  AND2_X1 U11372 ( .A1(n11298), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11892) );
  NAND2_X1 U11373 ( .A1(n21382), .A2(n17368), .ZN(n20747) );
  NAND2_X1 U11374 ( .A1(n21382), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14310) );
  INV_X2 U11375 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n19225) );
  NAND2_X1 U11376 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n21360) );
  AND2_X1 U11377 ( .A1(n12760), .A2(n12755), .ZN(n11386) );
  NAND2_X1 U11378 ( .A1(n11440), .A2(n11439), .ZN(n13252) );
  AOI21_X1 U11379 ( .B1(n17053), .B2(n17879), .A(n11289), .ZN(n12417) );
  OR2_X1 U11380 ( .A1(n14293), .A2(n17859), .ZN(n14301) );
  OAI21_X1 U11381 ( .B1(n16893), .B2(n17138), .A(n11365), .ZN(n12811) );
  AOI21_X1 U11382 ( .B1(n22685), .B2(n12758), .A(n11335), .ZN(n11334) );
  OAI21_X1 U11383 ( .B1(n12779), .B2(n12780), .A(n12435), .ZN(n12441) );
  NAND2_X1 U11384 ( .A1(n11368), .A2(n11366), .ZN(n16893) );
  AND2_X1 U11385 ( .A1(n13243), .A2(n11441), .ZN(n16271) );
  AND2_X1 U11386 ( .A1(n16308), .A2(n11442), .ZN(n11441) );
  NOR2_X1 U11387 ( .A1(n12778), .A2(n12791), .ZN(n12756) );
  XNOR2_X1 U11388 ( .A(n13831), .B(n13830), .ZN(n15990) );
  INV_X1 U11389 ( .A(n13242), .ZN(n16334) );
  OAI21_X1 U11390 ( .B1(n16060), .B2(n16061), .A(n16049), .ZN(n16293) );
  AND2_X1 U11391 ( .A1(n16160), .A2(n16159), .ZN(n22263) );
  OR2_X1 U11392 ( .A1(n16160), .A2(n16097), .ZN(n16095) );
  NAND2_X1 U11393 ( .A1(n16932), .A2(n12803), .ZN(n16922) );
  NAND2_X1 U11394 ( .A1(n11464), .A2(n11465), .ZN(n13242) );
  NAND2_X1 U11395 ( .A1(n13240), .A2(n16345), .ZN(n11464) );
  AOI21_X1 U11396 ( .B1(n16678), .B2(n16676), .A(n16675), .ZN(n14288) );
  NAND3_X1 U11397 ( .A1(n17307), .A2(n12408), .A3(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11340) );
  OAI211_X1 U11398 ( .C1(n16683), .C2(n16692), .A(n16685), .B(n16689), .ZN(
        n16678) );
  NOR2_X1 U11399 ( .A1(n14251), .A2(n14250), .ZN(n16683) );
  NAND2_X1 U11400 ( .A1(n11449), .A2(n11447), .ZN(n13238) );
  NAND2_X1 U11401 ( .A1(n16977), .A2(n12799), .ZN(n16969) );
  OR2_X1 U11402 ( .A1(n17051), .A2(n11336), .ZN(n11335) );
  OR2_X1 U11403 ( .A1(n12363), .A2(n12362), .ZN(n11289) );
  NOR2_X1 U11404 ( .A1(n16697), .A2(n11650), .ZN(n14251) );
  AOI21_X1 U11405 ( .B1(n11445), .B2(n11448), .A(n11444), .ZN(n11443) );
  NOR2_X1 U11406 ( .A1(n16699), .A2(n16698), .ZN(n16697) );
  XNOR2_X1 U11407 ( .A(n14215), .B(n11641), .ZN(n16699) );
  AND2_X1 U11408 ( .A1(n11578), .A2(n12394), .ZN(n11576) );
  INV_X1 U11409 ( .A(n13237), .ZN(n11448) );
  OAI21_X1 U11410 ( .B1(n16710), .B2(n11487), .A(n11486), .ZN(n14215) );
  XNOR2_X1 U11411 ( .A(n16679), .B(n12793), .ZN(n16829) );
  XNOR2_X1 U11412 ( .A(n12708), .B(n12707), .ZN(n19161) );
  NAND2_X1 U11413 ( .A1(n16710), .A2(n11259), .ZN(n11486) );
  NAND2_X1 U11414 ( .A1(n16712), .A2(n16711), .ZN(n16710) );
  INV_X1 U11415 ( .A(n12387), .ZN(n12382) );
  AOI211_X1 U11416 ( .C1(n14629), .C2(n18748), .A(n14628), .B(n14627), .ZN(
        n14630) );
  NAND2_X1 U11417 ( .A1(n11490), .A2(n11275), .ZN(n16712) );
  AND2_X1 U11418 ( .A1(n21296), .A2(n11208), .ZN(n21281) );
  AND2_X1 U11419 ( .A1(n16877), .A2(n11610), .ZN(n11608) );
  OR2_X1 U11420 ( .A1(n12401), .A2(n12430), .ZN(n12409) );
  NOR2_X1 U11421 ( .A1(n21273), .A2(n21274), .ZN(n21296) );
  OR2_X1 U11422 ( .A1(n12331), .A2(n16724), .ZN(n16726) );
  NAND2_X1 U11423 ( .A1(n12787), .A2(n12786), .ZN(n16017) );
  OR2_X1 U11424 ( .A1(n19012), .A2(n12430), .ZN(n16911) );
  OR2_X1 U11425 ( .A1(n15053), .A2(n15402), .ZN(n15404) );
  AND2_X1 U11426 ( .A1(n12002), .A2(n12001), .ZN(n12023) );
  XNOR2_X1 U11427 ( .A(n13134), .B(n21937), .ZN(n15218) );
  XNOR2_X1 U11428 ( .A(n12213), .B(n12214), .ZN(n19052) );
  AND2_X1 U11429 ( .A1(n12165), .A2(n12803), .ZN(n16930) );
  OR2_X1 U11430 ( .A1(n16794), .A2(n16795), .ZN(n16796) );
  AND2_X1 U11431 ( .A1(n22104), .A2(n15244), .ZN(n22260) );
  NAND2_X1 U11432 ( .A1(n15212), .A2(n13105), .ZN(n13134) );
  NAND2_X1 U11433 ( .A1(n21653), .A2(n14613), .ZN(n18589) );
  INV_X1 U11434 ( .A(n14613), .ZN(n18757) );
  NAND2_X1 U11435 ( .A1(n15210), .A2(n15209), .ZN(n15212) );
  OAI21_X1 U11436 ( .B1(n14999), .B2(n13471), .A(n13329), .ZN(n13330) );
  OR2_X1 U11437 ( .A1(n21871), .A2(n20741), .ZN(n18758) );
  OAI21_X2 U11438 ( .B1(n20674), .B2(P3_STATE2_REG_0__SCAN_IN), .A(n21871), 
        .ZN(n18753) );
  NOR2_X2 U11439 ( .A1(n17814), .A2(n15232), .ZN(n22236) );
  OAI22_X1 U11440 ( .A1(n12092), .A2(n12091), .B1(n12093), .B2(n12094), .ZN(
        n11305) );
  CLKBUF_X1 U11441 ( .A(n15993), .Z(n16256) );
  OAI21_X1 U11442 ( .B1(n14889), .B2(n14888), .A(n14031), .ZN(n14985) );
  AND2_X1 U11443 ( .A1(n11192), .A2(n11873), .ZN(n19754) );
  NAND2_X1 U11444 ( .A1(n13123), .A2(n13122), .ZN(n15031) );
  AND2_X1 U11445 ( .A1(n11321), .A2(n21845), .ZN(n21196) );
  AND2_X1 U11446 ( .A1(n12142), .A2(n11393), .ZN(n12166) );
  NAND2_X1 U11447 ( .A1(n11611), .A2(n13094), .ZN(n13096) );
  INV_X1 U11448 ( .A(n12178), .ZN(n12142) );
  NAND2_X1 U11449 ( .A1(n13067), .A2(n13216), .ZN(n13332) );
  OR2_X1 U11450 ( .A1(n13080), .A2(n13079), .ZN(n11612) );
  XNOR2_X1 U11451 ( .A(n13065), .B(n13064), .ZN(n13337) );
  NAND2_X1 U11452 ( .A1(n13080), .A2(n13079), .ZN(n14885) );
  NAND2_X1 U11453 ( .A1(n18688), .A2(n14414), .ZN(n18401) );
  NOR2_X2 U11454 ( .A1(n12736), .A2(n12711), .ZN(n19202) );
  AND2_X1 U11455 ( .A1(n11525), .A2(n11522), .ZN(n15817) );
  INV_X2 U11456 ( .A(n16727), .ZN(n11141) );
  NAND2_X1 U11457 ( .A1(n11838), .A2(n11574), .ZN(n11836) );
  NAND2_X1 U11458 ( .A1(n11573), .A2(n11572), .ZN(n11838) );
  AND2_X1 U11459 ( .A1(n12270), .A2(n11848), .ZN(n12271) );
  NAND2_X1 U11460 ( .A1(n11851), .A2(n11831), .ZN(n18858) );
  AND2_X1 U11461 ( .A1(n11504), .A2(n15022), .ZN(n11503) );
  OR2_X1 U11462 ( .A1(n12519), .A2(n12515), .ZN(n15202) );
  INV_X2 U11463 ( .A(n20683), .ZN(n20734) );
  OR3_X2 U11464 ( .A1(n15963), .A2(n20682), .A3(n11320), .ZN(n14564) );
  AOI211_X2 U11465 ( .C1(n14559), .C2(n14558), .A(n14557), .B(n14556), .ZN(
        n21377) );
  AOI21_X1 U11466 ( .B1(n15013), .B2(n11649), .A(n12514), .ZN(n12519) );
  AND2_X1 U11467 ( .A1(n14546), .A2(n20679), .ZN(n21816) );
  NAND2_X1 U11468 ( .A1(n11799), .A2(n11798), .ZN(n11587) );
  NOR2_X2 U11469 ( .A1(n14384), .A2(n21653), .ZN(n18548) );
  OR3_X1 U11470 ( .A1(n14562), .A2(n21231), .A3(n20736), .ZN(n20679) );
  AND2_X1 U11471 ( .A1(n14820), .A2(n14821), .ZN(n12510) );
  AND2_X1 U11472 ( .A1(n12728), .A2(n11756), .ZN(n11807) );
  NAND2_X1 U11473 ( .A1(n12689), .A2(n11768), .ZN(n11802) );
  NOR2_X1 U11474 ( .A1(n12113), .A2(n12052), .ZN(n11391) );
  INV_X1 U11475 ( .A(n11794), .ZN(n12722) );
  MUX2_X1 U11476 ( .A(n12045), .B(P2_EBX_REG_3__SCAN_IN), .S(n20020), .Z(
        n12052) );
  NAND2_X2 U11477 ( .A1(n15697), .A2(n12532), .ZN(n12516) );
  NAND2_X1 U11478 ( .A1(n12532), .A2(n12493), .ZN(n12653) );
  NAND2_X1 U11479 ( .A1(n11248), .A2(n12961), .ZN(n12970) );
  NAND2_X1 U11480 ( .A1(n11434), .A2(n11433), .ZN(n14403) );
  NAND3_X1 U11481 ( .A1(n11727), .A2(n11726), .A3(n11789), .ZN(n11778) );
  INV_X1 U11482 ( .A(n11793), .ZN(n11768) );
  INV_X1 U11483 ( .A(n14858), .ZN(n16026) );
  OR2_X1 U11484 ( .A1(n14833), .A2(n12989), .ZN(n14919) );
  AND2_X1 U11485 ( .A1(n11763), .A2(n20155), .ZN(n11725) );
  NAND2_X1 U11486 ( .A1(n11766), .A2(n11765), .ZN(n11780) );
  NAND2_X1 U11487 ( .A1(n20247), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11793) );
  INV_X1 U11488 ( .A(n12720), .ZN(n12726) );
  NAND2_X1 U11489 ( .A1(n11920), .A2(n11383), .ZN(n12040) );
  INV_X2 U11490 ( .A(n11771), .ZN(n13896) );
  NAND2_X1 U11491 ( .A1(n13047), .A2(n13009), .ZN(n14833) );
  CLKBUF_X1 U11492 ( .A(n12974), .Z(n12975) );
  NAND2_X1 U11493 ( .A1(n12494), .A2(n12717), .ZN(n11789) );
  AND2_X1 U11494 ( .A1(n16022), .A2(n13915), .ZN(n16192) );
  AND2_X2 U11495 ( .A1(n14899), .A2(n12962), .ZN(n14858) );
  INV_X2 U11496 ( .A(n12964), .ZN(n16021) );
  OR2_X2 U11497 ( .A1(n20662), .A2(n20601), .ZN(n20648) );
  OR2_X1 U11498 ( .A1(n12905), .A2(n12904), .ZN(n12962) );
  NAND2_X1 U11499 ( .A1(n11755), .A2(n11754), .ZN(n14235) );
  NAND2_X2 U11500 ( .A1(n11328), .A2(n11326), .ZN(n11762) );
  NAND2_X1 U11501 ( .A1(n11691), .A2(n11690), .ZN(n11769) );
  NAND2_X2 U11502 ( .A1(n11711), .A2(n11710), .ZN(n19758) );
  OR2_X1 U11503 ( .A1(n12865), .A2(n12864), .ZN(n12955) );
  AND4_X1 U11504 ( .A1(n12013), .A2(n12012), .A3(n12011), .A4(n12010), .ZN(
        n12020) );
  INV_X2 U11505 ( .A(U212), .ZN(n20663) );
  INV_X2 U11506 ( .A(U214), .ZN(n20662) );
  AND4_X1 U11507 ( .A1(n12910), .A2(n12909), .A3(n12908), .A4(n12907), .ZN(
        n12919) );
  AND4_X1 U11508 ( .A1(n12940), .A2(n12939), .A3(n12938), .A4(n12937), .ZN(
        n12941) );
  AND4_X1 U11509 ( .A1(n12853), .A2(n12852), .A3(n12851), .A4(n12850), .ZN(
        n12854) );
  AND4_X1 U11510 ( .A1(n12936), .A2(n12935), .A3(n12934), .A4(n12933), .ZN(
        n12942) );
  AND4_X1 U11511 ( .A1(n12932), .A2(n12931), .A3(n12930), .A4(n12929), .ZN(
        n12943) );
  AND4_X1 U11512 ( .A1(n12928), .A2(n12927), .A3(n12926), .A4(n12925), .ZN(
        n12944) );
  AND4_X1 U11513 ( .A1(n12914), .A2(n12913), .A3(n12912), .A4(n12911), .ZN(
        n12918) );
  AND3_X1 U11514 ( .A1(n11683), .A2(n11682), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11225) );
  AND2_X1 U11515 ( .A1(n11693), .A2(n11694), .ZN(n11329) );
  CLKBUF_X3 U11516 ( .A(n18101), .Z(n18332) );
  CLKBUF_X3 U11517 ( .A(n14349), .Z(n18350) );
  INV_X1 U11518 ( .A(n11190), .ZN(n11163) );
  BUF_X2 U11519 ( .A(n14390), .Z(n18055) );
  INV_X2 U11520 ( .A(n11190), .ZN(n11164) );
  CLKBUF_X2 U11521 ( .A(n18824), .Z(n21805) );
  CLKBUF_X1 U11522 ( .A(n11668), .Z(n11185) );
  CLKBUF_X1 U11523 ( .A(n13809), .Z(n13697) );
  BUF_X2 U11524 ( .A(n13032), .Z(n11176) );
  INV_X2 U11525 ( .A(n14606), .ZN(n11142) );
  BUF_X2 U11526 ( .A(n14389), .Z(n18234) );
  BUF_X4 U11527 ( .A(n14445), .Z(n11143) );
  NOR2_X1 U11528 ( .A1(n14309), .A2(n14307), .ZN(n18101) );
  BUF_X4 U11529 ( .A(n14395), .Z(n11144) );
  BUF_X4 U11530 ( .A(n14352), .Z(n11145) );
  CLKBUF_X3 U11531 ( .A(n11660), .Z(n11187) );
  INV_X1 U11532 ( .A(n19267), .ZN(n19127) );
  AND2_X2 U11533 ( .A1(n12848), .A2(n16603), .ZN(n13082) );
  NOR2_X1 U11534 ( .A1(n14309), .A2(n21360), .ZN(n14349) );
  INV_X2 U11535 ( .A(n18843), .ZN(n22303) );
  INV_X4 U11536 ( .A(n18103), .ZN(n18326) );
  INV_X2 U11537 ( .A(n20359), .ZN(n20410) );
  INV_X2 U11538 ( .A(n17988), .ZN(n17987) );
  INV_X2 U11539 ( .A(n14374), .ZN(n11147) );
  NOR2_X1 U11540 ( .A1(n21354), .A2(n18754), .ZN(n18824) );
  AND2_X2 U11541 ( .A1(n11890), .A2(n14137), .ZN(n11962) );
  OR2_X1 U11542 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n17747), .ZN(
        n18103) );
  NAND2_X1 U11543 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n21388), .ZN(
        n21383) );
  AND2_X2 U11544 ( .A1(n11438), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12847) );
  AND2_X2 U11545 ( .A1(n12840), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12848) );
  NAND2_X1 U11546 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n17368), .ZN(
        n14307) );
  INV_X2 U11547 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n21388) );
  INV_X1 U11548 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12840) );
  AND2_X2 U11549 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14872) );
  INV_X1 U11550 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12838) );
  INV_X1 U11551 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11438) );
  NOR2_X1 U11552 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14137) );
  NAND2_X1 U11553 ( .A1(n11589), .A2(n18900), .ZN(n12115) );
  INV_X2 U11554 ( .A(n15556), .ZN(n13375) );
  NOR2_X2 U11555 ( .A1(n15330), .A2(n15329), .ZN(n15328) );
  NAND2_X1 U11556 ( .A1(n12115), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17022) );
  NAND2_X2 U11557 ( .A1(n12053), .A2(n15638), .ZN(n17843) );
  NOR2_X2 U11558 ( .A1(n16377), .A2(n13235), .ZN(n20574) );
  NAND3_X1 U11559 ( .A1(n11956), .A2(n11957), .A3(n12030), .ZN(n11148) );
  NOR2_X1 U11560 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11299) );
  AND2_X1 U11561 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11890) );
  NAND2_X1 U11562 ( .A1(n15827), .A2(n15826), .ZN(n11149) );
  OR2_X1 U11563 ( .A1(n20551), .A2(n11160), .ZN(n11150) );
  NAND2_X1 U11564 ( .A1(n11150), .A2(n11151), .ZN(n15825) );
  AND2_X1 U11565 ( .A1(n15826), .A2(n11158), .ZN(n11151) );
  NAND2_X1 U11566 ( .A1(n13069), .A2(n13072), .ZN(n13080) );
  NAND2_X1 U11567 ( .A1(n13124), .A2(n15031), .ZN(n13156) );
  OR2_X1 U11568 ( .A1(n16412), .A2(n11152), .ZN(n16398) );
  AND2_X1 U11569 ( .A1(n21993), .A2(n16414), .ZN(n11152) );
  NAND2_X2 U11570 ( .A1(n12114), .A2(n18912), .ZN(n17021) );
  AND2_X2 U11571 ( .A1(n15813), .A2(n15812), .ZN(n15811) );
  OR2_X1 U11572 ( .A1(n16880), .A2(n11153), .ZN(n12778) );
  OR2_X1 U11573 ( .A1(n11343), .A2(n11583), .ZN(n11153) );
  XNOR2_X1 U11575 ( .A(n13218), .B(n13206), .ZN(n13318) );
  OR2_X1 U11576 ( .A1(n16860), .A2(n11583), .ZN(n11155) );
  OR2_X2 U11577 ( .A1(n16880), .A2(n11343), .ZN(n16860) );
  NAND2_X1 U11578 ( .A1(n11283), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11282) );
  AND2_X1 U11579 ( .A1(n11767), .A2(n11780), .ZN(n12689) );
  NAND2_X1 U11580 ( .A1(n11282), .A2(n11802), .ZN(n11156) );
  NAND2_X1 U11581 ( .A1(n11741), .A2(n12474), .ZN(n11727) );
  NAND2_X2 U11582 ( .A1(n11436), .A2(n11435), .ZN(n18216) );
  NOR2_X2 U11583 ( .A1(n14565), .A2(n21604), .ZN(n21809) );
  INV_X1 U11584 ( .A(n19245), .ZN(n11157) );
  INV_X1 U11585 ( .A(n12692), .ZN(n11774) );
  OAI22_X2 U11586 ( .A1(n11867), .A2(n11977), .B1(n11979), .B2(n11866), .ZN(
        n11868) );
  NAND2_X1 U11587 ( .A1(n20544), .A2(n11161), .ZN(n11158) );
  AND2_X1 U11588 ( .A1(n11158), .A2(n11159), .ZN(n15827) );
  OR2_X1 U11589 ( .A1(n11160), .A2(n20551), .ZN(n11159) );
  INV_X1 U11590 ( .A(n13214), .ZN(n11160) );
  AND2_X1 U11591 ( .A1(n13203), .A2(n13214), .ZN(n11161) );
  INV_X1 U11592 ( .A(n17799), .ZN(n11162) );
  OR2_X1 U11593 ( .A1(n14293), .A2(n19178), .ZN(n11387) );
  OAI21_X2 U11594 ( .B1(n16888), .B2(n11308), .A(n11307), .ZN(n16875) );
  NAND2_X2 U11595 ( .A1(n12212), .A2(n12211), .ZN(n16888) );
  AOI21_X2 U11596 ( .B1(n16051), .B2(n16049), .A(n16050), .ZN(n16285) );
  OR2_X2 U11597 ( .A1(n16070), .A2(n11628), .ZN(n16049) );
  NAND2_X2 U11598 ( .A1(n14894), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14893) );
  NOR2_X2 U11599 ( .A1(n12924), .A2(n11640), .ZN(n12964) );
  OR3_X1 U11600 ( .A1(n21371), .A2(n21388), .A3(n14310), .ZN(n11190) );
  AND2_X2 U11601 ( .A1(n11890), .A2(n19225), .ZN(n14278) );
  AND2_X2 U11602 ( .A1(n11890), .A2(n19225), .ZN(n11170) );
  CLKBUF_X1 U11603 ( .A(n11884), .Z(n11180) );
  NOR2_X2 U11604 ( .A1(n15934), .A2(n11620), .ZN(n16123) );
  OAI221_X2 U11605 ( .B1(n14564), .B2(n21358), .C1(n14564), .C2(n21357), .A(
        n21377), .ZN(n21576) );
  INV_X1 U11606 ( .A(n16605), .ZN(n11165) );
  INV_X2 U11607 ( .A(n16605), .ZN(n11166) );
  INV_X1 U11608 ( .A(n11166), .ZN(n11167) );
  AND2_X1 U11609 ( .A1(n12847), .A2(n12849), .ZN(n11168) );
  NAND2_X2 U11610 ( .A1(n11839), .A2(n11838), .ZN(n12269) );
  AND2_X1 U11611 ( .A1(n12848), .A2(n16603), .ZN(n11169) );
  AND2_X2 U11612 ( .A1(n12722), .A2(n11795), .ZN(n12732) );
  AND2_X1 U11613 ( .A1(n11789), .A2(n11788), .ZN(n11790) );
  AND2_X1 U11614 ( .A1(n12847), .A2(n12841), .ZN(n11171) );
  AND2_X1 U11615 ( .A1(n12847), .A2(n12841), .ZN(n12894) );
  AND3_X4 U11616 ( .A1(n19225), .A2(n11298), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11668) );
  AND2_X1 U11617 ( .A1(n12846), .A2(n12847), .ZN(n11172) );
  NOR2_X1 U11618 ( .A1(n12924), .A2(n11640), .ZN(n11173) );
  NAND2_X1 U11619 ( .A1(n11766), .A2(n11764), .ZN(n12260) );
  INV_X1 U11620 ( .A(n11824), .ZN(n11174) );
  INV_X1 U11621 ( .A(n11824), .ZN(n12272) );
  AND2_X4 U11622 ( .A1(n12732), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11824) );
  NOR2_X1 U11623 ( .A1(n16880), .A2(n11342), .ZN(n16850) );
  OR2_X4 U11624 ( .A1(n16894), .A2(n11580), .ZN(n16880) );
  XNOR2_X1 U11625 ( .A(n11478), .B(n11836), .ZN(n11854) );
  AND2_X2 U11626 ( .A1(n11770), .A2(n11769), .ZN(n12720) );
  INV_X1 U11627 ( .A(n11762), .ZN(n11757) );
  AND4_X1 U11628 ( .A1(n11762), .A2(n19758), .A3(n12442), .A4(n11182), .ZN(
        n11726) );
  NOR2_X2 U11629 ( .A1(n16110), .A2(n11613), .ZN(n16084) );
  INV_X2 U11630 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12054) );
  NAND2_X1 U11631 ( .A1(n12482), .A2(n11813), .ZN(n12335) );
  AOI21_X2 U11632 ( .B1(n12422), .B2(n11592), .A(n11590), .ZN(n16840) );
  NAND2_X2 U11633 ( .A1(n11631), .A2(n12231), .ZN(n12422) );
  NOR2_X2 U11634 ( .A1(n21380), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11175) );
  NOR2_X1 U11635 ( .A1(n21380), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14390) );
  OR2_X2 U11636 ( .A1(n12372), .A2(n15432), .ZN(n15430) );
  OAI21_X2 U11637 ( .B1(n14968), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n13008), 
        .ZN(n13062) );
  AND2_X2 U11638 ( .A1(n15437), .A2(n11861), .ZN(n11972) );
  AND2_X1 U11639 ( .A1(n11853), .A2(n15437), .ZN(n19904) );
  NOR2_X2 U11640 ( .A1(n15437), .A2(n11860), .ZN(n19837) );
  NAND2_X2 U11641 ( .A1(n11181), .A2(n11784), .ZN(n12494) );
  NAND2_X2 U11642 ( .A1(n11832), .A2(n11831), .ZN(n11830) );
  XNOR2_X2 U11643 ( .A(n11586), .B(n11587), .ZN(n11832) );
  AOI211_X1 U11644 ( .C1(n11972), .C2(n19933), .A(n19932), .B(n20338), .ZN(
        n19934) );
  OR2_X1 U11645 ( .A1(n11829), .A2(n11828), .ZN(n11851) );
  AND2_X1 U11646 ( .A1(n16907), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17014) );
  NAND3_X2 U11647 ( .A1(n11339), .A2(n11340), .A3(n11341), .ZN(n16907) );
  OR2_X2 U11648 ( .A1(n11872), .A2(n11865), .ZN(n11979) );
  NAND2_X1 U11649 ( .A1(n11681), .A2(n11680), .ZN(n11181) );
  NAND2_X1 U11650 ( .A1(n11681), .A2(n11680), .ZN(n11182) );
  AND2_X4 U11651 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12255) );
  XNOR2_X2 U11652 ( .A(n12269), .B(n12271), .ZN(n11855) );
  AOI21_X2 U11653 ( .B1(n16875), .B2(n11605), .A(n11603), .ZN(n11631) );
  NOR2_X2 U11654 ( .A1(n11860), .A2(n15441), .ZN(n11971) );
  CLKBUF_X3 U11655 ( .A(n11855), .Z(n15441) );
  AND4_X1 U11656 ( .A1(n11762), .A2(n11769), .A3(n19758), .A4(n12717), .ZN(
        n11766) );
  INV_X1 U11657 ( .A(n16036), .ZN(n16029) );
  INV_X1 U11658 ( .A(n12430), .ZN(n12438) );
  NAND2_X1 U11659 ( .A1(n16840), .A2(n16842), .ZN(n12779) );
  NAND2_X1 U11660 ( .A1(n12492), .A2(n18854), .ZN(n12736) );
  INV_X1 U11661 ( .A(n21224), .ZN(n14567) );
  NAND2_X1 U11662 ( .A1(n11757), .A2(n19758), .ZN(n12474) );
  INV_X1 U11663 ( .A(n11763), .ZN(n11764) );
  NAND2_X1 U11664 ( .A1(n14567), .A2(n21337), .ZN(n11434) );
  INV_X1 U11665 ( .A(n16164), .ZN(n11614) );
  NAND2_X1 U11666 ( .A1(n13918), .A2(n14002), .ZN(n13997) );
  NAND2_X1 U11667 ( .A1(n14828), .A2(n16021), .ZN(n14693) );
  INV_X1 U11668 ( .A(n16813), .ZN(n11548) );
  NAND2_X1 U11669 ( .A1(n11512), .A2(n11510), .ZN(n11509) );
  INV_X1 U11670 ( .A(n15561), .ZN(n11510) );
  XNOR2_X1 U11671 ( .A(n12436), .B(n12428), .ZN(n12429) );
  OR2_X1 U11672 ( .A1(n11544), .A2(n11543), .ZN(n11542) );
  INV_X1 U11673 ( .A(n15727), .ZN(n11543) );
  AOI21_X1 U11674 ( .B1(n14812), .B2(n11648), .A(n11556), .ZN(n11555) );
  INV_X1 U11675 ( .A(n14818), .ZN(n11556) );
  NAND2_X1 U11676 ( .A1(n13896), .A2(n19916), .ZN(n12541) );
  NOR2_X1 U11677 ( .A1(n20682), .A2(n15964), .ZN(n17757) );
  NOR2_X1 U11678 ( .A1(n14309), .A2(n14310), .ZN(n14445) );
  NAND3_X1 U11679 ( .A1(n18521), .A2(n11424), .A3(n11423), .ZN(n14426) );
  NOR2_X1 U11680 ( .A1(n18447), .A2(n11425), .ZN(n11424) );
  INV_X1 U11681 ( .A(n18471), .ZN(n11423) );
  NAND2_X1 U11682 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n11426), .ZN(
        n11425) );
  AOI21_X1 U11683 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n21838), .A(
        n14441), .ZN(n14469) );
  AND2_X1 U11684 ( .A1(n16021), .A2(n15229), .ZN(n13918) );
  CLKBUF_X1 U11685 ( .A(n14693), .Z(n16038) );
  AND2_X1 U11686 ( .A1(n14906), .A2(n16042), .ZN(n14923) );
  INV_X1 U11687 ( .A(n22283), .ZN(n16042) );
  NOR2_X1 U11688 ( .A1(n15838), .A2(n11551), .ZN(n11550) );
  INV_X1 U11689 ( .A(n15878), .ZN(n11551) );
  NAND2_X1 U11690 ( .A1(n16742), .A2(n12785), .ZN(n12787) );
  AOI21_X1 U11691 ( .B1(n15817), .B2(n15818), .A(n12538), .ZN(n14814) );
  XNOR2_X1 U11692 ( .A(n13845), .B(n13844), .ZN(n14296) );
  NAND2_X1 U11693 ( .A1(n13885), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13845) );
  NOR2_X1 U11694 ( .A1(n11594), .A2(n11593), .ZN(n11592) );
  INV_X1 U11695 ( .A(n12421), .ZN(n11594) );
  OR2_X1 U11696 ( .A1(n11582), .A2(n11343), .ZN(n11342) );
  INV_X1 U11697 ( .A(n12764), .ZN(n12768) );
  OR2_X1 U11698 ( .A1(n11309), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11307) );
  AND2_X1 U11699 ( .A1(n11309), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11308) );
  NOR2_X1 U11700 ( .A1(n20736), .A2(n20745), .ZN(n20742) );
  NAND2_X1 U11701 ( .A1(n18534), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11421) );
  NAND2_X1 U11702 ( .A1(n19553), .A2(n20741), .ZN(n14565) );
  NAND2_X1 U11703 ( .A1(n19243), .A2(n18854), .ZN(n19290) );
  AOI21_X1 U11704 ( .B1(n19161), .B2(n19202), .A(n11635), .ZN(n12753) );
  NAND2_X1 U11705 ( .A1(n11535), .A2(n11223), .ZN(n11336) );
  NAND2_X1 U11706 ( .A1(n17062), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11535) );
  INV_X1 U11707 ( .A(n12095), .ZN(n11306) );
  INV_X1 U11708 ( .A(n11305), .ZN(n11304) );
  NAND2_X1 U11709 ( .A1(n12038), .A2(n12027), .ZN(n12043) );
  OR2_X1 U11710 ( .A1(n13007), .A2(n13006), .ZN(n13057) );
  AND2_X2 U11711 ( .A1(n12847), .A2(n16603), .ZN(n13185) );
  NOR2_X1 U11712 ( .A1(n12955), .A2(n22274), .ZN(n13066) );
  INV_X1 U11713 ( .A(n13302), .ZN(n13270) );
  NAND2_X1 U11714 ( .A1(n13270), .A2(n13010), .ZN(n13303) );
  NAND2_X1 U11715 ( .A1(n12955), .A2(n16021), .ZN(n13081) );
  NOR2_X1 U11716 ( .A1(n12177), .A2(n11244), .ZN(n11395) );
  AOI21_X1 U11717 ( .B1(n11780), .B2(n20247), .A(n12451), .ZN(n11781) );
  AOI22_X1 U11718 ( .A1(n11188), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11140), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14143) );
  AND2_X1 U11719 ( .A1(n12809), .A2(n12191), .ZN(n12193) );
  NAND2_X1 U11720 ( .A1(n12400), .A2(n12399), .ZN(n12401) );
  NAND2_X1 U11721 ( .A1(n12389), .A2(n12382), .ZN(n12390) );
  NAND2_X1 U11722 ( .A1(n11840), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11777) );
  NOR2_X1 U11723 ( .A1(n11385), .A2(n11384), .ZN(n11383) );
  NAND2_X1 U11724 ( .A1(n11918), .A2(n11219), .ZN(n11385) );
  NAND2_X1 U11725 ( .A1(n16061), .A2(n11629), .ZN(n11628) );
  INV_X1 U11726 ( .A(n16071), .ZN(n11629) );
  NAND2_X1 U11727 ( .A1(n13707), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13716) );
  OR2_X1 U11728 ( .A1(n13716), .A2(n13715), .ZN(n13747) );
  INV_X1 U11729 ( .A(n16110), .ZN(n11615) );
  NAND2_X1 U11730 ( .A1(n14902), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13794) );
  NOR2_X1 U11731 ( .A1(n16259), .A2(n15936), .ZN(n11621) );
  INV_X1 U11732 ( .A(n15934), .ZN(n11622) );
  OR2_X1 U11733 ( .A1(n13911), .A2(n15575), .ZN(n13471) );
  OR2_X1 U11734 ( .A1(n13915), .A2(n15575), .ZN(n13822) );
  AND3_X1 U11735 ( .A1(n11463), .A2(n11465), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13245) );
  AND2_X1 U11736 ( .A1(n11193), .A2(n11452), .ZN(n11445) );
  INV_X1 U11737 ( .A(n13225), .ZN(n11451) );
  OAI21_X1 U11738 ( .B1(n12995), .B2(n12979), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n12980) );
  AND2_X1 U11739 ( .A1(n22670), .A2(n13107), .ZN(n15785) );
  AND2_X1 U11740 ( .A1(n15095), .A2(n13076), .ZN(n15547) );
  OR2_X1 U11741 ( .A1(n15337), .A2(n15248), .ZN(n22428) );
  INV_X1 U11742 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n22374) );
  OR2_X1 U11743 ( .A1(n13303), .A2(n14691), .ZN(n13309) );
  AND2_X1 U11744 ( .A1(n13081), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13286) );
  AND3_X1 U11745 ( .A1(n12480), .A2(n12479), .A3(n12716), .ZN(n12714) );
  NOR2_X1 U11746 ( .A1(n12220), .A2(n11396), .ZN(n12235) );
  NAND2_X1 U11747 ( .A1(n11397), .A2(n12233), .ZN(n11396) );
  AND2_X1 U11748 ( .A1(n12122), .A2(n12131), .ZN(n11388) );
  INV_X1 U11749 ( .A(n12061), .ZN(n11392) );
  NOR2_X1 U11750 ( .A1(n11254), .A2(n11499), .ZN(n11498) );
  INV_X1 U11751 ( .A(n15876), .ZN(n11499) );
  NAND2_X1 U11752 ( .A1(n11743), .A2(n11742), .ZN(n11794) );
  INV_X1 U11753 ( .A(n11741), .ZN(n11743) );
  NAND2_X1 U11754 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11538) );
  INV_X1 U11755 ( .A(n17021), .ZN(n11290) );
  NAND2_X1 U11756 ( .A1(n17022), .A2(n11297), .ZN(n11292) );
  AND2_X1 U11757 ( .A1(n16694), .A2(n12353), .ZN(n11521) );
  AND2_X1 U11758 ( .A1(n16876), .A2(n16877), .ZN(n11601) );
  INV_X1 U11759 ( .A(n11596), .ZN(n11595) );
  OAI21_X1 U11760 ( .B1(n11602), .B2(n11217), .A(n11604), .ZN(n11596) );
  NAND2_X1 U11761 ( .A1(n11608), .A2(n16876), .ZN(n11604) );
  INV_X1 U11762 ( .A(n11598), .ZN(n11597) );
  INV_X1 U11763 ( .A(n11608), .ZN(n11599) );
  INV_X1 U11764 ( .A(n15907), .ZN(n11517) );
  NOR2_X1 U11765 ( .A1(n11373), .A2(n12807), .ZN(n11370) );
  NOR2_X1 U11766 ( .A1(n15897), .A2(n11519), .ZN(n11518) );
  INV_X1 U11767 ( .A(n15832), .ZN(n11519) );
  NAND2_X1 U11768 ( .A1(n11545), .A2(n12626), .ZN(n11544) );
  INV_X1 U11769 ( .A(n15847), .ZN(n11545) );
  INV_X1 U11770 ( .A(n14891), .ZN(n11552) );
  NOR2_X1 U11771 ( .A1(n14210), .A2(n20243), .ZN(n14030) );
  NAND2_X1 U11772 ( .A1(n11229), .A2(n18879), .ZN(n11849) );
  AND2_X2 U11773 ( .A1(n11667), .A2(n11666), .ZN(n11784) );
  NOR2_X1 U11774 ( .A1(n21027), .A2(n21040), .ZN(n11349) );
  NOR2_X1 U11775 ( .A1(n14308), .A2(n21360), .ZN(n14352) );
  NAND2_X1 U11776 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n21371), .ZN(
        n14309) );
  NOR2_X1 U11777 ( .A1(n21383), .A2(n20747), .ZN(n14447) );
  NOR2_X1 U11778 ( .A1(n14307), .A2(n21383), .ZN(n14389) );
  AND2_X1 U11779 ( .A1(n14598), .A2(n11261), .ZN(n11413) );
  NOR2_X1 U11780 ( .A1(n18693), .A2(n14591), .ZN(n14594) );
  NOR2_X1 U11781 ( .A1(n18723), .A2(n14581), .ZN(n14582) );
  NAND2_X1 U11782 ( .A1(n14577), .A2(n21224), .ZN(n11433) );
  NOR2_X1 U11783 ( .A1(n17368), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n14468) );
  NOR2_X1 U11784 ( .A1(n14549), .A2(n21358), .ZN(n15950) );
  NOR2_X1 U11785 ( .A1(n21232), .A2(n19430), .ZN(n17367) );
  INV_X1 U11786 ( .A(n14564), .ZN(n14561) );
  NOR3_X1 U11787 ( .A1(n14555), .A2(n14551), .A3(n14559), .ZN(n21374) );
  INV_X1 U11788 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21827) );
  NAND2_X1 U11789 ( .A1(n11475), .A2(n13922), .ZN(n11476) );
  NAND2_X1 U11790 ( .A1(n14861), .A2(n14860), .ZN(n14931) );
  AND3_X1 U11791 ( .A1(n12948), .A2(n16042), .A3(n16029), .ZN(n15378) );
  INV_X1 U11792 ( .A(n13822), .ZN(n13828) );
  NAND2_X1 U11793 ( .A1(n13772), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13835) );
  NAND2_X1 U11794 ( .A1(n11201), .A2(n16220), .ZN(n11613) );
  AND2_X1 U11795 ( .A1(n13366), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13368) );
  INV_X1 U11796 ( .A(n12989), .ZN(n14838) );
  AND2_X1 U11797 ( .A1(n22004), .A2(n21907), .ZN(n22019) );
  INV_X1 U11798 ( .A(n20525), .ZN(n11455) );
  NOR2_X1 U11799 ( .A1(n15374), .A2(n20525), .ZN(n11456) );
  OR2_X1 U11800 ( .A1(n11458), .A2(n15374), .ZN(n20526) );
  INV_X1 U11801 ( .A(n11457), .ZN(n11458) );
  NOR2_X1 U11802 ( .A1(n15374), .A2(n15373), .ZN(n15397) );
  AND2_X1 U11803 ( .A1(n16439), .A2(n22062), .ZN(n22002) );
  NAND2_X1 U11804 ( .A1(n11476), .A2(n11474), .ZN(n15082) );
  OR2_X1 U11805 ( .A1(n14914), .A2(n15972), .ZN(n11474) );
  CLKBUF_X1 U11806 ( .A(n14968), .Z(n14969) );
  AND2_X1 U11807 ( .A1(n15287), .A2(n14966), .ZN(n15087) );
  NOR2_X1 U11808 ( .A1(n22430), .A2(n15782), .ZN(n22419) );
  INV_X1 U11809 ( .A(n13096), .ZN(n13098) );
  INV_X1 U11810 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n22415) );
  NOR2_X1 U11811 ( .A1(n22412), .A2(n15782), .ZN(n22439) );
  INV_X1 U11812 ( .A(n13338), .ZN(n15568) );
  AND2_X1 U11813 ( .A1(n15452), .A2(n15451), .ZN(n15453) );
  AOI21_X1 U11814 ( .B1(n22415), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n15782), 
        .ZN(n22387) );
  INV_X1 U11815 ( .A(n15124), .ZN(n15782) );
  OR2_X1 U11816 ( .A1(n15228), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n17814) );
  AND2_X1 U11817 ( .A1(n13843), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13885) );
  INV_X1 U11818 ( .A(n12425), .ZN(n12427) );
  NOR2_X1 U11819 ( .A1(n11398), .A2(n12228), .ZN(n11397) );
  INV_X1 U11820 ( .A(n11400), .ZN(n11398) );
  NOR2_X1 U11821 ( .A1(n12219), .A2(n11401), .ZN(n11400) );
  INV_X1 U11822 ( .A(n12223), .ZN(n11401) );
  INV_X1 U11823 ( .A(n12220), .ZN(n11399) );
  NAND2_X1 U11824 ( .A1(n12150), .A2(n11402), .ZN(n12213) );
  NOR2_X1 U11825 ( .A1(n11404), .A2(n12195), .ZN(n11402) );
  AND2_X1 U11826 ( .A1(n12661), .A2(n12660), .ZN(n16813) );
  INV_X1 U11827 ( .A(n15839), .ZN(n11549) );
  NAND2_X1 U11828 ( .A1(n11508), .A2(n12314), .ZN(n11507) );
  INV_X1 U11829 ( .A(n15707), .ZN(n12314) );
  INV_X1 U11830 ( .A(n11509), .ZN(n11508) );
  INV_X1 U11831 ( .A(n15628), .ZN(n11493) );
  AND2_X1 U11832 ( .A1(n11495), .A2(n15360), .ZN(n11494) );
  NAND2_X1 U11833 ( .A1(n11549), .A2(n11255), .ZN(n17133) );
  AND2_X1 U11834 ( .A1(n12540), .A2(n12539), .ZN(n14812) );
  NOR2_X1 U11835 ( .A1(n20060), .A2(n14816), .ZN(n15694) );
  AND2_X1 U11836 ( .A1(n12720), .A2(n19168), .ZN(n14809) );
  NOR2_X1 U11837 ( .A1(n13883), .A2(n19120), .ZN(n13882) );
  OR2_X1 U11838 ( .A1(n13879), .A2(n12773), .ZN(n13883) );
  NOR2_X1 U11839 ( .A1(n11236), .A2(n12359), .ZN(n13847) );
  OR3_X1 U11840 ( .A1(n12202), .A2(n12430), .A3(n12319), .ZN(n16919) );
  OR3_X1 U11841 ( .A1(n13902), .A2(n12430), .A3(n12791), .ZN(n12781) );
  AND2_X1 U11842 ( .A1(n12770), .A2(n11257), .ZN(n16679) );
  AND2_X1 U11843 ( .A1(n12657), .A2(n12656), .ZN(n15838) );
  NAND2_X1 U11844 ( .A1(n15108), .A2(n15695), .ZN(n15839) );
  NOR2_X1 U11845 ( .A1(n12798), .A2(n11381), .ZN(n11380) );
  INV_X1 U11846 ( .A(n17010), .ZN(n11381) );
  NOR2_X1 U11847 ( .A1(n12407), .A2(n11231), .ZN(n11339) );
  AND2_X1 U11848 ( .A1(n11524), .A2(n11523), .ZN(n11522) );
  INV_X1 U11849 ( .A(n15592), .ZN(n11523) );
  AND2_X1 U11850 ( .A1(n12469), .A2(n12478), .ZN(n19235) );
  INV_X1 U11851 ( .A(n12736), .ZN(n12757) );
  NAND2_X1 U11852 ( .A1(n14029), .A2(n14028), .ZN(n14803) );
  AOI22_X1 U11853 ( .A1(n14027), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19932), .B2(n19927), .ZN(n14028) );
  OR2_X1 U11854 ( .A1(n18858), .A2(n19259), .ZN(n14029) );
  XNOR2_X1 U11855 ( .A(n14803), .B(n14030), .ZN(n14881) );
  OAI21_X1 U11856 ( .B1(n17336), .B2(n19259), .A(n14026), .ZN(n14882) );
  NAND2_X1 U11857 ( .A1(n12467), .A2(n12466), .ZN(n19242) );
  NAND2_X1 U11858 ( .A1(n14015), .A2(n11479), .ZN(n14018) );
  NOR2_X1 U11859 ( .A1(n14017), .A2(n11480), .ZN(n11479) );
  INV_X1 U11860 ( .A(n14014), .ZN(n11480) );
  INV_X1 U11862 ( .A(n19914), .ZN(n19896) );
  INV_X1 U11863 ( .A(n11977), .ZN(n19889) );
  BUF_X1 U11864 ( .A(n11970), .Z(n19813) );
  OR2_X1 U11865 ( .A1(n19751), .A2(n19942), .ZN(n19944) );
  INV_X1 U11866 ( .A(n19751), .ZN(n19919) );
  NOR2_X1 U11867 ( .A1(n19820), .A2(n19925), .ZN(n19881) );
  INV_X1 U11868 ( .A(n19942), .ZN(n19932) );
  INV_X1 U11869 ( .A(n19919), .ZN(n20244) );
  NOR2_X1 U11870 ( .A1(n19820), .A2(n19915), .ZN(n19895) );
  NAND2_X1 U11871 ( .A1(n19270), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19259) );
  NOR2_X1 U11872 ( .A1(n21129), .A2(n21128), .ZN(n21144) );
  OAI21_X1 U11873 ( .B1(n21103), .B2(n11353), .A(n11352), .ZN(n21129) );
  NAND2_X1 U11874 ( .A1(n11354), .A2(n21101), .ZN(n11353) );
  NAND2_X1 U11875 ( .A1(n21128), .A2(n11354), .ZN(n11352) );
  INV_X1 U11876 ( .A(n21118), .ZN(n11354) );
  NOR2_X1 U11877 ( .A1(n21102), .A2(n21128), .ZN(n21103) );
  NOR2_X1 U11878 ( .A1(n21103), .A2(n21104), .ZN(n21116) );
  OR2_X1 U11879 ( .A1(n21167), .A2(n11322), .ZN(n11321) );
  AND2_X1 U11880 ( .A1(n21165), .A2(n21166), .ZN(n11322) );
  NOR2_X1 U11881 ( .A1(n20679), .A2(n14565), .ZN(n20682) );
  NOR2_X1 U11882 ( .A1(n21868), .A2(n21817), .ZN(n20681) );
  AND2_X1 U11883 ( .A1(n18561), .A2(n11360), .ZN(n18591) );
  AND2_X1 U11884 ( .A1(n11361), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11360) );
  AND2_X1 U11885 ( .A1(n11644), .A2(n20966), .ZN(n11364) );
  AND2_X1 U11886 ( .A1(n18478), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n18451) );
  NOR2_X1 U11887 ( .A1(n18411), .A2(n20955), .ZN(n20966) );
  NOR2_X1 U11888 ( .A1(n20738), .A2(n21871), .ZN(n14613) );
  AOI21_X2 U11889 ( .B1(n18556), .B2(n21668), .A(n11638), .ZN(n14430) );
  NOR2_X1 U11890 ( .A1(n11421), .A2(n21598), .ZN(n11420) );
  NAND3_X1 U11891 ( .A1(n14421), .A2(n11432), .A3(n21750), .ZN(n18604) );
  INV_X1 U11892 ( .A(n18548), .ZN(n21668) );
  NAND2_X1 U11893 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21876) );
  AND2_X1 U11894 ( .A1(n22104), .A2(n15226), .ZN(n22262) );
  AND2_X1 U11895 ( .A1(n15243), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n15244) );
  XNOR2_X1 U11896 ( .A(n15975), .B(n15974), .ZN(n16429) );
  AND2_X1 U11897 ( .A1(n16465), .A2(n20528), .ZN(n14007) );
  INV_X1 U11898 ( .A(n16265), .ZN(n16252) );
  XNOR2_X1 U11899 ( .A(n16050), .B(n13910), .ZN(n16277) );
  INV_X1 U11900 ( .A(n13909), .ZN(n13910) );
  AND2_X1 U11901 ( .A1(n22019), .A2(n22002), .ZN(n16545) );
  OR2_X1 U11902 ( .A1(n13838), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n22049) );
  AND2_X1 U11903 ( .A1(n14923), .A2(n14911), .ZN(n22053) );
  INV_X1 U11904 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n15570) );
  OR3_X1 U11905 ( .A1(n18852), .A2(n13906), .A3(n13905), .ZN(n19098) );
  AOI21_X1 U11906 ( .B1(n16661), .B2(n11532), .A(n11530), .ZN(n11529) );
  OAI21_X1 U11907 ( .B1(n11531), .B2(n19029), .A(n19029), .ZN(n11530) );
  INV_X1 U11908 ( .A(n11532), .ZN(n11531) );
  NAND2_X1 U11909 ( .A1(n13886), .A2(n16825), .ZN(n19164) );
  AND2_X1 U11910 ( .A1(n11211), .A2(n12221), .ZN(n19078) );
  OR2_X1 U11911 ( .A1(n12785), .A2(n16742), .ZN(n12786) );
  NAND2_X1 U11912 ( .A1(n16666), .A2(n16665), .ZN(n17050) );
  INV_X1 U11913 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n19120) );
  INV_X1 U11914 ( .A(n17850), .ZN(n17883) );
  INV_X1 U11915 ( .A(n17865), .ZN(n17878) );
  OR2_X1 U11916 ( .A1(n19290), .A2(n14673), .ZN(n17859) );
  NAND2_X1 U11917 ( .A1(n19290), .A2(n12356), .ZN(n17029) );
  XNOR2_X1 U11918 ( .A(n12441), .B(n12440), .ZN(n14293) );
  AOI21_X1 U11919 ( .B1(n16850), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16834) );
  OAI211_X1 U11920 ( .C1(n16846), .C2(n11287), .A(n11286), .B(n11285), .ZN(
        n17053) );
  NAND2_X1 U11921 ( .A1(n16847), .A2(n11288), .ZN(n11287) );
  OAI21_X1 U11922 ( .B1(n16847), .B2(n12247), .A(n11284), .ZN(n11286) );
  OAI21_X1 U11923 ( .B1(n12769), .B2(n12768), .A(n12767), .ZN(n17074) );
  AND2_X1 U11924 ( .A1(n12422), .A2(n12766), .ZN(n12767) );
  NOR2_X1 U11925 ( .A1(n12736), .A2(n12733), .ZN(n17174) );
  INV_X1 U11926 ( .A(n19178), .ZN(n19211) );
  INV_X1 U11927 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19833) );
  INV_X1 U11928 ( .A(n19915), .ZN(n19925) );
  NAND2_X1 U11929 ( .A1(n19833), .A2(n19916), .ZN(n19942) );
  INV_X1 U11930 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19916) );
  NAND2_X1 U11931 ( .A1(n20681), .A2(n21807), .ZN(n20745) );
  OAI22_X1 U11932 ( .A1(n21133), .A2(P3_EBX_REG_30__SCAN_IN), .B1(n21132), 
        .B2(n21131), .ZN(n21137) );
  NOR2_X1 U11933 ( .A1(n14529), .A2(n11324), .ZN(n11323) );
  NAND2_X1 U11934 ( .A1(n21296), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n21295) );
  INV_X1 U11935 ( .A(n21306), .ZN(n21312) );
  NAND2_X1 U11936 ( .A1(n11319), .A2(n11317), .ZN(n21326) );
  NOR2_X1 U11937 ( .A1(n21230), .A2(n11318), .ZN(n11317) );
  INV_X1 U11938 ( .A(n21332), .ZN(n11319) );
  AND3_X1 U11939 ( .A1(n14383), .A2(n14382), .A3(n14381), .ZN(n21653) );
  NAND2_X1 U11940 ( .A1(n21267), .A2(n21196), .ZN(n21333) );
  NOR2_X1 U11941 ( .A1(n21171), .A2(n21344), .ZN(n21338) );
  INV_X1 U11942 ( .A(n21338), .ZN(n21349) );
  XNOR2_X1 U11943 ( .A(n11409), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14629) );
  NAND2_X1 U11944 ( .A1(n21626), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11409) );
  INV_X1 U11945 ( .A(n18758), .ZN(n18748) );
  NAND2_X1 U11946 ( .A1(n11408), .A2(n11405), .ZN(n14608) );
  NAND2_X1 U11947 ( .A1(n14629), .A2(n21656), .ZN(n11408) );
  INV_X1 U11948 ( .A(n11406), .ZN(n11405) );
  OAI21_X1 U11949 ( .B1(n14614), .B2(n21731), .A(n11407), .ZN(n11406) );
  NOR2_X2 U11950 ( .A1(n21653), .A2(n21489), .ZN(n21801) );
  NAND2_X1 U11951 ( .A1(n11142), .A2(n21693), .ZN(n21680) );
  AOI21_X1 U11952 ( .B1(n14542), .B2(n14541), .A(n21868), .ZN(n21739) );
  OR3_X1 U11953 ( .A1(n14565), .A2(n21808), .A3(n14548), .ZN(n14541) );
  NAND2_X1 U11954 ( .A1(n21793), .A2(n21809), .ZN(n21489) );
  NAND2_X1 U11955 ( .A1(n11794), .A2(n12719), .ZN(n11806) );
  NOR2_X1 U11956 ( .A1(n11303), .A2(n12096), .ZN(n11302) );
  NAND2_X1 U11957 ( .A1(n11917), .A2(n11919), .ZN(n11384) );
  CLKBUF_X1 U11958 ( .A(n13433), .Z(n13802) );
  INV_X1 U11959 ( .A(n13286), .ZN(n13283) );
  OR2_X1 U11960 ( .A1(n13024), .A2(n13023), .ZN(n13031) );
  INV_X1 U11961 ( .A(n12971), .ZN(n12951) );
  OR2_X1 U11962 ( .A1(n13093), .A2(n13092), .ZN(n13100) );
  NOR2_X1 U11963 ( .A1(n11651), .A2(n11652), .ZN(n12915) );
  OR2_X1 U11964 ( .A1(n13121), .A2(n13120), .ZN(n13148) );
  NAND2_X1 U11965 ( .A1(n13046), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13302) );
  MUX2_X1 U11966 ( .A(n12044), .B(n12443), .S(n13906), .Z(n12261) );
  AOI21_X1 U11967 ( .B1(n11187), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A(
        n11271), .ZN(n14227) );
  AOI21_X1 U11968 ( .B1(n11188), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A(
        n11270), .ZN(n14221) );
  INV_X1 U11969 ( .A(n16705), .ZN(n11489) );
  AOI21_X1 U11970 ( .B1(n11188), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A(
        n11269), .ZN(n14207) );
  AOI21_X1 U11971 ( .B1(n11186), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A(
        n11268), .ZN(n14201) );
  AOI22_X1 U11972 ( .A1(n11186), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11140), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14186) );
  AOI22_X1 U11973 ( .A1(n11187), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11180), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14180) );
  AOI22_X1 U11974 ( .A1(n11187), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11140), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14168) );
  AOI22_X1 U11975 ( .A1(n11188), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11180), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14162) );
  NAND2_X1 U11976 ( .A1(n11772), .A2(n11762), .ZN(n11741) );
  INV_X1 U11977 ( .A(n16877), .ZN(n11607) );
  NOR2_X1 U11978 ( .A1(n11793), .A2(n11771), .ZN(n11813) );
  AND2_X1 U11979 ( .A1(n12194), .A2(n17873), .ZN(n11301) );
  NOR2_X1 U11980 ( .A1(n11394), .A2(n12143), .ZN(n11393) );
  INV_X1 U11981 ( .A(n12169), .ZN(n12143) );
  INV_X1 U11982 ( .A(n11395), .ZN(n11394) );
  OAI22_X1 U11983 ( .A1(n11935), .A2(n11977), .B1(n11979), .B2(n11934), .ZN(
        n11938) );
  INV_X1 U11984 ( .A(n11575), .ZN(n11573) );
  AOI21_X1 U11985 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19809), .A(
        n12029), .ZN(n12249) );
  NOR2_X1 U11986 ( .A1(n12028), .A2(n12042), .ZN(n12029) );
  AND2_X1 U11987 ( .A1(n19927), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12250) );
  INV_X1 U11988 ( .A(n11427), .ZN(n11426) );
  AOI21_X1 U11989 ( .B1(n21337), .B2(n14573), .A(n14567), .ZN(n14572) );
  NAND2_X1 U11990 ( .A1(n11311), .A2(n11313), .ZN(n11312) );
  AND2_X1 U11991 ( .A1(n14692), .A2(n14691), .ZN(n16028) );
  NAND2_X1 U11992 ( .A1(n11626), .A2(n11627), .ZN(n11625) );
  INV_X1 U11993 ( .A(n11628), .ZN(n11627) );
  INV_X1 U11994 ( .A(n16051), .ZN(n11626) );
  INV_X1 U11995 ( .A(n16112), .ZN(n11616) );
  AND2_X1 U11996 ( .A1(n13579), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13580) );
  NOR2_X1 U11997 ( .A1(n13545), .A2(n13544), .ZN(n13579) );
  INV_X1 U11998 ( .A(n13827), .ZN(n13539) );
  INV_X1 U11999 ( .A(n16062), .ZN(n11467) );
  NOR2_X1 U12000 ( .A1(n16073), .A2(n11469), .ZN(n11468) );
  INV_X1 U12001 ( .A(n16082), .ZN(n11469) );
  NOR2_X1 U12002 ( .A1(n16127), .A2(n11473), .ZN(n11472) );
  INV_X1 U12003 ( .A(n16176), .ZN(n11473) );
  NAND2_X1 U12004 ( .A1(n13947), .A2(n11462), .ZN(n11461) );
  INV_X1 U12005 ( .A(n15888), .ZN(n11462) );
  AND2_X1 U12006 ( .A1(n11453), .A2(n15396), .ZN(n11457) );
  INV_X1 U12007 ( .A(n15373), .ZN(n11453) );
  AND2_X1 U12008 ( .A1(n15146), .A2(n12962), .ZN(n13101) );
  INV_X1 U12009 ( .A(n13031), .ZN(n13052) );
  NOR2_X1 U12010 ( .A1(n11437), .A2(n12957), .ZN(n14686) );
  NAND2_X1 U12011 ( .A1(n12956), .A2(n12964), .ZN(n12957) );
  INV_X1 U12012 ( .A(n14833), .ZN(n12956) );
  OR2_X1 U12013 ( .A1(n12984), .A2(n13071), .ZN(n13072) );
  NAND2_X1 U12014 ( .A1(n13078), .A2(n13077), .ZN(n13079) );
  AOI21_X1 U12015 ( .B1(n14960), .B2(n22273), .A(n22277), .ZN(n15099) );
  NOR2_X1 U12016 ( .A1(n19076), .A2(n11568), .ZN(n11567) );
  INV_X1 U12017 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11568) );
  NAND2_X1 U12018 ( .A1(n12145), .A2(n11637), .ZN(n12162) );
  INV_X1 U12019 ( .A(n12174), .ZN(n12145) );
  NAND2_X1 U12020 ( .A1(n12142), .A2(n11395), .ZN(n12172) );
  INV_X1 U12021 ( .A(n12135), .ZN(n12133) );
  NAND2_X1 U12022 ( .A1(n11382), .A2(n12447), .ZN(n12041) );
  NAND2_X1 U12023 ( .A1(n12040), .A2(n12451), .ZN(n11382) );
  AOI21_X1 U12024 ( .B1(n14277), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n11279), .ZN(n14280) );
  AOI22_X1 U12025 ( .A1(n11186), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11180), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14265) );
  AOI21_X1 U12026 ( .B1(n14277), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n11278), .ZN(n14259) );
  AOI21_X1 U12027 ( .B1(n11186), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A(
        n11273), .ZN(n14247) );
  AOI21_X1 U12028 ( .B1(n11187), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n11272), .ZN(n14241) );
  INV_X1 U12029 ( .A(n16718), .ZN(n11491) );
  AOI22_X1 U12030 ( .A1(n11180), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_7__0__SCAN_IN), .B2(n11170), .ZN(n14149) );
  INV_X1 U12031 ( .A(n16735), .ZN(n11492) );
  INV_X1 U12032 ( .A(n15834), .ZN(n11500) );
  NOR2_X1 U12033 ( .A1(n11502), .A2(n15709), .ZN(n11501) );
  INV_X1 U12034 ( .A(n15693), .ZN(n11502) );
  NAND2_X1 U12035 ( .A1(n14016), .A2(n19970), .ZN(n14210) );
  AND2_X1 U12036 ( .A1(n13896), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14016) );
  NOR2_X1 U12037 ( .A1(n16965), .A2(n11564), .ZN(n11563) );
  INV_X1 U12038 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11564) );
  INV_X1 U12039 ( .A(n15625), .ZN(n11513) );
  INV_X1 U12040 ( .A(n15009), .ZN(n12287) );
  NOR2_X1 U12041 ( .A1(n13853), .A2(n11571), .ZN(n11570) );
  INV_X1 U12042 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11571) );
  NOR2_X1 U12043 ( .A1(n12061), .A2(n12052), .ZN(n12066) );
  NAND2_X1 U12044 ( .A1(n11390), .A2(n11389), .ZN(n12421) );
  NAND2_X1 U12045 ( .A1(n17058), .A2(n12420), .ZN(n11389) );
  INV_X1 U12046 ( .A(n16680), .ZN(n11520) );
  NAND2_X1 U12047 ( .A1(n11559), .A2(n16767), .ZN(n11558) );
  NOR2_X1 U12048 ( .A1(n16796), .A2(n11557), .ZN(n16663) );
  OR3_X1 U12049 ( .A1(n16777), .A2(n11558), .A3(n16757), .ZN(n11557) );
  NAND2_X1 U12050 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11343) );
  NAND2_X1 U12051 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11584) );
  NOR3_X1 U12052 ( .A1(n16796), .A2(n16777), .A3(n16786), .ZN(n16776) );
  NOR2_X1 U12053 ( .A1(n12805), .A2(n11377), .ZN(n11376) );
  AND2_X1 U12054 ( .A1(n12804), .A2(n16920), .ZN(n11377) );
  NOR2_X1 U12055 ( .A1(n11371), .A2(n12807), .ZN(n11369) );
  NAND2_X1 U12056 ( .A1(n16922), .A2(n11374), .ZN(n11373) );
  AND2_X1 U12057 ( .A1(n11378), .A2(n16920), .ZN(n11374) );
  AND2_X1 U12058 ( .A1(n15430), .A2(n12374), .ZN(n12376) );
  INV_X1 U12059 ( .A(n14989), .ZN(n11504) );
  NAND2_X1 U12060 ( .A1(n11830), .A2(n11820), .ZN(n11478) );
  NAND2_X1 U12061 ( .A1(n11586), .A2(n11585), .ZN(n11820) );
  INV_X1 U12062 ( .A(n11587), .ZN(n11585) );
  INV_X1 U12063 ( .A(n12040), .ZN(n12511) );
  NAND2_X1 U12064 ( .A1(n13887), .A2(n12471), .ZN(n12692) );
  AND2_X1 U12065 ( .A1(n11528), .A2(n15409), .ZN(n11524) );
  AND3_X1 U12066 ( .A1(n11790), .A2(n11791), .A3(n12725), .ZN(n12690) );
  AND2_X1 U12067 ( .A1(n11772), .A2(n15697), .ZN(n11773) );
  OAI21_X1 U12068 ( .B1(n16014), .B2(n19259), .A(n14022), .ZN(n14024) );
  NOR2_X1 U12069 ( .A1(n14210), .A2(n20194), .ZN(n14023) );
  NAND2_X1 U12070 ( .A1(n14024), .A2(n14023), .ZN(n14031) );
  NAND2_X1 U12071 ( .A1(n11717), .A2(n11716), .ZN(n11724) );
  NAND2_X1 U12072 ( .A1(n11722), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11723) );
  AND2_X1 U12073 ( .A1(n11699), .A2(n11698), .ZN(n11327) );
  NOR2_X1 U12074 ( .A1(n22321), .A2(n22332), .ZN(n19247) );
  NOR2_X1 U12075 ( .A1(n17368), .A2(n21388), .ZN(n11419) );
  NOR2_X1 U12076 ( .A1(n21388), .A2(n21371), .ZN(n11435) );
  INV_X1 U12077 ( .A(n20747), .ZN(n11436) );
  NOR2_X1 U12078 ( .A1(n11363), .A2(n11362), .ZN(n11361) );
  INV_X1 U12079 ( .A(n18531), .ZN(n11363) );
  INV_X1 U12080 ( .A(n14422), .ZN(n18445) );
  NAND2_X1 U12081 ( .A1(n18604), .A2(n21668), .ZN(n14422) );
  NOR2_X1 U12082 ( .A1(n18700), .A2(n14587), .ZN(n14589) );
  NAND2_X1 U12083 ( .A1(n18707), .A2(n14409), .ZN(n14412) );
  NAND2_X1 U12084 ( .A1(n18737), .A2(n14405), .ZN(n14406) );
  INV_X1 U12085 ( .A(n14403), .ZN(n14404) );
  INV_X1 U12086 ( .A(n11434), .ZN(n14574) );
  NOR2_X1 U12087 ( .A1(n14562), .A2(n21359), .ZN(n15951) );
  AND2_X1 U12088 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n21376) );
  NOR2_X1 U12089 ( .A1(n17757), .A2(n15965), .ZN(n21167) );
  CLKBUF_X1 U12090 ( .A(n12967), .Z(n16037) );
  NAND2_X1 U12091 ( .A1(n15225), .A2(n15224), .ZN(n22104) );
  AOI211_X1 U12092 ( .C1(P1_STATE2_REG_0__SCAN_IN), .C2(n15222), .A(n22052), 
        .B(n21874), .ZN(n15225) );
  AND2_X1 U12093 ( .A1(n14871), .A2(n13918), .ZN(n16030) );
  NOR2_X1 U12094 ( .A1(n16192), .A2(n14937), .ZN(n14938) );
  AND2_X1 U12095 ( .A1(n15065), .A2(n16040), .ZN(n20414) );
  NAND2_X1 U12096 ( .A1(n15535), .A2(n15064), .ZN(n15065) );
  AND2_X1 U12097 ( .A1(n11624), .A2(n13909), .ZN(n11623) );
  INV_X1 U12098 ( .A(n11625), .ZN(n11624) );
  NAND2_X1 U12099 ( .A1(n13748), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13750) );
  OR2_X1 U12100 ( .A1(n16303), .A2(n13668), .ZN(n13752) );
  NAND2_X1 U12101 ( .A1(n13664), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13666) );
  NAND2_X1 U12102 ( .A1(n13618), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13619) );
  NOR2_X1 U12103 ( .A1(n13619), .A2(n22212), .ZN(n13664) );
  NAND2_X1 U12104 ( .A1(n11615), .A2(n11239), .ZN(n16163) );
  AND2_X1 U12105 ( .A1(n13586), .A2(n13585), .ZN(n16240) );
  NAND2_X1 U12106 ( .A1(n13528), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13545) );
  NOR2_X1 U12107 ( .A1(n13511), .A2(n22161), .ZN(n13528) );
  NAND2_X1 U12108 ( .A1(n16174), .A2(n11621), .ZN(n11620) );
  NAND2_X1 U12109 ( .A1(n13494), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13511) );
  INV_X1 U12110 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n22161) );
  AND2_X1 U12111 ( .A1(n13478), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13494) );
  NAND2_X1 U12112 ( .A1(n11622), .A2(n13493), .ZN(n16260) );
  AND2_X1 U12113 ( .A1(n13423), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13424) );
  NOR2_X1 U12114 ( .A1(n13407), .A2(n15869), .ZN(n13423) );
  AND2_X1 U12115 ( .A1(n11260), .A2(n15885), .ZN(n11618) );
  NAND2_X1 U12116 ( .A1(n13392), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13407) );
  AND4_X1 U12117 ( .A1(n13391), .A2(n13390), .A3(n13389), .A4(n13388), .ZN(
        n15704) );
  AOI21_X1 U12118 ( .B1(n13372), .B2(n13503), .A(n13371), .ZN(n15557) );
  NOR2_X1 U12119 ( .A1(n13359), .A2(n13313), .ZN(n13366) );
  AND2_X1 U12120 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13320) );
  NAND2_X1 U12121 ( .A1(n13319), .A2(n13503), .ZN(n13325) );
  INV_X1 U12122 ( .A(n16271), .ZN(n11439) );
  NAND2_X1 U12123 ( .A1(n16104), .A2(n11466), .ZN(n16052) );
  AND2_X1 U12124 ( .A1(n11206), .A2(n16053), .ZN(n11466) );
  NAND2_X1 U12125 ( .A1(n16104), .A2(n11468), .ZN(n16075) );
  AND2_X1 U12126 ( .A1(n16156), .A2(n16106), .ZN(n16104) );
  AND2_X1 U12127 ( .A1(n13989), .A2(n13988), .ZN(n16155) );
  NOR2_X1 U12128 ( .A1(n16527), .A2(n16155), .ZN(n16156) );
  OR2_X1 U12129 ( .A1(n16525), .A2(n16524), .ZN(n16527) );
  NAND2_X1 U12130 ( .A1(n16560), .A2(n16161), .ZN(n16525) );
  NAND2_X1 U12131 ( .A1(n11446), .A2(n11443), .ZN(n16343) );
  NOR2_X1 U12132 ( .A1(n20578), .A2(n11281), .ZN(n11444) );
  AND2_X1 U12133 ( .A1(n13982), .A2(n13981), .ZN(n16558) );
  AND2_X1 U12134 ( .A1(n16115), .A2(n16558), .ZN(n16560) );
  AND2_X1 U12135 ( .A1(n20522), .A2(n16117), .ZN(n16115) );
  NOR2_X1 U12136 ( .A1(n20520), .A2(n20519), .ZN(n20522) );
  NAND2_X1 U12137 ( .A1(n11448), .A2(n11193), .ZN(n11447) );
  NAND2_X1 U12138 ( .A1(n11450), .A2(n16411), .ZN(n11449) );
  AND2_X1 U12139 ( .A1(n13972), .A2(n13971), .ZN(n16168) );
  NAND2_X1 U12140 ( .A1(n20509), .A2(n11470), .ZN(n20520) );
  AND2_X1 U12141 ( .A1(n11472), .A2(n11471), .ZN(n11470) );
  INV_X1 U12142 ( .A(n16168), .ZN(n11471) );
  NAND2_X1 U12143 ( .A1(n20509), .A2(n11472), .ZN(n16169) );
  NAND2_X1 U12144 ( .A1(n20509), .A2(n16176), .ZN(n16178) );
  AND2_X1 U12145 ( .A1(n20507), .A2(n20506), .ZN(n20509) );
  AND2_X1 U12146 ( .A1(n13962), .A2(n13961), .ZN(n15939) );
  NOR2_X1 U12147 ( .A1(n16139), .A2(n15939), .ZN(n20507) );
  NAND2_X1 U12148 ( .A1(n16188), .A2(n15948), .ZN(n16137) );
  OR2_X1 U12149 ( .A1(n16137), .A2(n16136), .ZN(n16139) );
  NOR2_X1 U12150 ( .A1(n15866), .A2(n11459), .ZN(n16188) );
  OR2_X1 U12151 ( .A1(n11461), .A2(n13952), .ZN(n11459) );
  NOR2_X1 U12152 ( .A1(n15866), .A2(n11461), .ZN(n16186) );
  NAND2_X1 U12153 ( .A1(n11460), .A2(n13947), .ZN(n15889) );
  INV_X1 U12154 ( .A(n15866), .ZN(n11460) );
  AND2_X1 U12155 ( .A1(n21888), .A2(n21892), .ZN(n22004) );
  INV_X1 U12156 ( .A(n22004), .ZN(n21909) );
  INV_X1 U12157 ( .A(n22007), .ZN(n21907) );
  NAND2_X1 U12158 ( .A1(n13930), .A2(n13929), .ZN(n15374) );
  NAND2_X1 U12159 ( .A1(n13936), .A2(n14002), .ZN(n15973) );
  INV_X1 U12160 ( .A(n13028), .ZN(n13029) );
  NAND2_X1 U12161 ( .A1(n13111), .A2(n13110), .ZN(n15092) );
  INV_X1 U12162 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14866) );
  INV_X1 U12163 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16595) );
  AND2_X1 U12164 ( .A1(n16032), .A2(n15229), .ZN(n16613) );
  NAND2_X1 U12165 ( .A1(n15030), .A2(n14999), .ZN(n22370) );
  AND2_X1 U12166 ( .A1(n15287), .A2(n15451), .ZN(n15291) );
  OR2_X1 U12167 ( .A1(n15030), .A2(n15333), .ZN(n15572) );
  INV_X2 U12168 ( .A(n12963), .ZN(n15379) );
  INV_X1 U12169 ( .A(n12962), .ZN(n15167) );
  NAND2_X1 U12170 ( .A1(n15987), .A2(n20555), .ZN(n15161) );
  OR3_X1 U12171 ( .A1(n22435), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n15099), 
        .ZN(n15168) );
  NAND2_X1 U12172 ( .A1(n13311), .A2(n13310), .ZN(n16036) );
  NAND2_X1 U12173 ( .A1(n13286), .A2(n13269), .ZN(n13311) );
  NAND2_X1 U12174 ( .A1(n13309), .A2(n13308), .ZN(n13310) );
  AND2_X1 U12175 ( .A1(n16023), .A2(n13047), .ZN(n12906) );
  NAND2_X1 U12176 ( .A1(n12714), .A2(n12713), .ZN(n19241) );
  AOI21_X1 U12177 ( .B1(n19029), .B2(n11533), .A(n16836), .ZN(n11532) );
  INV_X1 U12178 ( .A(n16660), .ZN(n11533) );
  NAND2_X1 U12179 ( .A1(n12243), .A2(n12242), .ZN(n12425) );
  NAND2_X1 U12180 ( .A1(n12150), .A2(n11403), .ZN(n12196) );
  NAND2_X1 U12181 ( .A1(n12150), .A2(n12151), .ZN(n12155) );
  NOR2_X1 U12182 ( .A1(n13870), .A2(n12358), .ZN(n13872) );
  OR2_X1 U12183 ( .A1(n19248), .A2(n19287), .ZN(n14659) );
  AND2_X1 U12184 ( .A1(n14037), .A2(n11496), .ZN(n11495) );
  INV_X1 U12185 ( .A(n15405), .ZN(n11496) );
  AND2_X1 U12186 ( .A1(n16662), .A2(n16744), .ZN(n16742) );
  AOI21_X1 U12187 ( .B1(n14277), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A(
        n11280), .ZN(n14272) );
  AND2_X1 U12188 ( .A1(n12663), .A2(n12662), .ZN(n17132) );
  NOR2_X1 U12189 ( .A1(n15839), .A2(n11546), .ZN(n17135) );
  NAND2_X1 U12190 ( .A1(n11255), .A2(n11547), .ZN(n11546) );
  INV_X1 U12191 ( .A(n17132), .ZN(n11547) );
  AND2_X1 U12192 ( .A1(n11786), .A2(n19758), .ZN(n15697) );
  OR2_X1 U12193 ( .A1(n14067), .A2(n14066), .ZN(n15876) );
  NAND2_X1 U12194 ( .A1(n14983), .A2(n14034), .ZN(n14976) );
  AND2_X1 U12195 ( .A1(n14790), .A2(n14789), .ZN(n17918) );
  NOR2_X1 U12196 ( .A1(n14659), .A2(n13887), .ZN(n14675) );
  NAND2_X1 U12197 ( .A1(n13847), .A2(n11566), .ZN(n13879) );
  AND2_X1 U12198 ( .A1(n11205), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11566) );
  NAND2_X1 U12199 ( .A1(n13847), .A2(n11205), .ZN(n13881) );
  NAND2_X1 U12200 ( .A1(n13847), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13877) );
  OR2_X1 U12201 ( .A1(n11538), .A2(n11537), .ZN(n11536) );
  INV_X1 U12202 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11537) );
  NOR3_X1 U12203 ( .A1(n13870), .A2(n11539), .A3(n11538), .ZN(n13875) );
  NAND2_X1 U12204 ( .A1(n13871), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13870) );
  AND2_X1 U12205 ( .A1(n13864), .A2(n11560), .ZN(n13871) );
  NOR2_X1 U12206 ( .A1(n11565), .A2(n11562), .ZN(n11560) );
  INV_X1 U12207 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11565) );
  NAND2_X1 U12208 ( .A1(n13864), .A2(n11563), .ZN(n13868) );
  AND2_X1 U12209 ( .A1(n13850), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13864) );
  NAND2_X1 U12210 ( .A1(n13864), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13866) );
  INV_X1 U12211 ( .A(n15041), .ZN(n12298) );
  NOR2_X1 U12212 ( .A1(n13859), .A2(n18933), .ZN(n13861) );
  NAND3_X1 U12213 ( .A1(n11569), .A2(n11200), .A3(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13859) );
  NAND2_X1 U12214 ( .A1(n11296), .A2(n15811), .ZN(n11295) );
  NAND2_X1 U12215 ( .A1(n15735), .A2(n12438), .ZN(n17875) );
  AND2_X1 U12216 ( .A1(n11569), .A2(n11200), .ZN(n13860) );
  NAND2_X1 U12217 ( .A1(n11569), .A2(n11570), .ZN(n13857) );
  INV_X1 U12218 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n13853) );
  NOR2_X1 U12219 ( .A1(n13855), .A2(n13853), .ZN(n13858) );
  NAND2_X1 U12220 ( .A1(n13856), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13855) );
  INV_X1 U12221 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n15433) );
  NOR2_X1 U12222 ( .A1(n13854), .A2(n15433), .ZN(n13856) );
  NOR2_X1 U12223 ( .A1(n12434), .A2(n12433), .ZN(n12435) );
  INV_X1 U12224 ( .A(n12781), .ZN(n12434) );
  INV_X1 U12225 ( .A(n12247), .ZN(n11288) );
  NAND2_X1 U12226 ( .A1(n11595), .A2(n11600), .ZN(n11603) );
  NAND2_X1 U12227 ( .A1(n11601), .A2(n16869), .ZN(n11600) );
  NAND2_X1 U12228 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11581) );
  AND2_X1 U12229 ( .A1(n11242), .A2(n16736), .ZN(n11516) );
  AND2_X1 U12230 ( .A1(n15713), .A2(n11242), .ZN(n16737) );
  NAND2_X1 U12231 ( .A1(n11375), .A2(n16920), .ZN(n16901) );
  NAND2_X1 U12232 ( .A1(n15713), .A2(n11518), .ZN(n15908) );
  OR2_X1 U12233 ( .A1(n11542), .A2(n11541), .ZN(n11540) );
  INV_X1 U12234 ( .A(n15110), .ZN(n11541) );
  AND3_X1 U12235 ( .A1(n12625), .A2(n12624), .A3(n12623), .ZN(n15039) );
  NOR2_X1 U12236 ( .A1(n15404), .A2(n15356), .ZN(n15626) );
  AND2_X1 U12237 ( .A1(n16989), .A2(n12184), .ZN(n16976) );
  NAND2_X1 U12238 ( .A1(n17012), .A2(n11379), .ZN(n16977) );
  AND2_X1 U12239 ( .A1(n11380), .A2(n16990), .ZN(n11379) );
  NAND2_X1 U12240 ( .A1(n17014), .A2(n17242), .ZN(n16987) );
  AND3_X1 U12241 ( .A1(n12585), .A2(n12584), .A3(n12583), .ZN(n15768) );
  AND3_X1 U12242 ( .A1(n12555), .A2(n12554), .A3(n12553), .ZN(n14891) );
  AND2_X1 U12243 ( .A1(n11553), .A2(n11197), .ZN(n14926) );
  NAND2_X1 U12244 ( .A1(n12385), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15814) );
  AND3_X1 U12245 ( .A1(n12529), .A2(n12528), .A3(n12527), .ZN(n15592) );
  NOR2_X1 U12246 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14661), .ZN(n17016) );
  INV_X1 U12247 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n15820) );
  CLKBUF_X1 U12248 ( .A(n11771), .Z(n14673) );
  AND2_X1 U12249 ( .A1(n12720), .A2(n12451), .ZN(n11795) );
  INV_X1 U12250 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n16001) );
  CLKBUF_X1 U12251 ( .A(n12692), .Z(n19245) );
  XNOR2_X1 U12252 ( .A(n12510), .B(n12504), .ZN(n15015) );
  INV_X1 U12253 ( .A(n12519), .ZN(n11528) );
  INV_X1 U12254 ( .A(n15203), .ZN(n11526) );
  OAI21_X1 U12255 ( .B1(n14024), .B2(n14023), .A(n14031), .ZN(n14889) );
  OAI22_X1 U12256 ( .A1(n14882), .A2(n14881), .B1(n14030), .B2(n14803), .ZN(
        n14888) );
  NOR2_X1 U12257 ( .A1(n19914), .A2(n19913), .ZN(n19929) );
  AND2_X1 U12258 ( .A1(n19880), .A2(n17899), .ZN(n19866) );
  INV_X1 U12259 ( .A(n11978), .ZN(n19794) );
  AND2_X1 U12260 ( .A1(n14013), .A2(n19755), .ZN(n19786) );
  INV_X1 U12261 ( .A(n11980), .ZN(n19778) );
  NAND3_X1 U12262 ( .A1(n15700), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19902), 
        .ZN(n19765) );
  NAND3_X1 U12263 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19752), .A3(n19902), 
        .ZN(n19764) );
  NAND2_X1 U12264 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19919), .ZN(n20154) );
  INV_X1 U12265 ( .A(n19765), .ZN(n20250) );
  INV_X1 U12266 ( .A(n19764), .ZN(n20251) );
  INV_X1 U12267 ( .A(n20154), .ZN(n20246) );
  NAND2_X1 U12268 ( .A1(n21128), .A2(n21080), .ZN(n11355) );
  NOR2_X1 U12269 ( .A1(n21083), .A2(n21062), .ZN(n11357) );
  NAND2_X1 U12270 ( .A1(n21128), .A2(n11347), .ZN(n11346) );
  INV_X1 U12271 ( .A(n21040), .ZN(n11347) );
  NOR2_X1 U12272 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n20807), .ZN(n20826) );
  AOI22_X1 U12273 ( .A1(n11145), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14531) );
  AOI22_X1 U12274 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18288), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14530) );
  NAND2_X1 U12275 ( .A1(n18130), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11325) );
  INV_X1 U12276 ( .A(n17367), .ZN(n21171) );
  INV_X1 U12277 ( .A(n18806), .ZN(n18808) );
  NOR2_X1 U12278 ( .A1(n20680), .A2(n21846), .ZN(n20683) );
  AND2_X1 U12279 ( .A1(n11202), .A2(n11251), .ZN(n11344) );
  NAND2_X1 U12280 ( .A1(n18561), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n18560) );
  NAND2_X1 U12281 ( .A1(n18451), .A2(n11199), .ZN(n18485) );
  NAND2_X1 U12282 ( .A1(n11314), .A2(n19551), .ZN(n18549) );
  NAND2_X1 U12283 ( .A1(n18562), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11314) );
  NAND2_X1 U12284 ( .A1(n18399), .A2(n11364), .ZN(n18601) );
  INV_X1 U12285 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18411) );
  INV_X1 U12286 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n20893) );
  NAND2_X1 U12287 ( .A1(n11415), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11418) );
  INV_X1 U12288 ( .A(n18671), .ZN(n11415) );
  AND2_X1 U12289 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18716) );
  AOI21_X1 U12290 ( .B1(n14602), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n11243), .ZN(n11407) );
  NOR2_X1 U12291 ( .A1(n21605), .A2(n21644), .ZN(n21626) );
  AND2_X1 U12292 ( .A1(n18538), .A2(n18536), .ZN(n18586) );
  NAND2_X1 U12293 ( .A1(n18537), .A2(n14428), .ZN(n21654) );
  NAND2_X1 U12294 ( .A1(n21652), .A2(n21809), .ZN(n21667) );
  AOI21_X1 U12295 ( .B1(n14426), .B2(n14425), .A(n18511), .ZN(n18557) );
  NAND2_X1 U12296 ( .A1(n18557), .A2(n21599), .ZN(n18556) );
  NAND2_X1 U12297 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11427) );
  NOR2_X1 U12298 ( .A1(n11422), .A2(n14600), .ZN(n21683) );
  INV_X1 U12299 ( .A(n21509), .ZN(n21732) );
  NAND2_X1 U12300 ( .A1(n11414), .A2(n11412), .ZN(n18611) );
  NAND2_X1 U12301 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18402), .ZN(
        n21509) );
  NAND2_X1 U12302 ( .A1(n18681), .A2(n14417), .ZN(n18665) );
  XNOR2_X1 U12303 ( .A(n18401), .B(n14416), .ZN(n18682) );
  INV_X1 U12304 ( .A(n14415), .ZN(n14416) );
  NAND2_X1 U12305 ( .A1(n18682), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18681) );
  XNOR2_X1 U12306 ( .A(n14589), .B(n14590), .ZN(n18694) );
  NOR2_X1 U12307 ( .A1(n18694), .A2(n21787), .ZN(n18693) );
  NOR2_X1 U12308 ( .A1(n18710), .A2(n14585), .ZN(n18702) );
  XNOR2_X1 U12309 ( .A(n14412), .B(n14411), .ZN(n18699) );
  INV_X1 U12310 ( .A(n14410), .ZN(n14411) );
  XNOR2_X1 U12311 ( .A(n14582), .B(n21463), .ZN(n18712) );
  NOR2_X1 U12312 ( .A1(n18712), .A2(n18711), .ZN(n18710) );
  XNOR2_X1 U12313 ( .A(n14403), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n18739) );
  NAND2_X1 U12314 ( .A1(n18738), .A2(n18739), .ZN(n18737) );
  OAI21_X1 U12315 ( .B1(n14471), .B2(n14470), .A(n14469), .ZN(n21817) );
  INV_X1 U12316 ( .A(n11313), .ZN(n14544) );
  AND2_X1 U12317 ( .A1(n14547), .A2(n15950), .ZN(n11320) );
  NAND2_X1 U12318 ( .A1(n21790), .A2(n21812), .ZN(n21625) );
  NAND2_X1 U12319 ( .A1(n15951), .A2(n20671), .ZN(n21812) );
  INV_X1 U12320 ( .A(n21812), .ZN(n21736) );
  NAND2_X1 U12321 ( .A1(n21376), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n21380) );
  INV_X1 U12322 ( .A(n14532), .ZN(n19553) );
  NOR2_X1 U12323 ( .A1(n14523), .A2(n14522), .ZN(n19511) );
  INV_X1 U12324 ( .A(n21231), .ZN(n19430) );
  NAND3_X1 U12325 ( .A1(n14512), .A2(n14511), .A3(n14510), .ZN(n21232) );
  INV_X1 U12326 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n20744) );
  OAI22_X1 U12327 ( .A1(n14611), .A2(n21811), .B1(n21808), .B2(n21457), .ZN(
        n21844) );
  NOR2_X1 U12328 ( .A1(n21857), .A2(n20744), .ZN(n21845) );
  OR2_X1 U12329 ( .A1(n20741), .A2(n20679), .ZN(n21846) );
  NAND2_X1 U12330 ( .A1(n22312), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n22304) );
  NAND2_X1 U12331 ( .A1(n14783), .A2(n14782), .ZN(n21874) );
  AND2_X1 U12332 ( .A1(n22236), .A2(n15980), .ZN(n22258) );
  INV_X1 U12333 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n22212) );
  AND2_X1 U12334 ( .A1(n13918), .A2(n15235), .ZN(n22199) );
  INV_X1 U12335 ( .A(n22166), .ZN(n22177) );
  NOR2_X1 U12336 ( .A1(n15938), .A2(n15937), .ZN(n22167) );
  INV_X1 U12337 ( .A(n22199), .ZN(n22267) );
  AND2_X1 U12338 ( .A1(n22104), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n22244) );
  AND2_X1 U12339 ( .A1(n17814), .A2(n15231), .ZN(n22235) );
  INV_X1 U12340 ( .A(n16191), .ZN(n16253) );
  NAND2_X1 U12341 ( .A1(n14936), .A2(n14935), .ZN(n16265) );
  NAND2_X1 U12342 ( .A1(n14931), .A2(n16042), .ZN(n14936) );
  OR2_X1 U12343 ( .A1(n16252), .A2(n14938), .ZN(n16268) );
  NOR2_X1 U12344 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n22273), .ZN(n20425) );
  CLKBUF_X1 U12345 ( .A(n15529), .Z(n15535) );
  XNOR2_X1 U12346 ( .A(n13837), .B(n13836), .ZN(n15243) );
  OR2_X1 U12347 ( .A1(n13835), .A2(n16275), .ZN(n13837) );
  INV_X1 U12348 ( .A(n20594), .ZN(n20584) );
  OR2_X1 U12349 ( .A1(n20588), .A2(n14944), .ZN(n20594) );
  INV_X1 U12350 ( .A(n22268), .ZN(n20591) );
  AND2_X1 U12351 ( .A1(n16537), .A2(n22013), .ZN(n21899) );
  NAND2_X1 U12352 ( .A1(n21909), .A2(n22050), .ZN(n22012) );
  INV_X1 U12353 ( .A(n21933), .ZN(n21956) );
  INV_X2 U12354 ( .A(n22049), .ZN(n22052) );
  NAND2_X1 U12355 ( .A1(n14923), .A2(n16613), .ZN(n21892) );
  AND2_X1 U12356 ( .A1(n14923), .A2(n14912), .ZN(n22056) );
  CLKBUF_X1 U12357 ( .A(n13340), .Z(n13341) );
  INV_X1 U12358 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n17795) );
  INV_X1 U12359 ( .A(n14999), .ZN(n15333) );
  NOR2_X1 U12360 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n16596) );
  OR2_X1 U12361 ( .A1(n22370), .A2(n22369), .ZN(n22592) );
  OAI21_X1 U12362 ( .B1(n22392), .B2(n22391), .A(n22390), .ZN(n22634) );
  AND2_X1 U12363 ( .A1(n15087), .A2(n13338), .ZN(n22642) );
  OAI211_X1 U12364 ( .C1(n22529), .C2(n22435), .A(n15783), .B(n22419), .ZN(
        n22532) );
  OAI21_X1 U12365 ( .B1(n15336), .B2(n22414), .A(n22387), .ZN(n22543) );
  NOR2_X1 U12366 ( .A1(n15572), .A2(n15655), .ZN(n22663) );
  AOI22_X1 U12367 ( .A1(n22431), .A2(n22440), .B1(n22430), .B2(n22429), .ZN(
        n22668) );
  INV_X1 U12368 ( .A(n22674), .ZN(n22667) );
  AND2_X1 U12369 ( .A1(n15453), .A2(n13338), .ZN(n22661) );
  NOR2_X1 U12370 ( .A1(n15782), .A2(n15481), .ZN(n16628) );
  NOR2_X1 U12371 ( .A1(n15782), .A2(n15494), .ZN(n16633) );
  NOR2_X1 U12372 ( .A1(n15782), .A2(n15492), .ZN(n16643) );
  NOR2_X1 U12373 ( .A1(n15168), .A2(n12961), .ZN(n22554) );
  OAI211_X1 U12374 ( .C1(n15546), .C2(n22553), .A(n22416), .B(n22439), .ZN(
        n22557) );
  INV_X1 U12375 ( .A(n22680), .ZN(n16653) );
  AND2_X1 U12376 ( .A1(n15453), .A2(n15568), .ZN(n22556) );
  INV_X1 U12377 ( .A(n22433), .ZN(n22400) );
  INV_X1 U12378 ( .A(n22464), .ZN(n22459) );
  INV_X1 U12379 ( .A(n16633), .ZN(n22469) );
  INV_X1 U12380 ( .A(n16638), .ZN(n22492) );
  INV_X1 U12381 ( .A(n22487), .ZN(n22482) );
  INV_X1 U12382 ( .A(n22511), .ZN(n22506) );
  INV_X1 U12383 ( .A(n16643), .ZN(n22516) );
  INV_X1 U12384 ( .A(n22578), .ZN(n22573) );
  INV_X1 U12385 ( .A(n22608), .ZN(n22601) );
  OR2_X1 U12386 ( .A1(n15458), .A2(n15655), .ZN(n22615) );
  NOR2_X1 U12387 ( .A1(n15782), .A2(n15649), .ZN(n22674) );
  NAND2_X1 U12388 ( .A1(n13312), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n22283) );
  NOR2_X1 U12389 ( .A1(n16036), .A2(n22435), .ZN(n22277) );
  NAND2_X1 U12390 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n22273) );
  NAND2_X1 U12391 ( .A1(n16659), .A2(n19029), .ZN(n19142) );
  OAI21_X1 U12392 ( .B1(n16661), .B2(n19015), .A(n11532), .ZN(n19141) );
  NAND2_X1 U12393 ( .A1(n19128), .A2(n19129), .ZN(n19126) );
  NAND2_X1 U12394 ( .A1(n19112), .A2(n19113), .ZN(n19111) );
  NAND2_X1 U12395 ( .A1(n11399), .A2(n11397), .ZN(n12234) );
  NAND2_X1 U12396 ( .A1(n11399), .A2(n11400), .ZN(n12230) );
  NAND2_X1 U12397 ( .A1(n19102), .A2(n19103), .ZN(n19101) );
  NAND2_X1 U12398 ( .A1(n19090), .A2(n19091), .ZN(n19089) );
  NAND2_X1 U12399 ( .A1(n19080), .A2(n19081), .ZN(n19079) );
  NAND2_X1 U12400 ( .A1(n19029), .A2(n19045), .ZN(n19057) );
  NAND2_X1 U12401 ( .A1(n19057), .A2(n19058), .ZN(n19056) );
  NAND2_X1 U12402 ( .A1(n11549), .A2(n11550), .ZN(n16814) );
  AND2_X1 U12403 ( .A1(n19151), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19157) );
  INV_X1 U12404 ( .A(n19098), .ZN(n19160) );
  OR2_X1 U12405 ( .A1(n12636), .A2(n12635), .ZN(n15565) );
  OR2_X1 U12406 ( .A1(n12607), .A2(n12606), .ZN(n15360) );
  OR2_X1 U12407 ( .A1(n12581), .A2(n12580), .ZN(n15058) );
  OR2_X1 U12408 ( .A1(n12566), .A2(n12565), .ZN(n15056) );
  NAND2_X1 U12409 ( .A1(n16703), .A2(n16705), .ZN(n16704) );
  XNOR2_X1 U12410 ( .A(n16710), .B(n14191), .ZN(n16703) );
  AND2_X1 U12411 ( .A1(n15701), .A2(n19752), .ZN(n20064) );
  AND2_X1 U12412 ( .A1(n15701), .A2(n15700), .ZN(n20063) );
  NAND2_X1 U12413 ( .A1(n11554), .A2(n11648), .ZN(n14819) );
  OR2_X1 U12414 ( .A1(n14814), .A2(n14812), .ZN(n11554) );
  AND2_X1 U12415 ( .A1(n20012), .A2(n16818), .ZN(n20018) );
  INV_X1 U12416 ( .A(n20012), .ZN(n20068) );
  INV_X1 U12417 ( .A(n16818), .ZN(n20067) );
  NAND2_X1 U12418 ( .A1(n14811), .A2(n18854), .ZN(n20060) );
  NOR2_X1 U12419 ( .A1(n17918), .A2(n17949), .ZN(n17928) );
  BUF_X1 U12421 ( .A(n17937), .Z(n17949) );
  NAND2_X1 U12422 ( .A1(n14675), .A2(n14673), .ZN(n14788) );
  INV_X1 U12423 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n18933) );
  AND3_X1 U12424 ( .A1(n11340), .A2(n11341), .A3(n12406), .ZN(n17869) );
  AND2_X1 U12425 ( .A1(n11506), .A2(n12270), .ZN(n14979) );
  NAND2_X1 U12426 ( .A1(n17029), .A2(n17766), .ZN(n17865) );
  INV_X1 U12427 ( .A(n17029), .ZN(n17866) );
  INV_X1 U12428 ( .A(n17859), .ZN(n17879) );
  OAI211_X1 U12429 ( .C1(n16017), .C2(n19180), .A(n12788), .B(n11634), .ZN(
        n12789) );
  XNOR2_X1 U12430 ( .A(n12784), .B(n12783), .ZN(n16831) );
  OR2_X1 U12431 ( .A1(n16875), .A2(n16876), .ZN(n11609) );
  OR2_X1 U12432 ( .A1(n11581), .A2(n17110), .ZN(n11580) );
  AND2_X1 U12433 ( .A1(n17012), .A2(n11380), .ZN(n16992) );
  NAND2_X1 U12434 ( .A1(n17012), .A2(n17010), .ZN(n17001) );
  CLKBUF_X1 U12435 ( .A(n17016), .Z(n19213) );
  INV_X1 U12436 ( .A(n19202), .ZN(n17283) );
  NAND2_X1 U12437 ( .A1(n16002), .A2(n12734), .ZN(n19183) );
  INV_X1 U12438 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19927) );
  INV_X1 U12439 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19926) );
  INV_X1 U12440 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19832) );
  INV_X1 U12441 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17769) );
  INV_X1 U12442 ( .A(n17365), .ZN(n19279) );
  NOR2_X1 U12443 ( .A1(n14803), .A2(n14802), .ZN(n19915) );
  INV_X1 U12444 ( .A(n14881), .ZN(n14883) );
  XNOR2_X1 U12445 ( .A(n14889), .B(n14888), .ZN(n19879) );
  NAND2_X1 U12446 ( .A1(n14983), .A2(n14986), .ZN(n19880) );
  OR2_X1 U12447 ( .A1(n14984), .A2(n14985), .ZN(n14986) );
  AOI21_X1 U12448 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n19269), .A(n15764), .ZN(
        n19166) );
  OAI21_X1 U12449 ( .B1(n19921), .B2(n19920), .A(n19919), .ZN(n20333) );
  OAI21_X1 U12450 ( .B1(n19892), .B2(n19888), .A(n19887), .ZN(n20321) );
  INV_X1 U12451 ( .A(n19882), .ZN(n20319) );
  OAI21_X1 U12452 ( .B1(n20293), .B2(n19835), .A(n19919), .ZN(n20295) );
  INV_X1 U12453 ( .A(n20214), .ZN(n20288) );
  OAI21_X1 U12454 ( .B1(n19816), .B2(n19812), .A(n19811), .ZN(n20283) );
  INV_X1 U12455 ( .A(n20274), .ZN(n20277) );
  INV_X1 U12456 ( .A(n20184), .ZN(n20189) );
  INV_X1 U12457 ( .A(n20145), .ZN(n20149) );
  AOI22_X1 U12458 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20251), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n20250), .ZN(n20052) );
  INV_X1 U12459 ( .A(n20045), .ZN(n20056) );
  OR2_X1 U12460 ( .A1(n19783), .A2(n19925), .ZN(n20267) );
  AOI22_X1 U12461 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n20250), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n20251), .ZN(n20345) );
  INV_X1 U12462 ( .A(n20337), .ZN(n20352) );
  AND2_X1 U12463 ( .A1(n20247), .A2(n20246), .ZN(n20347) );
  INV_X1 U12464 ( .A(n20227), .ZN(n20238) );
  AND2_X1 U12465 ( .A1(n13896), .A2(n20246), .ZN(n20237) );
  INV_X1 U12466 ( .A(n20187), .ZN(n20191) );
  AOI22_X1 U12467 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20251), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n20250), .ZN(n20184) );
  INV_X1 U12468 ( .A(n20138), .ZN(n20147) );
  AOI22_X1 U12469 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20251), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n20250), .ZN(n20145) );
  INV_X1 U12470 ( .A(n20100), .ZN(n20107) );
  INV_X1 U12471 ( .A(n20052), .ZN(n20054) );
  AOI22_X1 U12472 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n20250), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n20251), .ZN(n20045) );
  INV_X1 U12473 ( .A(n20261), .ZN(n20196) );
  INV_X1 U12474 ( .A(n19997), .ZN(n20004) );
  INV_X1 U12475 ( .A(n20199), .ZN(n20348) );
  INV_X1 U12476 ( .A(n19924), .ZN(n19956) );
  AND2_X1 U12477 ( .A1(n19758), .A2(n20246), .ZN(n19951) );
  NAND2_X1 U12478 ( .A1(n19768), .A2(n19895), .ZN(n20261) );
  NAND3_X1 U12479 ( .A1(n19256), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n19287) );
  NAND2_X1 U12480 ( .A1(n17954), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n17988) );
  NAND2_X1 U12481 ( .A1(n21844), .A2(n21845), .ZN(n21871) );
  NOR2_X1 U12482 ( .A1(n21116), .A2(n21128), .ZN(n21117) );
  AND2_X1 U12483 ( .A1(n11359), .A2(n11358), .ZN(n21081) );
  OR2_X1 U12484 ( .A1(n21060), .A2(n21128), .ZN(n11359) );
  NOR2_X1 U12485 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n21050), .ZN(n21069) );
  NOR2_X1 U12486 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n21024), .ZN(n21046) );
  OR2_X1 U12487 ( .A1(n21025), .A2(n21128), .ZN(n11351) );
  NOR2_X1 U12488 ( .A1(n20984), .A2(n21128), .ZN(n20985) );
  NOR2_X1 U12489 ( .A1(n20933), .A2(n20949), .ZN(n20936) );
  NOR2_X1 U12490 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n20917), .ZN(n20931) );
  NAND4_X1 U12491 ( .A1(n20742), .A2(P3_EBX_REG_31__SCAN_IN), .A3(n20741), 
        .A4(n20740), .ZN(n21135) );
  INV_X1 U12492 ( .A(n21076), .ZN(n21075) );
  NOR2_X1 U12493 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n20837), .ZN(n20855) );
  INV_X1 U12494 ( .A(n20933), .ZN(n20817) );
  NAND2_X1 U12495 ( .A1(n20737), .A2(n20742), .ZN(n21076) );
  INV_X1 U12496 ( .A(n21135), .ZN(n21160) );
  INV_X1 U12497 ( .A(n21132), .ZN(n21161) );
  NOR2_X1 U12498 ( .A1(n21068), .A2(n18263), .ZN(n18267) );
  INV_X1 U12499 ( .A(n21267), .ZN(n21197) );
  INV_X1 U12500 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18048) );
  NOR2_X1 U12501 ( .A1(n18365), .A2(n17990), .ZN(n17998) );
  NOR2_X2 U12502 ( .A1(n21197), .A2(n18365), .ZN(n18366) );
  INV_X1 U12503 ( .A(n21301), .ZN(n21268) );
  NAND2_X1 U12504 ( .A1(n21268), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n21273) );
  NOR2_X1 U12505 ( .A1(n21267), .A2(n21307), .ZN(n21302) );
  NOR3_X1 U12506 ( .A1(n21314), .A2(n21266), .A3(n21265), .ZN(n21308) );
  NAND2_X1 U12507 ( .A1(n21323), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n21314) );
  NOR2_X1 U12508 ( .A1(n21326), .A2(n21325), .ZN(n21323) );
  NOR2_X1 U12509 ( .A1(n21190), .A2(n21189), .ZN(n21194) );
  NOR2_X1 U12510 ( .A1(n21340), .A2(n21168), .ZN(n21169) );
  NOR2_X1 U12511 ( .A1(n14326), .A2(n14325), .ZN(n21213) );
  NOR2_X1 U12512 ( .A1(n14336), .A2(n14335), .ZN(n21224) );
  NOR2_X1 U12513 ( .A1(n21222), .A2(n21221), .ZN(n21226) );
  INV_X1 U12514 ( .A(n21345), .ZN(n21227) );
  NAND2_X1 U12515 ( .A1(n21196), .A2(P3_EAX_REG_1__SCAN_IN), .ZN(n21340) );
  INV_X1 U12516 ( .A(n21196), .ZN(n21344) );
  NOR2_X1 U12517 ( .A1(n21170), .A2(n21344), .ZN(n21345) );
  CLKBUF_X1 U12518 ( .A(n20731), .Z(n20728) );
  NOR2_X1 U12519 ( .A1(n20732), .A2(n20683), .ZN(n20731) );
  NAND2_X1 U12520 ( .A1(n18539), .A2(n21673), .ZN(n21652) );
  INV_X1 U12521 ( .A(n18562), .ZN(n18529) );
  AND3_X1 U12522 ( .A1(n18399), .A2(n11364), .A3(n11250), .ZN(n18478) );
  AND2_X1 U12523 ( .A1(n18753), .A2(n11315), .ZN(n18562) );
  INV_X1 U12524 ( .A(n19551), .ZN(n19639) );
  INV_X1 U12525 ( .A(n18416), .ZN(n18607) );
  INV_X1 U12526 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n20955) );
  NAND3_X1 U12527 ( .A1(n22296), .A2(n18753), .A3(P3_STATE2_REG_1__SCAN_IN), 
        .ZN(n18571) );
  NOR2_X1 U12528 ( .A1(n20893), .A2(n18443), .ZN(n20900) );
  INV_X1 U12529 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18443) );
  OR2_X1 U12530 ( .A1(n18758), .A2(n21397), .ZN(n11316) );
  INV_X1 U12531 ( .A(n18589), .ZN(n18672) );
  NAND3_X1 U12532 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20795) );
  INV_X1 U12533 ( .A(n18753), .ZN(n18730) );
  INV_X1 U12534 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20793) );
  INV_X1 U12535 ( .A(n18716), .ZN(n18717) );
  NAND2_X1 U12536 ( .A1(n19640), .A2(n19355), .ZN(n19551) );
  INV_X1 U12537 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n21354) );
  AOI21_X1 U12538 ( .B1(n11431), .B2(n21654), .A(n11430), .ZN(n21664) );
  AND2_X1 U12539 ( .A1(n21655), .A2(n21656), .ZN(n11430) );
  OAI21_X1 U12540 ( .B1(n21667), .B2(n21653), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11431) );
  NOR2_X1 U12541 ( .A1(n11422), .A2(n11421), .ZN(n18502) );
  OR3_X1 U12542 ( .A1(n11428), .A2(n11429), .A3(n11427), .ZN(n18512) );
  AND2_X1 U12543 ( .A1(n11432), .A2(n14421), .ZN(n18605) );
  NOR2_X1 U12544 ( .A1(n21544), .A2(n18612), .ZN(n21565) );
  INV_X1 U12545 ( .A(n21592), .ZN(n21606) );
  INV_X1 U12546 ( .A(n21693), .ZN(n21793) );
  INV_X1 U12547 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21508) );
  INV_X1 U12548 ( .A(n21680), .ZN(n21744) );
  NOR2_X1 U12549 ( .A1(n18370), .A2(n22296), .ZN(n19355) );
  INV_X1 U12550 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21838) );
  INV_X1 U12551 ( .A(n21845), .ZN(n21868) );
  NAND2_X1 U12552 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n22352) );
  NAND2_X1 U12553 ( .A1(n22345), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18843) );
  CLKBUF_X1 U12554 ( .A(n19636), .Z(n19593) );
  INV_X1 U12555 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20360) );
  NAND2_X1 U12556 ( .A1(n16277), .A2(n13916), .ZN(n14009) );
  NOR4_X1 U12557 ( .A1(n16454), .A2(n16453), .A3(n16452), .A4(n16451), .ZN(
        n16455) );
  AOI21_X1 U12558 ( .B1(n13904), .B2(n19159), .A(n13903), .ZN(n13907) );
  AND2_X1 U12559 ( .A1(n14299), .A2(n14298), .ZN(n14300) );
  NAND2_X1 U12560 ( .A1(n17055), .A2(n12415), .ZN(n16856) );
  AOI21_X1 U12561 ( .B1(n19110), .B2(n17878), .A(n12776), .ZN(n12777) );
  NAND2_X1 U12562 ( .A1(n11387), .A2(n11386), .ZN(P2_U3015) );
  NAND2_X1 U12563 ( .A1(n11337), .A2(n11334), .ZN(P2_U3018) );
  NAND2_X1 U12564 ( .A1(n17053), .A2(n19211), .ZN(n11337) );
  OAI21_X1 U12565 ( .B1(n12834), .B2(n19187), .A(n12833), .ZN(n12835) );
  OAI21_X1 U12566 ( .B1(n21139), .B2(n21851), .A(n21138), .ZN(n21140) );
  INV_X1 U12567 ( .A(n21281), .ZN(n21285) );
  NOR2_X1 U12568 ( .A1(n14614), .A2(n18589), .ZN(n14628) );
  AOI21_X1 U12569 ( .B1(n14608), .B2(n21739), .A(n14607), .ZN(n14609) );
  OAI21_X1 U12570 ( .B1(n21680), .B2(n21353), .A(n14618), .ZN(n14607) );
  AND2_X1 U12571 ( .A1(n12424), .A2(n16857), .ZN(n11189) );
  NAND2_X1 U12572 ( .A1(n11497), .A2(n11501), .ZN(n15692) );
  NOR2_X1 U12573 ( .A1(n16880), .A2(n17100), .ZN(n16867) );
  AND2_X1 U12574 ( .A1(n15910), .A2(n11204), .ZN(n11191) );
  AND2_X1 U12575 ( .A1(n11855), .A2(n17838), .ZN(n11192) );
  NAND2_X1 U12576 ( .A1(n12761), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12762) );
  INV_X1 U12577 ( .A(n12516), .ZN(n12678) );
  NOR2_X1 U12578 ( .A1(n14309), .A2(n20747), .ZN(n14395) );
  AND2_X1 U12579 ( .A1(n14156), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11921) );
  NAND2_X1 U12580 ( .A1(n20572), .A2(n13232), .ZN(n11193) );
  INV_X1 U12581 ( .A(n16869), .ZN(n11606) );
  NOR2_X1 U12582 ( .A1(n15564), .A2(n11254), .ZN(n15833) );
  AND3_X1 U12583 ( .A1(n13376), .A2(n13375), .A3(n11619), .ZN(n11194) );
  OR2_X1 U12584 ( .A1(n16894), .A2(n11581), .ZN(n12812) );
  AND2_X1 U12585 ( .A1(n15040), .A2(n11495), .ZN(n15358) );
  NAND2_X1 U12586 ( .A1(n11681), .A2(n11680), .ZN(n12031) );
  AND2_X1 U12587 ( .A1(n12974), .A2(n16022), .ZN(n11195) );
  AND2_X1 U12588 ( .A1(n11830), .A2(n11835), .ZN(n17336) );
  INV_X1 U12589 ( .A(n16412), .ZN(n20578) );
  AND2_X1 U12590 ( .A1(n11622), .A2(n11621), .ZN(n11196) );
  INV_X1 U12592 ( .A(n11189), .ZN(n11593) );
  INV_X1 U12593 ( .A(n12177), .ZN(n12141) );
  AND2_X1 U12594 ( .A1(n11555), .A2(n11552), .ZN(n11197) );
  OR3_X1 U12595 ( .A1(n16796), .A2(n16777), .A3(n11558), .ZN(n11198) );
  NAND2_X1 U12596 ( .A1(n12963), .A2(n12962), .ZN(n12989) );
  NAND2_X1 U12597 ( .A1(n12269), .A2(n12271), .ZN(n11506) );
  NAND2_X1 U12598 ( .A1(n11506), .A2(n11505), .ZN(n14980) );
  AND2_X1 U12599 ( .A1(n11645), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11199) );
  AND2_X1 U12600 ( .A1(n11570), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11200) );
  AND2_X1 U12601 ( .A1(n11239), .A2(n11614), .ZN(n11201) );
  INV_X1 U12602 ( .A(n11617), .ZN(n15860) );
  AND2_X1 U12603 ( .A1(n11199), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11202) );
  NAND2_X1 U12604 ( .A1(n11456), .A2(n11457), .ZN(n11203) );
  NOR2_X1 U12605 ( .A1(n16731), .A2(n11492), .ZN(n11204) );
  AND2_X1 U12606 ( .A1(n11567), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11205) );
  AND2_X1 U12607 ( .A1(n11468), .A2(n11467), .ZN(n11206) );
  AND2_X1 U12608 ( .A1(n11204), .A2(n16723), .ZN(n11207) );
  INV_X1 U12609 ( .A(n18754), .ZN(n11315) );
  AND3_X1 U12610 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(P3_EAX_REG_28__SCAN_IN), 
        .A3(P3_EAX_REG_27__SCAN_IN), .ZN(n11208) );
  OR2_X2 U12611 ( .A1(n14308), .A2(n20747), .ZN(n11209) );
  AND2_X1 U12612 ( .A1(n16104), .A2(n11206), .ZN(n11210) );
  OR2_X1 U12613 ( .A1(n12220), .A2(n12219), .ZN(n11211) );
  OR2_X1 U12614 ( .A1(n11847), .A2(n11846), .ZN(n12270) );
  NOR2_X1 U12615 ( .A1(n16110), .A2(n16112), .ZN(n16111) );
  NAND2_X1 U12616 ( .A1(n21376), .A2(n11419), .ZN(n14374) );
  AND4_X1 U12617 ( .A1(n12873), .A2(n12872), .A3(n12871), .A4(n12870), .ZN(
        n11212) );
  NAND2_X1 U12618 ( .A1(n11418), .A2(n11417), .ZN(n11416) );
  NAND2_X1 U12619 ( .A1(n18522), .A2(n21696), .ZN(n18521) );
  BUF_X1 U12620 ( .A(n11854), .Z(n16014) );
  INV_X1 U12621 ( .A(n11854), .ZN(n17838) );
  AND2_X1 U12622 ( .A1(n11373), .A2(n11371), .ZN(n11213) );
  AND2_X1 U12623 ( .A1(n11615), .A2(n11201), .ZN(n11214) );
  AND2_X1 U12624 ( .A1(n12054), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11893) );
  NOR2_X1 U12625 ( .A1(n16124), .A2(n16172), .ZN(n16171) );
  NAND2_X1 U12626 ( .A1(n12142), .A2(n12141), .ZN(n12170) );
  AND3_X1 U12627 ( .A1(n11697), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n11696), .ZN(n11215) );
  AND3_X1 U12628 ( .A1(n11695), .A2(n11716), .A3(n11692), .ZN(n11216) );
  NAND2_X1 U12630 ( .A1(n11609), .A2(n16877), .ZN(n16868) );
  AND2_X1 U12631 ( .A1(n11192), .A2(n11875), .ZN(n11978) );
  NAND2_X1 U12632 ( .A1(n13243), .A2(n16308), .ZN(n16300) );
  AND2_X1 U12633 ( .A1(n11607), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11217) );
  OAI21_X1 U12634 ( .B1(n18639), .B2(n14419), .A(n21668), .ZN(n14421) );
  AND4_X1 U12635 ( .A1(n14528), .A2(n14527), .A3(n14526), .A4(n14525), .ZN(
        n11218) );
  AND4_X1 U12636 ( .A1(n11925), .A2(n11924), .A3(n11923), .A4(n11922), .ZN(
        n11219) );
  AND2_X1 U12637 ( .A1(n11192), .A2(n11877), .ZN(n11982) );
  AND2_X1 U12638 ( .A1(n16846), .A2(n17058), .ZN(n11220) );
  AND2_X1 U12639 ( .A1(n12247), .A2(n17058), .ZN(n11221) );
  NAND2_X1 U12640 ( .A1(n11282), .A2(n11802), .ZN(n11840) );
  NAND2_X1 U12642 ( .A1(n16658), .A2(n12438), .ZN(n12423) );
  INV_X1 U12643 ( .A(n12423), .ZN(n11390) );
  NAND2_X1 U12644 ( .A1(n11724), .A2(n11723), .ZN(n12717) );
  OR2_X1 U12645 ( .A1(n12247), .A2(n17058), .ZN(n11222) );
  OR2_X1 U12646 ( .A1(n17052), .A2(n17283), .ZN(n11223) );
  AND3_X1 U12647 ( .A1(n12917), .A2(n12916), .A3(n12915), .ZN(n11224) );
  AND3_X1 U12648 ( .A1(n11687), .A2(n11716), .A3(n11686), .ZN(n11226) );
  NOR2_X1 U12649 ( .A1(n21295), .A2(n21290), .ZN(n11227) );
  OR2_X1 U12650 ( .A1(n11390), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11228) );
  AND2_X1 U12651 ( .A1(n11854), .A2(n18858), .ZN(n11229) );
  NAND2_X1 U12652 ( .A1(n12209), .A2(n12808), .ZN(n11230) );
  AND2_X1 U12653 ( .A1(n12410), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11231) );
  NOR2_X1 U12654 ( .A1(n16894), .A2(n17138), .ZN(n11232) );
  NOR2_X1 U12655 ( .A1(n21197), .A2(n19511), .ZN(n14545) );
  AND2_X1 U12656 ( .A1(n11579), .A2(n12390), .ZN(n11233) );
  NAND2_X1 U12657 ( .A1(n12193), .A2(n12192), .ZN(n11234) );
  AND2_X1 U12658 ( .A1(n11274), .A2(n11455), .ZN(n11235) );
  INV_X1 U12659 ( .A(n12406), .ZN(n12407) );
  OR2_X1 U12660 ( .A1(n12405), .A2(n17867), .ZN(n12406) );
  AND2_X2 U12661 ( .A1(n11892), .A2(n14137), .ZN(n11907) );
  OR3_X1 U12662 ( .A1(n13870), .A2(n11536), .A3(n11539), .ZN(n11236) );
  OR2_X1 U12663 ( .A1(n19758), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11237) );
  NAND2_X1 U12664 ( .A1(n14984), .A2(n14985), .ZN(n14983) );
  INV_X1 U12665 ( .A(n13855), .ZN(n11569) );
  NOR2_X1 U12666 ( .A1(n11515), .A2(n12771), .ZN(n12770) );
  NAND2_X1 U12667 ( .A1(n18665), .A2(n18666), .ZN(n18425) );
  NAND2_X1 U12668 ( .A1(n15910), .A2(n16735), .ZN(n16730) );
  NOR2_X1 U12669 ( .A1(n15564), .A2(n15709), .ZN(n15691) );
  NAND2_X1 U12670 ( .A1(n16104), .A2(n16082), .ZN(n16072) );
  OR3_X1 U12671 ( .A1(n16726), .A2(n16720), .A3(n11514), .ZN(n11238) );
  AND2_X1 U12672 ( .A1(n13624), .A2(n11616), .ZN(n11239) );
  AND2_X1 U12673 ( .A1(n13861), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13850) );
  NAND2_X1 U12674 ( .A1(n11783), .A2(n13906), .ZN(n12725) );
  AND2_X1 U12675 ( .A1(n13864), .A2(n11561), .ZN(n11240) );
  NOR2_X1 U12676 ( .A1(n15839), .A2(n15838), .ZN(n15877) );
  XNOR2_X1 U12677 ( .A(n18570), .B(n21147), .ZN(n20933) );
  NAND2_X1 U12678 ( .A1(n12123), .A2(n12122), .ZN(n12130) );
  NAND2_X1 U12679 ( .A1(n12066), .A2(n12067), .ZN(n12112) );
  NAND2_X1 U12680 ( .A1(n11333), .A2(n11331), .ZN(n17847) );
  AND2_X1 U12681 ( .A1(n17135), .A2(n12827), .ZN(n12826) );
  NAND2_X1 U12682 ( .A1(n15910), .A2(n11207), .ZN(n16717) );
  OR2_X1 U12683 ( .A1(n15404), .A2(n11509), .ZN(n11241) );
  NAND2_X1 U12684 ( .A1(n19169), .A2(n11785), .ZN(n12471) );
  NOR2_X1 U12685 ( .A1(n15404), .A2(n11507), .ZN(n15706) );
  NOR2_X1 U12686 ( .A1(n14993), .A2(n11540), .ZN(n15108) );
  AND2_X1 U12687 ( .A1(n14018), .A2(n14033), .ZN(n14984) );
  AND2_X1 U12688 ( .A1(n16663), .A2(n12681), .ZN(n16662) );
  XNOR2_X1 U12689 ( .A(n12031), .B(n11784), .ZN(n12477) );
  NAND2_X1 U12690 ( .A1(n15713), .A2(n15832), .ZN(n15831) );
  AND2_X1 U12691 ( .A1(n18399), .A2(n11644), .ZN(n18398) );
  AND2_X1 U12692 ( .A1(n11518), .A2(n11517), .ZN(n11242) );
  AND3_X1 U12693 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n21604), .A3(
        n21648), .ZN(n11243) );
  INV_X1 U12694 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n19256) );
  AND2_X1 U12695 ( .A1(n20020), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11244) );
  OR2_X1 U12696 ( .A1(n16796), .A2(n16786), .ZN(n11245) );
  INV_X1 U12697 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n21041) );
  INV_X1 U12698 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n13867) );
  INV_X1 U12699 ( .A(n12030), .ZN(n12526) );
  OR2_X1 U12700 ( .A1(n11968), .A2(n11967), .ZN(n12030) );
  AND2_X1 U12701 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n11246) );
  AND2_X1 U12702 ( .A1(n13670), .A2(n13669), .ZN(n16220) );
  INV_X1 U12703 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17030) );
  NAND2_X1 U12704 ( .A1(n15563), .A2(n15565), .ZN(n15564) );
  INV_X1 U12705 ( .A(n11562), .ZN(n11561) );
  NAND2_X1 U12706 ( .A1(n11563), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11562) );
  INV_X1 U12707 ( .A(n11485), .ZN(n11484) );
  NAND2_X1 U12708 ( .A1(n14975), .A2(n11276), .ZN(n11485) );
  NAND2_X1 U12709 ( .A1(n15713), .A2(n11516), .ZN(n12813) );
  INV_X1 U12710 ( .A(n11512), .ZN(n11511) );
  NOR2_X1 U12711 ( .A1(n15356), .A2(n11513), .ZN(n11512) );
  OR2_X1 U12712 ( .A1(n15404), .A2(n11511), .ZN(n11247) );
  AND2_X1 U12713 ( .A1(n12960), .A2(n13915), .ZN(n11248) );
  INV_X1 U12714 ( .A(n11372), .ZN(n11371) );
  NOR2_X1 U12715 ( .A1(n11376), .A2(n12806), .ZN(n11372) );
  AND2_X1 U12716 ( .A1(n11197), .A2(n14925), .ZN(n11249) );
  AND2_X1 U12717 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n14615), .ZN(
        n11250) );
  AND2_X1 U12718 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11251) );
  INV_X1 U12719 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n19270) );
  AND2_X1 U12720 ( .A1(n11452), .A2(n13246), .ZN(n11252) );
  INV_X1 U12721 ( .A(n19208), .ZN(n19180) );
  NAND2_X1 U12722 ( .A1(n14976), .A2(n14975), .ZN(n14974) );
  NAND2_X1 U12723 ( .A1(n11482), .A2(n11483), .ZN(n15006) );
  NAND2_X1 U12724 ( .A1(n11527), .A2(n11526), .ZN(n11525) );
  AND2_X1 U12725 ( .A1(n15006), .A2(n14036), .ZN(n15040) );
  AND2_X1 U12726 ( .A1(n14978), .A2(n12270), .ZN(n11505) );
  AND2_X1 U12727 ( .A1(n12673), .A2(n12672), .ZN(n16777) );
  NAND2_X1 U12728 ( .A1(n14814), .A2(n11648), .ZN(n11553) );
  NAND2_X1 U12729 ( .A1(n11553), .A2(n11555), .ZN(n14817) );
  NAND2_X1 U12730 ( .A1(n15040), .A2(n14037), .ZN(n15057) );
  NAND2_X1 U12731 ( .A1(n11525), .A2(n11524), .ZN(n15410) );
  NAND2_X1 U12732 ( .A1(n15040), .A2(n11494), .ZN(n15359) );
  OR3_X1 U12733 ( .A1(n13870), .A2(n11539), .A3(n12358), .ZN(n11253) );
  NAND2_X1 U12734 ( .A1(n11501), .A2(n11500), .ZN(n11254) );
  INV_X1 U12735 ( .A(n19029), .ZN(n19015) );
  NOR2_X1 U12736 ( .A1(n15652), .A2(n15651), .ZN(n15650) );
  AND2_X1 U12737 ( .A1(n11550), .A2(n11548), .ZN(n11255) );
  AND2_X1 U12738 ( .A1(n13882), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13843) );
  NOR2_X1 U12739 ( .A1(n14993), .A2(n11542), .ZN(n15107) );
  NOR2_X1 U12740 ( .A1(n15007), .A2(n15074), .ZN(n15042) );
  NOR2_X1 U12741 ( .A1(n15767), .A2(n15768), .ZN(n14994) );
  AND2_X1 U12742 ( .A1(n13847), .A2(n11567), .ZN(n11256) );
  AND3_X1 U12743 ( .A1(n18399), .A2(n11364), .A3(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18378) );
  AND2_X1 U12744 ( .A1(n18451), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18449) );
  AND2_X1 U12745 ( .A1(n11520), .A2(n11521), .ZN(n11257) );
  NAND2_X1 U12746 ( .A1(n12482), .A2(n20247), .ZN(n13887) );
  OR3_X1 U12747 ( .A1(n16720), .A2(n11514), .A3(n16706), .ZN(n11258) );
  NOR2_X1 U12748 ( .A1(n14993), .A2(n11544), .ZN(n15038) );
  AND2_X1 U12749 ( .A1(n14191), .A2(n16705), .ZN(n11259) );
  AND2_X1 U12750 ( .A1(n11619), .A2(n15861), .ZN(n11260) );
  NOR2_X1 U12751 ( .A1(n21538), .A2(n21495), .ZN(n11261) );
  NOR2_X1 U12752 ( .A1(n14993), .A2(n15847), .ZN(n15037) );
  INV_X1 U12753 ( .A(n11404), .ZN(n11403) );
  NAND2_X1 U12754 ( .A1(n12148), .A2(n12151), .ZN(n11404) );
  INV_X1 U12755 ( .A(n20738), .ZN(n20741) );
  NOR2_X1 U12756 ( .A1(n14481), .A2(n14480), .ZN(n20738) );
  AND2_X1 U12757 ( .A1(n11257), .A2(n12793), .ZN(n11262) );
  AND3_X1 U12758 ( .A1(n11506), .A2(n11505), .A3(n11504), .ZN(n11263) );
  AND2_X1 U12759 ( .A1(n11494), .A2(n11493), .ZN(n11264) );
  AND2_X1 U12760 ( .A1(n11351), .A2(n11350), .ZN(n11265) );
  AND2_X1 U12761 ( .A1(n11207), .A2(n11491), .ZN(n11266) );
  INV_X1 U12762 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n18592) );
  INV_X1 U12763 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n22274) );
  AND2_X1 U12764 ( .A1(n11525), .A2(n11528), .ZN(n11267) );
  INV_X1 U12765 ( .A(n15700), .ZN(n19752) );
  NAND2_X1 U12766 ( .A1(n18618), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18627) );
  AND2_X1 U12767 ( .A1(n11180), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11268) );
  AND2_X1 U12768 ( .A1(n11140), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n11269) );
  AND2_X1 U12769 ( .A1(n11180), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11270) );
  AND2_X1 U12770 ( .A1(n11140), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11271) );
  AND2_X1 U12771 ( .A1(n11180), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11272) );
  AND2_X1 U12772 ( .A1(n11140), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11273) );
  INV_X1 U12773 ( .A(n16786), .ZN(n11559) );
  NAND2_X1 U12774 ( .A1(n13941), .A2(n13940), .ZN(n11274) );
  XNOR2_X1 U12775 ( .A(n11476), .B(n14914), .ZN(n15028) );
  NAND2_X1 U12776 ( .A1(n18561), .A2(n11361), .ZN(n14619) );
  INV_X1 U12777 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11539) );
  OR2_X1 U12778 ( .A1(n14171), .A2(n13896), .ZN(n11275) );
  AND2_X1 U12779 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11276) );
  NAND2_X1 U12780 ( .A1(n18451), .A2(n11202), .ZN(n11345) );
  INV_X1 U12781 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11298) );
  INV_X1 U12782 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11362) );
  NOR2_X1 U12783 ( .A1(n18627), .A2(n18619), .ZN(n18399) );
  NAND2_X1 U12784 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11277) );
  AND2_X1 U12785 ( .A1(n11140), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11278) );
  AND2_X1 U12786 ( .A1(n11140), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11279) );
  AND2_X1 U12787 ( .A1(n11140), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11280) );
  NOR2_X1 U12788 ( .A1(n20795), .A2(n20793), .ZN(n18618) );
  INV_X1 U12789 ( .A(n14616), .ZN(n18561) );
  NAND2_X1 U12790 ( .A1(n18451), .A2(n11344), .ZN(n14616) );
  INV_X1 U12791 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21495) );
  NOR2_X1 U12792 ( .A1(n16547), .A2(n22022), .ZN(n11281) );
  INV_X1 U12793 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11610) );
  INV_X1 U12794 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11297) );
  INV_X1 U12795 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17138) );
  NOR2_X1 U12796 ( .A1(n14600), .A2(n21567), .ZN(n21682) );
  OAI21_X2 U12797 ( .B1(n15164), .B2(n15089), .A(n15088), .ZN(n22675) );
  OR2_X1 U12798 ( .A1(n15987), .A2(n16428), .ZN(n15164) );
  NAND2_X1 U12799 ( .A1(n11807), .A2(n11761), .ZN(n11283) );
  NAND2_X1 U12800 ( .A1(n16847), .A2(n11222), .ZN(n11284) );
  NAND2_X1 U12801 ( .A1(n16846), .A2(n11221), .ZN(n11285) );
  NAND2_X1 U12802 ( .A1(n11290), .A2(n11297), .ZN(n11296) );
  NAND2_X1 U12803 ( .A1(n17021), .A2(n11292), .ZN(n11291) );
  INV_X1 U12804 ( .A(n12120), .ZN(n11293) );
  NAND2_X2 U12805 ( .A1(n11295), .A2(n11294), .ZN(n17874) );
  XNOR2_X1 U12806 ( .A(n12115), .B(n12384), .ZN(n15813) );
  NOR2_X1 U12807 ( .A1(n12255), .A2(n11299), .ZN(n17345) );
  AND3_X2 U12808 ( .A1(n12129), .A2(n12128), .A3(n17873), .ZN(n17012) );
  NAND3_X1 U12809 ( .A1(n12129), .A2(n12128), .A3(n11301), .ZN(n11300) );
  NAND3_X1 U12810 ( .A1(n12099), .A2(n11302), .A3(n12098), .ZN(n12111) );
  NAND3_X1 U12811 ( .A1(n11306), .A2(n12097), .A3(n11304), .ZN(n11303) );
  INV_X1 U12812 ( .A(n16886), .ZN(n11309) );
  INV_X2 U12813 ( .A(n11855), .ZN(n15437) );
  NAND2_X1 U12814 ( .A1(n19470), .A2(n19553), .ZN(n14543) );
  INV_X1 U12815 ( .A(n14543), .ZN(n11310) );
  NAND2_X1 U12816 ( .A1(n11310), .A2(n14548), .ZN(n11311) );
  INV_X1 U12817 ( .A(n11312), .ZN(n14552) );
  NAND2_X1 U12818 ( .A1(n11312), .A2(n14545), .ZN(n14562) );
  OR2_X1 U12819 ( .A1(n19430), .A2(n14532), .ZN(n11313) );
  NAND3_X1 U12820 ( .A1(n14464), .A2(n14466), .A3(n14465), .ZN(n14532) );
  INV_X2 U12821 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n21371) );
  AND2_X2 U12822 ( .A1(n21756), .A2(n20738), .ZN(n21656) );
  NAND3_X1 U12823 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .A3(P3_EAX_REG_11__SCAN_IN), .ZN(n11318) );
  NAND2_X1 U12824 ( .A1(n14561), .A2(n21377), .ZN(n21373) );
  NAND2_X2 U12825 ( .A1(n11323), .A2(n11218), .ZN(n21267) );
  NAND3_X1 U12826 ( .A1(n14531), .A2(n14530), .A3(n11325), .ZN(n11324) );
  AND2_X4 U12827 ( .A1(n11892), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11884) );
  INV_X1 U12828 ( .A(n12375), .ZN(n11330) );
  NAND3_X1 U12829 ( .A1(n15430), .A2(n11330), .A3(n12374), .ZN(n11333) );
  NAND2_X1 U12830 ( .A1(n11332), .A2(n12375), .ZN(n11331) );
  NAND2_X1 U12831 ( .A1(n15430), .A2(n12374), .ZN(n11332) );
  NAND2_X1 U12832 ( .A1(n12387), .A2(n12388), .ZN(n11579) );
  INV_X1 U12833 ( .A(n12398), .ZN(n11338) );
  NAND2_X1 U12834 ( .A1(n11338), .A2(n12408), .ZN(n11341) );
  NAND2_X1 U12835 ( .A1(n17306), .A2(n12398), .ZN(n17027) );
  NAND2_X1 U12836 ( .A1(n17307), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17306) );
  INV_X1 U12837 ( .A(n11345), .ZN(n18516) );
  AOI21_X1 U12838 ( .B1(n21025), .B2(n11350), .A(n21128), .ZN(n21039) );
  NAND2_X1 U12839 ( .A1(n11348), .A2(n11346), .ZN(n21051) );
  NAND2_X1 U12840 ( .A1(n21025), .A2(n11349), .ZN(n11348) );
  INV_X1 U12841 ( .A(n11351), .ZN(n21026) );
  INV_X1 U12842 ( .A(n21027), .ZN(n11350) );
  AOI21_X1 U12843 ( .B1(n21060), .B2(n11358), .A(n21128), .ZN(n21082) );
  NAND2_X1 U12844 ( .A1(n11356), .A2(n11355), .ZN(n21090) );
  NAND2_X1 U12845 ( .A1(n21060), .A2(n11357), .ZN(n11356) );
  INV_X1 U12846 ( .A(n11359), .ZN(n21061) );
  INV_X1 U12847 ( .A(n21062), .ZN(n11358) );
  NAND3_X1 U12848 ( .A1(n12379), .A2(n12380), .A3(n12430), .ZN(n11589) );
  NAND2_X1 U12849 ( .A1(n12024), .A2(n11148), .ZN(n12380) );
  NAND2_X2 U12850 ( .A1(n11139), .A2(n12023), .ZN(n12379) );
  OR2_X1 U12851 ( .A1(n16922), .A2(n12804), .ZN(n11375) );
  NAND2_X1 U12852 ( .A1(n11373), .A2(n11367), .ZN(n11366) );
  NOR2_X1 U12853 ( .A1(n11372), .A2(n12198), .ZN(n11367) );
  NOR2_X1 U12854 ( .A1(n11370), .A2(n11369), .ZN(n11368) );
  INV_X1 U12855 ( .A(n12806), .ZN(n11378) );
  AND2_X2 U12856 ( .A1(n11180), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14068) );
  AND2_X2 U12857 ( .A1(n11140), .A2(n11716), .ZN(n14126) );
  NAND2_X1 U12858 ( .A1(n12123), .A2(n11388), .ZN(n12136) );
  INV_X1 U12859 ( .A(n12136), .ZN(n12134) );
  NAND4_X1 U12860 ( .A1(n12418), .A2(n12421), .A3(n11189), .A4(n17058), .ZN(
        n11591) );
  NAND3_X1 U12861 ( .A1(n11392), .A2(n12067), .A3(n11391), .ZN(n12116) );
  AOI21_X1 U12862 ( .B1(n14599), .B2(n21541), .A(n11410), .ZN(n11412) );
  AND2_X1 U12863 ( .A1(n14597), .A2(n11413), .ZN(n11410) );
  INV_X1 U12864 ( .A(n14599), .ZN(n11417) );
  NOR2_X1 U12865 ( .A1(n14596), .A2(n11411), .ZN(n18671) );
  AND2_X1 U12866 ( .A1(n14597), .A2(n14598), .ZN(n11411) );
  NAND2_X1 U12867 ( .A1(n14596), .A2(n11261), .ZN(n11414) );
  INV_X1 U12868 ( .A(n11418), .ZN(n18670) );
  INV_X1 U12869 ( .A(n11416), .ZN(n21397) );
  NAND3_X1 U12870 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n17747) );
  INV_X1 U12871 ( .A(n21729), .ZN(n11422) );
  NAND2_X1 U12872 ( .A1(n21729), .A2(n11420), .ZN(n18501) );
  OR2_X1 U12873 ( .A1(n18471), .A2(n18447), .ZN(n11429) );
  INV_X1 U12874 ( .A(n18521), .ZN(n11428) );
  INV_X1 U12875 ( .A(n14426), .ZN(n14427) );
  AOI22_X2 U12876 ( .A1(n14420), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(
        n18548), .B2(n21752), .ZN(n11432) );
  OR2_X2 U12877 ( .A1(n14348), .A2(n14347), .ZN(n21337) );
  OAI21_X1 U12878 ( .B1(n11437), .B2(n12968), .A(n12946), .ZN(n14840) );
  NAND2_X1 U12879 ( .A1(n12954), .A2(n12953), .ZN(n11437) );
  NOR2_X1 U12880 ( .A1(n16269), .A2(n11252), .ZN(n11440) );
  NOR2_X1 U12881 ( .A1(n16269), .A2(n16271), .ZN(n16280) );
  INV_X1 U12882 ( .A(n16476), .ZN(n11442) );
  NAND3_X1 U12883 ( .A1(n16411), .A2(n11450), .A3(n11452), .ZN(n11446) );
  NAND2_X1 U12884 ( .A1(n16411), .A2(n13225), .ZN(n16375) );
  NOR2_X2 U12885 ( .A1(n13237), .A2(n11451), .ZN(n11450) );
  INV_X1 U12886 ( .A(n15374), .ZN(n11454) );
  NAND3_X1 U12887 ( .A1(n11454), .A2(n11457), .A3(n11235), .ZN(n15652) );
  NAND2_X1 U12888 ( .A1(n12971), .A2(n12962), .ZN(n12990) );
  NAND2_X1 U12889 ( .A1(n11464), .A2(n16493), .ZN(n11463) );
  NAND2_X2 U12890 ( .A1(n13240), .A2(n11452), .ZN(n11465) );
  NAND2_X1 U12891 ( .A1(n11477), .A2(n13919), .ZN(n11475) );
  INV_X1 U12892 ( .A(n13925), .ZN(n11477) );
  NAND2_X1 U12893 ( .A1(n11837), .A2(n11478), .ZN(n11839) );
  NAND2_X1 U12894 ( .A1(n14015), .A2(n14014), .ZN(n11481) );
  NAND2_X1 U12895 ( .A1(n11481), .A2(n14017), .ZN(n14033) );
  NAND3_X1 U12896 ( .A1(n14984), .A2(n11484), .A3(n14985), .ZN(n11483) );
  INV_X1 U12897 ( .A(n11488), .ZN(n11487) );
  OAI21_X1 U12898 ( .B1(n14191), .B2(n11489), .A(n14193), .ZN(n11488) );
  NAND2_X1 U12899 ( .A1(n15910), .A2(n11266), .ZN(n11490) );
  INV_X1 U12900 ( .A(n15564), .ZN(n11497) );
  NAND2_X1 U12901 ( .A1(n11497), .A2(n11498), .ZN(n15875) );
  NAND4_X1 U12902 ( .A1(n11790), .A2(n12725), .A3(n11791), .A4(n12720), .ZN(
        n11816) );
  NAND3_X1 U12903 ( .A1(n11506), .A2(n11505), .A3(n11503), .ZN(n15008) );
  NOR2_X1 U12904 ( .A1(n16726), .A2(n16720), .ZN(n16719) );
  INV_X1 U12905 ( .A(n16713), .ZN(n11514) );
  NAND2_X1 U12906 ( .A1(n12770), .A2(n11262), .ZN(n12708) );
  NAND2_X1 U12907 ( .A1(n12770), .A2(n11521), .ZN(n12699) );
  AND2_X1 U12908 ( .A1(n12770), .A2(n16694), .ZN(n12352) );
  INV_X1 U12909 ( .A(n15202), .ZN(n11527) );
  INV_X1 U12910 ( .A(n11529), .ZN(n13886) );
  NAND2_X1 U12911 ( .A1(n16661), .A2(n16660), .ZN(n16659) );
  NAND2_X1 U12912 ( .A1(n11553), .A2(n11249), .ZN(n15767) );
  INV_X1 U12913 ( .A(n11827), .ZN(n11572) );
  NAND2_X1 U12914 ( .A1(n11822), .A2(n11821), .ZN(n11575) );
  INV_X1 U12915 ( .A(n11836), .ZN(n11837) );
  NAND2_X1 U12916 ( .A1(n11827), .A2(n11575), .ZN(n11574) );
  NAND2_X1 U12917 ( .A1(n15814), .A2(n11233), .ZN(n11577) );
  NAND3_X1 U12918 ( .A1(n11579), .A2(n12390), .A3(n12382), .ZN(n11578) );
  OR2_X1 U12919 ( .A1(n11584), .A2(n17079), .ZN(n11582) );
  OR3_X1 U12920 ( .A1(n11584), .A2(n17079), .A3(n11277), .ZN(n11583) );
  NAND2_X1 U12921 ( .A1(n11806), .A2(n11785), .ZN(n11756) );
  AND2_X2 U12922 ( .A1(n11777), .A2(n11776), .ZN(n11586) );
  NAND2_X1 U12923 ( .A1(n11957), .A2(n11956), .ZN(n11588) );
  NAND2_X1 U12924 ( .A1(n11588), .A2(n12526), .ZN(n12364) );
  OAI21_X1 U12925 ( .B1(n11228), .B2(n11593), .A(n11591), .ZN(n11590) );
  NAND2_X1 U12926 ( .A1(n11600), .A2(n11597), .ZN(n11605) );
  OAI21_X1 U12927 ( .B1(n11606), .B2(n11217), .A(n11599), .ZN(n11598) );
  NAND2_X1 U12928 ( .A1(n16869), .A2(n11610), .ZN(n11602) );
  NAND3_X1 U12929 ( .A1(n11612), .A2(n22274), .A3(n14885), .ZN(n11611) );
  NAND2_X1 U12930 ( .A1(n11612), .A2(n14885), .ZN(n15337) );
  NAND3_X1 U12931 ( .A1(n13376), .A2(n11618), .A3(n13375), .ZN(n15884) );
  NAND3_X1 U12932 ( .A1(n13376), .A2(n13375), .A3(n11260), .ZN(n11617) );
  NAND2_X1 U12933 ( .A1(n13376), .A2(n13375), .ZN(n15646) );
  INV_X1 U12934 ( .A(n15704), .ZN(n11619) );
  NOR2_X1 U12935 ( .A1(n16070), .A2(n11625), .ZN(n16050) );
  NAND2_X1 U12936 ( .A1(n16085), .A2(n11623), .ZN(n13831) );
  NOR2_X1 U12937 ( .A1(n16070), .A2(n16071), .ZN(n16060) );
  INV_X1 U12938 ( .A(n16324), .ZN(n13240) );
  INV_X1 U12939 ( .A(n15082), .ZN(n13930) );
  AOI22_X1 U12940 ( .A1(n11668), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11734) );
  AOI22_X1 U12941 ( .A1(n11668), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11701) );
  XNOR2_X1 U12942 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12449) );
  INV_X1 U12943 ( .A(n19857), .ZN(n19851) );
  AOI22_X1 U12944 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n14156), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11712) );
  CLKBUF_X1 U12945 ( .A(n16894), .Z(n17154) );
  NAND2_X1 U12946 ( .A1(n16084), .A2(n11643), .ZN(n16070) );
  AND2_X2 U12947 ( .A1(n12846), .A2(n14872), .ZN(n13083) );
  AND4_X1 U12948 ( .A1(n11859), .A2(n11858), .A3(n11857), .A4(n11856), .ZN(
        n11882) );
  OAI22_X1 U12949 ( .A1(n11936), .A2(n19857), .B1(n11980), .B2(n14070), .ZN(
        n11937) );
  AND2_X2 U12950 ( .A1(n15441), .A2(n11861), .ZN(n19825) );
  AND2_X2 U12951 ( .A1(n15441), .A2(n11853), .ZN(n19800) );
  AND2_X1 U12952 ( .A1(n12754), .A2(n12753), .ZN(n12755) );
  NAND2_X1 U12953 ( .A1(n17847), .A2(n19204), .ZN(n12378) );
  AOI22_X1 U12954 ( .A1(n13185), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13083), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12898) );
  AOI22_X1 U12955 ( .A1(n11886), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11664) );
  NAND2_X1 U12957 ( .A1(n11192), .A2(n11870), .ZN(n11980) );
  AND2_X4 U12958 ( .A1(n11893), .A2(n19225), .ZN(n11886) );
  NAND2_X1 U12959 ( .A1(n11794), .A2(n11770), .ZN(n11758) );
  AOI21_X1 U12960 ( .B1(n12948), .B2(n11639), .A(n12947), .ZN(n12958) );
  CLKBUF_X1 U12961 ( .A(n14686), .Z(n16032) );
  NAND2_X1 U12962 ( .A1(n15047), .A2(n13350), .ZN(n15207) );
  AND4_X1 U12963 ( .A1(n12845), .A2(n12844), .A3(n12843), .A4(n12842), .ZN(
        n12855) );
  AOI22_X1 U12964 ( .A1(n19837), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11971), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11931) );
  AND2_X4 U12965 ( .A1(n12847), .A2(n12849), .ZN(n13013) );
  OR2_X1 U12966 ( .A1(n16621), .A2(n15177), .ZN(n22382) );
  NAND2_X1 U12967 ( .A1(n16621), .A2(n22274), .ZN(n13123) );
  AND2_X1 U12968 ( .A1(n13248), .A2(n13247), .ZN(n11630) );
  INV_X1 U12969 ( .A(n12022), .ZN(n12430) );
  NAND2_X1 U12970 ( .A1(n14809), .A2(n11773), .ZN(n11779) );
  OR2_X1 U12971 ( .A1(n16829), .A2(n19098), .ZN(n11632) );
  AND2_X1 U12972 ( .A1(n12797), .A2(n12796), .ZN(n11633) );
  OR3_X1 U12973 ( .A1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n17035), .A3(
        n17036), .ZN(n11634) );
  OR2_X1 U12974 ( .A1(n12752), .A2(n12751), .ZN(n11635) );
  NOR2_X1 U12975 ( .A1(n22372), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11636) );
  OR2_X1 U12976 ( .A1(n12493), .A2(n12144), .ZN(n11637) );
  INV_X2 U12977 ( .A(n18366), .ZN(n18362) );
  INV_X1 U12978 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12358) );
  INV_X1 U12979 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n13544) );
  AND2_X1 U12980 ( .A1(n14427), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11638) );
  OR2_X1 U12981 ( .A1(n15229), .A2(n14847), .ZN(n11639) );
  NAND4_X1 U12982 ( .A1(n12923), .A2(n12922), .A3(n12921), .A4(n12920), .ZN(
        n11640) );
  INV_X1 U12983 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14746) );
  INV_X1 U12984 ( .A(n11870), .ZN(n11871) );
  AND2_X1 U12985 ( .A1(n14212), .A2(n14230), .ZN(n11641) );
  OR2_X1 U12986 ( .A1(n17074), .A2(n17859), .ZN(n11642) );
  INV_X1 U12987 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13246) );
  AOI21_X1 U12988 ( .B1(n11792), .B2(n11816), .A(n19270), .ZN(n11823) );
  INV_X1 U12989 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n19172) );
  NAND2_X1 U12990 ( .A1(n20524), .A2(n16033), .ZN(n20510) );
  OR2_X1 U12991 ( .A1(n12232), .A2(n17079), .ZN(n16857) );
  INV_X1 U12992 ( .A(n16857), .ZN(n12765) );
  INV_X1 U12993 ( .A(n17860), .ZN(n12415) );
  INV_X1 U12994 ( .A(n12391), .ZN(n12381) );
  AND2_X1 U12995 ( .A1(n13728), .A2(n16158), .ZN(n11643) );
  NAND2_X1 U12996 ( .A1(n13009), .A2(n15229), .ZN(n13215) );
  INV_X1 U12997 ( .A(n13215), .ZN(n13010) );
  INV_X1 U12998 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n13443) );
  INV_X1 U12999 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12359) );
  INV_X1 U13000 ( .A(n19187), .ZN(n12758) );
  INV_X1 U13001 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n15869) );
  NAND2_X2 U13002 ( .A1(n13914), .A2(n13913), .ZN(n20524) );
  AND2_X1 U13003 ( .A1(n20900), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11644) );
  AND2_X1 U13004 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11645) );
  OR2_X1 U13005 ( .A1(n21135), .A2(n21134), .ZN(n11646) );
  AND4_X1 U13006 ( .A1(n11897), .A2(n11896), .A3(n11895), .A4(n11894), .ZN(
        n11647) );
  NOR2_X1 U13007 ( .A1(n14310), .A2(n14308), .ZN(n14372) );
  INV_X1 U13008 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n15575) );
  INV_X1 U13009 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n22435) );
  INV_X1 U13010 ( .A(n15786), .ZN(n22424) );
  AND2_X2 U13011 ( .A1(n22268), .A2(n13832), .ZN(n20588) );
  NAND2_X2 U13012 ( .A1(n16265), .A2(n14938), .ZN(n16238) );
  INV_X1 U13013 ( .A(n15532), .ZN(n15381) );
  NAND2_X2 U13014 ( .A1(n15378), .A2(n15377), .ZN(n15532) );
  OR2_X1 U13015 ( .A1(n12430), .A2(n12653), .ZN(n11648) );
  OR2_X1 U13016 ( .A1(n12510), .A2(n12509), .ZN(n11649) );
  AND2_X1 U13017 ( .A1(n14215), .A2(n11641), .ZN(n11650) );
  INV_X1 U13018 ( .A(n20555), .ZN(n16428) );
  AND2_X2 U13019 ( .A1(n17821), .A2(n15786), .ZN(n20555) );
  INV_X1 U13020 ( .A(n13668), .ZN(n13791) );
  INV_X1 U13021 ( .A(n16111), .ZN(n16229) );
  AND2_X1 U13022 ( .A1(n13433), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11651) );
  NAND2_X1 U13023 ( .A1(n20524), .A2(n13915), .ZN(n16189) );
  INV_X1 U13024 ( .A(n16189), .ZN(n13916) );
  AND2_X1 U13025 ( .A1(n13083), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11652) );
  AND4_X1 U13026 ( .A1(n12869), .A2(n12868), .A3(n12867), .A4(n12866), .ZN(
        n11653) );
  INV_X1 U13027 ( .A(n12955), .ZN(n13047) );
  AND2_X1 U13028 ( .A1(n12955), .A2(n13915), .ZN(n11654) );
  INV_X1 U13029 ( .A(n19754), .ZN(n12076) );
  AND2_X1 U13030 ( .A1(n12976), .A2(n14834), .ZN(n12977) );
  NAND2_X1 U13031 ( .A1(n12978), .A2(n12977), .ZN(n12979) );
  AND4_X1 U13032 ( .A1(n11976), .A2(n11975), .A3(n11974), .A4(n11973), .ZN(
        n11990) );
  AND2_X1 U13033 ( .A1(n22415), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13277) );
  OR2_X1 U13034 ( .A1(n13168), .A2(n13167), .ZN(n13197) );
  INV_X1 U13035 ( .A(n11947), .ZN(n11948) );
  INV_X1 U13036 ( .A(n12418), .ZN(n12419) );
  AND2_X1 U13037 ( .A1(n17827), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13267) );
  OR2_X1 U13038 ( .A1(n13146), .A2(n13145), .ZN(n13150) );
  INV_X1 U13039 ( .A(n13725), .ZN(n13707) );
  INV_X1 U13040 ( .A(n15927), .ZN(n13441) );
  OAI22_X1 U13041 ( .A1(n13302), .A2(n13170), .B1(n13283), .B2(n13169), .ZN(
        n13179) );
  NAND2_X1 U13042 ( .A1(n12984), .A2(n12980), .ZN(n13073) );
  AOI22_X1 U13043 ( .A1(n13082), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13018), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12868) );
  AOI22_X1 U13044 ( .A1(n13185), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11165), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12888) );
  INV_X1 U13045 ( .A(n12043), .ZN(n12028) );
  NOR2_X1 U13046 ( .A1(n11949), .A2(n11948), .ZN(n11951) );
  AND2_X1 U13047 ( .A1(n12111), .A2(n12110), .ZN(n12399) );
  OAI22_X1 U13048 ( .A1(n11237), .A2(n12500), .B1(n12541), .B2(n14746), .ZN(
        n12501) );
  XNOR2_X1 U13049 ( .A(n11716), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12042) );
  AOI22_X1 U13050 ( .A1(n11668), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11170), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11719) );
  OR2_X1 U13051 ( .A1(n13295), .A2(n13267), .ZN(n13268) );
  INV_X1 U13052 ( .A(n13150), .ZN(n13171) );
  INV_X1 U13053 ( .A(n13747), .ZN(n13748) );
  NAND2_X1 U13054 ( .A1(n13427), .A2(n13441), .ZN(n13442) );
  OR2_X1 U13055 ( .A1(n13042), .A2(n13041), .ZN(n13219) );
  OR2_X1 U13056 ( .A1(n13191), .A2(n13190), .ZN(n13208) );
  INV_X1 U13057 ( .A(n13194), .ZN(n13192) );
  INV_X1 U13058 ( .A(n13081), .ZN(n13046) );
  AND4_X1 U13059 ( .A1(n12017), .A2(n12016), .A3(n12015), .A4(n12014), .ZN(
        n12019) );
  AND2_X1 U13060 ( .A1(n12671), .A2(n12670), .ZN(n16786) );
  INV_X1 U13061 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12384) );
  NAND2_X1 U13062 ( .A1(n11148), .A2(n12364), .ZN(n12375) );
  NAND2_X1 U13063 ( .A1(n14815), .A2(n12650), .ZN(n12512) );
  OR2_X1 U13064 ( .A1(n14437), .A2(n14438), .ZN(n14433) );
  NAND2_X1 U13065 ( .A1(n13268), .A2(n13294), .ZN(n14691) );
  NAND2_X1 U13066 ( .A1(n14838), .A2(n13918), .ZN(n13925) );
  NOR2_X1 U13067 ( .A1(n13771), .A2(n13770), .ZN(n13772) );
  INV_X1 U13068 ( .A(n16228), .ZN(n13624) );
  AND2_X1 U13069 ( .A1(n16134), .A2(n15929), .ZN(n13476) );
  INV_X1 U13070 ( .A(n15922), .ZN(n13426) );
  AND2_X1 U13071 ( .A1(n15575), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13827) );
  NAND2_X1 U13072 ( .A1(n15093), .A2(n12996), .ZN(n15454) );
  INV_X1 U13073 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17802) );
  NOR2_X1 U13074 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17769), .ZN(
        n12248) );
  NOR2_X1 U13075 ( .A1(n12493), .A2(n12146), .ZN(n12161) );
  INV_X1 U13076 ( .A(n15055), .ZN(n12297) );
  INV_X1 U13077 ( .A(n15039), .ZN(n12626) );
  AND2_X1 U13078 ( .A1(n16976), .A2(n16974), .ZN(n12799) );
  AND2_X1 U13079 ( .A1(n12049), .A2(n12531), .ZN(n12113) );
  AND3_X1 U13080 ( .A1(n15013), .A2(n11649), .A3(n12514), .ZN(n12515) );
  OAI211_X1 U13081 ( .C1(n14667), .C2(n12653), .A(n12512), .B(n12495), .ZN(
        n14820) );
  INV_X1 U13082 ( .A(n11887), .ZN(n11888) );
  AND2_X1 U13083 ( .A1(n17768), .A2(n19282), .ZN(n19760) );
  OAI21_X1 U13084 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n21371), .A(
        n14433), .ZN(n14434) );
  AOI21_X1 U13085 ( .B1(n21827), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n14432), .ZN(n14438) );
  AND2_X1 U13086 ( .A1(n18548), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14428) );
  OR2_X1 U13087 ( .A1(n18548), .A2(n21495), .ZN(n14418) );
  INV_X2 U13088 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17368) );
  INV_X1 U13089 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18281) );
  INV_X1 U13090 ( .A(n15238), .ZN(n15233) );
  INV_X1 U13091 ( .A(n15865), .ZN(n13947) );
  INV_X1 U13092 ( .A(n15936), .ZN(n13493) );
  OR2_X1 U13093 ( .A1(n13750), .A2(n13749), .ZN(n13771) );
  AND2_X1 U13094 ( .A1(n13727), .A2(n13726), .ZN(n16158) );
  OR2_X1 U13095 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n13668) );
  INV_X1 U13096 ( .A(n13471), .ZN(n13503) );
  OAI21_X1 U13097 ( .B1(n13302), .B2(n13051), .A(n13050), .ZN(n13064) );
  AOI221_X1 U13098 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n12249), 
        .C1(n19172), .C2(n12249), .A(n12248), .ZN(n12465) );
  AND2_X1 U13099 ( .A1(n15058), .A2(n15056), .ZN(n14037) );
  NAND2_X1 U13100 ( .A1(n14011), .A2(n19916), .ZN(n14027) );
  OR2_X1 U13101 ( .A1(n14211), .A2(n14213), .ZN(n14230) );
  NOR2_X1 U13102 ( .A1(n12736), .A2(n19241), .ZN(n17171) );
  INV_X1 U13103 ( .A(n14235), .ZN(n11771) );
  INV_X1 U13104 ( .A(n11979), .ZN(n19842) );
  AOI21_X1 U13105 ( .B1(n19279), .B2(n19270), .A(n19760), .ZN(n19751) );
  NOR2_X1 U13106 ( .A1(n11646), .A2(n21131), .ZN(n21136) );
  OR2_X1 U13107 ( .A1(n21204), .A2(n14385), .ZN(n14384) );
  INV_X1 U13108 ( .A(n21232), .ZN(n14548) );
  INV_X1 U13109 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n13665) );
  INV_X1 U13110 ( .A(n22235), .ZN(n22254) );
  INV_X1 U13111 ( .A(n22244), .ZN(n22256) );
  AND2_X1 U13112 ( .A1(n13950), .A2(n13949), .ZN(n15888) );
  OR2_X1 U13113 ( .A1(n21878), .A2(n21876), .ZN(n15377) );
  AND2_X1 U13114 ( .A1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n13580), .ZN(
        n13618) );
  NOR2_X1 U13115 ( .A1(n13459), .A2(n13443), .ZN(n13478) );
  AND2_X1 U13116 ( .A1(n16437), .A2(n16436), .ZN(n16531) );
  INV_X1 U13117 ( .A(n15081), .ZN(n13929) );
  INV_X1 U13118 ( .A(n16620), .ZN(n16607) );
  NAND2_X1 U13119 ( .A1(n15291), .A2(n15568), .ZN(n22640) );
  INV_X1 U13120 ( .A(n22671), .ZN(n22639) );
  INV_X1 U13121 ( .A(n22554), .ZN(n22535) );
  INV_X1 U13122 ( .A(n17343), .ZN(n19239) );
  NAND2_X1 U13123 ( .A1(n18852), .A2(n13893), .ZN(n19151) );
  INV_X1 U13124 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13846) );
  XNOR2_X1 U13125 ( .A(n12787), .B(n12688), .ZN(n19158) );
  OR2_X1 U13126 ( .A1(n14136), .A2(n14135), .ZN(n14155) );
  INV_X1 U13127 ( .A(n20062), .ZN(n16819) );
  INV_X1 U13128 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n19076) );
  INV_X1 U13129 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16965) );
  OR2_X1 U13130 ( .A1(n17309), .A2(n12739), .ZN(n17211) );
  AND3_X1 U13131 ( .A1(n12611), .A2(n12610), .A3(n12609), .ZN(n15847) );
  OR2_X1 U13132 ( .A1(n15850), .A2(n12185), .ZN(n16974) );
  INV_X1 U13133 ( .A(n12260), .ZN(n12469) );
  AND2_X1 U13134 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19897) );
  INV_X1 U13135 ( .A(n19944), .ZN(n19902) );
  INV_X1 U13136 ( .A(n19879), .ZN(n17899) );
  NAND2_X1 U13137 ( .A1(n19270), .A2(n19256), .ZN(n19261) );
  NOR2_X1 U13138 ( .A1(n21137), .A2(n21136), .ZN(n21138) );
  NOR2_X1 U13139 ( .A1(n21010), .A2(n21128), .ZN(n21013) );
  NOR2_X1 U13140 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n20942), .ZN(n20957) );
  NOR2_X1 U13141 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n20891), .ZN(n20904) );
  OR4_X1 U13142 ( .A1(n15954), .A2(n20825), .A3(n18031), .A4(n15953), .ZN(
        n15955) );
  INV_X1 U13143 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n20825) );
  NOR2_X1 U13144 ( .A1(n14617), .A2(n21093), .ZN(n18531) );
  INV_X1 U13145 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n21064) );
  NOR2_X1 U13146 ( .A1(n18405), .A2(n21555), .ZN(n21729) );
  OR2_X1 U13147 ( .A1(n18665), .A2(n18548), .ZN(n18402) );
  OR4_X1 U13148 ( .A1(n18394), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18446) );
  NOR2_X1 U13149 ( .A1(n14579), .A2(n18734), .ZN(n18725) );
  NOR2_X1 U13150 ( .A1(n14502), .A2(n14501), .ZN(n20736) );
  AOI211_X1 U13151 ( .C1(n11143), .C2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n14509), .B(n14508), .ZN(n14510) );
  INV_X1 U13152 ( .A(n21809), .ZN(n21457) );
  OR2_X1 U13153 ( .A1(n16039), .A2(n22283), .ZN(n14782) );
  OR3_X1 U13154 ( .A1(n16101), .A2(n16310), .A3(n20464), .ZN(n16092) );
  OR2_X1 U13155 ( .A1(n13666), .A2(n13665), .ZN(n13725) );
  NAND2_X1 U13156 ( .A1(n13424), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13459) );
  INV_X1 U13157 ( .A(n22092), .ZN(n22197) );
  INV_X1 U13158 ( .A(n22236), .ZN(n22220) );
  NOR2_X1 U13159 ( .A1(n20524), .A2(n16043), .ZN(n14006) );
  AND2_X1 U13160 ( .A1(n13992), .A2(n13991), .ZN(n16106) );
  INV_X1 U13161 ( .A(n20510), .ZN(n20528) );
  AOI21_X1 U13162 ( .B1(n15378), .B2(n14934), .A(n14933), .ZN(n14935) );
  NOR2_X2 U13163 ( .A1(n15532), .A2(n15379), .ZN(n15522) );
  AND2_X1 U13164 ( .A1(n13368), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13392) );
  NAND2_X1 U13165 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n13320), .ZN(
        n13359) );
  NOR2_X1 U13166 ( .A1(n16036), .A2(n22283), .ZN(n15063) );
  NAND2_X1 U13167 ( .A1(n16596), .A2(n22274), .ZN(n13838) );
  OR2_X1 U13168 ( .A1(n21944), .A2(n21925), .ZN(n21933) );
  AND2_X1 U13169 ( .A1(n14923), .A2(n16030), .ZN(n22007) );
  AND2_X1 U13170 ( .A1(n14966), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n15335) );
  OR2_X1 U13171 ( .A1(n14862), .A2(n14931), .ZN(n17803) );
  INV_X1 U13172 ( .A(n22623), .ZN(n22589) );
  INV_X1 U13173 ( .A(n22592), .ZN(n22633) );
  OAI21_X1 U13174 ( .B1(n15658), .B2(n15662), .A(n22439), .ZN(n15684) );
  AND2_X1 U13175 ( .A1(n15291), .A2(n13338), .ZN(n15688) );
  OAI211_X1 U13176 ( .C1(n15786), .C2(n22398), .A(n15104), .B(n22387), .ZN(
        n15172) );
  AND2_X1 U13177 ( .A1(n15087), .A2(n15568), .ZN(n22531) );
  INV_X1 U13178 ( .A(n22652), .ZN(n15780) );
  NOR2_X1 U13179 ( .A1(n15572), .A2(n14966), .ZN(n15569) );
  NOR2_X2 U13180 ( .A1(n15572), .A2(n22369), .ZN(n22654) );
  NOR2_X1 U13181 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15099), .ZN(n15124) );
  OAI211_X1 U13182 ( .C1(n15786), .C2(n15460), .A(n22387), .B(n15459), .ZN(
        n15539) );
  NOR2_X1 U13183 ( .A1(n15782), .A2(n15496), .ZN(n16638) );
  NOR2_X1 U13184 ( .A1(n15782), .A2(n15559), .ZN(n16648) );
  NOR2_X1 U13185 ( .A1(n15168), .A2(n16033), .ZN(n22671) );
  AND2_X1 U13186 ( .A1(n17825), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13312) );
  INV_X1 U13187 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n22311) );
  INV_X1 U13188 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n22312) );
  INV_X1 U13189 ( .A(n20466), .ZN(n20470) );
  OAI21_X1 U13190 ( .B1(n13902), .B2(n19149), .A(n13901), .ZN(n13903) );
  AND2_X1 U13191 ( .A1(n14675), .A2(n13897), .ZN(n19135) );
  INV_X1 U13192 ( .A(n19151), .ZN(n19134) );
  INV_X1 U13193 ( .A(n19149), .ZN(n19136) );
  NOR2_X1 U13194 ( .A1(n14659), .A2(n19257), .ZN(n19159) );
  INV_X1 U13195 ( .A(n19287), .ZN(n18854) );
  OR2_X1 U13196 ( .A1(n14125), .A2(n14124), .ZN(n16723) );
  INV_X1 U13197 ( .A(n16740), .ZN(n16732) );
  OR2_X1 U13198 ( .A1(n14047), .A2(n14046), .ZN(n15693) );
  INV_X1 U13199 ( .A(n14788), .ZN(n14775) );
  NAND2_X1 U13200 ( .A1(n19161), .A2(n17878), .ZN(n14299) );
  OAI21_X1 U13201 ( .B1(n12834), .B2(n17860), .A(n12818), .ZN(n12819) );
  AND2_X1 U13202 ( .A1(n17029), .A2(n14670), .ZN(n17850) );
  AND2_X1 U13203 ( .A1(n16726), .A2(n16725), .ZN(n19065) );
  NOR2_X1 U13204 ( .A1(n16987), .A2(n17228), .ZN(n16980) );
  AND2_X1 U13205 ( .A1(n15594), .A2(n15593), .ZN(n19207) );
  INV_X1 U13206 ( .A(n12365), .ZN(n14667) );
  NAND2_X1 U13207 ( .A1(n19242), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17365) );
  INV_X1 U13208 ( .A(n20344), .ZN(n20353) );
  AND2_X1 U13209 ( .A1(n19929), .A2(n19915), .ZN(n20340) );
  INV_X1 U13210 ( .A(n20324), .ZN(n20326) );
  OAI21_X1 U13211 ( .B1(n19892), .B2(n19891), .A(n19890), .ZN(n20320) );
  INV_X1 U13212 ( .A(n20317), .ZN(n20308) );
  AND2_X1 U13213 ( .A1(n19866), .A2(n19895), .ZN(n20220) );
  INV_X1 U13214 ( .A(n20219), .ZN(n20301) );
  INV_X1 U13215 ( .A(n20298), .ZN(n20211) );
  OAI21_X1 U13216 ( .B1(n19816), .B2(n19815), .A(n19814), .ZN(n20282) );
  AND2_X1 U13217 ( .A1(n19819), .A2(n19895), .ZN(n20208) );
  NOR2_X1 U13218 ( .A1(n19880), .A2(n17899), .ZN(n19819) );
  INV_X1 U13219 ( .A(n20345), .ZN(n20349) );
  AOI21_X1 U13220 ( .B1(n20255), .B2(n19919), .A(n19772), .ZN(n20258) );
  NOR2_X1 U13221 ( .A1(n19880), .A2(n19879), .ZN(n19768) );
  NAND2_X1 U13222 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n17768) );
  INV_X1 U13223 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n22328) );
  XOR2_X1 U13224 ( .A(n20738), .B(n18807), .Z(n20671) );
  AOI211_X1 U13225 ( .C1(n14444), .C2(n14443), .A(n14539), .B(n14442), .ZN(
        n21813) );
  NOR2_X1 U13226 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n21079), .ZN(n21097) );
  AND2_X1 U13227 ( .A1(n21075), .A2(n21078), .ZN(n21089) );
  NOR2_X1 U13228 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n21004), .ZN(n21019) );
  NOR2_X1 U13229 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n20977), .ZN(n20993) );
  NOR2_X1 U13230 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n20862), .ZN(n20882) );
  NOR2_X1 U13231 ( .A1(n21803), .A2(n20859), .ZN(n20886) );
  INV_X1 U13232 ( .A(n21146), .ZN(n21127) );
  OAI211_X2 U13233 ( .C1(n21857), .C2(n21856), .A(n20746), .B(n20745), .ZN(
        n21077) );
  NOR2_X1 U13234 ( .A1(n21267), .A2(n18241), .ZN(n18279) );
  INV_X1 U13235 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n20992) );
  NAND2_X1 U13236 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n18128), .ZN(n18127) );
  INV_X1 U13237 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n20798) );
  NAND4_X1 U13238 ( .A1(n21845), .A2(n18807), .A3(n20741), .A4(n21165), .ZN(
        n18365) );
  NOR2_X1 U13239 ( .A1(n21255), .A2(n21260), .ZN(n21254) );
  NOR2_X1 U13240 ( .A1(n21267), .A2(n21314), .ZN(n21261) );
  INV_X1 U13241 ( .A(n20736), .ZN(n18807) );
  NOR2_X1 U13242 ( .A1(n17756), .A2(n20735), .ZN(n17755) );
  INV_X1 U13243 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n21093) );
  NAND2_X1 U13244 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21565), .ZN(
        n21567) );
  NOR2_X2 U13245 ( .A1(n21653), .A2(n18757), .ZN(n18661) );
  NOR2_X1 U13246 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19317), .ZN(n19640) );
  NAND2_X1 U13247 ( .A1(n21670), .A2(n18535), .ZN(n21671) );
  AND2_X1 U13248 ( .A1(n21725), .A2(n21799), .ZN(n21753) );
  INV_X1 U13249 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n21763) );
  NAND2_X1 U13250 ( .A1(n18699), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18698) );
  NOR2_X1 U13251 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n17758), .ZN(n14606) );
  INV_X1 U13252 ( .A(n19640), .ZN(n19552) );
  NOR2_X1 U13253 ( .A1(n21855), .A2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n21367) );
  INV_X1 U13254 ( .A(n19620), .ZN(n19717) );
  INV_X1 U13255 ( .A(n19679), .ZN(n19692) );
  INV_X1 U13256 ( .A(n19609), .ZN(n19686) );
  INV_X1 U13257 ( .A(n19341), .ZN(n19342) );
  INV_X1 U13258 ( .A(n19656), .ZN(n19669) );
  INV_X1 U13259 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n22301) );
  INV_X1 U13260 ( .A(n22352), .ZN(n22341) );
  NOR2_X1 U13261 ( .A1(n22301), .A2(n18843), .ZN(n18837) );
  INV_X1 U13262 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n22345) );
  NOR2_X1 U13263 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n14656), .ZN(n19636)
         );
  INV_X1 U13264 ( .A(n15378), .ZN(n14783) );
  INV_X1 U13265 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n22286) );
  INV_X1 U13266 ( .A(n22262), .ZN(n22246) );
  NOR2_X1 U13267 ( .A1(n14007), .A2(n14006), .ZN(n14008) );
  INV_X1 U13268 ( .A(n16277), .ZN(n16197) );
  INV_X1 U13269 ( .A(n22263), .ZN(n16219) );
  OR2_X1 U13270 ( .A1(n16135), .A2(n15931), .ZN(n22159) );
  AND2_X1 U13271 ( .A1(n15091), .A2(n15090), .ZN(n15649) );
  AND2_X1 U13272 ( .A1(n15052), .A2(n15051), .ZN(n15496) );
  NAND2_X1 U13273 ( .A1(n20414), .A2(n16021), .ZN(n15623) );
  INV_X1 U13274 ( .A(n20414), .ZN(n20437) );
  NAND2_X1 U13275 ( .A1(n15378), .A2(n15379), .ZN(n15529) );
  INV_X1 U13276 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21949) );
  INV_X1 U13277 ( .A(n22056), .ZN(n22033) );
  INV_X1 U13278 ( .A(n22053), .ZN(n22031) );
  INV_X1 U13279 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17827) );
  AOI22_X1 U13280 ( .A1(n22359), .A2(n22364), .B1(n22358), .B2(n22412), .ZN(
        n22621) );
  AOI22_X1 U13281 ( .A1(n22373), .A2(n22377), .B1(n22412), .B2(n11636), .ZN(
        n22628) );
  AOI22_X1 U13282 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n22388), .B1(n22386), 
        .B2(n22391), .ZN(n22637) );
  OR2_X1 U13283 ( .A1(n22370), .A2(n15655), .ZN(n22631) );
  AOI21_X1 U13284 ( .B1(n15657), .B2(n15290), .A(n15289), .ZN(n15327) );
  AOI22_X1 U13285 ( .A1(n22397), .A2(n22405), .B1(n22430), .B2(n11636), .ZN(
        n22646) );
  INV_X1 U13286 ( .A(n22642), .ZN(n15175) );
  NAND2_X1 U13287 ( .A1(n15569), .A2(n15568), .ZN(n22604) );
  AOI22_X1 U13288 ( .A1(n22413), .A2(n22420), .B1(n22412), .B2(n22411), .ZN(
        n22659) );
  INV_X1 U13289 ( .A(n22663), .ZN(n22546) );
  INV_X1 U13290 ( .A(n16628), .ZN(n22445) );
  INV_X1 U13291 ( .A(n16648), .ZN(n22613) );
  INV_X1 U13292 ( .A(n22556), .ZN(n15542) );
  INV_X1 U13293 ( .A(n22547), .ZN(n22560) );
  OR2_X1 U13294 ( .A1(n15458), .A2(n22369), .ZN(n22680) );
  INV_X1 U13295 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n17825) );
  INV_X1 U13296 ( .A(n22287), .ZN(n22289) );
  NAND2_X1 U13297 ( .A1(n13890), .A2(n19245), .ZN(n18852) );
  INV_X1 U13298 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n22292) );
  OR3_X1 U13299 ( .A1(n18852), .A2(n13906), .A3(n13891), .ZN(n19149) );
  INV_X1 U13300 ( .A(n19157), .ZN(n19121) );
  INV_X1 U13301 ( .A(n19159), .ZN(n19133) );
  AND2_X1 U13302 ( .A1(n14290), .A2(n18854), .ZN(n16727) );
  NAND2_X1 U13303 ( .A1(n16727), .A2(n19758), .ZN(n16740) );
  INV_X1 U13304 ( .A(n20060), .ZN(n16817) );
  NAND2_X1 U13305 ( .A1(n16817), .A2(n14816), .ZN(n16818) );
  NAND2_X1 U13306 ( .A1(n17918), .A2(n11768), .ZN(n14959) );
  INV_X1 U13307 ( .A(n17918), .ZN(n17951) );
  OAI21_X1 U13308 ( .B1(n14674), .B2(n22321), .A(n14788), .ZN(n14749) );
  CLKBUF_X1 U13309 ( .A(n14749), .Z(n14780) );
  NAND2_X1 U13310 ( .A1(n22685), .A2(n12415), .ZN(n12416) );
  NOR2_X1 U13311 ( .A1(n16938), .A2(n17177), .ZN(n17179) );
  OR2_X1 U13312 ( .A1(n19290), .A2(n13896), .ZN(n17860) );
  INV_X1 U13313 ( .A(n12835), .ZN(n12836) );
  OR2_X1 U13314 ( .A1(n17305), .A2(n17304), .ZN(n17858) );
  NAND2_X1 U13315 ( .A1(n12757), .A2(n19233), .ZN(n19178) );
  NAND2_X1 U13316 ( .A1(n12757), .A2(n19235), .ZN(n19187) );
  INV_X1 U13317 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19809) );
  INV_X1 U13318 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n20243) );
  AOI21_X1 U13319 ( .B1(n19950), .B2(n19949), .A(n20244), .ZN(n20357) );
  INV_X1 U13320 ( .A(n20340), .ZN(n20235) );
  NAND2_X1 U13321 ( .A1(n19896), .A2(n19895), .ZN(n20336) );
  NAND2_X1 U13322 ( .A1(n19896), .A2(n19881), .ZN(n20324) );
  NAND2_X1 U13323 ( .A1(n19866), .A2(n19855), .ZN(n20317) );
  INV_X1 U13324 ( .A(n20220), .ZN(n20311) );
  NAND2_X1 U13325 ( .A1(n19866), .A2(n19881), .ZN(n20219) );
  NAND2_X1 U13326 ( .A1(n19819), .A2(n19865), .ZN(n20298) );
  NAND2_X1 U13327 ( .A1(n19819), .A2(n19855), .ZN(n20214) );
  INV_X1 U13328 ( .A(n20208), .ZN(n20286) );
  AOI22_X1 U13329 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n20250), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n20251), .ZN(n20187) );
  NAND2_X1 U13330 ( .A1(n19881), .A2(n19819), .ZN(n20274) );
  AOI22_X1 U13331 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20251), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n20250), .ZN(n20337) );
  AOI22_X1 U13332 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n20250), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n20251), .ZN(n20138) );
  AOI22_X1 U13333 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20251), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n20250), .ZN(n19924) );
  AOI22_X1 U13334 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20251), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n20250), .ZN(n20105) );
  INV_X1 U13335 ( .A(n22295), .ZN(n17765) );
  AND2_X1 U13336 ( .A1(n17984), .A2(n17953), .ZN(n22332) );
  NAND2_X1 U13337 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n21354), .ZN(n21857) );
  INV_X1 U13338 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n22296) );
  INV_X1 U13339 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n21058) );
  INV_X1 U13340 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n20973) );
  NAND2_X1 U13341 ( .A1(n21077), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n21146) );
  AND2_X1 U13342 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n18267), .ZN(n18262) );
  NOR2_X1 U13343 ( .A1(n20992), .A2(n18324), .ZN(n18340) );
  AND2_X1 U13344 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17999), .ZN(n18128) );
  INV_X1 U13345 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18184) );
  INV_X1 U13346 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18195) );
  INV_X1 U13347 ( .A(n21333), .ZN(n21324) );
  NOR2_X1 U13348 ( .A1(n21179), .A2(n21186), .ZN(n21183) );
  NOR2_X1 U13349 ( .A1(n14316), .A2(n14315), .ZN(n21204) );
  NAND2_X1 U13350 ( .A1(n18808), .A2(n18807), .ZN(n18826) );
  NAND2_X1 U13351 ( .A1(n17755), .A2(n20681), .ZN(n18806) );
  NOR2_X1 U13352 ( .A1(n18562), .A2(n18593), .ZN(n18740) );
  INV_X1 U13353 ( .A(n21739), .ZN(n21693) );
  INV_X1 U13354 ( .A(n21801), .ZN(n21770) );
  INV_X1 U13355 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21825) );
  INV_X1 U13356 ( .A(n19724), .ZN(n19715) );
  INV_X1 U13357 ( .A(n19704), .ZN(n19696) );
  INV_X1 U13358 ( .A(n19698), .ZN(n19690) );
  INV_X1 U13359 ( .A(n19681), .ZN(n19673) );
  INV_X1 U13360 ( .A(n19663), .ZN(n19650) );
  INV_X1 U13361 ( .A(n19583), .ZN(n19592) );
  INV_X1 U13362 ( .A(n19658), .ZN(n19556) );
  INV_X1 U13363 ( .A(n20970), .ZN(n21851) );
  NAND2_X1 U13364 ( .A1(n18843), .A2(n18827), .ZN(n17752) );
  INV_X1 U13365 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n21440) );
  INV_X1 U13366 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n21464) );
  AND2_X2 U13367 ( .A1(n14644), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n15987)
         );
  OAI211_X1 U13368 ( .C1(n17860), .C2(n17077), .A(n11642), .B(n12777), .ZN(
        P2_U2988) );
  AOI22_X1 U13369 ( .A1(n11188), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11658) );
  AND2_X4 U13370 ( .A1(n11891), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14139) );
  AOI22_X1 U13371 ( .A1(n11884), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14139), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11657) );
  AOI22_X1 U13372 ( .A1(n11886), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11170), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11656) );
  AND2_X4 U13373 ( .A1(n12255), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11883) );
  AND2_X4 U13374 ( .A1(n12255), .A2(n12054), .ZN(n14156) );
  AOI22_X1 U13375 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n14156), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11655) );
  NAND4_X1 U13376 ( .A1(n11658), .A2(n11657), .A3(n11656), .A4(n11655), .ZN(
        n11659) );
  NAND2_X1 U13377 ( .A1(n11659), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11667) );
  AOI22_X1 U13378 ( .A1(n11186), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14139), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11663) );
  AOI22_X1 U13379 ( .A1(n11884), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11662) );
  AOI22_X1 U13380 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n14156), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11661) );
  NAND4_X1 U13381 ( .A1(n11664), .A2(n11663), .A3(n11662), .A4(n11661), .ZN(
        n11665) );
  NAND2_X1 U13382 ( .A1(n11665), .A2(n11716), .ZN(n11666) );
  INV_X2 U13383 ( .A(n11784), .ZN(n11772) );
  AOI22_X1 U13384 ( .A1(n11668), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11670) );
  AOI22_X1 U13385 ( .A1(n11884), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11886), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11669) );
  NAND2_X1 U13386 ( .A1(n11670), .A2(n11669), .ZN(n11674) );
  AOI22_X1 U13387 ( .A1(n11188), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14139), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11672) );
  AOI22_X1 U13388 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n14156), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11671) );
  NAND2_X1 U13389 ( .A1(n11672), .A2(n11671), .ZN(n11673) );
  OAI21_X2 U13390 ( .B1(n11674), .B2(n11673), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11681) );
  AOI22_X1 U13391 ( .A1(n11884), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11886), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11678) );
  AOI22_X1 U13392 ( .A1(n11668), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11170), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11677) );
  AOI22_X1 U13393 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14156), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11676) );
  AOI22_X1 U13394 ( .A1(n11186), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14139), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11675) );
  NAND4_X1 U13395 ( .A1(n11678), .A2(n11677), .A3(n11676), .A4(n11675), .ZN(
        n11679) );
  NAND2_X1 U13396 ( .A1(n11679), .A2(n11716), .ZN(n11680) );
  NAND2_X1 U13397 ( .A1(n11772), .A2(n11182), .ZN(n11763) );
  AOI22_X1 U13398 ( .A1(n11884), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11886), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11683) );
  AOI22_X1 U13399 ( .A1(n11668), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11170), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11682) );
  AOI22_X1 U13400 ( .A1(n11186), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14139), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11685) );
  AOI22_X1 U13401 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n14156), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11684) );
  NAND3_X1 U13402 ( .A1(n11225), .A2(n11685), .A3(n11684), .ZN(n11691) );
  AOI22_X1 U13403 ( .A1(n11186), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14139), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11687) );
  AOI22_X1 U13404 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n14156), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11686) );
  AOI22_X1 U13405 ( .A1(n11668), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11689) );
  AOI22_X1 U13406 ( .A1(n11884), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11886), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11688) );
  NAND3_X1 U13407 ( .A1(n11226), .A2(n11689), .A3(n11688), .ZN(n11690) );
  AOI22_X1 U13408 ( .A1(n11884), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11886), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11695) );
  AOI22_X1 U13409 ( .A1(n11188), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n14139), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11694) );
  AOI22_X1 U13410 ( .A1(n11668), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11170), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11693) );
  AOI22_X1 U13411 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14156), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11692) );
  AOI22_X1 U13412 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n14156), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11696) );
  AOI22_X1 U13413 ( .A1(n11668), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11170), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11699) );
  AOI22_X1 U13414 ( .A1(n11187), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14139), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11698) );
  AOI22_X1 U13415 ( .A1(n11884), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11886), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11697) );
  AOI22_X1 U13416 ( .A1(n11884), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11886), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11703) );
  AOI22_X1 U13417 ( .A1(n11187), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14139), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11702) );
  AOI22_X1 U13418 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n14156), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11700) );
  NAND4_X1 U13419 ( .A1(n11703), .A2(n11702), .A3(n11701), .A4(n11700), .ZN(
        n11704) );
  NAND2_X1 U13420 ( .A1(n11704), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11711) );
  AOI22_X1 U13421 ( .A1(n11884), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11886), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11708) );
  AOI22_X1 U13422 ( .A1(n11187), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n14139), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11707) );
  AOI22_X1 U13423 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n14156), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11706) );
  AOI22_X1 U13424 ( .A1(n11668), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11705) );
  NAND4_X1 U13425 ( .A1(n11708), .A2(n11707), .A3(n11706), .A4(n11705), .ZN(
        n11709) );
  NAND2_X1 U13426 ( .A1(n11709), .A2(n11716), .ZN(n11710) );
  AOI22_X1 U13427 ( .A1(n11884), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11886), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11715) );
  AOI22_X1 U13428 ( .A1(n11187), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n14139), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11714) );
  AOI22_X1 U13429 ( .A1(n11668), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11713) );
  NAND4_X1 U13430 ( .A1(n11715), .A2(n11714), .A3(n11713), .A4(n11712), .ZN(
        n11717) );
  AOI22_X1 U13431 ( .A1(n11884), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11886), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11721) );
  AOI22_X1 U13432 ( .A1(n11186), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14139), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11720) );
  AOI22_X1 U13433 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n14156), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11718) );
  NAND4_X1 U13434 ( .A1(n11721), .A2(n11720), .A3(n11719), .A4(n11718), .ZN(
        n11722) );
  NAND3_X1 U13435 ( .A1(n11725), .A2(n11727), .A3(n11789), .ZN(n11740) );
  AOI22_X1 U13436 ( .A1(n11884), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11886), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11731) );
  AOI22_X1 U13437 ( .A1(n11188), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14139), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11730) );
  AOI22_X1 U13438 ( .A1(n11668), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11729) );
  AOI22_X1 U13439 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14156), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11728) );
  NAND4_X1 U13440 ( .A1(n11731), .A2(n11730), .A3(n11729), .A4(n11728), .ZN(
        n11732) );
  NAND2_X1 U13441 ( .A1(n11732), .A2(n11716), .ZN(n11739) );
  AOI22_X1 U13442 ( .A1(n11884), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11886), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11736) );
  AOI22_X1 U13443 ( .A1(n11188), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14139), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11735) );
  AOI22_X1 U13444 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n14156), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11733) );
  NAND4_X1 U13445 ( .A1(n11736), .A2(n11735), .A3(n11734), .A4(n11733), .ZN(
        n11737) );
  NAND2_X1 U13446 ( .A1(n11737), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11738) );
  NAND3_X1 U13447 ( .A1(n11740), .A2(n11778), .A3(n11785), .ZN(n12728) );
  NOR2_X1 U13448 ( .A1(n19758), .A2(n11182), .ZN(n11742) );
  AOI22_X1 U13449 ( .A1(n11884), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11886), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11747) );
  AOI22_X1 U13450 ( .A1(n11187), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14139), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11746) );
  AOI22_X1 U13451 ( .A1(n11668), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11745) );
  AOI22_X1 U13452 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n14156), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11744) );
  NAND4_X1 U13453 ( .A1(n11747), .A2(n11746), .A3(n11745), .A4(n11744), .ZN(
        n11748) );
  NAND2_X1 U13454 ( .A1(n11748), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11755) );
  AOI22_X1 U13455 ( .A1(n11884), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11886), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11752) );
  AOI22_X1 U13456 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n11186), .B1(
        n14139), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11751) );
  AOI22_X1 U13457 ( .A1(n11668), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11750) );
  AOI22_X1 U13458 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n14156), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11749) );
  NAND4_X1 U13459 ( .A1(n11752), .A2(n11751), .A3(n11750), .A4(n11749), .ZN(
        n11753) );
  NAND2_X1 U13460 ( .A1(n11753), .A2(n11716), .ZN(n11754) );
  AND2_X1 U13461 ( .A1(n12494), .A2(n11771), .ZN(n12719) );
  NAND2_X1 U13462 ( .A1(n12477), .A2(n11762), .ZN(n12476) );
  NAND2_X1 U13463 ( .A1(n12494), .A2(n11757), .ZN(n12472) );
  NAND3_X1 U13464 ( .A1(n12476), .A2(n19758), .A3(n12472), .ZN(n12715) );
  NAND2_X1 U13465 ( .A1(n12715), .A2(n12717), .ZN(n11759) );
  NAND2_X1 U13466 ( .A1(n11759), .A2(n11758), .ZN(n11805) );
  NAND2_X1 U13467 ( .A1(n11805), .A2(n12451), .ZN(n11761) );
  NAND3_X1 U13468 ( .A1(n12260), .A2(n20155), .A3(n13896), .ZN(n11767) );
  NOR2_X1 U13469 ( .A1(n12031), .A2(n11772), .ZN(n11765) );
  INV_X1 U13471 ( .A(n11778), .ZN(n19169) );
  INV_X1 U13472 ( .A(n12031), .ZN(n11786) );
  NAND2_X2 U13473 ( .A1(n11774), .A2(n11779), .ZN(n12709) );
  NOR2_X1 U13474 ( .A1(n19261), .A2(n19926), .ZN(n11775) );
  NAND3_X1 U13475 ( .A1(n11779), .A2(n11785), .A3(n11778), .ZN(n11782) );
  NAND2_X1 U13476 ( .A1(n11782), .A2(n11781), .ZN(n11792) );
  INV_X1 U13477 ( .A(n19168), .ZN(n11783) );
  NAND3_X1 U13478 ( .A1(n11786), .A2(n19970), .A3(n11785), .ZN(n11787) );
  NAND2_X1 U13479 ( .A1(n11787), .A2(n11770), .ZN(n11791) );
  INV_X1 U13480 ( .A(n12474), .ZN(n11788) );
  NAND2_X1 U13481 ( .A1(n11823), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11799) );
  AOI21_X1 U13482 ( .B1(n11843), .B2(P2_REIP_REG_1__SCAN_IN), .A(n11246), .ZN(
        n11797) );
  NAND2_X1 U13483 ( .A1(n11824), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n11796) );
  AND2_X1 U13484 ( .A1(n11797), .A2(n11796), .ZN(n11798) );
  INV_X1 U13485 ( .A(n11823), .ZN(n11812) );
  INV_X1 U13486 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n18862) );
  INV_X2 U13487 ( .A(n12335), .ZN(n11843) );
  NAND2_X1 U13488 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11800) );
  NAND2_X1 U13489 ( .A1(n19261), .A2(n11800), .ZN(n11801) );
  AOI21_X1 U13490 ( .B1(n11843), .B2(P2_REIP_REG_0__SCAN_IN), .A(n11801), .ZN(
        n11803) );
  INV_X1 U13491 ( .A(n11804), .ZN(n11811) );
  NAND2_X1 U13492 ( .A1(n11805), .A2(n11806), .ZN(n11808) );
  NAND2_X1 U13493 ( .A1(n11808), .A2(n11807), .ZN(n11809) );
  NAND2_X1 U13494 ( .A1(n11809), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11810) );
  OAI211_X2 U13495 ( .C1(n11812), .C2(n19184), .A(n11811), .B(n11810), .ZN(
        n11828) );
  INV_X1 U13496 ( .A(n11813), .ZN(n11814) );
  NOR2_X1 U13497 ( .A1(n11814), .A2(n12726), .ZN(n11815) );
  OAI22_X1 U13498 ( .A1(n11840), .A2(n11815), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n11824), .ZN(n11819) );
  INV_X1 U13499 ( .A(n11816), .ZN(n12710) );
  NOR2_X1 U13500 ( .A1(n19261), .A2(n19927), .ZN(n11817) );
  AOI21_X1 U13501 ( .B1(n12710), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n11817), 
        .ZN(n11818) );
  NAND2_X1 U13502 ( .A1(n11819), .A2(n11818), .ZN(n11829) );
  NAND2_X2 U13503 ( .A1(n11828), .A2(n11829), .ZN(n11831) );
  NAND2_X1 U13504 ( .A1(n11156), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11822) );
  AOI21_X1 U13505 ( .B1(n19270), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n11821) );
  AOI22_X1 U13506 ( .A1(n11843), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11826) );
  NAND2_X1 U13507 ( .A1(n11824), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n11825) );
  OAI211_X1 U13508 ( .C1(n11812), .C2(n16001), .A(n11826), .B(n11825), .ZN(
        n11827) );
  INV_X1 U13509 ( .A(n11831), .ZN(n11834) );
  BUF_X1 U13510 ( .A(n11832), .Z(n11850) );
  INV_X1 U13511 ( .A(n11850), .ZN(n11833) );
  NAND2_X1 U13512 ( .A1(n11834), .A2(n11833), .ZN(n11835) );
  NAND2_X1 U13513 ( .A1(n11229), .A2(n17336), .ZN(n11860) );
  NAND2_X1 U13514 ( .A1(n11156), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11842) );
  OR2_X1 U13515 ( .A1(n19261), .A2(n19809), .ZN(n11841) );
  NAND2_X1 U13516 ( .A1(n11842), .A2(n11841), .ZN(n11847) );
  CLKBUF_X3 U13517 ( .A(n11843), .Z(n12703) );
  AOI22_X1 U13518 ( .A1(n12703), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11845) );
  NAND2_X1 U13519 ( .A1(n12700), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n11844) );
  OAI211_X1 U13520 ( .C1(n11812), .C2(n15820), .A(n11845), .B(n11844), .ZN(
        n11846) );
  NAND2_X1 U13521 ( .A1(n11847), .A2(n11846), .ZN(n11848) );
  NOR2_X1 U13522 ( .A1(n15437), .A2(n11849), .ZN(n11970) );
  AOI22_X1 U13523 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n11971), .B1(
        n11970), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11859) );
  NOR2_X2 U13524 ( .A1(n15441), .A2(n11849), .ZN(n11969) );
  NOR2_X1 U13525 ( .A1(n18858), .A2(n11850), .ZN(n11870) );
  AND2_X1 U13526 ( .A1(n16014), .A2(n11870), .ZN(n11861) );
  AOI22_X1 U13527 ( .A1(n11969), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n11972), .ZN(n11858) );
  INV_X1 U13528 ( .A(n11851), .ZN(n11852) );
  NOR2_X1 U13529 ( .A1(n11830), .A2(n11852), .ZN(n11873) );
  AND2_X1 U13530 ( .A1(n16014), .A2(n11873), .ZN(n11853) );
  AOI22_X1 U13531 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19904), .B1(
        n19800), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11857) );
  NAND2_X1 U13532 ( .A1(n19778), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11856) );
  NAND2_X2 U13533 ( .A1(n15437), .A2(n17838), .ZN(n11872) );
  INV_X1 U13534 ( .A(n17336), .ZN(n18879) );
  NAND2_X1 U13535 ( .A1(n18879), .A2(n18858), .ZN(n11876) );
  INV_X1 U13536 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11864) );
  NAND2_X1 U13537 ( .A1(n19837), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11863) );
  AOI21_X1 U13538 ( .B1(n19825), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A(
        n14673), .ZN(n11862) );
  OAI211_X1 U13539 ( .C1(n19857), .C2(n11864), .A(n11863), .B(n11862), .ZN(
        n11869) );
  INV_X1 U13540 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11867) );
  NAND2_X1 U13541 ( .A1(n17336), .A2(n18858), .ZN(n11874) );
  INV_X1 U13542 ( .A(n11873), .ZN(n11865) );
  INV_X1 U13543 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11866) );
  NOR2_X1 U13544 ( .A1(n11869), .A2(n11868), .ZN(n11881) );
  NOR2_X2 U13545 ( .A1(n11872), .A2(n11871), .ZN(n19873) );
  AOI22_X1 U13546 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19873), .B1(
        n19754), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11879) );
  INV_X1 U13547 ( .A(n11874), .ZN(n11875) );
  INV_X1 U13548 ( .A(n11876), .ZN(n11877) );
  AOI22_X1 U13549 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n11978), .B1(
        n11982), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11878) );
  AND2_X1 U13550 ( .A1(n11879), .A2(n11878), .ZN(n11880) );
  NAND3_X1 U13551 ( .A1(n11882), .A2(n11881), .A3(n11880), .ZN(n11927) );
  INV_X1 U13552 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n20356) );
  NAND2_X1 U13553 ( .A1(n11883), .A2(n11716), .ZN(n12007) );
  AOI22_X1 U13554 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17363), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11900) );
  AOI22_X1 U13555 ( .A1(n14126), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11942), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11899) );
  AOI22_X1 U13556 ( .A1(n14071), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14072), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11885) );
  INV_X1 U13557 ( .A(n11885), .ZN(n11889) );
  AND2_X2 U13558 ( .A1(n14277), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14069) );
  AOI22_X1 U13559 ( .A1(n14068), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14069), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11887) );
  NOR2_X1 U13560 ( .A1(n11889), .A2(n11888), .ZN(n11898) );
  AND2_X1 U13561 ( .A1(n14139), .A2(n11716), .ZN(n11901) );
  AOI22_X1 U13562 ( .A1(n11909), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11901), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11897) );
  AND2_X2 U13563 ( .A1(n14156), .A2(n11716), .ZN(n14104) );
  AOI22_X1 U13564 ( .A1(n14104), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11921), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11896) );
  AOI22_X1 U13565 ( .A1(n11962), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11906), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11895) );
  AND2_X1 U13566 ( .A1(n11893), .A2(n14137), .ZN(n11908) );
  AOI22_X1 U13567 ( .A1(n11907), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11908), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11894) );
  NAND4_X1 U13568 ( .A1(n11900), .A2(n11899), .A3(n11898), .A4(n11647), .ZN(
        n12365) );
  AOI22_X1 U13569 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n14104), .B1(
        n11942), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11905) );
  AOI22_X1 U13570 ( .A1(n11901), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12556), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11904) );
  AOI22_X1 U13571 ( .A1(n14072), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11921), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11903) );
  AOI22_X1 U13572 ( .A1(n14068), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17363), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11902) );
  NAND4_X1 U13573 ( .A1(n11905), .A2(n11904), .A3(n11903), .A4(n11902), .ZN(
        n11915) );
  AOI22_X1 U13574 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n11962), .B1(
        n11906), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11913) );
  AOI22_X1 U13575 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n11907), .B1(
        n11908), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11912) );
  AOI22_X1 U13576 ( .A1(n14126), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11911) );
  AOI22_X1 U13577 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n14069), .B1(
        n14071), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11910) );
  NAND4_X1 U13578 ( .A1(n11913), .A2(n11912), .A3(n11911), .A4(n11910), .ZN(
        n11914) );
  NOR2_X1 U13579 ( .A1(n11915), .A2(n11914), .ZN(n12505) );
  NOR2_X1 U13580 ( .A1(n14667), .A2(n12505), .ZN(n11916) );
  NAND2_X1 U13581 ( .A1(n14673), .A2(n11916), .ZN(n12369) );
  AOI22_X1 U13582 ( .A1(n14068), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14069), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11920) );
  AOI22_X1 U13583 ( .A1(n14071), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14072), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11919) );
  AOI22_X1 U13584 ( .A1(n14126), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11942), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11918) );
  AOI22_X1 U13585 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17363), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11917) );
  AOI22_X1 U13586 ( .A1(n11909), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11901), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11925) );
  AOI22_X1 U13587 ( .A1(n14104), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11921), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11924) );
  AOI22_X1 U13588 ( .A1(n11962), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11906), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11923) );
  AOI22_X1 U13589 ( .A1(n11907), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11908), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11922) );
  NAND2_X1 U13590 ( .A1(n12369), .A2(n12511), .ZN(n11926) );
  NAND2_X1 U13591 ( .A1(n11927), .A2(n11926), .ZN(n12050) );
  INV_X1 U13592 ( .A(n12050), .ZN(n11957) );
  AOI22_X1 U13593 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n11969), .B1(
        n11970), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11930) );
  AOI22_X1 U13594 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19904), .B1(
        n19800), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11929) );
  AOI22_X1 U13595 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n11972), .B1(
        n19825), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11928) );
  AND4_X1 U13596 ( .A1(n11931), .A2(n11930), .A3(n11929), .A4(n11928), .ZN(
        n11941) );
  AOI22_X1 U13597 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19873), .B1(
        n19754), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11933) );
  AOI22_X1 U13598 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n11978), .B1(
        n11982), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11932) );
  AND2_X1 U13599 ( .A1(n11933), .A2(n11932), .ZN(n11940) );
  INV_X1 U13600 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11935) );
  INV_X1 U13601 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11934) );
  INV_X1 U13602 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11936) );
  INV_X1 U13603 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14070) );
  NOR2_X1 U13604 ( .A1(n11938), .A2(n11937), .ZN(n11939) );
  NAND3_X1 U13605 ( .A1(n11941), .A2(n11940), .A3(n11939), .ZN(n11955) );
  AOI22_X1 U13606 ( .A1(n14126), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11942), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11953) );
  AOI22_X1 U13607 ( .A1(n14068), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14069), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11952) );
  AOI22_X1 U13608 ( .A1(n11909), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11901), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11946) );
  AOI22_X1 U13609 ( .A1(n14104), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11921), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11945) );
  AOI22_X1 U13610 ( .A1(n11962), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11906), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11944) );
  AOI22_X1 U13611 ( .A1(n11907), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11908), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11943) );
  NAND4_X1 U13612 ( .A1(n11946), .A2(n11945), .A3(n11944), .A4(n11943), .ZN(
        n11949) );
  AOI22_X1 U13613 ( .A1(n14071), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14072), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11947) );
  AOI22_X1 U13614 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17363), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11950) );
  NAND4_X1 U13615 ( .A1(n11953), .A2(n11952), .A3(n11951), .A4(n11950), .ZN(
        n12044) );
  INV_X1 U13616 ( .A(n12044), .ZN(n12522) );
  NAND2_X1 U13617 ( .A1(n12522), .A2(n14673), .ZN(n11954) );
  NAND2_X1 U13618 ( .A1(n11955), .A2(n11954), .ZN(n12051) );
  INV_X1 U13619 ( .A(n12051), .ZN(n11956) );
  AOI22_X1 U13620 ( .A1(n14068), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14069), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11961) );
  AOI22_X1 U13621 ( .A1(n14071), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14072), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11960) );
  AOI22_X1 U13622 ( .A1(n14126), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11942), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11959) );
  AOI22_X1 U13623 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17363), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11958) );
  NAND4_X1 U13624 ( .A1(n11961), .A2(n11960), .A3(n11959), .A4(n11958), .ZN(
        n11968) );
  AOI22_X1 U13625 ( .A1(n11909), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11901), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11966) );
  AOI22_X1 U13626 ( .A1(n14104), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11921), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11965) );
  AOI22_X1 U13627 ( .A1(n11962), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11906), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11964) );
  AOI22_X1 U13628 ( .A1(n11907), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11908), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11963) );
  NAND4_X1 U13629 ( .A1(n11966), .A2(n11965), .A3(n11964), .A4(n11963), .ZN(
        n11967) );
  AOI22_X1 U13630 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n11969), .B1(
        n19813), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11976) );
  AOI22_X1 U13631 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n11971), .B1(
        n19837), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11975) );
  AOI22_X1 U13632 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19904), .B1(
        n19825), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11974) );
  AOI22_X1 U13633 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n11972), .B1(
        n19800), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11973) );
  AOI22_X1 U13634 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19889), .B1(
        n11978), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11989) );
  AOI22_X1 U13635 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19842), .B1(
        n19851), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11988) );
  INV_X1 U13636 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14097) );
  INV_X1 U13637 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11981) );
  OAI22_X1 U13638 ( .A1(n14097), .A2(n11980), .B1(n12076), .B2(n11981), .ZN(
        n11986) );
  INV_X1 U13639 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11984) );
  INV_X1 U13640 ( .A(n19873), .ZN(n19870) );
  INV_X1 U13641 ( .A(n11982), .ZN(n12079) );
  INV_X1 U13642 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11983) );
  OAI22_X1 U13643 ( .A1(n11984), .A2(n19870), .B1(n12079), .B2(n11983), .ZN(
        n11985) );
  NOR2_X1 U13644 ( .A1(n11986), .A2(n11985), .ZN(n11987) );
  NAND4_X1 U13645 ( .A1(n11990), .A2(n11989), .A3(n11988), .A4(n11987), .ZN(
        n12002) );
  AOI22_X1 U13646 ( .A1(n14069), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14126), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11994) );
  AOI22_X1 U13647 ( .A1(n14071), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11942), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11993) );
  AOI22_X1 U13648 ( .A1(n14068), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14072), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11992) );
  AOI22_X1 U13649 ( .A1(n11921), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17363), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11991) );
  NAND4_X1 U13650 ( .A1(n11994), .A2(n11993), .A3(n11992), .A4(n11991), .ZN(
        n12000) );
  AOI22_X1 U13651 ( .A1(n11909), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11901), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11998) );
  AOI22_X1 U13652 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14104), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11997) );
  AOI22_X1 U13653 ( .A1(n11907), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11962), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11996) );
  AOI22_X1 U13654 ( .A1(n11908), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11906), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11995) );
  NAND4_X1 U13655 ( .A1(n11998), .A2(n11997), .A3(n11996), .A4(n11995), .ZN(
        n11999) );
  NOR2_X1 U13656 ( .A1(n12000), .A2(n11999), .ZN(n12047) );
  NAND2_X1 U13657 ( .A1(n12047), .A2(n14673), .ZN(n12001) );
  INV_X1 U13658 ( .A(n14126), .ZN(n12006) );
  INV_X1 U13659 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12005) );
  INV_X1 U13660 ( .A(n11942), .ZN(n12004) );
  INV_X1 U13661 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12003) );
  OAI22_X1 U13662 ( .A1(n12006), .A2(n12005), .B1(n12004), .B2(n12003), .ZN(
        n12009) );
  INV_X1 U13663 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n19960) );
  INV_X1 U13664 ( .A(n12556), .ZN(n14077) );
  INV_X1 U13665 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14273) );
  OAI22_X1 U13666 ( .A1(n19960), .A2(n14077), .B1(n12007), .B2(n14273), .ZN(
        n12008) );
  NOR2_X1 U13667 ( .A1(n12009), .A2(n12008), .ZN(n12021) );
  NAND2_X1 U13668 ( .A1(n14068), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12013) );
  NAND2_X1 U13669 ( .A1(n14069), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n12012) );
  NAND2_X1 U13670 ( .A1(n14072), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12011) );
  NAND2_X1 U13671 ( .A1(n14071), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n12010) );
  AOI22_X1 U13672 ( .A1(n11907), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11908), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12017) );
  AOI22_X1 U13673 ( .A1(n11962), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11906), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12016) );
  NAND2_X1 U13674 ( .A1(n11909), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n12015) );
  NAND2_X1 U13675 ( .A1(n11901), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12014) );
  AOI22_X1 U13676 ( .A1(n14104), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11921), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12018) );
  NAND4_X1 U13677 ( .A1(n12021), .A2(n12020), .A3(n12019), .A4(n12018), .ZN(
        n12022) );
  INV_X1 U13678 ( .A(n12023), .ZN(n12024) );
  INV_X1 U13679 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n12275) );
  NAND2_X1 U13680 ( .A1(n12449), .A2(n12250), .ZN(n12026) );
  NAND2_X1 U13681 ( .A1(n19926), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12025) );
  NAND2_X1 U13682 ( .A1(n12026), .A2(n12025), .ZN(n12034) );
  XNOR2_X1 U13683 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12035) );
  NAND2_X1 U13684 ( .A1(n12034), .A2(n12035), .ZN(n12038) );
  NAND2_X1 U13685 ( .A1(n19832), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12027) );
  NAND3_X1 U13686 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12249), .A3(
        n19172), .ZN(n12444) );
  MUX2_X1 U13687 ( .A(n12444), .B(n12030), .S(n12451), .Z(n12262) );
  MUX2_X1 U13688 ( .A(n12275), .B(n12262), .S(n12493), .Z(n12067) );
  OR2_X1 U13689 ( .A1(n12505), .A2(n20020), .ZN(n12033) );
  NOR2_X1 U13690 ( .A1(n12493), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n12057) );
  INV_X1 U13691 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n18871) );
  NAND2_X1 U13692 ( .A1(n12057), .A2(n18871), .ZN(n12032) );
  NAND2_X1 U13693 ( .A1(n12033), .A2(n12032), .ZN(n12063) );
  INV_X1 U13694 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n15746) );
  INV_X1 U13695 ( .A(n12034), .ZN(n12037) );
  INV_X1 U13696 ( .A(n12035), .ZN(n12036) );
  NAND2_X1 U13697 ( .A1(n12037), .A2(n12036), .ZN(n12039) );
  AND2_X1 U13698 ( .A1(n12039), .A2(n12038), .ZN(n12448) );
  AND2_X1 U13699 ( .A1(n13906), .A2(n12448), .ZN(n12263) );
  INV_X1 U13700 ( .A(n12263), .ZN(n12447) );
  MUX2_X1 U13701 ( .A(n15746), .B(n12041), .S(n12493), .Z(n12062) );
  NAND2_X1 U13702 ( .A1(n12063), .A2(n12062), .ZN(n12061) );
  XNOR2_X1 U13703 ( .A(n12043), .B(n12042), .ZN(n12443) );
  INV_X1 U13704 ( .A(n12261), .ZN(n12045) );
  INV_X1 U13705 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n12046) );
  NAND2_X1 U13706 ( .A1(n20020), .A2(n12046), .ZN(n12049) );
  INV_X1 U13707 ( .A(n12047), .ZN(n12048) );
  NAND2_X1 U13708 ( .A1(n12048), .A2(n12493), .ZN(n12531) );
  XNOR2_X1 U13709 ( .A(n12112), .B(n12113), .ZN(n18900) );
  XNOR2_X1 U13710 ( .A(n12051), .B(n12050), .ZN(n12372) );
  BUF_X1 U13711 ( .A(n12372), .Z(n15431) );
  OR2_X1 U13712 ( .A1(n15431), .A2(n12022), .ZN(n12053) );
  XNOR2_X1 U13713 ( .A(n12052), .B(n12061), .ZN(n15638) );
  INV_X1 U13714 ( .A(n12250), .ZN(n12056) );
  NAND2_X1 U13715 ( .A1(n12054), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12055) );
  NAND2_X1 U13716 ( .A1(n12056), .A2(n12055), .ZN(n12252) );
  INV_X1 U13717 ( .A(n12252), .ZN(n12454) );
  MUX2_X1 U13718 ( .A(n12365), .B(n12454), .S(n13906), .Z(n12264) );
  INV_X1 U13719 ( .A(n12264), .ZN(n12058) );
  AOI21_X1 U13720 ( .B1(n12058), .B2(n12493), .A(n12057), .ZN(n18859) );
  NAND2_X1 U13721 ( .A1(n18859), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14665) );
  INV_X1 U13722 ( .A(n12063), .ZN(n12060) );
  NAND3_X1 U13723 ( .A1(n20020), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n12059) );
  NAND2_X1 U13724 ( .A1(n12060), .A2(n12059), .ZN(n18872) );
  NAND2_X1 U13725 ( .A1(n14665), .A2(n18872), .ZN(n14744) );
  OR2_X1 U13726 ( .A1(n14665), .A2(n18872), .ZN(n14745) );
  NAND2_X1 U13727 ( .A1(n14746), .A2(n14745), .ZN(n14742) );
  AND2_X1 U13728 ( .A1(n14744), .A2(n14742), .ZN(n16000) );
  OAI21_X1 U13729 ( .B1(n12063), .B2(n12062), .A(n12061), .ZN(n15747) );
  XNOR2_X1 U13730 ( .A(n15747), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n15999) );
  NAND2_X1 U13731 ( .A1(n16000), .A2(n15999), .ZN(n15998) );
  INV_X1 U13732 ( .A(n15747), .ZN(n12064) );
  NAND2_X1 U13733 ( .A1(n12064), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12065) );
  AND2_X1 U13734 ( .A1(n15998), .A2(n12065), .ZN(n15428) );
  XNOR2_X1 U13735 ( .A(n12067), .B(n12066), .ZN(n17844) );
  INV_X1 U13736 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19204) );
  AND2_X1 U13737 ( .A1(n17844), .A2(n19204), .ZN(n12069) );
  AOI21_X1 U13738 ( .B1(n15428), .B2(n15820), .A(n12069), .ZN(n12068) );
  NAND2_X1 U13739 ( .A1(n17843), .A2(n12068), .ZN(n12074) );
  INV_X1 U13740 ( .A(n15428), .ZN(n12072) );
  INV_X1 U13741 ( .A(n12069), .ZN(n12070) );
  AND2_X1 U13742 ( .A1(n12070), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12071) );
  INV_X1 U13743 ( .A(n17844), .ZN(n18885) );
  AOI22_X1 U13744 ( .A1(n12072), .A2(n12071), .B1(n18885), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12073) );
  NAND2_X1 U13745 ( .A1(n12074), .A2(n12073), .ZN(n15812) );
  INV_X1 U13746 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12077) );
  INV_X1 U13747 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12075) );
  OAI22_X1 U13748 ( .A1(n12077), .A2(n11980), .B1(n12076), .B2(n12075), .ZN(
        n12082) );
  INV_X1 U13749 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12080) );
  INV_X1 U13750 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12078) );
  OAI22_X1 U13751 ( .A1(n12080), .A2(n19794), .B1(n12079), .B2(n12078), .ZN(
        n12081) );
  NOR2_X1 U13752 ( .A1(n12082), .A2(n12081), .ZN(n12099) );
  NAND2_X1 U13753 ( .A1(n11969), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n12086) );
  NAND2_X1 U13754 ( .A1(n19813), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12085) );
  NAND2_X1 U13755 ( .A1(n19837), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n12084) );
  NAND2_X1 U13756 ( .A1(n11971), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12083) );
  NAND4_X1 U13757 ( .A1(n12086), .A2(n12085), .A3(n12084), .A4(n12083), .ZN(
        n12096) );
  INV_X1 U13758 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12090) );
  INV_X1 U13759 ( .A(n19825), .ZN(n12089) );
  INV_X1 U13760 ( .A(n19800), .ZN(n12088) );
  INV_X1 U13761 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12087) );
  OAI22_X1 U13762 ( .A1(n12090), .A2(n12089), .B1(n12088), .B2(n12087), .ZN(
        n12095) );
  INV_X1 U13763 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12094) );
  INV_X1 U13764 ( .A(n11972), .ZN(n12093) );
  INV_X1 U13765 ( .A(n19904), .ZN(n12092) );
  INV_X1 U13766 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12091) );
  AOI22_X1 U13767 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19842), .B1(
        n19851), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12098) );
  AOI22_X1 U13768 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19889), .B1(
        n19873), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12097) );
  AOI22_X1 U13769 ( .A1(n14068), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n14069), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12103) );
  AOI22_X1 U13770 ( .A1(n14071), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14072), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12102) );
  AOI22_X1 U13771 ( .A1(n14126), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11942), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12101) );
  AOI22_X1 U13772 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17363), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12100) );
  NAND4_X1 U13773 ( .A1(n12103), .A2(n12102), .A3(n12101), .A4(n12100), .ZN(
        n12109) );
  AOI22_X1 U13774 ( .A1(n11909), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11901), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12107) );
  AOI22_X1 U13775 ( .A1(n14104), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11921), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12106) );
  AOI22_X1 U13776 ( .A1(n11962), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11906), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12105) );
  AOI22_X1 U13777 ( .A1(n11907), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11908), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12104) );
  NAND4_X1 U13778 ( .A1(n12107), .A2(n12106), .A3(n12105), .A4(n12104), .ZN(
        n12108) );
  NOR2_X1 U13779 ( .A1(n12109), .A2(n12108), .ZN(n12537) );
  NAND2_X1 U13780 ( .A1(n12537), .A2(n14673), .ZN(n12110) );
  XNOR2_X1 U13781 ( .A(n12379), .B(n12399), .ZN(n12386) );
  NAND2_X1 U13782 ( .A1(n12386), .A2(n12430), .ZN(n12114) );
  MUX2_X1 U13783 ( .A(P2_EBX_REG_6__SCAN_IN), .B(n12537), .S(n12493), .Z(
        n12117) );
  XNOR2_X1 U13784 ( .A(n12116), .B(n12117), .ZN(n18912) );
  INV_X1 U13785 ( .A(n12116), .ZN(n12119) );
  INV_X1 U13786 ( .A(n12117), .ZN(n12118) );
  NAND2_X1 U13787 ( .A1(n12119), .A2(n12118), .ZN(n12121) );
  INV_X1 U13788 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n12285) );
  MUX2_X1 U13789 ( .A(n12285), .B(n12022), .S(n12493), .Z(n12122) );
  XNOR2_X1 U13790 ( .A(n12121), .B(n12122), .ZN(n18925) );
  NAND2_X1 U13791 ( .A1(n18925), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17024) );
  OAI21_X1 U13792 ( .B1(n17022), .B2(n11297), .A(n17024), .ZN(n12120) );
  NAND2_X1 U13793 ( .A1(n17874), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12124) );
  INV_X1 U13794 ( .A(n12121), .ZN(n12123) );
  NAND2_X1 U13795 ( .A1(n20020), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12131) );
  XNOR2_X1 U13796 ( .A(n12130), .B(n12131), .ZN(n15735) );
  NAND2_X1 U13797 ( .A1(n12124), .A2(n17875), .ZN(n12129) );
  INV_X1 U13798 ( .A(n17874), .ZN(n12126) );
  INV_X1 U13799 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12125) );
  NAND2_X1 U13800 ( .A1(n12126), .A2(n12125), .ZN(n12128) );
  INV_X1 U13801 ( .A(n18925), .ZN(n12127) );
  INV_X1 U13802 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n19196) );
  NAND2_X1 U13803 ( .A1(n12127), .A2(n19196), .ZN(n17873) );
  INV_X1 U13804 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n12132) );
  NOR2_X1 U13805 ( .A1(n12493), .A2(n12132), .ZN(n12135) );
  NAND2_X1 U13806 ( .A1(n12134), .A2(n12133), .ZN(n12138) );
  NAND2_X1 U13807 ( .A1(n12136), .A2(n12135), .ZN(n12137) );
  NAND2_X1 U13808 ( .A1(n12138), .A2(n12137), .ZN(n18934) );
  INV_X1 U13809 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17279) );
  OAI21_X1 U13810 ( .B1(n18934), .B2(n12430), .A(n17279), .ZN(n17010) );
  INV_X1 U13811 ( .A(n12138), .ZN(n12139) );
  NAND2_X1 U13812 ( .A1(n20020), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n12182) );
  NAND2_X1 U13813 ( .A1(n12139), .A2(n12182), .ZN(n12178) );
  INV_X1 U13814 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n12140) );
  NOR2_X1 U13815 ( .A1(n12493), .A2(n12140), .ZN(n12177) );
  NAND2_X1 U13816 ( .A1(n20020), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n12169) );
  NAND2_X1 U13817 ( .A1(n20020), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n12167) );
  NAND2_X1 U13818 ( .A1(n12166), .A2(n12167), .ZN(n12174) );
  INV_X1 U13819 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n12144) );
  INV_X1 U13820 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n12146) );
  NOR2_X2 U13821 ( .A1(n12162), .A2(n12161), .ZN(n12157) );
  NAND2_X1 U13822 ( .A1(n20020), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n12158) );
  AND2_X2 U13823 ( .A1(n12157), .A2(n12158), .ZN(n12150) );
  NAND2_X1 U13824 ( .A1(n20020), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12151) );
  NAND2_X1 U13825 ( .A1(n20020), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n12148) );
  INV_X1 U13826 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n19039) );
  NOR2_X1 U13827 ( .A1(n12493), .A2(n19039), .ZN(n12195) );
  NAND2_X1 U13828 ( .A1(n20020), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12214) );
  NAND2_X1 U13829 ( .A1(n19052), .A2(n12438), .ZN(n12147) );
  INV_X1 U13830 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12825) );
  NAND2_X1 U13831 ( .A1(n12147), .A2(n12825), .ZN(n12809) );
  NAND2_X1 U13832 ( .A1(n19024), .A2(n12438), .ZN(n12149) );
  INV_X1 U13833 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17148) );
  NAND2_X1 U13834 ( .A1(n12149), .A2(n17148), .ZN(n16900) );
  INV_X1 U13835 ( .A(n12150), .ZN(n12153) );
  INV_X1 U13836 ( .A(n12151), .ZN(n12152) );
  NAND2_X1 U13837 ( .A1(n12153), .A2(n12152), .ZN(n12154) );
  NAND2_X1 U13838 ( .A1(n12155), .A2(n12154), .ZN(n19012) );
  INV_X1 U13839 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17159) );
  NAND2_X1 U13840 ( .A1(n16911), .A2(n17159), .ZN(n12156) );
  NAND2_X1 U13841 ( .A1(n16900), .A2(n12156), .ZN(n12806) );
  INV_X1 U13842 ( .A(n12157), .ZN(n12159) );
  XNOR2_X1 U13843 ( .A(n12159), .B(n12158), .ZN(n19004) );
  NAND2_X1 U13844 ( .A1(n19004), .A2(n12438), .ZN(n12160) );
  INV_X1 U13845 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12319) );
  NAND2_X1 U13846 ( .A1(n12160), .A2(n12319), .ZN(n16920) );
  XNOR2_X1 U13847 ( .A(n12162), .B(n12161), .ZN(n12163) );
  INV_X1 U13848 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17177) );
  OAI21_X1 U13849 ( .B1(n12163), .B2(n12430), .A(n17177), .ZN(n12165) );
  INV_X1 U13850 ( .A(n12163), .ZN(n18987) );
  AND2_X1 U13851 ( .A1(n12022), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12164) );
  NAND2_X1 U13852 ( .A1(n18987), .A2(n12164), .ZN(n12803) );
  INV_X1 U13853 ( .A(n12166), .ZN(n12168) );
  XNOR2_X1 U13854 ( .A(n12168), .B(n12167), .ZN(n15721) );
  AOI21_X1 U13855 ( .B1(n15721), .B2(n12438), .A(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16943) );
  XNOR2_X1 U13856 ( .A(n12172), .B(n12169), .ZN(n18965) );
  NAND2_X1 U13857 ( .A1(n18965), .A2(n12438), .ZN(n12205) );
  INV_X1 U13858 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17233) );
  NAND2_X1 U13859 ( .A1(n12205), .A2(n17233), .ZN(n16967) );
  NAND2_X1 U13860 ( .A1(n12170), .A2(n11244), .ZN(n12171) );
  NAND2_X1 U13861 ( .A1(n12172), .A2(n12171), .ZN(n15850) );
  OR2_X1 U13862 ( .A1(n15850), .A2(n12430), .ZN(n12173) );
  INV_X1 U13863 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17228) );
  NAND2_X1 U13864 ( .A1(n12173), .A2(n17228), .ZN(n16975) );
  NAND2_X1 U13865 ( .A1(n16967), .A2(n16975), .ZN(n16939) );
  NOR2_X1 U13866 ( .A1(n16943), .A2(n16939), .ZN(n12176) );
  XNOR2_X1 U13867 ( .A(n12174), .B(n11637), .ZN(n18975) );
  NAND2_X1 U13868 ( .A1(n18975), .A2(n12438), .ZN(n12175) );
  INV_X1 U13869 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12412) );
  NAND2_X1 U13870 ( .A1(n12175), .A2(n12412), .ZN(n16945) );
  AND2_X1 U13871 ( .A1(n12176), .A2(n16945), .ZN(n12800) );
  NAND2_X1 U13872 ( .A1(n12178), .A2(n12177), .ZN(n12179) );
  AND2_X1 U13873 ( .A1(n12170), .A2(n12179), .ZN(n12186) );
  AND2_X1 U13874 ( .A1(n12022), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12180) );
  NAND2_X1 U13875 ( .A1(n12186), .A2(n12180), .ZN(n16989) );
  INV_X1 U13876 ( .A(n18934), .ZN(n12181) );
  NAND3_X1 U13877 ( .A1(n12181), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n12022), .ZN(n17011) );
  XNOR2_X1 U13878 ( .A(n12138), .B(n12182), .ZN(n15773) );
  NAND2_X1 U13879 ( .A1(n15773), .A2(n12438), .ZN(n12187) );
  INV_X1 U13880 ( .A(n12187), .ZN(n12183) );
  NAND2_X1 U13881 ( .A1(n12183), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17000) );
  NAND2_X1 U13882 ( .A1(n17011), .A2(n17000), .ZN(n16991) );
  INV_X1 U13883 ( .A(n16991), .ZN(n12184) );
  NAND2_X1 U13884 ( .A1(n12022), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12185) );
  INV_X1 U13885 ( .A(n12186), .ZN(n18953) );
  INV_X1 U13886 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17254) );
  OAI21_X1 U13887 ( .B1(n18953), .B2(n12430), .A(n17254), .ZN(n16990) );
  INV_X1 U13888 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17270) );
  NAND2_X1 U13889 ( .A1(n12187), .A2(n17270), .ZN(n16999) );
  NAND2_X1 U13890 ( .A1(n16990), .A2(n16999), .ZN(n12188) );
  NAND2_X1 U13891 ( .A1(n12799), .A2(n12188), .ZN(n12189) );
  NAND4_X1 U13892 ( .A1(n16920), .A2(n16930), .A3(n12800), .A4(n12189), .ZN(
        n12190) );
  NOR2_X1 U13893 ( .A1(n12806), .A2(n12190), .ZN(n12191) );
  AND2_X1 U13894 ( .A1(n17010), .A2(n12193), .ZN(n12194) );
  INV_X1 U13895 ( .A(n12799), .ZN(n12192) );
  NAND2_X1 U13896 ( .A1(n12200), .A2(n17138), .ZN(n12199) );
  NAND2_X1 U13897 ( .A1(n12196), .A2(n12195), .ZN(n12197) );
  AND2_X1 U13898 ( .A1(n12213), .A2(n12197), .ZN(n19037) );
  NAND2_X1 U13899 ( .A1(n19037), .A2(n12438), .ZN(n12807) );
  INV_X1 U13900 ( .A(n12807), .ZN(n12198) );
  NAND2_X1 U13901 ( .A1(n12199), .A2(n12198), .ZN(n12212) );
  INV_X1 U13902 ( .A(n12200), .ZN(n12210) );
  INV_X1 U13903 ( .A(n19024), .ZN(n12201) );
  OR3_X1 U13904 ( .A1(n12201), .A2(n12430), .A3(n17148), .ZN(n16899) );
  OAI21_X1 U13905 ( .B1(n16911), .B2(n17159), .A(n16899), .ZN(n12805) );
  INV_X1 U13906 ( .A(n19004), .ZN(n12202) );
  AND2_X1 U13907 ( .A1(n12022), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12203) );
  NAND2_X1 U13908 ( .A1(n18975), .A2(n12203), .ZN(n16944) );
  AND2_X1 U13909 ( .A1(n12022), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12204) );
  NAND2_X1 U13910 ( .A1(n15721), .A2(n12204), .ZN(n16941) );
  OR2_X1 U13911 ( .A1(n12205), .A2(n17233), .ZN(n16968) );
  AND2_X1 U13912 ( .A1(n16941), .A2(n16968), .ZN(n12206) );
  AND2_X1 U13913 ( .A1(n16944), .A2(n12206), .ZN(n12801) );
  NAND3_X1 U13914 ( .A1(n16919), .A2(n12801), .A3(n12803), .ZN(n12207) );
  NOR2_X1 U13915 ( .A1(n12805), .A2(n12207), .ZN(n12209) );
  AND2_X1 U13916 ( .A1(n12022), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12208) );
  NAND2_X1 U13917 ( .A1(n19052), .A2(n12208), .ZN(n12808) );
  AOI21_X1 U13918 ( .B1(n12210), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n11230), .ZN(n12211) );
  INV_X1 U13919 ( .A(n12213), .ZN(n12215) );
  NAND2_X1 U13920 ( .A1(n12215), .A2(n12214), .ZN(n12216) );
  NAND2_X1 U13921 ( .A1(n20020), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12217) );
  XNOR2_X1 U13922 ( .A(n12216), .B(n12217), .ZN(n19063) );
  NAND2_X1 U13923 ( .A1(n19063), .A2(n12438), .ZN(n16886) );
  INV_X1 U13924 ( .A(n12216), .ZN(n12218) );
  NAND2_X1 U13925 ( .A1(n12218), .A2(n12217), .ZN(n12220) );
  INV_X1 U13926 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n12338) );
  NOR2_X1 U13927 ( .A1(n12493), .A2(n12338), .ZN(n12219) );
  NAND2_X1 U13928 ( .A1(n12220), .A2(n12219), .ZN(n12221) );
  AOI21_X1 U13929 ( .B1(n19078), .B2(n12438), .A(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16876) );
  AND2_X1 U13930 ( .A1(n12022), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12222) );
  NAND2_X1 U13931 ( .A1(n19078), .A2(n12222), .ZN(n16877) );
  NAND2_X1 U13932 ( .A1(n20020), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12223) );
  XNOR2_X1 U13933 ( .A(n11211), .B(n12223), .ZN(n19085) );
  NAND2_X1 U13934 ( .A1(n19085), .A2(n12438), .ZN(n16869) );
  INV_X1 U13935 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n12224) );
  NOR2_X1 U13936 ( .A1(n12493), .A2(n12224), .ZN(n12228) );
  NAND2_X1 U13937 ( .A1(n20020), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n12233) );
  XNOR2_X1 U13938 ( .A(n12234), .B(n12233), .ZN(n19108) );
  NAND2_X1 U13939 ( .A1(n19108), .A2(n12438), .ZN(n12225) );
  INV_X1 U13940 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17066) );
  NAND2_X1 U13941 ( .A1(n12225), .A2(n17066), .ZN(n12227) );
  AND2_X1 U13942 ( .A1(n12022), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12226) );
  NAND2_X1 U13943 ( .A1(n19108), .A2(n12226), .ZN(n12424) );
  NAND2_X1 U13944 ( .A1(n12227), .A2(n12424), .ZN(n12764) );
  INV_X1 U13945 ( .A(n12228), .ZN(n12229) );
  XNOR2_X1 U13946 ( .A(n12230), .B(n12229), .ZN(n19096) );
  NAND2_X1 U13947 ( .A1(n19096), .A2(n12438), .ZN(n12232) );
  INV_X1 U13948 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17079) );
  AND2_X1 U13949 ( .A1(n12232), .A2(n17079), .ZN(n16858) );
  NOR2_X1 U13950 ( .A1(n12764), .A2(n16858), .ZN(n12231) );
  NAND3_X1 U13951 ( .A1(n12422), .A2(n17066), .A3(n16857), .ZN(n12240) );
  NAND2_X1 U13952 ( .A1(n20020), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12236) );
  NAND2_X1 U13953 ( .A1(n12235), .A2(n12236), .ZN(n12245) );
  INV_X1 U13954 ( .A(n12235), .ZN(n12238) );
  INV_X1 U13955 ( .A(n12236), .ZN(n12237) );
  NAND2_X1 U13956 ( .A1(n12238), .A2(n12237), .ZN(n12239) );
  NAND2_X1 U13957 ( .A1(n12245), .A2(n12239), .ZN(n19122) );
  OR2_X1 U13958 ( .A1(n19122), .A2(n12430), .ZN(n12418) );
  NAND2_X1 U13959 ( .A1(n12240), .A2(n12419), .ZN(n16846) );
  INV_X1 U13960 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17058) );
  NAND2_X1 U13961 ( .A1(n12422), .A2(n12418), .ZN(n16847) );
  INV_X1 U13962 ( .A(n12245), .ZN(n12243) );
  INV_X1 U13963 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n12241) );
  NOR2_X1 U13964 ( .A1(n12493), .A2(n12241), .ZN(n12244) );
  INV_X1 U13965 ( .A(n12244), .ZN(n12242) );
  NAND2_X1 U13966 ( .A1(n12245), .A2(n12244), .ZN(n12246) );
  AND2_X1 U13967 ( .A1(n12425), .A2(n12246), .ZN(n16658) );
  XNOR2_X1 U13968 ( .A(n12423), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12247) );
  NAND3_X1 U13969 ( .A1(n12444), .A2(n12448), .A3(n12443), .ZN(n12253) );
  XNOR2_X1 U13970 ( .A(n12449), .B(n12250), .ZN(n12452) );
  NOR2_X1 U13971 ( .A1(n12253), .A2(n12452), .ZN(n12251) );
  OR2_X1 U13972 ( .A1(n12465), .A2(n12251), .ZN(n19248) );
  OAI21_X1 U13973 ( .B1(n12253), .B2(n12252), .A(n19256), .ZN(n12254) );
  OR2_X1 U13974 ( .A1(n19248), .A2(n12254), .ZN(n12259) );
  NAND2_X1 U13975 ( .A1(n12255), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12256) );
  NAND2_X1 U13976 ( .A1(n12256), .A2(n19172), .ZN(n19167) );
  INV_X1 U13977 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n12257) );
  OAI21_X1 U13978 ( .B1(n14068), .B2(n19167), .A(n12257), .ZN(n12258) );
  NAND2_X1 U13979 ( .A1(n12258), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n17885) );
  NAND2_X1 U13980 ( .A1(n12259), .A2(n17885), .ZN(n19272) );
  AND2_X1 U13981 ( .A1(n12469), .A2(n12451), .ZN(n19233) );
  NAND2_X1 U13982 ( .A1(n19272), .A2(n19233), .ZN(n12268) );
  NAND2_X1 U13983 ( .A1(n12262), .A2(n12261), .ZN(n12462) );
  AOI21_X1 U13984 ( .B1(n12264), .B2(n12449), .A(n12263), .ZN(n12265) );
  NOR2_X1 U13985 ( .A1(n12462), .A2(n12265), .ZN(n12266) );
  OR2_X1 U13986 ( .A1(n12266), .A2(n12465), .ZN(n19234) );
  INV_X1 U13987 ( .A(n19234), .ZN(n12267) );
  AND2_X1 U13988 ( .A1(n14673), .A2(n20247), .ZN(n12478) );
  NAND2_X1 U13989 ( .A1(n12267), .A2(n19235), .ZN(n12486) );
  NAND2_X1 U13990 ( .A1(n12268), .A2(n12486), .ZN(n19243) );
  INV_X2 U13991 ( .A(n12706), .ZN(n12698) );
  NAND2_X1 U13992 ( .A1(n12698), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12274) );
  AOI22_X1 U13993 ( .A1(n12703), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12273) );
  OAI211_X1 U13994 ( .C1(n12275), .C2(n12272), .A(n12274), .B(n12273), .ZN(
        n14978) );
  AOI22_X1 U13995 ( .A1(n12703), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12277) );
  NAND2_X1 U13996 ( .A1(n12700), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n12276) );
  NAND2_X1 U13997 ( .A1(n12277), .A2(n12276), .ZN(n12278) );
  AOI21_X1 U13998 ( .B1(n12698), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n12278), .ZN(n14989) );
  NAND2_X1 U13999 ( .A1(n12698), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12282) );
  AOI22_X1 U14000 ( .A1(n12703), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12280) );
  NAND2_X1 U14001 ( .A1(n12700), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n12279) );
  AND2_X1 U14002 ( .A1(n12280), .A2(n12279), .ZN(n12281) );
  NAND2_X1 U14003 ( .A1(n12282), .A2(n12281), .ZN(n15022) );
  INV_X1 U14004 ( .A(n15008), .ZN(n12288) );
  NAND2_X1 U14005 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12284) );
  NAND2_X1 U14006 ( .A1(n12703), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n12283) );
  OAI211_X1 U14007 ( .C1(n12272), .C2(n12285), .A(n12284), .B(n12283), .ZN(
        n12286) );
  AOI21_X1 U14008 ( .B1(n12698), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n12286), .ZN(n15009) );
  NAND2_X1 U14009 ( .A1(n12288), .A2(n12287), .ZN(n15007) );
  INV_X1 U14010 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n15739) );
  NAND2_X1 U14011 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12290) );
  NAND2_X1 U14012 ( .A1(n12703), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n12289) );
  OAI211_X1 U14013 ( .C1(n12272), .C2(n15739), .A(n12290), .B(n12289), .ZN(
        n12291) );
  AOI21_X1 U14014 ( .B1(n12698), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n12291), .ZN(n15074) );
  AOI22_X1 U14015 ( .A1(n12703), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12293) );
  NAND2_X1 U14016 ( .A1(n12700), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12292) );
  OAI211_X1 U14017 ( .C1(n12706), .C2(n17279), .A(n12293), .B(n12292), .ZN(
        n15043) );
  NAND2_X1 U14018 ( .A1(n15042), .A2(n15043), .ZN(n15041) );
  INV_X1 U14019 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n15772) );
  NAND2_X1 U14020 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12295) );
  NAND2_X1 U14021 ( .A1(n12703), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n12294) );
  OAI211_X1 U14022 ( .C1(n12272), .C2(n15772), .A(n12295), .B(n12294), .ZN(
        n12296) );
  AOI21_X1 U14023 ( .B1(n12698), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n12296), .ZN(n15055) );
  NAND2_X1 U14024 ( .A1(n12298), .A2(n12297), .ZN(n15053) );
  AOI22_X1 U14025 ( .A1(n12703), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n12300) );
  NAND2_X1 U14026 ( .A1(n12700), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n12299) );
  NAND2_X1 U14027 ( .A1(n12300), .A2(n12299), .ZN(n12301) );
  AOI21_X1 U14028 ( .B1(n12698), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n12301), .ZN(n15402) );
  INV_X1 U14029 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n12304) );
  NAND2_X1 U14030 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12303) );
  INV_X1 U14031 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n17965) );
  OR2_X1 U14032 ( .A1(n12335), .A2(n17965), .ZN(n12302) );
  OAI211_X1 U14033 ( .C1(n12272), .C2(n12304), .A(n12303), .B(n12302), .ZN(
        n12305) );
  AOI21_X1 U14034 ( .B1(n12698), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n12305), .ZN(n15356) );
  AOI22_X1 U14035 ( .A1(n12703), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n12307) );
  NAND2_X1 U14036 ( .A1(n12700), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n12306) );
  OAI211_X1 U14037 ( .C1(n12706), .C2(n17233), .A(n12307), .B(n12306), .ZN(
        n15625) );
  INV_X1 U14038 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n15726) );
  NAND2_X1 U14039 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12309) );
  INV_X1 U14040 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n17966) );
  OR2_X1 U14041 ( .A1(n12335), .A2(n17966), .ZN(n12308) );
  OAI211_X1 U14042 ( .C1(n12272), .C2(n15726), .A(n12309), .B(n12308), .ZN(
        n12310) );
  AOI21_X1 U14043 ( .B1(n12698), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n12310), .ZN(n15561) );
  AOI22_X1 U14044 ( .A1(n12703), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n12312) );
  NAND2_X1 U14045 ( .A1(n12700), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n12311) );
  NAND2_X1 U14046 ( .A1(n12312), .A2(n12311), .ZN(n12313) );
  AOI21_X1 U14047 ( .B1(n12698), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n12313), .ZN(n15707) );
  AOI22_X1 U14048 ( .A1(n12703), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n12316) );
  NAND2_X1 U14049 ( .A1(n12700), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12315) );
  OAI211_X1 U14050 ( .C1(n12706), .C2(n17177), .A(n12316), .B(n12315), .ZN(
        n15714) );
  AOI22_X1 U14051 ( .A1(n12703), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n12318) );
  NAND2_X1 U14052 ( .A1(n12700), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n12317) );
  OAI211_X1 U14053 ( .C1(n12706), .C2(n12319), .A(n12318), .B(n12317), .ZN(
        n15832) );
  AOI22_X1 U14054 ( .A1(n12703), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n12321) );
  NAND2_X1 U14055 ( .A1(n12700), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12320) );
  NAND2_X1 U14056 ( .A1(n12321), .A2(n12320), .ZN(n12322) );
  AOI21_X1 U14057 ( .B1(n12698), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n12322), .ZN(n15897) );
  AOI22_X1 U14058 ( .A1(n12703), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n12324) );
  NAND2_X1 U14059 ( .A1(n12700), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n12323) );
  NAND2_X1 U14060 ( .A1(n12324), .A2(n12323), .ZN(n12325) );
  AOI21_X1 U14061 ( .B1(n12698), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n12325), .ZN(n15907) );
  AOI22_X1 U14062 ( .A1(n12703), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n12327) );
  NAND2_X1 U14063 ( .A1(n12700), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12326) );
  OAI211_X1 U14064 ( .C1(n12706), .C2(n17138), .A(n12327), .B(n12326), .ZN(
        n16736) );
  AOI22_X1 U14065 ( .A1(n12703), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n12329) );
  NAND2_X1 U14066 ( .A1(n12700), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12328) );
  NAND2_X1 U14067 ( .A1(n12329), .A2(n12328), .ZN(n12330) );
  AOI21_X1 U14068 ( .B1(n12698), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n12330), .ZN(n12814) );
  AOI22_X1 U14069 ( .A1(n11843), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n12333) );
  NAND2_X1 U14070 ( .A1(n12700), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12332) );
  NAND2_X1 U14071 ( .A1(n12333), .A2(n12332), .ZN(n12334) );
  AOI21_X1 U14072 ( .B1(n12698), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n12334), .ZN(n16724) );
  NAND2_X1 U14073 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12337) );
  INV_X1 U14074 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n17973) );
  OR2_X1 U14075 ( .A1(n12335), .A2(n17973), .ZN(n12336) );
  OAI211_X1 U14076 ( .C1(n12272), .C2(n12338), .A(n12337), .B(n12336), .ZN(
        n12339) );
  AOI21_X1 U14077 ( .B1(n12698), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n12339), .ZN(n16720) );
  AOI22_X1 U14078 ( .A1(n12703), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n12341) );
  NAND2_X1 U14079 ( .A1(n12700), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12340) );
  OAI211_X1 U14080 ( .C1(n12706), .C2(n11610), .A(n12341), .B(n12340), .ZN(
        n16713) );
  AOI22_X1 U14081 ( .A1(n12703), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n12343) );
  NAND2_X1 U14082 ( .A1(n12700), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n12342) );
  NAND2_X1 U14083 ( .A1(n12343), .A2(n12342), .ZN(n12344) );
  AOI21_X1 U14084 ( .B1(n12698), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n12344), .ZN(n16706) );
  AOI22_X1 U14085 ( .A1(n12703), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n12346) );
  NAND2_X1 U14086 ( .A1(n12700), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n12345) );
  NAND2_X1 U14087 ( .A1(n12346), .A2(n12345), .ZN(n12347) );
  AOI21_X1 U14088 ( .B1(n12698), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n12347), .ZN(n12771) );
  AOI22_X1 U14089 ( .A1(n11843), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n12349) );
  NAND2_X1 U14090 ( .A1(n12700), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12348) );
  OAI211_X1 U14091 ( .C1(n12706), .C2(n17058), .A(n12349), .B(n12348), .ZN(
        n16694) );
  INV_X1 U14092 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12420) );
  AOI22_X1 U14093 ( .A1(n12703), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n12351) );
  NAND2_X1 U14094 ( .A1(n12700), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n12350) );
  OAI211_X1 U14095 ( .C1(n12706), .C2(n12420), .A(n12351), .B(n12350), .ZN(
        n12353) );
  OR2_X1 U14096 ( .A1(n12352), .A2(n12353), .ZN(n12354) );
  NAND2_X1 U14097 ( .A1(n12699), .A2(n12354), .ZN(n17052) );
  INV_X1 U14098 ( .A(n17768), .ZN(n12355) );
  NOR2_X1 U14099 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n12355), .ZN(n17884) );
  NAND2_X1 U14100 ( .A1(n17884), .A2(n19270), .ZN(n12356) );
  AND2_X1 U14101 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n17766) );
  NOR2_X1 U14102 ( .A1(n17052), .A2(n17865), .ZN(n12363) );
  NAND2_X1 U14103 ( .A1(n22292), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12357) );
  NAND2_X1 U14104 ( .A1(n19259), .A2(n12357), .ZN(n14670) );
  NAND2_X1 U14105 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13854) );
  INV_X1 U14106 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16861) );
  INV_X1 U14107 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12773) );
  NOR2_X1 U14108 ( .A1(n13882), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12360) );
  OR2_X1 U14109 ( .A1(n13843), .A2(n12360), .ZN(n16660) );
  NAND2_X1 U14110 ( .A1(n19256), .A2(n19916), .ZN(n19263) );
  INV_X1 U14111 ( .A(n19263), .ZN(n19170) );
  NAND2_X1 U14112 ( .A1(n19170), .A2(n19833), .ZN(n14661) );
  NAND2_X1 U14113 ( .A1(n19213), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n17049) );
  NAND2_X1 U14114 ( .A1(n17866), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12361) );
  OAI211_X1 U14115 ( .C1(n17883), .C2(n16660), .A(n17049), .B(n12361), .ZN(
        n12362) );
  INV_X1 U14116 ( .A(n12505), .ZN(n12366) );
  NAND2_X1 U14117 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n14667), .ZN(
        n14666) );
  NOR2_X1 U14118 ( .A1(n12505), .A2(n14666), .ZN(n12368) );
  NOR2_X1 U14119 ( .A1(n12365), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12367) );
  XOR2_X1 U14120 ( .A(n12367), .B(n12366), .Z(n14739) );
  NOR2_X1 U14121 ( .A1(n14746), .A2(n14739), .ZN(n14738) );
  NOR2_X1 U14122 ( .A1(n12368), .A2(n14738), .ZN(n12370) );
  XNOR2_X1 U14123 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n12370), .ZN(
        n16010) );
  XNOR2_X1 U14124 ( .A(n12369), .B(n12511), .ZN(n16009) );
  NAND2_X1 U14125 ( .A1(n16010), .A2(n16009), .ZN(n16008) );
  OR2_X1 U14126 ( .A1(n12370), .A2(n16001), .ZN(n12371) );
  NAND2_X1 U14127 ( .A1(n16008), .A2(n12371), .ZN(n12373) );
  XNOR2_X1 U14128 ( .A(n12373), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n15432) );
  NAND2_X1 U14129 ( .A1(n12373), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12374) );
  NAND2_X1 U14130 ( .A1(n12376), .A2(n12375), .ZN(n12377) );
  NAND2_X1 U14131 ( .A1(n12379), .A2(n12380), .ZN(n12391) );
  NAND2_X1 U14132 ( .A1(n12382), .A2(n12381), .ZN(n12395) );
  NAND2_X1 U14133 ( .A1(n12387), .A2(n12391), .ZN(n12383) );
  NAND2_X1 U14134 ( .A1(n12395), .A2(n12383), .ZN(n15816) );
  INV_X1 U14135 ( .A(n15816), .ZN(n12385) );
  INV_X1 U14136 ( .A(n12396), .ZN(n12388) );
  OAI21_X1 U14137 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n12381), .A(
        n12388), .ZN(n12389) );
  INV_X1 U14138 ( .A(n12399), .ZN(n12392) );
  MUX2_X1 U14139 ( .A(n12392), .B(n12384), .S(n12391), .Z(n12393) );
  OAI21_X1 U14140 ( .B1(n12396), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n12393), .ZN(n12394) );
  NAND2_X1 U14141 ( .A1(n15814), .A2(n12395), .ZN(n12397) );
  NAND2_X1 U14142 ( .A1(n12397), .A2(n12396), .ZN(n12398) );
  INV_X1 U14143 ( .A(n12379), .ZN(n12400) );
  NAND2_X1 U14144 ( .A1(n12401), .A2(n12430), .ZN(n12402) );
  NAND2_X1 U14145 ( .A1(n12409), .A2(n12402), .ZN(n12403) );
  XNOR2_X1 U14146 ( .A(n12403), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17028) );
  XNOR2_X1 U14147 ( .A(n12409), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17870) );
  AND2_X1 U14148 ( .A1(n17028), .A2(n17870), .ZN(n12408) );
  INV_X1 U14149 ( .A(n17870), .ZN(n12405) );
  INV_X1 U14150 ( .A(n12403), .ZN(n12404) );
  NAND2_X1 U14151 ( .A1(n12404), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17867) );
  INV_X1 U14152 ( .A(n12409), .ZN(n12410) );
  NAND3_X1 U14153 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12411) );
  NAND2_X1 U14154 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16937) );
  NOR2_X1 U14155 ( .A1(n12411), .A2(n16937), .ZN(n17216) );
  NAND2_X1 U14156 ( .A1(n17216), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17200) );
  OR2_X1 U14157 ( .A1(n17200), .A2(n12412), .ZN(n17173) );
  NAND3_X1 U14158 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12413) );
  NOR2_X1 U14159 ( .A1(n17173), .A2(n12413), .ZN(n17139) );
  AND2_X1 U14160 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17139), .ZN(
        n12414) );
  INV_X1 U14161 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17110) );
  INV_X1 U14162 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17100) );
  NAND2_X1 U14164 ( .A1(n12417), .A2(n12416), .ZN(P2_U2986) );
  NAND2_X1 U14165 ( .A1(n20020), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12426) );
  XOR2_X1 U14166 ( .A(n12426), .B(n12427), .Z(n19137) );
  NAND2_X1 U14167 ( .A1(n19137), .A2(n12438), .ZN(n12431) );
  INV_X1 U14168 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17039) );
  NAND2_X1 U14169 ( .A1(n12431), .A2(n17039), .ZN(n16842) );
  NAND2_X1 U14170 ( .A1(n12427), .A2(n12426), .ZN(n12436) );
  NAND2_X1 U14171 ( .A1(n20020), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12428) );
  AOI21_X1 U14172 ( .B1(n12429), .B2(n12438), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12780) );
  INV_X1 U14173 ( .A(n12429), .ZN(n13902) );
  INV_X1 U14174 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12791) );
  INV_X1 U14175 ( .A(n12431), .ZN(n12432) );
  NAND2_X1 U14176 ( .A1(n12432), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16841) );
  INV_X1 U14177 ( .A(n16841), .ZN(n12433) );
  NOR2_X1 U14178 ( .A1(n12436), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12437) );
  MUX2_X1 U14179 ( .A(n12437), .B(n12121), .S(n12493), .Z(n19148) );
  NAND2_X1 U14180 ( .A1(n19148), .A2(n12438), .ZN(n12439) );
  XNOR2_X1 U14181 ( .A(n12439), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12440) );
  NAND2_X1 U14182 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19281) );
  INV_X1 U14183 ( .A(n19281), .ZN(n22321) );
  INV_X1 U14184 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n17954) );
  NAND2_X2 U14185 ( .A1(n17987), .A2(n22328), .ZN(n17984) );
  NOR2_X1 U14186 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_0__SCAN_IN), 
        .ZN(n22322) );
  NAND2_X1 U14187 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n22322), .ZN(n17953) );
  NAND2_X1 U14188 ( .A1(n12442), .A2(n19247), .ZN(n12491) );
  AND2_X1 U14189 ( .A1(n12444), .A2(n12443), .ZN(n12461) );
  INV_X1 U14190 ( .A(n12448), .ZN(n12445) );
  OAI21_X1 U14191 ( .B1(n11768), .B2(n14673), .A(n12445), .ZN(n12446) );
  NAND2_X1 U14192 ( .A1(n12447), .A2(n12446), .ZN(n12459) );
  NAND2_X1 U14193 ( .A1(n19168), .A2(n12448), .ZN(n12457) );
  NAND2_X1 U14194 ( .A1(n12454), .A2(n12449), .ZN(n12450) );
  NAND2_X1 U14195 ( .A1(n12451), .A2(n12450), .ZN(n12456) );
  INV_X1 U14196 ( .A(n12452), .ZN(n12453) );
  OAI211_X1 U14197 ( .C1(n13896), .C2(n12454), .A(n11785), .B(n12453), .ZN(
        n12455) );
  NAND3_X1 U14198 ( .A1(n12457), .A2(n12456), .A3(n12455), .ZN(n12458) );
  NAND2_X1 U14199 ( .A1(n12459), .A2(n12458), .ZN(n12460) );
  AOI22_X1 U14200 ( .A1(n12462), .A2(n13906), .B1(n12461), .B2(n12460), .ZN(
        n12463) );
  OR2_X1 U14201 ( .A1(n12463), .A2(n12465), .ZN(n12464) );
  MUX2_X1 U14202 ( .A(n12464), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n19270), .Z(n12467) );
  NAND2_X1 U14203 ( .A1(n12465), .A2(n11768), .ZN(n12466) );
  NAND2_X1 U14204 ( .A1(n19242), .A2(n13896), .ZN(n12490) );
  AOI21_X1 U14205 ( .B1(n12467), .B2(n11785), .A(n11762), .ZN(n12468) );
  NAND2_X1 U14206 ( .A1(n12490), .A2(n12468), .ZN(n12489) );
  NAND3_X1 U14207 ( .A1(n19272), .A2(n12469), .A3(n13896), .ZN(n12487) );
  NAND2_X1 U14208 ( .A1(n12482), .A2(n19247), .ZN(n12470) );
  OR2_X1 U14209 ( .A1(n19248), .A2(n12470), .ZN(n12481) );
  NAND2_X1 U14210 ( .A1(n12472), .A2(n20155), .ZN(n12473) );
  NAND2_X1 U14211 ( .A1(n12471), .A2(n12473), .ZN(n12480) );
  INV_X1 U14212 ( .A(n19758), .ZN(n14816) );
  OR2_X1 U14213 ( .A1(n12474), .A2(n13896), .ZN(n12712) );
  OAI211_X1 U14214 ( .C1(n11785), .C2(n14816), .A(n12712), .B(n20155), .ZN(
        n12475) );
  AND3_X1 U14215 ( .A1(n12476), .A2(n12475), .A3(n12726), .ZN(n12479) );
  OAI21_X1 U14216 ( .B1(n12477), .B2(n14816), .A(n12478), .ZN(n12716) );
  AND2_X1 U14217 ( .A1(n12481), .A2(n12714), .ZN(n15762) );
  MUX2_X1 U14218 ( .A(n12482), .B(n12442), .S(n14673), .Z(n12483) );
  NAND2_X1 U14219 ( .A1(n12483), .A2(n19281), .ZN(n12484) );
  OR2_X1 U14220 ( .A1(n19248), .A2(n12484), .ZN(n12485) );
  AND4_X1 U14221 ( .A1(n12487), .A2(n15762), .A3(n12486), .A4(n12485), .ZN(
        n12488) );
  OAI211_X1 U14222 ( .C1(n12491), .C2(n12490), .A(n12489), .B(n12488), .ZN(
        n12492) );
  NOR2_X1 U14223 ( .A1(n13896), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12532) );
  INV_X1 U14224 ( .A(n12494), .ZN(n14815) );
  INV_X2 U14225 ( .A(n12541), .ZN(n12650) );
  MUX2_X1 U14226 ( .A(n19758), .B(n19927), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12495) );
  INV_X1 U14227 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18861) );
  OR2_X1 U14228 ( .A1(n12516), .A2(n18861), .ZN(n12499) );
  INV_X1 U14229 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n14822) );
  NAND2_X1 U14230 ( .A1(n13896), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12496) );
  OAI211_X1 U14231 ( .C1(n19758), .C2(n14822), .A(n12496), .B(n19916), .ZN(
        n12497) );
  INV_X1 U14232 ( .A(n12497), .ZN(n12498) );
  NAND2_X1 U14233 ( .A1(n12499), .A2(n12498), .ZN(n14821) );
  INV_X1 U14234 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n18870) );
  OR2_X1 U14235 ( .A1(n12516), .A2(n18870), .ZN(n12503) );
  INV_X1 U14236 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n12500) );
  INV_X1 U14237 ( .A(n12501), .ZN(n12502) );
  NAND2_X1 U14238 ( .A1(n12503), .A2(n12502), .ZN(n12509) );
  INV_X1 U14239 ( .A(n12509), .ZN(n12504) );
  OR2_X1 U14240 ( .A1(n12505), .A2(n12653), .ZN(n12508) );
  NAND2_X1 U14241 ( .A1(n12494), .A2(n19758), .ZN(n12506) );
  MUX2_X1 U14242 ( .A(n12506), .B(n19926), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12507) );
  AND2_X1 U14243 ( .A1(n12508), .A2(n12507), .ZN(n15014) );
  NAND2_X1 U14244 ( .A1(n15015), .A2(n15014), .ZN(n15013) );
  OR2_X1 U14245 ( .A1(n12653), .A2(n12511), .ZN(n12513) );
  OAI211_X1 U14246 ( .C1(n19916), .C2(n19832), .A(n12513), .B(n12512), .ZN(
        n12514) );
  INV_X1 U14247 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n17956) );
  OR2_X1 U14248 ( .A1(n12516), .A2(n17956), .ZN(n12518) );
  AOI22_X1 U14249 ( .A1(n12686), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n12650), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12517) );
  NAND2_X1 U14250 ( .A1(n12518), .A2(n12517), .ZN(n15203) );
  INV_X1 U14251 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n12520) );
  OAI22_X1 U14252 ( .A1(n12516), .A2(n12520), .B1(n15820), .B2(n12541), .ZN(
        n12524) );
  AOI22_X1 U14253 ( .A1(n12686), .A2(P2_EAX_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12521) );
  OAI21_X1 U14254 ( .B1(n12522), .B2(n12653), .A(n12521), .ZN(n12523) );
  OR2_X1 U14255 ( .A1(n12524), .A2(n12523), .ZN(n15409) );
  INV_X1 U14256 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n12525) );
  OR2_X1 U14257 ( .A1(n12516), .A2(n12525), .ZN(n12529) );
  AOI22_X1 U14258 ( .A1(n12686), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n12650), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12528) );
  OR2_X1 U14259 ( .A1(n12653), .A2(n12526), .ZN(n12527) );
  INV_X1 U14260 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n12536) );
  INV_X1 U14261 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n12530) );
  OR2_X1 U14262 ( .A1(n12516), .A2(n12530), .ZN(n12535) );
  INV_X1 U14263 ( .A(n12531), .ZN(n12533) );
  AOI22_X1 U14264 ( .A1(n12533), .A2(n12532), .B1(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n12650), .ZN(n12534) );
  OAI211_X1 U14265 ( .C1(n11237), .C2(n12536), .A(n12535), .B(n12534), .ZN(
        n15818) );
  NOR2_X1 U14266 ( .A1(n12653), .A2(n12537), .ZN(n12538) );
  INV_X1 U14267 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n17957) );
  OR2_X1 U14268 ( .A1(n12516), .A2(n17957), .ZN(n12540) );
  AOI22_X1 U14269 ( .A1(n12686), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n12650), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12539) );
  INV_X1 U14270 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n17932) );
  INV_X1 U14271 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n17958) );
  OAI222_X1 U14272 ( .A1(n12541), .A2(n19196), .B1(n11237), .B2(n17932), .C1(
        n12516), .C2(n17958), .ZN(n14818) );
  INV_X1 U14273 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n12542) );
  OR2_X1 U14274 ( .A1(n12516), .A2(n12542), .ZN(n12555) );
  AOI22_X1 U14275 ( .A1(n12686), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n12650), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12554) );
  AOI22_X1 U14276 ( .A1(n14068), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n14069), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12546) );
  AOI22_X1 U14277 ( .A1(n14071), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14072), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12545) );
  AOI22_X1 U14278 ( .A1(n14126), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11942), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12544) );
  AOI22_X1 U14279 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17363), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12543) );
  NAND4_X1 U14280 ( .A1(n12546), .A2(n12545), .A3(n12544), .A4(n12543), .ZN(
        n12552) );
  AOI22_X1 U14281 ( .A1(n11909), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11901), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12550) );
  AOI22_X1 U14282 ( .A1(n14104), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11921), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12549) );
  AOI22_X1 U14283 ( .A1(n11907), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11962), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12548) );
  AOI22_X1 U14284 ( .A1(n11908), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11906), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12547) );
  NAND4_X1 U14285 ( .A1(n12550), .A2(n12549), .A3(n12548), .A4(n12547), .ZN(
        n12551) );
  NOR2_X1 U14286 ( .A1(n12552), .A2(n12551), .ZN(n15077) );
  OR2_X1 U14287 ( .A1(n12653), .A2(n15077), .ZN(n12553) );
  INV_X1 U14288 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n17962) );
  AOI22_X1 U14289 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n14069), .B1(
        n14068), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12560) );
  AOI22_X1 U14290 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n14071), .B1(
        n14072), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12559) );
  AOI22_X1 U14291 ( .A1(n14126), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11942), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12558) );
  AOI22_X1 U14292 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n12556), .B1(
        n17363), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12557) );
  NAND4_X1 U14293 ( .A1(n12560), .A2(n12559), .A3(n12558), .A4(n12557), .ZN(
        n12566) );
  AOI22_X1 U14294 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11901), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12564) );
  AOI22_X1 U14295 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n11921), .B1(
        n14104), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12563) );
  AOI22_X1 U14296 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11962), .B1(
        n11906), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12562) );
  AOI22_X1 U14297 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n11908), .B1(
        n11907), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12561) );
  NAND4_X1 U14298 ( .A1(n12564), .A2(n12563), .A3(n12562), .A4(n12561), .ZN(
        n12565) );
  INV_X1 U14299 ( .A(n15056), .ZN(n12567) );
  OAI22_X1 U14300 ( .A1(n12516), .A2(n17962), .B1(n12653), .B2(n12567), .ZN(
        n12568) );
  INV_X1 U14301 ( .A(n12568), .ZN(n12570) );
  AOI22_X1 U14302 ( .A1(n12686), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n12650), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12569) );
  NAND2_X1 U14303 ( .A1(n12570), .A2(n12569), .ZN(n14925) );
  INV_X1 U14304 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n12571) );
  OR2_X1 U14305 ( .A1(n12516), .A2(n12571), .ZN(n12585) );
  AOI22_X1 U14306 ( .A1(n12686), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n12650), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12584) );
  AOI22_X1 U14307 ( .A1(n14068), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n14071), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12575) );
  AOI22_X1 U14308 ( .A1(n14069), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14072), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12574) );
  AOI22_X1 U14309 ( .A1(n14126), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11942), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12573) );
  AOI22_X1 U14310 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17363), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12572) );
  NAND4_X1 U14311 ( .A1(n12575), .A2(n12574), .A3(n12573), .A4(n12572), .ZN(
        n12581) );
  AOI22_X1 U14312 ( .A1(n11909), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11901), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12579) );
  AOI22_X1 U14313 ( .A1(n14104), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11921), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12578) );
  AOI22_X1 U14314 ( .A1(n11962), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11906), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12577) );
  AOI22_X1 U14315 ( .A1(n11907), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11908), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12576) );
  NAND4_X1 U14316 ( .A1(n12579), .A2(n12578), .A3(n12577), .A4(n12576), .ZN(
        n12580) );
  INV_X1 U14317 ( .A(n15058), .ZN(n12582) );
  OR2_X1 U14318 ( .A1(n12653), .A2(n12582), .ZN(n12583) );
  AOI22_X1 U14319 ( .A1(n14068), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n14069), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12589) );
  AOI22_X1 U14320 ( .A1(n14071), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n14072), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12588) );
  AOI22_X1 U14321 ( .A1(n14126), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11942), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12587) );
  AOI22_X1 U14322 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17363), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12586) );
  NAND4_X1 U14323 ( .A1(n12589), .A2(n12588), .A3(n12587), .A4(n12586), .ZN(
        n12595) );
  AOI22_X1 U14324 ( .A1(n11909), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11901), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12593) );
  AOI22_X1 U14325 ( .A1(n14104), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11921), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12592) );
  AOI22_X1 U14326 ( .A1(n11962), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11906), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12591) );
  AOI22_X1 U14327 ( .A1(n11907), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11908), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12590) );
  NAND4_X1 U14328 ( .A1(n12593), .A2(n12592), .A3(n12591), .A4(n12590), .ZN(
        n12594) );
  NOR2_X1 U14329 ( .A1(n12595), .A2(n12594), .ZN(n15405) );
  INV_X1 U14330 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n17964) );
  OR2_X1 U14331 ( .A1(n12516), .A2(n17964), .ZN(n12597) );
  AOI22_X1 U14332 ( .A1(n12686), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n12650), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12596) );
  OAI211_X1 U14333 ( .C1(n15405), .C2(n12653), .A(n12597), .B(n12596), .ZN(
        n14995) );
  OR2_X1 U14334 ( .A1(n12516), .A2(n17965), .ZN(n12611) );
  AOI22_X1 U14335 ( .A1(n12686), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n12650), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12610) );
  AOI22_X1 U14336 ( .A1(n14069), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14126), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12601) );
  AOI22_X1 U14337 ( .A1(n14068), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n14072), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12600) );
  AOI22_X1 U14338 ( .A1(n14071), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11942), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12599) );
  AOI22_X1 U14339 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11921), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12598) );
  NAND4_X1 U14340 ( .A1(n12601), .A2(n12600), .A3(n12599), .A4(n12598), .ZN(
        n12607) );
  AOI22_X1 U14341 ( .A1(n11909), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11901), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12605) );
  AOI22_X1 U14342 ( .A1(n14104), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17363), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12604) );
  AOI22_X1 U14343 ( .A1(n11962), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11906), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12603) );
  AOI22_X1 U14344 ( .A1(n11907), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11908), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12602) );
  NAND4_X1 U14345 ( .A1(n12605), .A2(n12604), .A3(n12603), .A4(n12602), .ZN(
        n12606) );
  INV_X1 U14346 ( .A(n15360), .ZN(n12608) );
  OR2_X1 U14347 ( .A1(n12653), .A2(n12608), .ZN(n12609) );
  INV_X1 U14348 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n12612) );
  OR2_X1 U14349 ( .A1(n12516), .A2(n12612), .ZN(n12625) );
  AOI22_X1 U14350 ( .A1(n12686), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n12650), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12624) );
  AOI22_X1 U14351 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n14069), .B1(
        n14068), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12616) );
  AOI22_X1 U14352 ( .A1(n14071), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14072), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12615) );
  AOI22_X1 U14353 ( .A1(n14126), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11942), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12614) );
  AOI22_X1 U14354 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17363), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12613) );
  NAND4_X1 U14355 ( .A1(n12616), .A2(n12615), .A3(n12614), .A4(n12613), .ZN(
        n12622) );
  AOI22_X1 U14356 ( .A1(n11909), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11901), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12620) );
  AOI22_X1 U14357 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n11921), .B1(
        n14104), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12619) );
  AOI22_X1 U14358 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n11962), .B1(
        n11906), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12618) );
  AOI22_X1 U14359 ( .A1(n11907), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11908), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12617) );
  NAND4_X1 U14360 ( .A1(n12620), .A2(n12619), .A3(n12618), .A4(n12617), .ZN(
        n12621) );
  NOR2_X1 U14361 ( .A1(n12622), .A2(n12621), .ZN(n15628) );
  OR2_X1 U14362 ( .A1(n12653), .A2(n15628), .ZN(n12623) );
  AOI22_X1 U14363 ( .A1(n14069), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14126), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12630) );
  AOI22_X1 U14364 ( .A1(n14068), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11942), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12629) );
  AOI22_X1 U14365 ( .A1(n14071), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14072), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12628) );
  AOI22_X1 U14366 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17363), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12627) );
  NAND4_X1 U14367 ( .A1(n12630), .A2(n12629), .A3(n12628), .A4(n12627), .ZN(
        n12636) );
  AOI22_X1 U14368 ( .A1(n11909), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11901), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12634) );
  AOI22_X1 U14369 ( .A1(n14104), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11921), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12633) );
  AOI22_X1 U14370 ( .A1(n11962), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11906), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12632) );
  AOI22_X1 U14371 ( .A1(n11907), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11908), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12631) );
  NAND4_X1 U14372 ( .A1(n12634), .A2(n12633), .A3(n12632), .A4(n12631), .ZN(
        n12635) );
  INV_X1 U14373 ( .A(n15565), .ZN(n12639) );
  OR2_X1 U14374 ( .A1(n12516), .A2(n17966), .ZN(n12638) );
  AOI22_X1 U14375 ( .A1(n12686), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n12650), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12637) );
  OAI211_X1 U14376 ( .C1(n12639), .C2(n12653), .A(n12638), .B(n12637), .ZN(
        n15727) );
  AOI22_X1 U14377 ( .A1(n14068), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n14069), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12643) );
  AOI22_X1 U14378 ( .A1(n14071), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n14072), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12642) );
  AOI22_X1 U14379 ( .A1(n14126), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11942), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12641) );
  AOI22_X1 U14380 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17363), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12640) );
  NAND4_X1 U14381 ( .A1(n12643), .A2(n12642), .A3(n12641), .A4(n12640), .ZN(
        n12649) );
  AOI22_X1 U14382 ( .A1(n11909), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11901), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12647) );
  AOI22_X1 U14383 ( .A1(n14104), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11921), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12646) );
  AOI22_X1 U14384 ( .A1(n11962), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11906), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12645) );
  AOI22_X1 U14385 ( .A1(n11907), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11908), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12644) );
  NAND4_X1 U14386 ( .A1(n12647), .A2(n12646), .A3(n12645), .A4(n12644), .ZN(
        n12648) );
  NOR2_X1 U14387 ( .A1(n12649), .A2(n12648), .ZN(n15709) );
  NAND2_X1 U14388 ( .A1(n12678), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n12652) );
  INV_X2 U14389 ( .A(n11237), .ZN(n12686) );
  AOI22_X1 U14390 ( .A1(n12686), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n12650), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12651) );
  OAI211_X1 U14391 ( .C1(n15709), .C2(n12653), .A(n12652), .B(n12651), .ZN(
        n15110) );
  INV_X1 U14392 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n18989) );
  OR2_X1 U14393 ( .A1(n12516), .A2(n18989), .ZN(n12655) );
  AOI22_X1 U14394 ( .A1(n12686), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n12650), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12654) );
  NAND2_X1 U14395 ( .A1(n12655), .A2(n12654), .ZN(n15695) );
  INV_X1 U14396 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n17969) );
  OR2_X1 U14397 ( .A1(n12516), .A2(n17969), .ZN(n12657) );
  AOI22_X1 U14398 ( .A1(n12686), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n12650), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12656) );
  INV_X1 U14399 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19011) );
  OR2_X1 U14400 ( .A1(n12516), .A2(n19011), .ZN(n12659) );
  AOI22_X1 U14401 ( .A1(n12686), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n12650), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12658) );
  NAND2_X1 U14402 ( .A1(n12659), .A2(n12658), .ZN(n15878) );
  INV_X1 U14403 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19026) );
  OR2_X1 U14404 ( .A1(n12516), .A2(n19026), .ZN(n12661) );
  AOI22_X1 U14405 ( .A1(n12686), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n12650), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12660) );
  INV_X1 U14406 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19040) );
  OR2_X1 U14407 ( .A1(n12516), .A2(n19040), .ZN(n12663) );
  AOI22_X1 U14408 ( .A1(n12686), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n12650), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12662) );
  INV_X1 U14409 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n17971) );
  OR2_X1 U14410 ( .A1(n12516), .A2(n17971), .ZN(n12665) );
  AOI22_X1 U14411 ( .A1(n12686), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n12650), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12664) );
  NAND2_X1 U14412 ( .A1(n12665), .A2(n12664), .ZN(n12827) );
  INV_X1 U14413 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n17972) );
  OR2_X1 U14414 ( .A1(n12516), .A2(n17972), .ZN(n12667) );
  AOI22_X1 U14415 ( .A1(n12686), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n12650), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12666) );
  NAND2_X1 U14416 ( .A1(n12667), .A2(n12666), .ZN(n17112) );
  NAND2_X1 U14417 ( .A1(n12826), .A2(n17112), .ZN(n16794) );
  OR2_X1 U14418 ( .A1(n12516), .A2(n17973), .ZN(n12669) );
  AOI22_X1 U14419 ( .A1(n12686), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n12650), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12668) );
  AND2_X1 U14420 ( .A1(n12669), .A2(n12668), .ZN(n16795) );
  INV_X1 U14421 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n17974) );
  OR2_X1 U14422 ( .A1(n12516), .A2(n17974), .ZN(n12671) );
  AOI22_X1 U14423 ( .A1(n12686), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n12650), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12670) );
  INV_X1 U14424 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n17976) );
  OR2_X1 U14425 ( .A1(n12516), .A2(n17976), .ZN(n12673) );
  AOI22_X1 U14426 ( .A1(n12686), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n12650), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12672) );
  INV_X1 U14427 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n17977) );
  OR2_X1 U14428 ( .A1(n12516), .A2(n17977), .ZN(n12675) );
  AOI22_X1 U14429 ( .A1(n12686), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n12650), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12674) );
  NAND2_X1 U14430 ( .A1(n12675), .A2(n12674), .ZN(n16767) );
  INV_X1 U14431 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n17979) );
  OR2_X1 U14432 ( .A1(n12516), .A2(n17979), .ZN(n12677) );
  AOI22_X1 U14433 ( .A1(n12686), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n12650), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12676) );
  AND2_X1 U14434 ( .A1(n12677), .A2(n12676), .ZN(n16757) );
  NAND2_X1 U14435 ( .A1(n12678), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12680) );
  AOI22_X1 U14436 ( .A1(n12686), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n12650), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12679) );
  AND2_X1 U14437 ( .A1(n12680), .A2(n12679), .ZN(n16664) );
  INV_X1 U14438 ( .A(n16664), .ZN(n12681) );
  INV_X1 U14439 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n17982) );
  OR2_X1 U14440 ( .A1(n12516), .A2(n17982), .ZN(n12683) );
  AOI22_X1 U14441 ( .A1(n12686), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n12650), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12682) );
  NAND2_X1 U14442 ( .A1(n12683), .A2(n12682), .ZN(n16744) );
  INV_X1 U14443 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n17983) );
  OR2_X1 U14444 ( .A1(n12516), .A2(n17983), .ZN(n12685) );
  AOI22_X1 U14445 ( .A1(n12686), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n12650), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12684) );
  NAND2_X1 U14446 ( .A1(n12685), .A2(n12684), .ZN(n12785) );
  INV_X1 U14447 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19152) );
  AOI22_X1 U14448 ( .A1(n12686), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n12650), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12687) );
  OAI21_X1 U14449 ( .B1(n12516), .B2(n19152), .A(n12687), .ZN(n12688) );
  INV_X1 U14450 ( .A(n12689), .ZN(n12691) );
  NAND2_X1 U14451 ( .A1(n12691), .A2(n12690), .ZN(n17343) );
  NAND2_X1 U14452 ( .A1(n19245), .A2(n13896), .ZN(n12693) );
  AND2_X1 U14453 ( .A1(n17343), .A2(n12693), .ZN(n12694) );
  NOR2_X2 U14454 ( .A1(n12736), .A2(n12694), .ZN(n19208) );
  NAND2_X1 U14455 ( .A1(n19158), .A2(n19208), .ZN(n12754) );
  AOI22_X1 U14456 ( .A1(n12703), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n12696) );
  NAND2_X1 U14457 ( .A1(n12700), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12695) );
  NAND2_X1 U14458 ( .A1(n12696), .A2(n12695), .ZN(n12697) );
  AOI21_X1 U14459 ( .B1(n12698), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n12697), .ZN(n16680) );
  AOI22_X1 U14460 ( .A1(n11843), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n12702) );
  NAND2_X1 U14461 ( .A1(n12700), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12701) );
  OAI211_X1 U14462 ( .C1(n12706), .C2(n12791), .A(n12702), .B(n12701), .ZN(
        n12793) );
  AOI22_X1 U14463 ( .A1(n12703), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n12705) );
  NAND2_X1 U14464 ( .A1(n12700), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n12704) );
  OAI211_X1 U14465 ( .C1(n12706), .C2(n13846), .A(n12705), .B(n12704), .ZN(
        n12707) );
  AOI21_X1 U14466 ( .B1(n12709), .B2(n14673), .A(n12710), .ZN(n12711) );
  NAND3_X1 U14467 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17036) );
  OR2_X1 U14468 ( .A1(n12791), .A2(n17036), .ZN(n12749) );
  INV_X1 U14469 ( .A(n12712), .ZN(n12713) );
  INV_X1 U14470 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19184) );
  NOR2_X1 U14471 ( .A1(n19184), .A2(n14746), .ZN(n17319) );
  NAND2_X1 U14472 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n17319), .ZN(
        n16004) );
  INV_X1 U14473 ( .A(n16004), .ZN(n15997) );
  INV_X1 U14474 ( .A(n17319), .ZN(n15996) );
  NAND2_X1 U14475 ( .A1(n16001), .A2(n15996), .ZN(n16003) );
  INV_X1 U14476 ( .A(n17171), .ZN(n16002) );
  NAND2_X1 U14477 ( .A1(n12715), .A2(n13896), .ZN(n15755) );
  NAND2_X1 U14478 ( .A1(n15755), .A2(n12716), .ZN(n12718) );
  NAND2_X1 U14479 ( .A1(n12718), .A2(n12717), .ZN(n12731) );
  INV_X1 U14480 ( .A(n12719), .ZN(n12721) );
  NAND2_X1 U14481 ( .A1(n12721), .A2(n12720), .ZN(n12724) );
  INV_X1 U14482 ( .A(n14809), .ZN(n12723) );
  MUX2_X1 U14483 ( .A(n12724), .B(n12723), .S(n12722), .Z(n12730) );
  INV_X1 U14484 ( .A(n12725), .ZN(n14664) );
  NAND2_X1 U14485 ( .A1(n12726), .A2(n11762), .ZN(n12727) );
  AOI22_X1 U14486 ( .A1(n14664), .A2(n12727), .B1(n20247), .B2(n12442), .ZN(
        n12729) );
  NAND4_X1 U14487 ( .A1(n12731), .A2(n12730), .A3(n12729), .A4(n12728), .ZN(
        n17364) );
  NOR2_X1 U14488 ( .A1(n17364), .A2(n12732), .ZN(n12733) );
  INV_X1 U14489 ( .A(n17174), .ZN(n12734) );
  OAI211_X1 U14490 ( .C1(n17171), .C2(n15997), .A(n16003), .B(n19183), .ZN(
        n17309) );
  NAND3_X1 U14491 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17308) );
  NOR2_X1 U14492 ( .A1(n11297), .A2(n17308), .ZN(n17291) );
  NAND3_X1 U14493 ( .A1(n17291), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12739) );
  INV_X1 U14494 ( .A(n17139), .ZN(n17125) );
  NOR2_X1 U14495 ( .A1(n17211), .A2(n17125), .ZN(n17131) );
  AND2_X1 U14496 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12742) );
  NAND2_X1 U14497 ( .A1(n17131), .A2(n12742), .ZN(n12824) );
  NOR2_X1 U14498 ( .A1(n12825), .A2(n12824), .ZN(n17101) );
  NAND3_X1 U14499 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n17101), .ZN(n12747) );
  NOR2_X1 U14500 ( .A1(n11610), .A2(n12747), .ZN(n17067) );
  NAND3_X1 U14501 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(n17067), .ZN(n17035) );
  NOR3_X1 U14502 ( .A1(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n12749), .A3(
        n17035), .ZN(n12752) );
  INV_X1 U14503 ( .A(n19183), .ZN(n17318) );
  NOR2_X1 U14504 ( .A1(n17066), .A2(n17079), .ZN(n12748) );
  INV_X1 U14505 ( .A(n16003), .ZN(n12735) );
  NAND2_X1 U14506 ( .A1(n17171), .A2(n12735), .ZN(n12737) );
  NAND2_X1 U14507 ( .A1(n12736), .A2(n18976), .ZN(n19176) );
  NAND2_X1 U14508 ( .A1(n12737), .A2(n19176), .ZN(n15442) );
  AND2_X1 U14509 ( .A1(n17171), .A2(n12739), .ZN(n12738) );
  NOR2_X1 U14510 ( .A1(n15442), .A2(n12738), .ZN(n17130) );
  INV_X1 U14511 ( .A(n12739), .ZN(n12740) );
  NAND2_X1 U14512 ( .A1(n12740), .A2(n15997), .ZN(n17124) );
  NAND2_X1 U14513 ( .A1(n17174), .A2(n17124), .ZN(n12741) );
  NAND2_X1 U14514 ( .A1(n17130), .A2(n12741), .ZN(n17286) );
  NAND3_X1 U14515 ( .A1(n17139), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n12742), .ZN(n12743) );
  AND2_X1 U14516 ( .A1(n19183), .A2(n12743), .ZN(n12744) );
  OR2_X1 U14517 ( .A1(n17286), .A2(n12744), .ZN(n12823) );
  OR2_X1 U14518 ( .A1(n17110), .A2(n17100), .ZN(n12745) );
  AND2_X1 U14519 ( .A1(n19183), .A2(n12745), .ZN(n12746) );
  OR2_X1 U14520 ( .A1(n12823), .A2(n12746), .ZN(n17092) );
  NOR2_X1 U14521 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n12747), .ZN(
        n17090) );
  NOR2_X1 U14522 ( .A1(n17092), .A2(n17090), .ZN(n17080) );
  OAI21_X1 U14523 ( .B1(n17318), .B2(n12748), .A(n17080), .ZN(n17062) );
  AOI21_X1 U14524 ( .B1(n12749), .B2(n19183), .A(n17062), .ZN(n12792) );
  INV_X2 U14525 ( .A(n19213), .ZN(n18976) );
  NOR2_X1 U14526 ( .A1(n18976), .A2(n19152), .ZN(n14294) );
  INV_X1 U14527 ( .A(n14294), .ZN(n12750) );
  OAI21_X1 U14528 ( .B1(n12792), .B2(n13846), .A(n12750), .ZN(n12751) );
  XNOR2_X1 U14529 ( .A(n12756), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14302) );
  INV_X1 U14530 ( .A(n14302), .ZN(n12759) );
  NAND2_X1 U14531 ( .A1(n12759), .A2(n12758), .ZN(n12760) );
  OAI21_X1 U14532 ( .B1(n11154), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n12762), .ZN(n17077) );
  INV_X1 U14533 ( .A(n11631), .ZN(n12763) );
  AOI21_X1 U14534 ( .B1(n12763), .B2(n16857), .A(n16858), .ZN(n12769) );
  NAND2_X1 U14535 ( .A1(n12768), .A2(n12765), .ZN(n12766) );
  AND2_X1 U14536 ( .A1(n11515), .A2(n12771), .ZN(n12772) );
  NOR2_X1 U14537 ( .A1(n12770), .A2(n12772), .ZN(n19110) );
  NAND2_X1 U14538 ( .A1(n13879), .A2(n12773), .ZN(n12774) );
  NAND2_X1 U14539 ( .A1(n13883), .A2(n12774), .ZN(n19113) );
  NOR2_X1 U14540 ( .A1(n18976), .A2(n17977), .ZN(n17068) );
  AOI21_X1 U14541 ( .B1(n17866), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n17068), .ZN(n12775) );
  OAI21_X1 U14542 ( .B1(n17883), .B2(n19113), .A(n12775), .ZN(n12776) );
  XOR2_X1 U14543 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n11155), .Z(
        n16833) );
  NAND2_X1 U14544 ( .A1(n12779), .A2(n16841), .ZN(n12784) );
  INV_X1 U14545 ( .A(n12780), .ZN(n12782) );
  NAND2_X1 U14546 ( .A1(n12782), .A2(n12781), .ZN(n12783) );
  NAND2_X1 U14547 ( .A1(n16831), .A2(n19211), .ZN(n12797) );
  NOR2_X1 U14548 ( .A1(n18976), .A2(n17983), .ZN(n16827) );
  INV_X1 U14549 ( .A(n16827), .ZN(n12788) );
  INV_X1 U14550 ( .A(n12789), .ZN(n12790) );
  OAI21_X1 U14551 ( .B1(n12792), .B2(n12791), .A(n12790), .ZN(n12795) );
  NOR2_X1 U14552 ( .A1(n16829), .A2(n17283), .ZN(n12794) );
  NOR2_X1 U14553 ( .A1(n12795), .A2(n12794), .ZN(n12796) );
  OAI21_X1 U14554 ( .B1(n16833), .B2(n19187), .A(n11633), .ZN(P2_U3016) );
  INV_X1 U14555 ( .A(n16999), .ZN(n12798) );
  NAND2_X1 U14556 ( .A1(n16969), .A2(n12800), .ZN(n12802) );
  NAND2_X1 U14557 ( .A1(n12802), .A2(n12801), .ZN(n16931) );
  NAND2_X1 U14558 ( .A1(n16931), .A2(n16930), .ZN(n16932) );
  INV_X1 U14559 ( .A(n16919), .ZN(n12804) );
  NAND2_X1 U14560 ( .A1(n12809), .A2(n12808), .ZN(n12810) );
  XNOR2_X1 U14561 ( .A(n12811), .B(n12810), .ZN(n12822) );
  NAND2_X1 U14562 ( .A1(n12822), .A2(n17879), .ZN(n12821) );
  OAI21_X1 U14563 ( .B1(n11232), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n12812), .ZN(n12834) );
  AOI21_X1 U14564 ( .B1(n11236), .B2(n12359), .A(n13847), .ZN(n13876) );
  NAND2_X1 U14565 ( .A1(n19213), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12829) );
  OAI21_X1 U14566 ( .B1(n17029), .B2(n12359), .A(n12829), .ZN(n12817) );
  NAND2_X1 U14567 ( .A1(n12813), .A2(n12814), .ZN(n12815) );
  NAND2_X1 U14568 ( .A1(n12331), .A2(n12815), .ZN(n19054) );
  NOR2_X1 U14569 ( .A1(n19054), .A2(n17865), .ZN(n12816) );
  AOI211_X1 U14570 ( .C1(n17850), .C2(n13876), .A(n12817), .B(n12816), .ZN(
        n12818) );
  INV_X1 U14571 ( .A(n12819), .ZN(n12820) );
  NAND2_X1 U14572 ( .A1(n12821), .A2(n12820), .ZN(P2_U2993) );
  NAND2_X1 U14573 ( .A1(n12822), .A2(n19211), .ZN(n12837) );
  INV_X1 U14574 ( .A(n19054), .ZN(n12832) );
  INV_X1 U14575 ( .A(n12823), .ZN(n17111) );
  AOI21_X1 U14576 ( .B1(n12825), .B2(n12824), .A(n17111), .ZN(n12831) );
  NOR2_X1 U14577 ( .A1(n17135), .A2(n12827), .ZN(n12828) );
  OR2_X1 U14578 ( .A1(n12826), .A2(n12828), .ZN(n19053) );
  OAI21_X1 U14579 ( .B1(n19180), .B2(n19053), .A(n12829), .ZN(n12830) );
  AOI211_X1 U14580 ( .C1(n12832), .C2(n19202), .A(n12831), .B(n12830), .ZN(
        n12833) );
  NAND2_X1 U14581 ( .A1(n12837), .A2(n12836), .ZN(P2_U3025) );
  INV_X1 U14582 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12839) );
  AND2_X2 U14583 ( .A1(n12839), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12846) );
  AOI22_X1 U14584 ( .A1(n13185), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13083), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12845) );
  NOR2_X4 U14585 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12841) );
  NOR2_X4 U14586 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14961) );
  AND2_X2 U14587 ( .A1(n14961), .A2(n12841), .ZN(n13444) );
  AOI22_X1 U14588 ( .A1(n11177), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13444), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12844) );
  AND2_X4 U14589 ( .A1(n12841), .A2(n14872), .ZN(n13433) );
  AOI22_X1 U14590 ( .A1(n12894), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13433), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12843) );
  AND2_X4 U14591 ( .A1(n12846), .A2(n14961), .ZN(n13809) );
  AOI22_X1 U14592 ( .A1(n13809), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11165), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12842) );
  AND2_X2 U14593 ( .A1(n16603), .A2(n14961), .ZN(n13012) );
  AOI22_X1 U14594 ( .A1(n13012), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11172), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12853) );
  AND2_X2 U14595 ( .A1(n16603), .A2(n14872), .ZN(n13018) );
  AOI22_X1 U14596 ( .A1(n11169), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13018), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12852) );
  AOI22_X1 U14597 ( .A1(n13136), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11168), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12851) );
  AOI22_X1 U14598 ( .A1(n13377), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12997), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12850) );
  NAND2_X1 U14599 ( .A1(n12855), .A2(n12854), .ZN(n12950) );
  AOI22_X1 U14600 ( .A1(n13377), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13012), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12859) );
  AOI22_X1 U14601 ( .A1(n12894), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13083), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12858) );
  AOI22_X1 U14602 ( .A1(n13013), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13433), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12857) );
  AOI22_X1 U14603 ( .A1(n13809), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11165), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12856) );
  NAND4_X1 U14604 ( .A1(n12859), .A2(n12858), .A3(n12857), .A4(n12856), .ZN(
        n12865) );
  AOI22_X1 U14605 ( .A1(n12899), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12997), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12863) );
  AOI22_X1 U14606 ( .A1(n13136), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13185), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12862) );
  AOI22_X1 U14607 ( .A1(n13082), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13018), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12861) );
  AOI22_X1 U14608 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13444), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12860) );
  NAND4_X1 U14609 ( .A1(n12863), .A2(n12862), .A3(n12861), .A4(n12860), .ZN(
        n12864) );
  AOI22_X1 U14610 ( .A1(n13136), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13083), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12869) );
  AOI22_X1 U14611 ( .A1(n13809), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13444), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12867) );
  AOI22_X1 U14612 ( .A1(n12899), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12997), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12866) );
  AOI22_X1 U14613 ( .A1(n13377), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13012), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12873) );
  AOI22_X1 U14614 ( .A1(n13185), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12894), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12872) );
  AOI22_X1 U14615 ( .A1(n13013), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13433), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12871) );
  AOI22_X1 U14616 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11165), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12870) );
  NAND2_X2 U14617 ( .A1(n11653), .A2(n11212), .ZN(n13009) );
  AOI22_X1 U14618 ( .A1(n13012), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12899), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12877) );
  AOI22_X1 U14619 ( .A1(n13082), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13018), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12876) );
  AOI22_X1 U14620 ( .A1(n13136), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13013), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12875) );
  AOI22_X1 U14621 ( .A1(n13377), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12997), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12874) );
  NAND4_X1 U14622 ( .A1(n12877), .A2(n12876), .A3(n12875), .A4(n12874), .ZN(
        n12883) );
  AOI22_X1 U14623 ( .A1(n13185), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13083), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12881) );
  AOI22_X1 U14624 ( .A1(n11177), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13444), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12880) );
  AOI22_X1 U14625 ( .A1(n11171), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13433), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12879) );
  AOI22_X1 U14626 ( .A1(n13809), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11165), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12878) );
  NAND4_X1 U14627 ( .A1(n12881), .A2(n12880), .A3(n12879), .A4(n12878), .ZN(
        n12882) );
  AOI22_X1 U14628 ( .A1(n13082), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13013), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12887) );
  AOI22_X1 U14629 ( .A1(n13083), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13809), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12886) );
  AOI22_X1 U14630 ( .A1(n12899), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12997), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12885) );
  AOI22_X1 U14631 ( .A1(n13136), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13433), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12884) );
  NAND4_X1 U14632 ( .A1(n12887), .A2(n12886), .A3(n12885), .A4(n12884), .ZN(
        n12893) );
  AOI22_X1 U14633 ( .A1(n13377), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13012), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12891) );
  AOI22_X1 U14634 ( .A1(n13018), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11171), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12890) );
  AOI22_X1 U14635 ( .A1(n11146), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13444), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12889) );
  NAND4_X1 U14636 ( .A1(n12891), .A2(n12890), .A3(n12889), .A4(n12888), .ZN(
        n12892) );
  AOI22_X1 U14637 ( .A1(n11146), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13444), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12897) );
  AOI22_X1 U14638 ( .A1(n11171), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13433), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12896) );
  AOI22_X1 U14639 ( .A1(n13809), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11165), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12895) );
  NAND4_X1 U14640 ( .A1(n12898), .A2(n12897), .A3(n12896), .A4(n12895), .ZN(
        n12905) );
  AOI22_X1 U14641 ( .A1(n13012), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12899), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12903) );
  AOI22_X1 U14642 ( .A1(n13082), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13018), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12902) );
  AOI22_X1 U14643 ( .A1(n13136), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13013), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12901) );
  AOI22_X1 U14644 ( .A1(n13377), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12997), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12900) );
  NAND4_X1 U14645 ( .A1(n12903), .A2(n12902), .A3(n12901), .A4(n12900), .ZN(
        n12904) );
  AND3_X2 U14646 ( .A1(n12906), .A2(n16192), .A3(n14858), .ZN(n14828) );
  NAND2_X1 U14647 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12910) );
  NAND2_X1 U14648 ( .A1(n13809), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12909) );
  NAND2_X1 U14649 ( .A1(n13444), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12908) );
  NAND2_X1 U14650 ( .A1(n11165), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12907) );
  NAND2_X1 U14651 ( .A1(n13377), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12914) );
  NAND2_X1 U14652 ( .A1(n13012), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12913) );
  NAND2_X1 U14653 ( .A1(n12899), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12912) );
  NAND2_X1 U14654 ( .A1(n12997), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12911) );
  NAND2_X1 U14655 ( .A1(n11171), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12917) );
  NAND2_X1 U14656 ( .A1(n13185), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12916) );
  NAND3_X1 U14657 ( .A1(n12919), .A2(n12918), .A3(n11224), .ZN(n12924) );
  NAND2_X1 U14658 ( .A1(n13082), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12923) );
  NAND2_X1 U14659 ( .A1(n13018), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12922) );
  NAND2_X1 U14660 ( .A1(n13136), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12921) );
  NAND2_X1 U14661 ( .A1(n13013), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12920) );
  INV_X1 U14662 ( .A(n14693), .ZN(n12948) );
  NAND2_X1 U14663 ( .A1(n13377), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12928) );
  NAND2_X1 U14664 ( .A1(n13012), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12927) );
  NAND2_X1 U14665 ( .A1(n12899), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12926) );
  NAND2_X1 U14666 ( .A1(n12997), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12925) );
  NAND2_X1 U14667 ( .A1(n13082), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12932) );
  NAND2_X1 U14668 ( .A1(n13018), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12931) );
  NAND2_X1 U14669 ( .A1(n13136), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12930) );
  NAND2_X1 U14670 ( .A1(n13013), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12929) );
  NAND2_X1 U14671 ( .A1(n11171), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12936) );
  NAND2_X1 U14672 ( .A1(n13185), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12935) );
  NAND2_X1 U14673 ( .A1(n13083), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12934) );
  NAND2_X1 U14674 ( .A1(n13433), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12933) );
  NAND2_X1 U14675 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12940) );
  NAND2_X1 U14676 ( .A1(n13809), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12939) );
  NAND2_X1 U14677 ( .A1(n13444), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12938) );
  NAND2_X1 U14678 ( .A1(n11165), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12937) );
  NAND2_X1 U14679 ( .A1(n22311), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n12945) );
  NAND2_X1 U14680 ( .A1(n22304), .A2(n12945), .ZN(n14847) );
  NAND2_X1 U14681 ( .A1(n15379), .A2(n11173), .ZN(n12967) );
  INV_X1 U14682 ( .A(n12967), .ZN(n12946) );
  NAND2_X1 U14683 ( .A1(n11195), .A2(n12946), .ZN(n14829) );
  NAND2_X1 U14684 ( .A1(n13915), .A2(n13911), .ZN(n15992) );
  OR2_X2 U14685 ( .A1(n14829), .A2(n15992), .ZN(n14908) );
  INV_X1 U14686 ( .A(n14908), .ZN(n12947) );
  NAND2_X1 U14687 ( .A1(n14899), .A2(n13009), .ZN(n12949) );
  MUX2_X1 U14688 ( .A(n12955), .B(n12949), .S(n13911), .Z(n12954) );
  INV_X2 U14689 ( .A(n12950), .ZN(n16023) );
  NAND2_X1 U14690 ( .A1(n11654), .A2(n12951), .ZN(n12973) );
  NAND2_X1 U14691 ( .A1(n15167), .A2(n13915), .ZN(n12952) );
  NAND2_X1 U14692 ( .A1(n12973), .A2(n12952), .ZN(n12953) );
  NAND2_X1 U14693 ( .A1(n14686), .A2(n15379), .ZN(n14827) );
  NAND2_X1 U14694 ( .A1(n12958), .A2(n14827), .ZN(n12959) );
  NAND2_X1 U14695 ( .A1(n12959), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12984) );
  AND2_X2 U14696 ( .A1(n15379), .A2(n16021), .ZN(n21878) );
  NAND2_X1 U14697 ( .A1(n16022), .A2(n13911), .ZN(n12960) );
  INV_X1 U14698 ( .A(n12955), .ZN(n12961) );
  NAND2_X1 U14699 ( .A1(n12964), .A2(n15229), .ZN(n15239) );
  NAND2_X1 U14700 ( .A1(n14919), .A2(n15239), .ZN(n12965) );
  AOI21_X1 U14701 ( .B1(n21878), .B2(n12970), .A(n12965), .ZN(n12969) );
  AND2_X1 U14702 ( .A1(n14833), .A2(n12966), .ZN(n12968) );
  NAND2_X1 U14703 ( .A1(n12969), .A2(n14840), .ZN(n12995) );
  INV_X1 U14704 ( .A(n12970), .ZN(n12972) );
  NAND2_X1 U14705 ( .A1(n12972), .A2(n12971), .ZN(n14842) );
  NAND2_X1 U14706 ( .A1(n14842), .A2(n16592), .ZN(n12978) );
  INV_X1 U14707 ( .A(n12975), .ZN(n12976) );
  NAND2_X1 U14708 ( .A1(n16026), .A2(n16021), .ZN(n14834) );
  NAND2_X1 U14709 ( .A1(n13073), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12983) );
  NAND2_X1 U14710 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n13075) );
  OAI21_X1 U14711 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n13075), .ZN(n22372) );
  INV_X1 U14712 ( .A(n13312), .ZN(n13108) );
  NAND2_X1 U14713 ( .A1(n13108), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n13070) );
  OAI21_X1 U14714 ( .B1(n13838), .B2(n22372), .A(n13070), .ZN(n12981) );
  INV_X1 U14715 ( .A(n12981), .ZN(n12982) );
  NAND2_X1 U14716 ( .A1(n12983), .A2(n12982), .ZN(n12986) );
  INV_X1 U14717 ( .A(n12984), .ZN(n12985) );
  XNOR2_X2 U14718 ( .A(n12986), .B(n12985), .ZN(n15093) );
  NAND2_X1 U14719 ( .A1(n13073), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12988) );
  MUX2_X1 U14720 ( .A(n13838), .B(n13312), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n12987) );
  NAND2_X1 U14721 ( .A1(n12988), .A2(n12987), .ZN(n13030) );
  NAND3_X1 U14722 ( .A1(n14842), .A2(n15229), .A3(n16592), .ZN(n12993) );
  NAND2_X1 U14723 ( .A1(n16596), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20598) );
  AOI21_X1 U14724 ( .B1(n12966), .B2(n16021), .A(n20598), .ZN(n12992) );
  AND2_X1 U14725 ( .A1(n16037), .A2(n12989), .ZN(n14786) );
  NAND2_X1 U14726 ( .A1(n14786), .A2(n12990), .ZN(n12991) );
  NAND2_X1 U14727 ( .A1(n12975), .A2(n16023), .ZN(n14918) );
  NAND4_X1 U14728 ( .A1(n12993), .A2(n12992), .A3(n12991), .A4(n14918), .ZN(
        n12994) );
  OR2_X1 U14729 ( .A1(n12995), .A2(n12994), .ZN(n13028) );
  NAND2_X1 U14730 ( .A1(n13030), .A2(n13028), .ZN(n12996) );
  OR2_X2 U14731 ( .A1(n15093), .A2(n12996), .ZN(n13069) );
  AOI22_X1 U14732 ( .A1(n13801), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13001) );
  AOI22_X1 U14733 ( .A1(n13804), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13809), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13000) );
  AOI22_X1 U14734 ( .A1(n11146), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12999) );
  AOI22_X1 U14735 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12998) );
  NAND4_X1 U14736 ( .A1(n13001), .A2(n13000), .A3(n12999), .A4(n12998), .ZN(
        n13007) );
  AOI22_X1 U14737 ( .A1(n13563), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12899), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13005) );
  AOI22_X1 U14738 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13013), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13004) );
  AOI22_X1 U14739 ( .A1(n13779), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13433), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13003) );
  AOI22_X1 U14740 ( .A1(n13778), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13002) );
  NAND4_X1 U14741 ( .A1(n13005), .A2(n13004), .A3(n13003), .A4(n13002), .ZN(
        n13006) );
  NAND2_X1 U14742 ( .A1(n13066), .A2(n13057), .ZN(n13008) );
  INV_X1 U14743 ( .A(n13062), .ZN(n13011) );
  NAND2_X1 U14744 ( .A1(n13011), .A2(n13010), .ZN(n13027) );
  AOI22_X1 U14745 ( .A1(n13563), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12899), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13017) );
  AOI22_X1 U14746 ( .A1(n13801), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13013), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13016) );
  AOI22_X1 U14747 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13015) );
  AOI22_X1 U14748 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n11146), .B1(
        n13433), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13014) );
  NAND4_X1 U14749 ( .A1(n13017), .A2(n13016), .A3(n13015), .A4(n13014), .ZN(
        n13024) );
  AOI22_X1 U14750 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n13810), .B1(
        n13731), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13022) );
  AOI22_X1 U14751 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n13804), .B1(
        n13779), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13021) );
  AOI22_X1 U14752 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n13809), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13020) );
  AOI22_X1 U14753 ( .A1(n13778), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13019) );
  NAND4_X1 U14754 ( .A1(n13022), .A2(n13021), .A3(n13020), .A4(n13019), .ZN(
        n13023) );
  NAND2_X1 U14755 ( .A1(n13057), .A2(n13031), .ZN(n13129) );
  OAI211_X1 U14756 ( .C1(n13057), .C2(n13031), .A(n21878), .B(n13129), .ZN(
        n13025) );
  AND3_X1 U14757 ( .A1(n13025), .A2(n14858), .A3(n13009), .ZN(n13026) );
  NAND2_X1 U14758 ( .A1(n13027), .A2(n13026), .ZN(n13054) );
  XNOR2_X1 U14759 ( .A(n13030), .B(n13029), .ZN(n13340) );
  NAND2_X1 U14760 ( .A1(n13340), .A2(n22274), .ZN(n13045) );
  AOI22_X1 U14761 ( .A1(n13801), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13013), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13036) );
  AOI22_X1 U14762 ( .A1(n13804), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13778), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13035) );
  AOI22_X1 U14763 ( .A1(n11146), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13809), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13034) );
  AOI22_X1 U14764 ( .A1(n13810), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13033) );
  NAND4_X1 U14765 ( .A1(n13036), .A2(n13035), .A3(n13034), .A4(n13033), .ZN(
        n13042) );
  AOI22_X1 U14766 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13563), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13040) );
  AOI22_X1 U14767 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12899), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13039) );
  AOI22_X1 U14768 ( .A1(n13779), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13433), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13038) );
  AOI22_X1 U14769 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13037) );
  NAND4_X1 U14770 ( .A1(n13040), .A2(n13039), .A3(n13038), .A4(n13037), .ZN(
        n13041) );
  XNOR2_X1 U14771 ( .A(n13052), .B(n13219), .ZN(n13043) );
  NAND2_X1 U14772 ( .A1(n13043), .A2(n13066), .ZN(n13044) );
  INV_X1 U14773 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13051) );
  NAND2_X1 U14774 ( .A1(n12961), .A2(n13219), .ZN(n13048) );
  OAI211_X1 U14775 ( .C1(n13052), .C2(n16021), .A(n13048), .B(
        P1_STATE2_REG_0__SCAN_IN), .ZN(n13049) );
  INV_X1 U14776 ( .A(n13049), .ZN(n13050) );
  AOI21_X1 U14777 ( .B1(n13052), .B2(n21878), .A(n13101), .ZN(n13053) );
  OAI21_X2 U14778 ( .B1(n13337), .B2(n13215), .A(n13053), .ZN(n14894) );
  NAND2_X1 U14779 ( .A1(n15070), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15071) );
  INV_X1 U14780 ( .A(n13054), .ZN(n13055) );
  OR2_X1 U14781 ( .A1(n13055), .A2(n14893), .ZN(n13056) );
  NAND2_X1 U14782 ( .A1(n15071), .A2(n13056), .ZN(n13104) );
  INV_X1 U14783 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n16433) );
  XNOR2_X1 U14784 ( .A(n13104), .B(n16433), .ZN(n15210) );
  INV_X1 U14785 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13060) );
  NAND3_X1 U14786 ( .A1(n15146), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n13057), 
        .ZN(n13059) );
  INV_X1 U14787 ( .A(n13219), .ZN(n13204) );
  NAND2_X1 U14788 ( .A1(n13066), .A2(n13204), .ZN(n13058) );
  OAI211_X1 U14789 ( .C1(n13302), .C2(n13060), .A(n13059), .B(n13058), .ZN(
        n13061) );
  OR2_X2 U14790 ( .A1(n13062), .A2(n13061), .ZN(n13068) );
  NAND2_X1 U14791 ( .A1(n13062), .A2(n13061), .ZN(n13063) );
  NAND2_X2 U14792 ( .A1(n13068), .A2(n13063), .ZN(n13331) );
  NAND2_X1 U14793 ( .A1(n13065), .A2(n13064), .ZN(n13067) );
  NAND2_X1 U14794 ( .A1(n13066), .A2(n13219), .ZN(n13216) );
  OAI21_X2 U14795 ( .B1(n13331), .B2(n13332), .A(n13068), .ZN(n13097) );
  INV_X1 U14796 ( .A(n13097), .ZN(n13095) );
  AND2_X1 U14797 ( .A1(n13070), .A2(n16595), .ZN(n13071) );
  NAND2_X1 U14798 ( .A1(n13073), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13078) );
  INV_X1 U14799 ( .A(n13075), .ZN(n13074) );
  NAND2_X1 U14800 ( .A1(n13074), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n15095) );
  NAND2_X1 U14801 ( .A1(n13075), .A2(n17795), .ZN(n13076) );
  INV_X1 U14802 ( .A(n13838), .ZN(n13109) );
  AOI22_X1 U14803 ( .A1(n15547), .A2(n13109), .B1(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n13108), .ZN(n13077) );
  AOI22_X1 U14804 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11172), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13087) );
  AOI22_X1 U14805 ( .A1(n13801), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13086) );
  AOI22_X1 U14806 ( .A1(n13013), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13779), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13085) );
  AOI22_X1 U14807 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13778), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13084) );
  NAND4_X1 U14808 ( .A1(n13087), .A2(n13086), .A3(n13085), .A4(n13084), .ZN(
        n13093) );
  AOI22_X1 U14809 ( .A1(n13563), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13091) );
  AOI22_X1 U14810 ( .A1(n13809), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13090) );
  AOI22_X1 U14811 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13433), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13089) );
  AOI22_X1 U14812 ( .A1(n13804), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13088) );
  NAND4_X1 U14813 ( .A1(n13091), .A2(n13090), .A3(n13089), .A4(n13088), .ZN(
        n13092) );
  AOI22_X1 U14814 ( .A1(n13270), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13286), .B2(n13100), .ZN(n13094) );
  NAND2_X2 U14815 ( .A1(n13095), .A2(n13096), .ZN(n13126) );
  NAND2_X1 U14816 ( .A1(n13097), .A2(n13098), .ZN(n13099) );
  NAND2_X2 U14817 ( .A1(n13126), .A2(n13099), .ZN(n14999) );
  INV_X1 U14818 ( .A(n13100), .ZN(n13128) );
  XNOR2_X1 U14819 ( .A(n13129), .B(n13128), .ZN(n13102) );
  AOI21_X1 U14820 ( .B1(n13102), .B2(n21878), .A(n13101), .ZN(n13103) );
  NAND2_X1 U14821 ( .A1(n13104), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13105) );
  INV_X1 U14822 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21937) );
  INV_X1 U14823 ( .A(n13126), .ZN(n13124) );
  NAND2_X1 U14824 ( .A1(n13073), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13111) );
  INV_X1 U14825 ( .A(n15095), .ZN(n13106) );
  NAND2_X1 U14826 ( .A1(n13106), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n22670) );
  NAND2_X1 U14827 ( .A1(n15095), .A2(n15570), .ZN(n13107) );
  AOI22_X1 U14828 ( .A1(n15785), .A2(n13109), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n13108), .ZN(n13110) );
  XNOR2_X2 U14829 ( .A(n14885), .B(n15092), .ZN(n16621) );
  AOI22_X1 U14830 ( .A1(n13563), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11172), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13115) );
  AOI22_X1 U14831 ( .A1(n13801), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13114) );
  AOI22_X1 U14832 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13013), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13113) );
  AOI22_X1 U14833 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13112) );
  NAND4_X1 U14834 ( .A1(n13115), .A2(n13114), .A3(n13113), .A4(n13112), .ZN(
        n13121) );
  AOI22_X1 U14835 ( .A1(n13804), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13778), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13119) );
  AOI22_X1 U14836 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13118) );
  AOI22_X1 U14837 ( .A1(n13779), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13433), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13117) );
  AOI22_X1 U14838 ( .A1(n13809), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13116) );
  NAND4_X1 U14839 ( .A1(n13119), .A2(n13118), .A3(n13117), .A4(n13116), .ZN(
        n13120) );
  AOI22_X1 U14840 ( .A1(n13270), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13286), .B2(n13148), .ZN(n13122) );
  INV_X1 U14841 ( .A(n15031), .ZN(n13125) );
  NAND2_X1 U14842 ( .A1(n13126), .A2(n13125), .ZN(n13127) );
  NAND2_X1 U14843 ( .A1(n13156), .A2(n13127), .ZN(n15030) );
  OR2_X1 U14844 ( .A1(n15030), .A2(n13215), .ZN(n13133) );
  NAND2_X1 U14845 ( .A1(n13129), .A2(n13128), .ZN(n13149) );
  INV_X1 U14846 ( .A(n13148), .ZN(n13130) );
  XNOR2_X1 U14847 ( .A(n13149), .B(n13130), .ZN(n13131) );
  NAND2_X1 U14848 ( .A1(n13131), .A2(n21878), .ZN(n13132) );
  NAND2_X1 U14849 ( .A1(n13133), .A2(n13132), .ZN(n15217) );
  NAND2_X1 U14850 ( .A1(n15218), .A2(n15217), .ZN(n15216) );
  NAND2_X1 U14851 ( .A1(n13134), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13135) );
  NAND2_X1 U14852 ( .A1(n15216), .A2(n13135), .ZN(n20533) );
  INV_X1 U14853 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13147) );
  AOI22_X1 U14854 ( .A1(n13563), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11172), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13140) );
  AOI22_X1 U14855 ( .A1(n13801), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13139) );
  AOI22_X1 U14856 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13013), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13138) );
  AOI22_X1 U14857 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13137) );
  NAND4_X1 U14858 ( .A1(n13140), .A2(n13139), .A3(n13138), .A4(n13137), .ZN(
        n13146) );
  AOI22_X1 U14859 ( .A1(n13804), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13778), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13144) );
  AOI22_X1 U14860 ( .A1(n11177), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13143) );
  AOI22_X1 U14861 ( .A1(n13779), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13433), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13142) );
  AOI22_X1 U14862 ( .A1(n13697), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13141) );
  NAND4_X1 U14863 ( .A1(n13144), .A2(n13143), .A3(n13142), .A4(n13141), .ZN(
        n13145) );
  OAI22_X1 U14864 ( .A1(n13302), .A2(n13147), .B1(n13283), .B2(n13171), .ZN(
        n13157) );
  XNOR2_X1 U14865 ( .A(n13156), .B(n13157), .ZN(n13357) );
  NAND2_X1 U14866 ( .A1(n13357), .A2(n13010), .ZN(n13153) );
  NAND2_X1 U14867 ( .A1(n13149), .A2(n13148), .ZN(n13172) );
  XNOR2_X1 U14868 ( .A(n13172), .B(n13150), .ZN(n13151) );
  NAND2_X1 U14869 ( .A1(n13151), .A2(n21878), .ZN(n13152) );
  NAND2_X1 U14870 ( .A1(n13153), .A2(n13152), .ZN(n13154) );
  INV_X1 U14871 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n21930) );
  XNOR2_X1 U14872 ( .A(n13154), .B(n21930), .ZN(n20532) );
  NAND2_X1 U14873 ( .A1(n20533), .A2(n20532), .ZN(n20531) );
  NAND2_X1 U14874 ( .A1(n13154), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13155) );
  NAND2_X1 U14875 ( .A1(n20531), .A2(n13155), .ZN(n20540) );
  INV_X1 U14876 ( .A(n13156), .ZN(n13158) );
  NAND2_X1 U14877 ( .A1(n13158), .A2(n13157), .ZN(n13178) );
  INV_X1 U14878 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13170) );
  AOI22_X1 U14879 ( .A1(n13801), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13563), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13162) );
  AOI22_X1 U14880 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13161) );
  AOI22_X1 U14881 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13013), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13160) );
  AOI22_X1 U14882 ( .A1(n13779), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13433), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13159) );
  NAND4_X1 U14883 ( .A1(n13162), .A2(n13161), .A3(n13160), .A4(n13159), .ZN(
        n13168) );
  AOI22_X1 U14884 ( .A1(n11146), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13778), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13166) );
  AOI22_X1 U14885 ( .A1(n13800), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13165) );
  AOI22_X1 U14886 ( .A1(n13810), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13164) );
  AOI22_X1 U14887 ( .A1(n13697), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13163) );
  NAND4_X1 U14888 ( .A1(n13166), .A2(n13165), .A3(n13164), .A4(n13163), .ZN(
        n13167) );
  INV_X1 U14889 ( .A(n13197), .ZN(n13169) );
  XNOR2_X1 U14890 ( .A(n13178), .B(n13179), .ZN(n13358) );
  NAND2_X1 U14891 ( .A1(n13358), .A2(n13010), .ZN(n13175) );
  OR2_X1 U14892 ( .A1(n13172), .A2(n13171), .ZN(n13196) );
  XNOR2_X1 U14893 ( .A(n13196), .B(n13197), .ZN(n13173) );
  NAND2_X1 U14894 ( .A1(n13173), .A2(n21878), .ZN(n13174) );
  NAND2_X1 U14895 ( .A1(n13175), .A2(n13174), .ZN(n13176) );
  INV_X1 U14896 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21939) );
  XNOR2_X1 U14897 ( .A(n13176), .B(n21939), .ZN(n20539) );
  NAND2_X1 U14898 ( .A1(n20540), .A2(n20539), .ZN(n20538) );
  NAND2_X1 U14899 ( .A1(n13176), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13177) );
  NAND2_X1 U14900 ( .A1(n20538), .A2(n13177), .ZN(n20546) );
  INV_X1 U14901 ( .A(n13178), .ZN(n13180) );
  NAND2_X1 U14902 ( .A1(n13180), .A2(n13179), .ZN(n13195) );
  INV_X1 U14903 ( .A(n13195), .ZN(n13193) );
  AOI22_X1 U14904 ( .A1(n13563), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13800), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13184) );
  AOI22_X1 U14905 ( .A1(n13801), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13183) );
  AOI22_X1 U14906 ( .A1(n13731), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13013), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13182) );
  AOI22_X1 U14907 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13181) );
  NAND4_X1 U14908 ( .A1(n13184), .A2(n13183), .A3(n13182), .A4(n13181), .ZN(
        n13191) );
  AOI22_X1 U14909 ( .A1(n13804), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13778), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13189) );
  AOI22_X1 U14910 ( .A1(n11146), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13188) );
  AOI22_X1 U14911 ( .A1(n13779), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13433), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13187) );
  AOI22_X1 U14912 ( .A1(n13697), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13186) );
  NAND4_X1 U14913 ( .A1(n13189), .A2(n13188), .A3(n13187), .A4(n13186), .ZN(
        n13190) );
  AOI22_X1 U14914 ( .A1(n13270), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13286), .B2(n13208), .ZN(n13194) );
  NAND2_X2 U14915 ( .A1(n13193), .A2(n13192), .ZN(n13218) );
  NAND2_X1 U14916 ( .A1(n13195), .A2(n13194), .ZN(n13372) );
  NAND3_X1 U14917 ( .A1(n13218), .A2(n13010), .A3(n13372), .ZN(n13201) );
  INV_X1 U14918 ( .A(n13196), .ZN(n13198) );
  NAND2_X1 U14919 ( .A1(n13198), .A2(n13197), .ZN(n13207) );
  XNOR2_X1 U14920 ( .A(n13207), .B(n13208), .ZN(n13199) );
  NAND2_X1 U14921 ( .A1(n13199), .A2(n21878), .ZN(n13200) );
  NAND2_X1 U14922 ( .A1(n13201), .A2(n13200), .ZN(n13202) );
  XNOR2_X1 U14923 ( .A(n13202), .B(n21949), .ZN(n20545) );
  NAND2_X1 U14924 ( .A1(n20546), .A2(n20545), .ZN(n20544) );
  NAND2_X1 U14925 ( .A1(n13202), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13203) );
  NAND2_X1 U14926 ( .A1(n20544), .A2(n13203), .ZN(n20552) );
  INV_X1 U14927 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13205) );
  OAI22_X1 U14928 ( .A1(n13302), .A2(n13205), .B1(n13283), .B2(n13204), .ZN(
        n13206) );
  NAND2_X1 U14929 ( .A1(n13318), .A2(n13010), .ZN(n13212) );
  INV_X1 U14930 ( .A(n13207), .ZN(n13209) );
  NAND2_X1 U14931 ( .A1(n13209), .A2(n13208), .ZN(n13221) );
  XNOR2_X1 U14932 ( .A(n13221), .B(n13219), .ZN(n13210) );
  NAND2_X1 U14933 ( .A1(n13210), .A2(n21878), .ZN(n13211) );
  NAND2_X1 U14934 ( .A1(n13212), .A2(n13211), .ZN(n13213) );
  INV_X1 U14935 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21965) );
  XNOR2_X1 U14936 ( .A(n13213), .B(n21965), .ZN(n20551) );
  NAND2_X1 U14937 ( .A1(n20552), .A2(n20551), .ZN(n20550) );
  NAND2_X1 U14938 ( .A1(n13213), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13214) );
  NOR2_X1 U14939 ( .A1(n13216), .A2(n13215), .ZN(n13217) );
  NAND2_X4 U14940 ( .A1(n13218), .A2(n13217), .ZN(n16412) );
  NAND2_X1 U14941 ( .A1(n21878), .A2(n13219), .ZN(n13220) );
  OR2_X1 U14942 ( .A1(n13221), .A2(n13220), .ZN(n13222) );
  NAND2_X1 U14943 ( .A1(n16412), .A2(n13222), .ZN(n13223) );
  INV_X1 U14944 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21966) );
  XNOR2_X1 U14945 ( .A(n13223), .B(n21966), .ZN(n15826) );
  NAND2_X1 U14946 ( .A1(n13223), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13224) );
  NAND2_X1 U14947 ( .A1(n15825), .A2(n13224), .ZN(n15915) );
  XNOR2_X1 U14948 ( .A(n11452), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15914) );
  NAND2_X2 U14949 ( .A1(n15915), .A2(n15914), .ZN(n16411) );
  INV_X2 U14950 ( .A(n16412), .ZN(n16352) );
  NAND2_X1 U14951 ( .A1(n16352), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13225) );
  NAND2_X1 U14952 ( .A1(n16352), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16388) );
  INV_X1 U14953 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n21901) );
  NAND2_X1 U14954 ( .A1(n16412), .A2(n21901), .ZN(n13226) );
  NAND2_X1 U14955 ( .A1(n16388), .A2(n13226), .ZN(n16403) );
  INV_X1 U14956 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16401) );
  NAND2_X1 U14957 ( .A1(n16412), .A2(n16401), .ZN(n20560) );
  NAND2_X1 U14958 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n13227) );
  NAND2_X1 U14959 ( .A1(n16412), .A2(n13227), .ZN(n16400) );
  NAND2_X1 U14960 ( .A1(n20560), .A2(n16400), .ZN(n13228) );
  NOR2_X1 U14961 ( .A1(n16403), .A2(n13228), .ZN(n16386) );
  INV_X1 U14962 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n13959) );
  NAND2_X1 U14963 ( .A1(n16412), .A2(n13959), .ZN(n13229) );
  NAND2_X1 U14964 ( .A1(n16386), .A2(n13229), .ZN(n16376) );
  NAND2_X1 U14965 ( .A1(n21901), .A2(n13959), .ZN(n13230) );
  NAND2_X1 U14966 ( .A1(n20578), .A2(n13230), .ZN(n13233) );
  NAND2_X1 U14967 ( .A1(n16376), .A2(n13233), .ZN(n20572) );
  AND2_X1 U14968 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n22028) );
  AND2_X1 U14969 ( .A1(n22028), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n22023) );
  INV_X1 U14970 ( .A(n22023), .ZN(n13231) );
  NAND2_X1 U14971 ( .A1(n16412), .A2(n13231), .ZN(n13232) );
  INV_X1 U14972 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n21993) );
  INV_X1 U14973 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16414) );
  NAND2_X1 U14974 ( .A1(n20578), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n20559) );
  NAND2_X1 U14975 ( .A1(n16398), .A2(n20559), .ZN(n16387) );
  INV_X1 U14976 ( .A(n13233), .ZN(n13234) );
  INV_X1 U14977 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n22015) );
  NOR2_X1 U14978 ( .A1(n16412), .A2(n22015), .ZN(n13235) );
  OAI21_X1 U14979 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n20578), .ZN(n13236) );
  NAND2_X1 U14980 ( .A1(n20574), .A2(n13236), .ZN(n13237) );
  AND2_X1 U14981 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16546) );
  NAND2_X1 U14982 ( .A1(n16546), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16547) );
  INV_X1 U14983 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n22022) );
  INV_X1 U14984 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16432) );
  NOR2_X2 U14985 ( .A1(n16343), .A2(n16432), .ZN(n16324) );
  NOR4_X1 U14986 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n13239) );
  AND2_X1 U14987 ( .A1(n13238), .A2(n13239), .ZN(n16345) );
  NOR2_X1 U14988 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16513) );
  NAND3_X1 U14989 ( .A1(n13242), .A2(n16513), .A3(n13990), .ZN(n13241) );
  NAND2_X1 U14990 ( .A1(n13241), .A2(n16352), .ZN(n16308) );
  AND2_X1 U14991 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16504) );
  NAND2_X1 U14992 ( .A1(n16504), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16493) );
  INV_X1 U14993 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16494) );
  INV_X1 U14994 ( .A(n13245), .ZN(n13243) );
  INV_X1 U14995 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16291) );
  INV_X1 U14996 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13244) );
  NAND2_X1 U14997 ( .A1(n16291), .A2(n13244), .ZN(n16476) );
  AND2_X1 U14998 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16458) );
  AOI21_X1 U14999 ( .B1(n13245), .B2(n16458), .A(n16352), .ZN(n16269) );
  INV_X1 U15000 ( .A(n13252), .ZN(n13249) );
  INV_X1 U15001 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16449) );
  XNOR2_X1 U15002 ( .A(n11452), .B(n16449), .ZN(n13251) );
  INV_X1 U15003 ( .A(n13251), .ZN(n13248) );
  INV_X1 U15004 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16448) );
  AND2_X1 U15005 ( .A1(n16412), .A2(n16448), .ZN(n13254) );
  INV_X1 U15006 ( .A(n13254), .ZN(n13247) );
  NAND2_X1 U15007 ( .A1(n13249), .A2(n11630), .ZN(n13258) );
  NAND2_X1 U15008 ( .A1(n16448), .A2(n13246), .ZN(n13250) );
  NAND2_X1 U15009 ( .A1(n16352), .A2(n13250), .ZN(n13253) );
  NAND3_X1 U15010 ( .A1(n13252), .A2(n13251), .A3(n13253), .ZN(n13257) );
  INV_X1 U15011 ( .A(n13253), .ZN(n13255) );
  OAI21_X1 U15012 ( .B1(n13255), .B2(n13254), .A(n16449), .ZN(n13256) );
  NAND3_X1 U15013 ( .A1(n13258), .A2(n13257), .A3(n13256), .ZN(n16456) );
  OR2_X1 U15014 ( .A1(n12971), .A2(n12955), .ZN(n13259) );
  AND2_X1 U15015 ( .A1(n11248), .A2(n13259), .ZN(n14832) );
  NAND2_X1 U15016 ( .A1(n16592), .A2(n15146), .ZN(n13260) );
  NAND3_X1 U15017 ( .A1(n14832), .A2(n14858), .A3(n13260), .ZN(n14849) );
  NOR2_X1 U15018 ( .A1(n14849), .A2(n14833), .ZN(n17804) );
  XNOR2_X1 U15019 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n13273) );
  NAND2_X1 U15020 ( .A1(n13277), .A2(n13273), .ZN(n13262) );
  NAND2_X1 U15021 ( .A1(n22374), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13261) );
  NAND2_X1 U15022 ( .A1(n13262), .A2(n13261), .ZN(n13272) );
  XNOR2_X1 U15023 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n13271) );
  NAND2_X1 U15024 ( .A1(n13272), .A2(n13271), .ZN(n13264) );
  NAND2_X1 U15025 ( .A1(n17795), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13263) );
  NAND2_X1 U15026 ( .A1(n13264), .A2(n13263), .ZN(n13298) );
  XNOR2_X1 U15027 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n13296) );
  NAND2_X1 U15028 ( .A1(n13298), .A2(n13296), .ZN(n13266) );
  NAND2_X1 U15029 ( .A1(n15570), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13265) );
  NAND2_X1 U15030 ( .A1(n13266), .A2(n13265), .ZN(n13295) );
  NAND2_X1 U15031 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n17802), .ZN(
        n13294) );
  INV_X1 U15032 ( .A(n14691), .ZN(n13269) );
  AOI21_X1 U15033 ( .B1(n15379), .B2(n13009), .A(n12946), .ZN(n13293) );
  XOR2_X1 U15034 ( .A(n13272), .B(n13271), .Z(n14688) );
  NAND2_X1 U15035 ( .A1(n13286), .A2(n14688), .ZN(n13292) );
  INV_X1 U15036 ( .A(n13273), .ZN(n13274) );
  XNOR2_X1 U15037 ( .A(n13274), .B(n13277), .ZN(n14687) );
  INV_X1 U15038 ( .A(n14687), .ZN(n13275) );
  NAND2_X1 U15039 ( .A1(n15379), .A2(n13275), .ZN(n13282) );
  NAND2_X1 U15040 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16022), .ZN(n13284) );
  OAI21_X1 U15041 ( .B1(n13302), .B2(n14687), .A(n13284), .ZN(n13288) );
  AND2_X1 U15042 ( .A1(n14866), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n13276) );
  NOR2_X1 U15043 ( .A1(n13277), .A2(n13276), .ZN(n13279) );
  INV_X1 U15044 ( .A(n13279), .ZN(n13278) );
  OAI21_X1 U15045 ( .B1(n13283), .B2(n13278), .A(n13303), .ZN(n13281) );
  OAI211_X1 U15046 ( .C1(n15146), .C2(n14833), .A(n13293), .B(n13279), .ZN(
        n13280) );
  OAI211_X1 U15047 ( .C1(n13282), .C2(n13288), .A(n13281), .B(n13280), .ZN(
        n13291) );
  NOR2_X1 U15048 ( .A1(n15379), .A2(n13283), .ZN(n13289) );
  INV_X1 U15049 ( .A(n13284), .ZN(n13285) );
  NOR3_X1 U15050 ( .A1(n13286), .A2(n15379), .A3(n13285), .ZN(n13287) );
  OAI22_X1 U15051 ( .A1(n13289), .A2(n13288), .B1(n13287), .B2(n14687), .ZN(
        n13290) );
  OAI211_X1 U15052 ( .C1(n13293), .C2(n13292), .A(n13291), .B(n13290), .ZN(
        n13306) );
  AND2_X1 U15053 ( .A1(n13293), .A2(n13292), .ZN(n13301) );
  OR2_X1 U15054 ( .A1(n13295), .A2(n13294), .ZN(n13300) );
  INV_X1 U15055 ( .A(n13296), .ZN(n13297) );
  XNOR2_X1 U15056 ( .A(n13298), .B(n13297), .ZN(n13299) );
  NAND2_X1 U15057 ( .A1(n13300), .A2(n13299), .ZN(n14690) );
  OAI22_X1 U15058 ( .A1(n14688), .A2(n13302), .B1(n13301), .B2(n14690), .ZN(
        n13305) );
  INV_X1 U15059 ( .A(n13303), .ZN(n13304) );
  AOI222_X1 U15060 ( .A1(n13306), .A2(n13305), .B1(n22274), .B2(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C1(n14690), .C2(n13304), .ZN(
        n13307) );
  INV_X1 U15061 ( .A(n13307), .ZN(n13308) );
  INV_X1 U15062 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n13316) );
  NAND2_X1 U15063 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n13313) );
  NOR2_X1 U15064 ( .A1(n13368), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13314) );
  OR2_X1 U15065 ( .A1(n13392), .A2(n13314), .ZN(n22126) );
  AOI22_X1 U15066 ( .A1(n22126), .A2(n13791), .B1(n13827), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n13315) );
  OAI21_X1 U15067 ( .B1(n13822), .B2(n13316), .A(n13315), .ZN(n13317) );
  AOI21_X1 U15068 ( .B1(n13318), .B2(n13503), .A(n13317), .ZN(n15648) );
  INV_X1 U15069 ( .A(n15648), .ZN(n13376) );
  INV_X1 U15070 ( .A(n15030), .ZN(n13319) );
  INV_X1 U15071 ( .A(n15992), .ZN(n14937) );
  AND2_X1 U15072 ( .A1(n14937), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13342) );
  INV_X1 U15073 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n13322) );
  OAI21_X1 U15074 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n13320), .A(
        n13359), .ZN(n15395) );
  AOI22_X1 U15075 ( .A1(n13791), .A2(n15395), .B1(n13827), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13321) );
  OAI21_X1 U15076 ( .B1(n13822), .B2(n13322), .A(n13321), .ZN(n13323) );
  AOI21_X1 U15077 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13342), .A(
        n13323), .ZN(n13324) );
  NAND2_X1 U15078 ( .A1(n13325), .A2(n13324), .ZN(n15208) );
  INV_X1 U15079 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n13327) );
  XNOR2_X1 U15080 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15286) );
  AOI21_X1 U15081 ( .B1(n13791), .B2(n15286), .A(n13827), .ZN(n13326) );
  OAI21_X1 U15082 ( .B1(n13822), .B2(n13327), .A(n13326), .ZN(n13328) );
  AOI21_X1 U15083 ( .B1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n13342), .A(
        n13328), .ZN(n13329) );
  NAND2_X1 U15084 ( .A1(n13827), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13350) );
  NAND2_X1 U15085 ( .A1(n13330), .A2(n13350), .ZN(n15050) );
  INV_X1 U15086 ( .A(n15050), .ZN(n13349) );
  XNOR2_X2 U15087 ( .A(n13331), .B(n13332), .ZN(n14966) );
  NAND2_X1 U15088 ( .A1(n14966), .A2(n13503), .ZN(n13336) );
  INV_X1 U15089 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n13333) );
  INV_X1 U15090 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n22071) );
  OAI22_X1 U15091 ( .A1(n13822), .A2(n13333), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n22071), .ZN(n13334) );
  AOI21_X1 U15092 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n13342), .A(
        n13334), .ZN(n13335) );
  NAND2_X1 U15093 ( .A1(n13336), .A2(n13335), .ZN(n15002) );
  NAND2_X1 U15095 ( .A1(n13338), .A2(n16023), .ZN(n13339) );
  NAND2_X1 U15096 ( .A1(n13339), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14927) );
  INV_X1 U15097 ( .A(n13342), .ZN(n13353) );
  NAND2_X1 U15098 ( .A1(n15575), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13344) );
  NAND2_X1 U15099 ( .A1(n13828), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n13343) );
  OAI211_X1 U15100 ( .C1(n13353), .C2(n14866), .A(n13344), .B(n13343), .ZN(
        n13345) );
  AOI21_X1 U15101 ( .B1(n13341), .B2(n13503), .A(n13345), .ZN(n13346) );
  OR2_X1 U15102 ( .A1(n14927), .A2(n13346), .ZN(n14928) );
  INV_X1 U15103 ( .A(n13346), .ZN(n14929) );
  OR2_X1 U15104 ( .A1(n14929), .A2(n13668), .ZN(n13347) );
  NAND2_X1 U15105 ( .A1(n14928), .A2(n13347), .ZN(n15001) );
  NAND2_X1 U15106 ( .A1(n15002), .A2(n15001), .ZN(n15049) );
  INV_X1 U15107 ( .A(n15049), .ZN(n13348) );
  NAND2_X1 U15108 ( .A1(n13349), .A2(n13348), .ZN(n15047) );
  NAND2_X1 U15109 ( .A1(n15208), .A2(n15207), .ZN(n15330) );
  NAND2_X1 U15110 ( .A1(n15575), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13352) );
  NAND2_X1 U15111 ( .A1(n13828), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n13351) );
  OAI211_X1 U15112 ( .C1(n13353), .C2(n17802), .A(n13352), .B(n13351), .ZN(
        n13355) );
  INV_X1 U15113 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n13354) );
  XNOR2_X1 U15114 ( .A(n13354), .B(n13359), .ZN(n22090) );
  MUX2_X1 U15115 ( .A(n13355), .B(n22090), .S(n13791), .Z(n13356) );
  AOI21_X1 U15116 ( .B1(n13357), .B2(n13503), .A(n13356), .ZN(n15329) );
  NAND2_X1 U15117 ( .A1(n13358), .A2(n13503), .ZN(n13365) );
  INV_X1 U15118 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n15426) );
  INV_X1 U15119 ( .A(n13359), .ZN(n13360) );
  AOI21_X1 U15120 ( .B1(n13360), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n13361) );
  OR2_X1 U15121 ( .A1(n13361), .A2(n13366), .ZN(n22103) );
  AOI22_X1 U15122 ( .A1(n22103), .A2(n13791), .B1(n13827), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n13362) );
  OAI21_X1 U15123 ( .B1(n13822), .B2(n15426), .A(n13362), .ZN(n13363) );
  INV_X1 U15124 ( .A(n13363), .ZN(n13364) );
  NAND2_X1 U15125 ( .A1(n13365), .A2(n13364), .ZN(n15423) );
  NAND2_X1 U15126 ( .A1(n15328), .A2(n15423), .ZN(n15422) );
  INV_X1 U15127 ( .A(n15422), .ZN(n13374) );
  INV_X1 U15128 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n13370) );
  NOR2_X1 U15129 ( .A1(n13366), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13367) );
  OR2_X1 U15130 ( .A1(n13368), .A2(n13367), .ZN(n22114) );
  AOI22_X1 U15131 ( .A1(n22114), .A2(n13791), .B1(n13827), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n13369) );
  OAI21_X1 U15132 ( .B1(n13822), .B2(n13370), .A(n13369), .ZN(n13371) );
  INV_X1 U15133 ( .A(n15557), .ZN(n13373) );
  NAND2_X1 U15134 ( .A1(n13374), .A2(n13373), .ZN(n15556) );
  AOI22_X1 U15135 ( .A1(n13800), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13013), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13381) );
  AOI22_X1 U15136 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n11179), .B1(
        n13778), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13380) );
  AOI22_X1 U15137 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13379) );
  AOI22_X1 U15138 ( .A1(n13779), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13433), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13378) );
  NAND4_X1 U15139 ( .A1(n13381), .A2(n13380), .A3(n13379), .A4(n13378), .ZN(
        n13387) );
  AOI22_X1 U15140 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n13810), .B1(
        n13563), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13385) );
  AOI22_X1 U15141 ( .A1(n13801), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13784), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13384) );
  AOI22_X1 U15142 ( .A1(n13804), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13383) );
  AOI22_X1 U15143 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n13809), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13382) );
  NAND4_X1 U15144 ( .A1(n13385), .A2(n13384), .A3(n13383), .A4(n13382), .ZN(
        n13386) );
  OAI21_X1 U15145 ( .B1(n13387), .B2(n13386), .A(n13503), .ZN(n13391) );
  NAND2_X1 U15146 ( .A1(n13828), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n13390) );
  XNOR2_X1 U15147 ( .A(n13392), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n22131) );
  NAND2_X1 U15148 ( .A1(n22131), .A2(n13791), .ZN(n13389) );
  NAND2_X1 U15149 ( .A1(n13827), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13388) );
  XOR2_X1 U15150 ( .A(n15869), .B(n13407), .Z(n15920) );
  AOI22_X1 U15151 ( .A1(n13563), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13396) );
  AOI22_X1 U15152 ( .A1(n13801), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13731), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13395) );
  AOI22_X1 U15153 ( .A1(n13779), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13778), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13394) );
  AOI22_X1 U15154 ( .A1(n13697), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13393) );
  NAND4_X1 U15155 ( .A1(n13396), .A2(n13395), .A3(n13394), .A4(n13393), .ZN(
        n13402) );
  AOI22_X1 U15156 ( .A1(n13800), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13013), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13400) );
  AOI22_X1 U15157 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13399) );
  AOI22_X1 U15158 ( .A1(n13804), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13433), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13398) );
  AOI22_X1 U15159 ( .A1(n11146), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13397) );
  NAND4_X1 U15160 ( .A1(n13400), .A2(n13399), .A3(n13398), .A4(n13397), .ZN(
        n13401) );
  NOR2_X1 U15161 ( .A1(n13402), .A2(n13401), .ZN(n13403) );
  OAI22_X1 U15162 ( .A1(n13471), .A2(n13403), .B1(n13539), .B2(n15869), .ZN(
        n13405) );
  INV_X1 U15163 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n15902) );
  NOR2_X1 U15164 ( .A1(n13822), .A2(n15902), .ZN(n13404) );
  NOR2_X1 U15165 ( .A1(n13405), .A2(n13404), .ZN(n13406) );
  OAI21_X1 U15166 ( .B1(n15920), .B2(n13668), .A(n13406), .ZN(n15861) );
  XNOR2_X1 U15167 ( .A(n13423), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16423) );
  NAND2_X1 U15168 ( .A1(n16423), .A2(n13791), .ZN(n13422) );
  INV_X1 U15169 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n15904) );
  INV_X1 U15170 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n15892) );
  OAI22_X1 U15171 ( .A1(n13822), .A2(n15904), .B1(n13539), .B2(n15892), .ZN(
        n13420) );
  AOI22_X1 U15172 ( .A1(n13731), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13411) );
  AOI22_X1 U15173 ( .A1(n13810), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13013), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13410) );
  AOI22_X1 U15174 ( .A1(n13800), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13409) );
  AOI22_X1 U15175 ( .A1(n13778), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13408) );
  NAND4_X1 U15176 ( .A1(n13411), .A2(n13410), .A3(n13409), .A4(n13408), .ZN(
        n13417) );
  AOI22_X1 U15177 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13563), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13415) );
  AOI22_X1 U15178 ( .A1(n13779), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13809), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13414) );
  AOI22_X1 U15179 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13413) );
  AOI22_X1 U15180 ( .A1(n13801), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13433), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13412) );
  NAND4_X1 U15181 ( .A1(n13415), .A2(n13414), .A3(n13413), .A4(n13412), .ZN(
        n13416) );
  NOR2_X1 U15182 ( .A1(n13417), .A2(n13416), .ZN(n13418) );
  NOR2_X1 U15183 ( .A1(n13471), .A2(n13418), .ZN(n13419) );
  NOR2_X1 U15184 ( .A1(n13420), .A2(n13419), .ZN(n13421) );
  NAND2_X1 U15185 ( .A1(n13422), .A2(n13421), .ZN(n15885) );
  INV_X1 U15186 ( .A(n15884), .ZN(n13427) );
  OAI21_X1 U15187 ( .B1(n13424), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n13459), .ZN(n22147) );
  INV_X1 U15188 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n15924) );
  INV_X1 U15189 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n22139) );
  OAI22_X1 U15190 ( .A1(n13822), .A2(n15924), .B1(n13539), .B2(n22139), .ZN(
        n13425) );
  AOI21_X1 U15191 ( .B1(n22147), .B2(n13791), .A(n13425), .ZN(n15922) );
  NAND2_X1 U15192 ( .A1(n13427), .A2(n13426), .ZN(n15926) );
  AOI22_X1 U15193 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13431) );
  AOI22_X1 U15194 ( .A1(n13801), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13013), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13430) );
  AOI22_X1 U15195 ( .A1(n13731), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13778), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13429) );
  AOI22_X1 U15196 ( .A1(n13697), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13428) );
  NAND4_X1 U15197 ( .A1(n13431), .A2(n13430), .A3(n13429), .A4(n13428), .ZN(
        n13439) );
  AOI22_X1 U15198 ( .A1(n13804), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13779), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13437) );
  AOI22_X1 U15199 ( .A1(n13563), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13436) );
  AOI22_X1 U15200 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13435) );
  AOI22_X1 U15201 ( .A1(n13800), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13802), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13434) );
  NAND4_X1 U15202 ( .A1(n13437), .A2(n13436), .A3(n13435), .A4(n13434), .ZN(
        n13438) );
  OR2_X1 U15203 ( .A1(n13439), .A2(n13438), .ZN(n13440) );
  NAND2_X1 U15204 ( .A1(n13503), .A2(n13440), .ZN(n15927) );
  NAND2_X1 U15205 ( .A1(n15926), .A2(n13442), .ZN(n13477) );
  XOR2_X1 U15206 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n13478), .Z(
        n16407) );
  AOI22_X1 U15207 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13448) );
  AOI22_X1 U15208 ( .A1(n13801), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13013), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13447) );
  AOI22_X1 U15209 ( .A1(n11146), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13446) );
  AOI22_X1 U15210 ( .A1(n13697), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13445) );
  NAND4_X1 U15211 ( .A1(n13448), .A2(n13447), .A3(n13446), .A4(n13445), .ZN(
        n13454) );
  AOI22_X1 U15212 ( .A1(n13563), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13800), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13452) );
  AOI22_X1 U15213 ( .A1(n13779), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13778), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13451) );
  AOI22_X1 U15214 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13450) );
  AOI22_X1 U15215 ( .A1(n13810), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13802), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13449) );
  NAND4_X1 U15216 ( .A1(n13452), .A2(n13451), .A3(n13450), .A4(n13449), .ZN(
        n13453) );
  NOR2_X1 U15217 ( .A1(n13454), .A2(n13453), .ZN(n13455) );
  INV_X1 U15218 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16404) );
  OAI22_X1 U15219 ( .A1(n13471), .A2(n13455), .B1(n13539), .B2(n16404), .ZN(
        n13457) );
  INV_X1 U15220 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n16266) );
  NOR2_X1 U15221 ( .A1(n13822), .A2(n16266), .ZN(n13456) );
  NOR2_X1 U15222 ( .A1(n13457), .A2(n13456), .ZN(n13458) );
  OAI21_X1 U15223 ( .B1(n16407), .B2(n13668), .A(n13458), .ZN(n16134) );
  XNOR2_X1 U15224 ( .A(n13459), .B(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n22156) );
  OR2_X1 U15225 ( .A1(n22156), .A2(n13668), .ZN(n13475) );
  AOI22_X1 U15226 ( .A1(n13804), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11146), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13463) );
  AOI22_X1 U15227 ( .A1(n13563), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13800), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13462) );
  AOI22_X1 U15228 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13461) );
  AOI22_X1 U15229 ( .A1(n13731), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13802), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13460) );
  NAND4_X1 U15230 ( .A1(n13463), .A2(n13462), .A3(n13461), .A4(n13460), .ZN(
        n13469) );
  AOI22_X1 U15231 ( .A1(n13801), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13467) );
  AOI22_X1 U15232 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13779), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13466) );
  AOI22_X1 U15233 ( .A1(n13697), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13465) );
  AOI22_X1 U15234 ( .A1(n13778), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13464) );
  NAND4_X1 U15235 ( .A1(n13467), .A2(n13466), .A3(n13465), .A4(n13464), .ZN(
        n13468) );
  NOR2_X1 U15236 ( .A1(n13469), .A2(n13468), .ZN(n13470) );
  OAI22_X1 U15237 ( .A1(n13471), .A2(n13470), .B1(n13539), .B2(n13443), .ZN(
        n13473) );
  INV_X1 U15238 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n15932) );
  NOR2_X1 U15239 ( .A1(n13822), .A2(n15932), .ZN(n13472) );
  NOR2_X1 U15240 ( .A1(n13473), .A2(n13472), .ZN(n13474) );
  NAND2_X1 U15241 ( .A1(n13475), .A2(n13474), .ZN(n15929) );
  XNOR2_X1 U15242 ( .A(n13494), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16393) );
  AOI22_X1 U15243 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13800), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13482) );
  AOI22_X1 U15244 ( .A1(n13810), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13013), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13481) );
  AOI22_X1 U15245 ( .A1(n13778), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13480) );
  AOI22_X1 U15246 ( .A1(n13731), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13802), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13479) );
  NAND4_X1 U15247 ( .A1(n13482), .A2(n13481), .A3(n13480), .A4(n13479), .ZN(
        n13488) );
  AOI22_X1 U15248 ( .A1(n13801), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13779), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13486) );
  AOI22_X1 U15249 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13809), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13485) );
  AOI22_X1 U15250 ( .A1(n13563), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13484) );
  AOI22_X1 U15251 ( .A1(n13804), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13483) );
  NAND4_X1 U15252 ( .A1(n13486), .A2(n13485), .A3(n13484), .A4(n13483), .ZN(
        n13487) );
  OAI21_X1 U15253 ( .B1(n13488), .B2(n13487), .A(n13503), .ZN(n13491) );
  NAND2_X1 U15254 ( .A1(n13828), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n13490) );
  NAND2_X1 U15255 ( .A1(n13827), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13489) );
  NAND3_X1 U15256 ( .A1(n13491), .A2(n13490), .A3(n13489), .ZN(n13492) );
  AOI21_X1 U15257 ( .B1(n16393), .B2(n13791), .A(n13492), .ZN(n15936) );
  XOR2_X1 U15258 ( .A(n22161), .B(n13511), .Z(n22164) );
  INV_X1 U15259 ( .A(n22164), .ZN(n13510) );
  AOI22_X1 U15260 ( .A1(n13810), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13779), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13498) );
  AOI22_X1 U15261 ( .A1(n13804), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13778), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13497) );
  AOI22_X1 U15262 ( .A1(n11177), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13496) );
  AOI22_X1 U15263 ( .A1(n13563), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13495) );
  NAND4_X1 U15264 ( .A1(n13498), .A2(n13497), .A3(n13496), .A4(n13495), .ZN(
        n13505) );
  AOI22_X1 U15265 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13800), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13502) );
  AOI22_X1 U15266 ( .A1(n13801), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11168), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13501) );
  AOI22_X1 U15267 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13802), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13500) );
  AOI22_X1 U15268 ( .A1(n13697), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13499) );
  NAND4_X1 U15269 ( .A1(n13502), .A2(n13501), .A3(n13500), .A4(n13499), .ZN(
        n13504) );
  OAI21_X1 U15270 ( .B1(n13505), .B2(n13504), .A(n13503), .ZN(n13508) );
  NAND2_X1 U15271 ( .A1(n13828), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n13507) );
  NAND2_X1 U15272 ( .A1(n13827), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13506) );
  NAND3_X1 U15273 ( .A1(n13508), .A2(n13507), .A3(n13506), .ZN(n13509) );
  AOI21_X1 U15274 ( .B1(n13510), .B2(n13791), .A(n13509), .ZN(n16259) );
  INV_X1 U15275 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n22172) );
  XNOR2_X1 U15276 ( .A(n13528), .B(n22172), .ZN(n22174) );
  INV_X1 U15277 ( .A(n16592), .ZN(n14902) );
  NAND2_X1 U15278 ( .A1(n13794), .A2(n13668), .ZN(n13597) );
  AOI22_X1 U15279 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n13801), .B1(
        n13778), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13517) );
  NAND2_X1 U15280 ( .A1(n13800), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n13513) );
  NAND2_X1 U15281 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n13512) );
  AND3_X1 U15282 ( .A1(n13513), .A2(n13512), .A3(n13668), .ZN(n13516) );
  AOI22_X1 U15283 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n13731), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13515) );
  AOI22_X1 U15284 ( .A1(n13779), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13514) );
  NAND4_X1 U15285 ( .A1(n13517), .A2(n13516), .A3(n13515), .A4(n13514), .ZN(
        n13523) );
  AOI22_X1 U15286 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13013), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13521) );
  AOI22_X1 U15287 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n13804), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13520) );
  AOI22_X1 U15288 ( .A1(n13563), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13809), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13519) );
  AOI22_X1 U15289 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n11176), .B1(
        n13802), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13518) );
  NAND4_X1 U15290 ( .A1(n13521), .A2(n13520), .A3(n13519), .A4(n13518), .ZN(
        n13522) );
  OR2_X1 U15291 ( .A1(n13523), .A2(n13522), .ZN(n13526) );
  INV_X1 U15292 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13524) );
  OAI22_X1 U15293 ( .A1(n13822), .A2(n13524), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n22172), .ZN(n13525) );
  AOI21_X1 U15294 ( .B1(n13597), .B2(n13526), .A(n13525), .ZN(n13527) );
  AOI21_X1 U15295 ( .B1(n22174), .B2(n13791), .A(n13527), .ZN(n16174) );
  XOR2_X1 U15296 ( .A(n13544), .B(n13545), .Z(n20583) );
  INV_X1 U15297 ( .A(n13794), .ZN(n13819) );
  AOI22_X1 U15298 ( .A1(n13801), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13532) );
  AOI22_X1 U15299 ( .A1(n13804), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13809), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13531) );
  AOI22_X1 U15300 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13530) );
  AOI22_X1 U15301 ( .A1(n13013), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13802), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13529) );
  NAND4_X1 U15302 ( .A1(n13532), .A2(n13531), .A3(n13530), .A4(n13529), .ZN(
        n13538) );
  AOI22_X1 U15303 ( .A1(n13563), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13800), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13536) );
  AOI22_X1 U15304 ( .A1(n13731), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13779), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13535) );
  AOI22_X1 U15305 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13534) );
  AOI22_X1 U15306 ( .A1(n13778), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13533) );
  NAND4_X1 U15307 ( .A1(n13536), .A2(n13535), .A3(n13534), .A4(n13533), .ZN(
        n13537) );
  OR2_X1 U15308 ( .A1(n13538), .A2(n13537), .ZN(n13542) );
  INV_X1 U15309 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13540) );
  OAI22_X1 U15310 ( .A1(n13822), .A2(n13540), .B1(n13539), .B2(n13544), .ZN(
        n13541) );
  AOI21_X1 U15311 ( .B1(n13819), .B2(n13542), .A(n13541), .ZN(n13543) );
  OAI21_X1 U15312 ( .B1(n20583), .B2(n13668), .A(n13543), .ZN(n16125) );
  NAND2_X1 U15313 ( .A1(n16123), .A2(n16125), .ZN(n16124) );
  INV_X1 U15314 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n22185) );
  XNOR2_X1 U15315 ( .A(n13579), .B(n22185), .ZN(n16370) );
  NAND2_X1 U15316 ( .A1(n16370), .A2(n13791), .ZN(n13562) );
  AOI22_X1 U15317 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13731), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13549) );
  AOI22_X1 U15318 ( .A1(n13563), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13809), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13548) );
  AOI22_X1 U15319 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13547) );
  AOI22_X1 U15320 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13802), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13546) );
  NAND4_X1 U15321 ( .A1(n13549), .A2(n13548), .A3(n13547), .A4(n13546), .ZN(
        n13557) );
  AOI22_X1 U15322 ( .A1(n13810), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13555) );
  NAND2_X1 U15323 ( .A1(n11146), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n13551) );
  NAND2_X1 U15324 ( .A1(n13800), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n13550) );
  AND3_X1 U15325 ( .A1(n13551), .A2(n13550), .A3(n13668), .ZN(n13554) );
  AOI22_X1 U15326 ( .A1(n13779), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13778), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13553) );
  AOI22_X1 U15327 ( .A1(n13801), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13552) );
  NAND4_X1 U15328 ( .A1(n13555), .A2(n13554), .A3(n13553), .A4(n13552), .ZN(
        n13556) );
  OAI21_X1 U15329 ( .B1(n13557), .B2(n13556), .A(n13597), .ZN(n13560) );
  NAND2_X1 U15330 ( .A1(n13828), .A2(P1_EAX_REG_18__SCAN_IN), .ZN(n13559) );
  NAND2_X1 U15331 ( .A1(n15575), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13558) );
  NAND3_X1 U15332 ( .A1(n13560), .A2(n13559), .A3(n13558), .ZN(n13561) );
  NAND2_X1 U15333 ( .A1(n13562), .A2(n13561), .ZN(n16172) );
  AOI22_X1 U15334 ( .A1(n13563), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13567) );
  AOI22_X1 U15335 ( .A1(n13801), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11168), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13566) );
  AOI22_X1 U15336 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13565) );
  AOI22_X1 U15337 ( .A1(n13804), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13802), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13564) );
  NAND4_X1 U15338 ( .A1(n13567), .A2(n13566), .A3(n13565), .A4(n13564), .ZN(
        n13573) );
  AOI22_X1 U15339 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13800), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13571) );
  AOI22_X1 U15340 ( .A1(n13779), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13778), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13570) );
  AOI22_X1 U15341 ( .A1(n11177), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13569) );
  AOI22_X1 U15342 ( .A1(n13697), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13568) );
  NAND4_X1 U15343 ( .A1(n13571), .A2(n13570), .A3(n13569), .A4(n13568), .ZN(
        n13572) );
  NOR2_X1 U15344 ( .A1(n13573), .A2(n13572), .ZN(n13578) );
  INV_X1 U15345 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13575) );
  NAND2_X1 U15346 ( .A1(n15575), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13574) );
  OAI211_X1 U15347 ( .C1(n13822), .C2(n13575), .A(n13668), .B(n13574), .ZN(
        n13576) );
  INV_X1 U15348 ( .A(n13576), .ZN(n13577) );
  OAI21_X1 U15349 ( .B1(n13794), .B2(n13578), .A(n13577), .ZN(n13586) );
  INV_X1 U15350 ( .A(n13618), .ZN(n13584) );
  INV_X1 U15351 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n13582) );
  INV_X1 U15352 ( .A(n13580), .ZN(n13581) );
  NAND2_X1 U15353 ( .A1(n13582), .A2(n13581), .ZN(n13583) );
  NAND2_X1 U15354 ( .A1(n13584), .A2(n13583), .ZN(n22195) );
  OR2_X1 U15355 ( .A1(n22195), .A2(n13668), .ZN(n13585) );
  NAND2_X1 U15356 ( .A1(n16171), .A2(n16240), .ZN(n16110) );
  AOI22_X1 U15357 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13784), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13590) );
  AOI22_X1 U15358 ( .A1(n13810), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13778), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13589) );
  AOI22_X1 U15359 ( .A1(n13804), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13809), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13588) );
  AOI22_X1 U15360 ( .A1(n13800), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13587) );
  NAND4_X1 U15361 ( .A1(n13590), .A2(n13589), .A3(n13588), .A4(n13587), .ZN(
        n13599) );
  AOI22_X1 U15362 ( .A1(n13801), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13779), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13596) );
  NAND2_X1 U15363 ( .A1(n13563), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n13592) );
  NAND2_X1 U15364 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n13591) );
  AND3_X1 U15365 ( .A1(n13592), .A2(n13668), .A3(n13591), .ZN(n13595) );
  AOI22_X1 U15366 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13594) );
  AOI22_X1 U15367 ( .A1(n11146), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13802), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13593) );
  NAND4_X1 U15368 ( .A1(n13596), .A2(n13595), .A3(n13594), .A4(n13593), .ZN(
        n13598) );
  OAI21_X1 U15369 ( .B1(n13599), .B2(n13598), .A(n13597), .ZN(n13602) );
  NAND2_X1 U15370 ( .A1(n13828), .A2(P1_EAX_REG_20__SCAN_IN), .ZN(n13601) );
  NAND2_X1 U15371 ( .A1(n15575), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13600) );
  NAND3_X1 U15372 ( .A1(n13602), .A2(n13601), .A3(n13600), .ZN(n13604) );
  INV_X1 U15373 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n16365) );
  XNOR2_X1 U15374 ( .A(n13618), .B(n16365), .ZN(n16363) );
  NAND2_X1 U15375 ( .A1(n16363), .A2(n13791), .ZN(n13603) );
  NAND2_X1 U15376 ( .A1(n13604), .A2(n13603), .ZN(n16112) );
  AOI22_X1 U15377 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13563), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13608) );
  AOI22_X1 U15378 ( .A1(n13810), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13731), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13607) );
  AOI22_X1 U15379 ( .A1(n13778), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13802), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13606) );
  AOI22_X1 U15380 ( .A1(n11177), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13605) );
  NAND4_X1 U15381 ( .A1(n13608), .A2(n13607), .A3(n13606), .A4(n13605), .ZN(
        n13614) );
  AOI22_X1 U15382 ( .A1(n13801), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11168), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13612) );
  AOI22_X1 U15383 ( .A1(n13804), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13779), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13611) );
  AOI22_X1 U15384 ( .A1(n13809), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13610) );
  AOI22_X1 U15385 ( .A1(n13800), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13609) );
  NAND4_X1 U15386 ( .A1(n13612), .A2(n13611), .A3(n13610), .A4(n13609), .ZN(
        n13613) );
  NOR2_X1 U15387 ( .A1(n13614), .A2(n13613), .ZN(n13617) );
  OAI21_X1 U15388 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n22286), .A(
        n15575), .ZN(n13616) );
  NAND2_X1 U15389 ( .A1(n13828), .A2(P1_EAX_REG_21__SCAN_IN), .ZN(n13615) );
  OAI211_X1 U15390 ( .C1(n13794), .C2(n13617), .A(n13616), .B(n13615), .ZN(
        n13623) );
  AND2_X1 U15391 ( .A1(n13619), .A2(n22212), .ZN(n13620) );
  OR2_X1 U15392 ( .A1(n13620), .A2(n13664), .ZN(n22219) );
  INV_X1 U15393 ( .A(n22219), .ZN(n13621) );
  NAND2_X1 U15394 ( .A1(n13621), .A2(n13791), .ZN(n13622) );
  NAND2_X1 U15395 ( .A1(n13623), .A2(n13622), .ZN(n16228) );
  AOI22_X1 U15396 ( .A1(n13563), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13800), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13628) );
  AOI22_X1 U15397 ( .A1(n13801), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13627) );
  AOI22_X1 U15398 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11168), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13626) );
  AOI22_X1 U15399 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13625) );
  NAND4_X1 U15400 ( .A1(n13628), .A2(n13627), .A3(n13626), .A4(n13625), .ZN(
        n13634) );
  AOI22_X1 U15401 ( .A1(n13804), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13778), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13632) );
  AOI22_X1 U15402 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13631) );
  AOI22_X1 U15403 ( .A1(n13779), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13802), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13630) );
  AOI22_X1 U15404 ( .A1(n13697), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13629) );
  NAND4_X1 U15405 ( .A1(n13632), .A2(n13631), .A3(n13630), .A4(n13629), .ZN(
        n13633) );
  NOR2_X1 U15406 ( .A1(n13634), .A2(n13633), .ZN(n13637) );
  NAND2_X1 U15407 ( .A1(n13828), .A2(P1_EAX_REG_22__SCAN_IN), .ZN(n13636) );
  OAI21_X1 U15408 ( .B1(n22286), .B2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15575), .ZN(n13635) );
  OAI211_X1 U15409 ( .C1(n13794), .C2(n13637), .A(n13636), .B(n13635), .ZN(
        n13640) );
  INV_X1 U15410 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n13638) );
  XNOR2_X1 U15411 ( .A(n13664), .B(n13638), .ZN(n16347) );
  NAND2_X1 U15412 ( .A1(n16347), .A2(n13791), .ZN(n13639) );
  NAND2_X1 U15413 ( .A1(n13640), .A2(n13639), .ZN(n16164) );
  AOI22_X1 U15414 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n13779), .B1(
        n13809), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13644) );
  AOI22_X1 U15415 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13643) );
  AOI22_X1 U15416 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n11176), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13642) );
  AOI22_X1 U15417 ( .A1(n13563), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13802), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13641) );
  NAND4_X1 U15418 ( .A1(n13644), .A2(n13643), .A3(n13642), .A4(n13641), .ZN(
        n13650) );
  AOI22_X1 U15419 ( .A1(n13810), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13800), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13648) );
  AOI22_X1 U15420 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n13784), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13647) );
  AOI22_X1 U15421 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n13801), .B1(
        n13013), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13646) );
  AOI22_X1 U15422 ( .A1(n13778), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13645) );
  NAND4_X1 U15423 ( .A1(n13648), .A2(n13647), .A3(n13646), .A4(n13645), .ZN(
        n13649) );
  NOR2_X1 U15424 ( .A1(n13650), .A2(n13649), .ZN(n13682) );
  AOI22_X1 U15425 ( .A1(n13013), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13778), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13654) );
  AOI22_X1 U15426 ( .A1(n11177), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13653) );
  AOI22_X1 U15427 ( .A1(n13800), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13652) );
  AOI22_X1 U15428 ( .A1(n13809), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13651) );
  NAND4_X1 U15429 ( .A1(n13654), .A2(n13653), .A3(n13652), .A4(n13651), .ZN(
        n13660) );
  AOI22_X1 U15430 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13563), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13658) );
  AOI22_X1 U15431 ( .A1(n13801), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13657) );
  AOI22_X1 U15432 ( .A1(n13804), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13779), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13656) );
  AOI22_X1 U15433 ( .A1(n13731), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13802), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13655) );
  NAND4_X1 U15434 ( .A1(n13658), .A2(n13657), .A3(n13656), .A4(n13655), .ZN(
        n13659) );
  NOR2_X1 U15435 ( .A1(n13660), .A2(n13659), .ZN(n13681) );
  XNOR2_X1 U15436 ( .A(n13682), .B(n13681), .ZN(n13663) );
  OAI21_X1 U15437 ( .B1(n22286), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n15575), .ZN(n13662) );
  NAND2_X1 U15438 ( .A1(n13828), .A2(P1_EAX_REG_23__SCAN_IN), .ZN(n13661) );
  OAI211_X1 U15439 ( .C1(n13794), .C2(n13663), .A(n13662), .B(n13661), .ZN(
        n13670) );
  NAND2_X1 U15440 ( .A1(n13666), .A2(n13665), .ZN(n13667) );
  NAND2_X1 U15441 ( .A1(n13725), .A2(n13667), .ZN(n22252) );
  OR2_X1 U15442 ( .A1(n22252), .A2(n13668), .ZN(n13669) );
  AOI22_X1 U15443 ( .A1(n13810), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13800), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13674) );
  AOI22_X1 U15444 ( .A1(n13731), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11168), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13673) );
  AOI22_X1 U15445 ( .A1(n11146), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13779), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13672) );
  AOI22_X1 U15446 ( .A1(n13563), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13671) );
  NAND4_X1 U15447 ( .A1(n13674), .A2(n13673), .A3(n13672), .A4(n13671), .ZN(
        n13680) );
  AOI22_X1 U15448 ( .A1(n13801), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13799), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13678) );
  AOI22_X1 U15449 ( .A1(n13804), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13802), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13677) );
  AOI22_X1 U15450 ( .A1(n13809), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13676) );
  AOI22_X1 U15451 ( .A1(n13778), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13675) );
  NAND4_X1 U15452 ( .A1(n13678), .A2(n13677), .A3(n13676), .A4(n13675), .ZN(
        n13679) );
  NOR2_X1 U15453 ( .A1(n13680), .A2(n13679), .ZN(n13711) );
  NOR2_X1 U15454 ( .A1(n13682), .A2(n13681), .ZN(n13721) );
  AOI22_X1 U15455 ( .A1(n13563), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13800), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13686) );
  AOI22_X1 U15456 ( .A1(n13801), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13685) );
  AOI22_X1 U15457 ( .A1(n13731), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13013), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13684) );
  AOI22_X1 U15458 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13683) );
  NAND4_X1 U15459 ( .A1(n13686), .A2(n13685), .A3(n13684), .A4(n13683), .ZN(
        n13692) );
  AOI22_X1 U15460 ( .A1(n13804), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13778), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13690) );
  AOI22_X1 U15461 ( .A1(n11146), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13689) );
  AOI22_X1 U15462 ( .A1(n13779), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13802), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13688) );
  AOI22_X1 U15463 ( .A1(n13809), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13687) );
  NAND4_X1 U15464 ( .A1(n13690), .A2(n13689), .A3(n13688), .A4(n13687), .ZN(
        n13691) );
  OR2_X1 U15465 ( .A1(n13692), .A2(n13691), .ZN(n13720) );
  NAND2_X1 U15466 ( .A1(n13721), .A2(n13720), .ZN(n13710) );
  NOR2_X1 U15467 ( .A1(n13711), .A2(n13710), .ZN(n13730) );
  AOI22_X1 U15468 ( .A1(n13563), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13800), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13696) );
  AOI22_X1 U15469 ( .A1(n13801), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13695) );
  AOI22_X1 U15470 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13013), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13694) );
  AOI22_X1 U15471 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13693) );
  NAND4_X1 U15472 ( .A1(n13696), .A2(n13695), .A3(n13694), .A4(n13693), .ZN(
        n13703) );
  AOI22_X1 U15473 ( .A1(n13804), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13778), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13701) );
  AOI22_X1 U15474 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13700) );
  AOI22_X1 U15475 ( .A1(n13779), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13802), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13699) );
  AOI22_X1 U15476 ( .A1(n13697), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13698) );
  NAND4_X1 U15477 ( .A1(n13701), .A2(n13700), .A3(n13699), .A4(n13698), .ZN(
        n13702) );
  OR2_X1 U15478 ( .A1(n13703), .A2(n13702), .ZN(n13729) );
  XNOR2_X1 U15479 ( .A(n13730), .B(n13729), .ZN(n13706) );
  NAND2_X1 U15480 ( .A1(n13828), .A2(P1_EAX_REG_26__SCAN_IN), .ZN(n13705) );
  OAI21_X1 U15481 ( .B1(n22286), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15575), .ZN(n13704) );
  OAI211_X1 U15482 ( .C1(n13706), .C2(n13794), .A(n13705), .B(n13704), .ZN(
        n13709) );
  INV_X1 U15483 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n13715) );
  XNOR2_X1 U15484 ( .A(n13747), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16088) );
  NAND2_X1 U15485 ( .A1(n16088), .A2(n13791), .ZN(n13708) );
  NAND2_X1 U15486 ( .A1(n13709), .A2(n13708), .ZN(n16086) );
  XNOR2_X1 U15487 ( .A(n13711), .B(n13710), .ZN(n13714) );
  OAI21_X1 U15488 ( .B1(n22286), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n15575), .ZN(n13713) );
  NAND2_X1 U15489 ( .A1(n13828), .A2(P1_EAX_REG_25__SCAN_IN), .ZN(n13712) );
  OAI211_X1 U15490 ( .C1(n13714), .C2(n13794), .A(n13713), .B(n13712), .ZN(
        n13719) );
  NAND2_X1 U15491 ( .A1(n13716), .A2(n13715), .ZN(n13717) );
  AND2_X1 U15492 ( .A1(n13747), .A2(n13717), .ZN(n16100) );
  NAND2_X1 U15493 ( .A1(n16100), .A2(n13791), .ZN(n13718) );
  NAND2_X1 U15494 ( .A1(n13719), .A2(n13718), .ZN(n16097) );
  NOR2_X1 U15495 ( .A1(n16086), .A2(n16097), .ZN(n13728) );
  XNOR2_X1 U15496 ( .A(n13721), .B(n13720), .ZN(n13724) );
  NAND2_X1 U15497 ( .A1(n13828), .A2(P1_EAX_REG_24__SCAN_IN), .ZN(n13723) );
  OAI21_X1 U15498 ( .B1(n22286), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15575), .ZN(n13722) );
  OAI211_X1 U15499 ( .C1(n13724), .C2(n13794), .A(n13723), .B(n13722), .ZN(
        n13727) );
  XNOR2_X1 U15500 ( .A(n13725), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n22261) );
  NAND2_X1 U15501 ( .A1(n22261), .A2(n13791), .ZN(n13726) );
  NAND2_X1 U15502 ( .A1(n13730), .A2(n13729), .ZN(n13764) );
  AOI22_X1 U15503 ( .A1(n13810), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13800), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13735) );
  AOI22_X1 U15504 ( .A1(n13801), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13731), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13734) );
  AOI22_X1 U15505 ( .A1(n11146), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13809), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13733) );
  AOI22_X1 U15506 ( .A1(n13779), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13732) );
  NAND4_X1 U15507 ( .A1(n13735), .A2(n13734), .A3(n13733), .A4(n13732), .ZN(
        n13741) );
  AOI22_X1 U15508 ( .A1(n13563), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11168), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13739) );
  AOI22_X1 U15509 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13738) );
  AOI22_X1 U15510 ( .A1(n13778), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13737) );
  AOI22_X1 U15511 ( .A1(n13804), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13802), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13736) );
  NAND4_X1 U15512 ( .A1(n13739), .A2(n13738), .A3(n13737), .A4(n13736), .ZN(
        n13740) );
  NOR2_X1 U15513 ( .A1(n13741), .A2(n13740), .ZN(n13765) );
  XNOR2_X1 U15514 ( .A(n13764), .B(n13765), .ZN(n13746) );
  INV_X1 U15515 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13743) );
  NAND2_X1 U15516 ( .A1(n15575), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13742) );
  OAI211_X1 U15517 ( .C1(n13822), .C2(n13743), .A(n13668), .B(n13742), .ZN(
        n13744) );
  INV_X1 U15518 ( .A(n13744), .ZN(n13745) );
  OAI21_X1 U15519 ( .B1(n13746), .B2(n13794), .A(n13745), .ZN(n13753) );
  INV_X1 U15520 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n13749) );
  NAND2_X1 U15521 ( .A1(n13750), .A2(n13749), .ZN(n13751) );
  NAND2_X1 U15522 ( .A1(n13771), .A2(n13751), .ZN(n16303) );
  NAND2_X1 U15523 ( .A1(n13753), .A2(n13752), .ZN(n16071) );
  XNOR2_X1 U15524 ( .A(n13771), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16063) );
  AOI22_X1 U15525 ( .A1(n13563), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13800), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13757) );
  AOI22_X1 U15526 ( .A1(n13801), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13756) );
  AOI22_X1 U15527 ( .A1(n13731), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13013), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13755) );
  AOI22_X1 U15528 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13754) );
  NAND4_X1 U15529 ( .A1(n13757), .A2(n13756), .A3(n13755), .A4(n13754), .ZN(
        n13763) );
  AOI22_X1 U15530 ( .A1(n13804), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13778), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13761) );
  AOI22_X1 U15531 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13760) );
  AOI22_X1 U15532 ( .A1(n13779), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13802), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13759) );
  AOI22_X1 U15533 ( .A1(n13809), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13758) );
  NAND4_X1 U15534 ( .A1(n13761), .A2(n13760), .A3(n13759), .A4(n13758), .ZN(
        n13762) );
  OR2_X1 U15535 ( .A1(n13763), .A2(n13762), .ZN(n13776) );
  NOR2_X1 U15536 ( .A1(n13765), .A2(n13764), .ZN(n13777) );
  XOR2_X1 U15537 ( .A(n13776), .B(n13777), .Z(n13768) );
  INV_X1 U15538 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n15621) );
  NOR2_X1 U15539 ( .A1(n22286), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13766) );
  OAI22_X1 U15540 ( .A1(n13822), .A2(n15621), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13766), .ZN(n13767) );
  AOI21_X1 U15541 ( .B1(n13768), .B2(n13819), .A(n13767), .ZN(n13769) );
  AOI21_X1 U15542 ( .B1(n13791), .B2(n16063), .A(n13769), .ZN(n16061) );
  INV_X1 U15543 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n13770) );
  INV_X1 U15544 ( .A(n13772), .ZN(n13774) );
  INV_X1 U15545 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n13773) );
  NAND2_X1 U15546 ( .A1(n13774), .A2(n13773), .ZN(n13775) );
  NAND2_X1 U15547 ( .A1(n13835), .A2(n13775), .ZN(n16283) );
  NAND2_X1 U15548 ( .A1(n13777), .A2(n13776), .ZN(n13797) );
  AOI22_X1 U15549 ( .A1(n13801), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13800), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13783) );
  AOI22_X1 U15550 ( .A1(n13779), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13778), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13782) );
  AOI22_X1 U15551 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13781) );
  AOI22_X1 U15552 ( .A1(n13563), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13780) );
  NAND4_X1 U15553 ( .A1(n13783), .A2(n13782), .A3(n13781), .A4(n13780), .ZN(
        n13790) );
  AOI22_X1 U15554 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13788) );
  AOI22_X1 U15555 ( .A1(n13731), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11168), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13787) );
  AOI22_X1 U15556 ( .A1(n13804), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13802), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13786) );
  AOI22_X1 U15557 ( .A1(n13809), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13785) );
  NAND4_X1 U15558 ( .A1(n13788), .A2(n13787), .A3(n13786), .A4(n13785), .ZN(
        n13789) );
  NOR2_X1 U15559 ( .A1(n13790), .A2(n13789), .ZN(n13798) );
  XNOR2_X1 U15560 ( .A(n13797), .B(n13798), .ZN(n13795) );
  AOI21_X1 U15561 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n15575), .A(
        n13791), .ZN(n13793) );
  NAND2_X1 U15562 ( .A1(n13828), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n13792) );
  OAI211_X1 U15563 ( .C1(n13795), .C2(n13794), .A(n13793), .B(n13792), .ZN(
        n13796) );
  OAI21_X1 U15564 ( .B1(n13668), .B2(n16283), .A(n13796), .ZN(n16051) );
  NOR2_X1 U15565 ( .A1(n13798), .A2(n13797), .ZN(n13818) );
  AOI22_X1 U15566 ( .A1(n13799), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13563), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13808) );
  AOI22_X1 U15567 ( .A1(n13801), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13800), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13807) );
  AOI22_X1 U15568 ( .A1(n13731), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13802), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13806) );
  AOI22_X1 U15569 ( .A1(n13804), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13805) );
  NAND4_X1 U15570 ( .A1(n13808), .A2(n13807), .A3(n13806), .A4(n13805), .ZN(
        n13816) );
  AOI22_X1 U15571 ( .A1(n13013), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13779), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13814) );
  AOI22_X1 U15572 ( .A1(n11146), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13809), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13813) );
  AOI22_X1 U15573 ( .A1(n13810), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13432), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13812) );
  AOI22_X1 U15574 ( .A1(n13778), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11166), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13811) );
  NAND4_X1 U15575 ( .A1(n13814), .A2(n13813), .A3(n13812), .A4(n13811), .ZN(
        n13815) );
  NOR2_X1 U15576 ( .A1(n13816), .A2(n13815), .ZN(n13817) );
  XNOR2_X1 U15577 ( .A(n13818), .B(n13817), .ZN(n13820) );
  NAND2_X1 U15578 ( .A1(n13820), .A2(n13819), .ZN(n13826) );
  INV_X1 U15579 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n15614) );
  OAI21_X1 U15580 ( .B1(n22286), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15575), .ZN(n13821) );
  OAI21_X1 U15581 ( .B1(n13822), .B2(n15614), .A(n13821), .ZN(n13823) );
  INV_X1 U15582 ( .A(n13823), .ZN(n13825) );
  XNOR2_X1 U15583 ( .A(n13835), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16273) );
  AND2_X1 U15584 ( .A1(n16273), .A2(n13791), .ZN(n13824) );
  AOI21_X1 U15585 ( .B1(n13826), .B2(n13825), .A(n13824), .ZN(n13909) );
  AOI22_X1 U15586 ( .A1(n13828), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n13827), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13829) );
  INV_X1 U15587 ( .A(n13829), .ZN(n13830) );
  AND3_X1 U15588 ( .A1(n22274), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n17821) );
  NOR2_X2 U15589 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15786) );
  NAND2_X1 U15590 ( .A1(n15990), .A2(n20555), .ZN(n13842) );
  NAND2_X1 U15591 ( .A1(n22424), .A2(n13838), .ZN(n21875) );
  NAND2_X1 U15592 ( .A1(n21875), .A2(n22274), .ZN(n13832) );
  NAND2_X1 U15593 ( .A1(n22274), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13834) );
  NAND2_X1 U15594 ( .A1(n22286), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13833) );
  AND2_X1 U15595 ( .A1(n13834), .A2(n13833), .ZN(n14944) );
  INV_X1 U15596 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16275) );
  INV_X1 U15597 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13836) );
  INV_X1 U15598 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n17628) );
  NOR2_X1 U15599 ( .A1(n22049), .A2(n17628), .ZN(n16452) );
  AOI21_X1 U15600 ( .B1(n20588), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n16452), .ZN(n13839) );
  OAI21_X1 U15601 ( .B1(n20594), .B2(n15243), .A(n13839), .ZN(n13840) );
  INV_X1 U15602 ( .A(n13840), .ZN(n13841) );
  OAI211_X1 U15603 ( .C1(n16456), .C2(n22268), .A(n13842), .B(n13841), .ZN(
        P1_U2968) );
  INV_X1 U15604 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13844) );
  AOI22_X4 U15605 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13846), .B1(n14296), 
        .B2(n19270), .ZN(n19029) );
  OAI21_X1 U15606 ( .B1(n13847), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n13877), .ZN(n19068) );
  INV_X1 U15607 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16904) );
  AOI21_X1 U15608 ( .B1(n16904), .B2(n11253), .A(n13875), .ZN(n19030) );
  AOI21_X1 U15609 ( .B1(n13870), .B2(n12358), .A(n13872), .ZN(n19001) );
  NOR2_X1 U15610 ( .A1(n11240), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13848) );
  OR2_X1 U15611 ( .A1(n13871), .A2(n13848), .ZN(n16950) );
  INV_X1 U15612 ( .A(n16950), .ZN(n18980) );
  INV_X1 U15613 ( .A(n13868), .ZN(n13849) );
  AOI21_X1 U15614 ( .B1(n16965), .B2(n13866), .A(n13849), .ZN(n18963) );
  NOR2_X1 U15615 ( .A1(n13850), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13851) );
  OR2_X1 U15616 ( .A1(n13864), .A2(n13851), .ZN(n18961) );
  INV_X1 U15617 ( .A(n18961), .ZN(n13863) );
  AND2_X1 U15618 ( .A1(n13859), .A2(n18933), .ZN(n13852) );
  NOR2_X1 U15619 ( .A1(n13861), .A2(n13852), .ZN(n18937) );
  AOI21_X1 U15620 ( .B1(n17030), .B2(n13857), .A(n13860), .ZN(n18923) );
  AOI21_X1 U15621 ( .B1(n13853), .B2(n13855), .A(n13858), .ZN(n18898) );
  AOI21_X1 U15622 ( .B1(n15433), .B2(n13854), .A(n13856), .ZN(n15634) );
  INV_X1 U15623 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n18865) );
  AOI22_X1 U15624 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19184), .B1(n18865), 
        .B2(n19270), .ZN(n18857) );
  AOI22_X1 U15625 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14746), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19270), .ZN(n17339) );
  NOR2_X1 U15626 ( .A1(n18857), .A2(n17339), .ZN(n17338) );
  OAI21_X1 U15627 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n13854), .ZN(n17836) );
  NAND2_X1 U15628 ( .A1(n17338), .A2(n17836), .ZN(n15632) );
  NOR2_X1 U15629 ( .A1(n15634), .A2(n15632), .ZN(n18889) );
  OAI21_X1 U15630 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n13856), .A(
        n13855), .ZN(n18888) );
  NAND2_X1 U15631 ( .A1(n18889), .A2(n18888), .ZN(n18897) );
  NOR2_X1 U15632 ( .A1(n18898), .A2(n18897), .ZN(n18909) );
  OAI21_X1 U15633 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n13858), .A(
        n13857), .ZN(n18911) );
  NAND2_X1 U15634 ( .A1(n18909), .A2(n18911), .ZN(n18922) );
  NOR2_X1 U15635 ( .A1(n18923), .A2(n18922), .ZN(n15733) );
  OAI21_X1 U15636 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n13860), .A(
        n13859), .ZN(n17882) );
  NAND2_X1 U15637 ( .A1(n15733), .A2(n17882), .ZN(n18938) );
  NOR2_X1 U15638 ( .A1(n18937), .A2(n18938), .ZN(n15769) );
  NOR2_X1 U15639 ( .A1(n13861), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13862) );
  OR2_X1 U15640 ( .A1(n13850), .A2(n13862), .ZN(n17005) );
  NAND2_X1 U15641 ( .A1(n15769), .A2(n17005), .ZN(n18956) );
  NOR2_X1 U15642 ( .A1(n13863), .A2(n18956), .ZN(n15853) );
  OR2_X1 U15643 ( .A1(n13864), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13865) );
  NAND2_X1 U15644 ( .A1(n13866), .A2(n13865), .ZN(n16982) );
  NAND2_X1 U15645 ( .A1(n15853), .A2(n16982), .ZN(n18962) );
  NOR2_X1 U15646 ( .A1(n18963), .A2(n18962), .ZN(n15719) );
  AND2_X1 U15647 ( .A1(n13868), .A2(n13867), .ZN(n13869) );
  OR2_X1 U15648 ( .A1(n13869), .A2(n11240), .ZN(n16958) );
  NAND2_X1 U15649 ( .A1(n15719), .A2(n16958), .ZN(n18979) );
  NOR2_X1 U15650 ( .A1(n18980), .A2(n18979), .ZN(n18991) );
  OAI21_X1 U15651 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n13871), .A(
        n13870), .ZN(n18992) );
  NAND2_X1 U15652 ( .A1(n18991), .A2(n18992), .ZN(n19000) );
  NOR2_X1 U15653 ( .A1(n19001), .A2(n19000), .ZN(n19014) );
  INV_X1 U15654 ( .A(n13872), .ZN(n13873) );
  NAND2_X1 U15655 ( .A1(n13873), .A2(n11539), .ZN(n13874) );
  NAND2_X1 U15656 ( .A1(n11253), .A2(n13874), .ZN(n19017) );
  NAND2_X1 U15657 ( .A1(n19014), .A2(n19017), .ZN(n19028) );
  NOR2_X1 U15658 ( .A1(n19030), .A2(n19028), .ZN(n19047) );
  OAI21_X1 U15659 ( .B1(n13875), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n11236), .ZN(n19051) );
  NAND2_X1 U15660 ( .A1(n19047), .A2(n19051), .ZN(n19045) );
  INV_X1 U15661 ( .A(n13876), .ZN(n19058) );
  NAND2_X1 U15662 ( .A1(n19056), .A2(n19029), .ZN(n19067) );
  NAND2_X1 U15663 ( .A1(n19068), .A2(n19067), .ZN(n19066) );
  NAND2_X1 U15664 ( .A1(n19029), .A2(n19066), .ZN(n19080) );
  AOI21_X1 U15665 ( .B1(n19076), .B2(n13877), .A(n11256), .ZN(n16881) );
  INV_X1 U15666 ( .A(n16881), .ZN(n19081) );
  NAND2_X1 U15667 ( .A1(n19029), .A2(n19079), .ZN(n19090) );
  OR2_X1 U15668 ( .A1(n11256), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13878) );
  NAND2_X1 U15669 ( .A1(n13881), .A2(n13878), .ZN(n19091) );
  NAND2_X1 U15670 ( .A1(n19029), .A2(n19089), .ZN(n19102) );
  INV_X1 U15671 ( .A(n13879), .ZN(n13880) );
  AOI21_X1 U15672 ( .B1(n16861), .B2(n13881), .A(n13880), .ZN(n16864) );
  INV_X1 U15673 ( .A(n16864), .ZN(n19103) );
  NAND2_X1 U15674 ( .A1(n19029), .A2(n19101), .ZN(n19112) );
  NAND2_X1 U15675 ( .A1(n19029), .A2(n19111), .ZN(n19128) );
  AOI21_X1 U15676 ( .B1(n19120), .B2(n13883), .A(n13882), .ZN(n16854) );
  INV_X1 U15677 ( .A(n16854), .ZN(n19129) );
  NAND2_X1 U15678 ( .A1(n19029), .A2(n19126), .ZN(n16661) );
  INV_X1 U15679 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16838) );
  INV_X1 U15680 ( .A(n13843), .ZN(n13884) );
  AOI21_X1 U15681 ( .B1(n16838), .B2(n13884), .A(n13885), .ZN(n16836) );
  INV_X1 U15682 ( .A(n16836), .ZN(n19143) );
  XNOR2_X1 U15683 ( .A(n13885), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16825) );
  NAND4_X1 U15684 ( .A1(n19270), .A2(n19833), .A3(n22292), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19267) );
  OAI211_X1 U15685 ( .C1(n13886), .C2(n16825), .A(n19127), .B(n19164), .ZN(
        n13908) );
  INV_X1 U15686 ( .A(n16017), .ZN(n13904) );
  INV_X1 U15687 ( .A(n19247), .ZN(n13888) );
  NOR2_X1 U15688 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n13888), .ZN(n13894) );
  NAND2_X1 U15689 ( .A1(n14673), .A2(n13894), .ZN(n13889) );
  OR2_X1 U15690 ( .A1(n13887), .A2(n13889), .ZN(n19257) );
  INV_X1 U15691 ( .A(n14659), .ZN(n13890) );
  NAND2_X1 U15692 ( .A1(n19281), .A2(n22292), .ZN(n13905) );
  NAND2_X1 U15693 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n13905), .ZN(n13891) );
  NAND2_X1 U15694 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19833), .ZN(n19273) );
  NOR3_X1 U15695 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n19916), .A3(n19273), 
        .ZN(n19277) );
  NAND2_X1 U15696 ( .A1(n19267), .A2(n18976), .ZN(n13892) );
  NOR2_X1 U15697 ( .A1(n19277), .A2(n13892), .ZN(n13893) );
  INV_X1 U15698 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13899) );
  INV_X1 U15699 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n19154) );
  NAND2_X1 U15700 ( .A1(n19154), .A2(n13905), .ZN(n13895) );
  AOI21_X1 U15701 ( .B1(n13896), .B2(n13895), .A(n13894), .ZN(n13897) );
  AOI22_X1 U15702 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(n19135), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19134), .ZN(n13898) );
  OAI21_X1 U15703 ( .B1(n19121), .B2(n13899), .A(n13898), .ZN(n13900) );
  INV_X1 U15704 ( .A(n13900), .ZN(n13901) );
  NAND3_X1 U15705 ( .A1(n13908), .A2(n13907), .A3(n11632), .ZN(P2_U2825) );
  NOR2_X1 U15706 ( .A1(n16026), .A2(n16592), .ZN(n14871) );
  NAND3_X1 U15707 ( .A1(n16030), .A2(n16042), .A3(n16036), .ZN(n13914) );
  INV_X1 U15708 ( .A(n13915), .ZN(n16033) );
  NAND4_X1 U15709 ( .A1(n16033), .A2(n12961), .A3(n16042), .A4(n13911), .ZN(
        n14932) );
  NOR2_X1 U15710 ( .A1(n14932), .A2(n15972), .ZN(n13912) );
  NAND2_X1 U15711 ( .A1(n11195), .A2(n13912), .ZN(n13913) );
  NAND2_X1 U15712 ( .A1(n15167), .A2(n16021), .ZN(n13936) );
  AND2_X1 U15713 ( .A1(n15972), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13917) );
  AOI21_X1 U15714 ( .B1(n15973), .B2(P1_EBX_REG_30__SCAN_IN), .A(n13917), .ZN(
        n15971) );
  INV_X1 U15715 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n22064) );
  NAND2_X1 U15716 ( .A1(n13936), .A2(n22064), .ZN(n13921) );
  INV_X1 U15717 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13919) );
  NAND2_X1 U15718 ( .A1(n13918), .A2(n13919), .ZN(n13920) );
  NAND3_X1 U15719 ( .A1(n13921), .A2(n12989), .A3(n13920), .ZN(n13922) );
  NAND2_X1 U15720 ( .A1(n13936), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n13924) );
  INV_X1 U15721 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n14988) );
  NAND2_X1 U15722 ( .A1(n12989), .A2(n14988), .ZN(n13923) );
  AND2_X1 U15723 ( .A1(n13924), .A2(n13923), .ZN(n14914) );
  OR2_X1 U15724 ( .A1(n13925), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n13928) );
  NAND2_X1 U15725 ( .A1(n13936), .A2(n16433), .ZN(n13926) );
  OAI211_X1 U15726 ( .C1(P1_EBX_REG_2__SCAN_IN), .C2(n15972), .A(n13926), .B(
        n14002), .ZN(n13927) );
  AND2_X1 U15727 ( .A1(n13928), .A2(n13927), .ZN(n15081) );
  MUX2_X1 U15728 ( .A(n13997), .B(n14002), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n13931) );
  OAI21_X1 U15729 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n15973), .A(
        n13931), .ZN(n15373) );
  OR2_X1 U15730 ( .A1(n13925), .A2(P1_EBX_REG_4__SCAN_IN), .ZN(n13935) );
  NAND2_X1 U15731 ( .A1(n13936), .A2(n21930), .ZN(n13933) );
  INV_X1 U15732 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n15399) );
  NAND2_X1 U15733 ( .A1(n13918), .A2(n15399), .ZN(n13932) );
  NAND3_X1 U15734 ( .A1(n13933), .A2(n14002), .A3(n13932), .ZN(n13934) );
  NAND2_X1 U15735 ( .A1(n13935), .A2(n13934), .ZN(n15396) );
  NAND2_X1 U15736 ( .A1(n14002), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13937) );
  OAI211_X1 U15737 ( .C1(P1_EBX_REG_5__SCAN_IN), .C2(n15972), .A(n13936), .B(
        n13937), .ZN(n13938) );
  OAI21_X1 U15738 ( .B1(n13997), .B2(P1_EBX_REG_5__SCAN_IN), .A(n13938), .ZN(
        n20525) );
  OR2_X1 U15739 ( .A1(n13925), .A2(P1_EBX_REG_6__SCAN_IN), .ZN(n13941) );
  NAND2_X1 U15740 ( .A1(n13936), .A2(n21949), .ZN(n13939) );
  OAI211_X1 U15741 ( .C1(P1_EBX_REG_6__SCAN_IN), .C2(n15972), .A(n13939), .B(
        n14002), .ZN(n13940) );
  MUX2_X1 U15742 ( .A(n13997), .B(n14002), .S(P1_EBX_REG_7__SCAN_IN), .Z(
        n13942) );
  OAI21_X1 U15743 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n15973), .A(
        n13942), .ZN(n15651) );
  OR2_X1 U15744 ( .A1(n13925), .A2(P1_EBX_REG_8__SCAN_IN), .ZN(n13945) );
  NAND2_X1 U15745 ( .A1(n13936), .A2(n21966), .ZN(n13943) );
  OAI211_X1 U15746 ( .C1(P1_EBX_REG_8__SCAN_IN), .C2(n15972), .A(n13943), .B(
        n14002), .ZN(n13944) );
  NAND2_X1 U15747 ( .A1(n13945), .A2(n13944), .ZN(n15857) );
  NAND2_X1 U15748 ( .A1(n15650), .A2(n15857), .ZN(n15866) );
  MUX2_X1 U15749 ( .A(n13997), .B(n14002), .S(P1_EBX_REG_9__SCAN_IN), .Z(
        n13946) );
  OAI21_X1 U15750 ( .B1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15973), .A(
        n13946), .ZN(n15865) );
  OR2_X1 U15751 ( .A1(n13925), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n13950) );
  NAND2_X1 U15752 ( .A1(n13936), .A2(n21993), .ZN(n13948) );
  OAI211_X1 U15753 ( .C1(P1_EBX_REG_10__SCAN_IN), .C2(n15972), .A(n13948), .B(
        n14002), .ZN(n13949) );
  MUX2_X1 U15754 ( .A(n13997), .B(n14002), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n13951) );
  OAI21_X1 U15755 ( .B1(n15973), .B2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n13951), .ZN(n13952) );
  INV_X1 U15756 ( .A(n13952), .ZN(n16185) );
  OR2_X1 U15757 ( .A1(n13925), .A2(P1_EBX_REG_12__SCAN_IN), .ZN(n13956) );
  NAND2_X1 U15758 ( .A1(n14002), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13953) );
  NAND2_X1 U15759 ( .A1(n13936), .A2(n13953), .ZN(n13954) );
  OAI21_X1 U15760 ( .B1(P1_EBX_REG_12__SCAN_IN), .B2(n15972), .A(n13954), .ZN(
        n13955) );
  NAND2_X1 U15761 ( .A1(n13956), .A2(n13955), .ZN(n15948) );
  NAND2_X1 U15762 ( .A1(n14002), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13957) );
  OAI211_X1 U15763 ( .C1(P1_EBX_REG_13__SCAN_IN), .C2(n15972), .A(n13936), .B(
        n13957), .ZN(n13958) );
  OAI21_X1 U15764 ( .B1(n13997), .B2(P1_EBX_REG_13__SCAN_IN), .A(n13958), .ZN(
        n16136) );
  OR2_X1 U15765 ( .A1(n13925), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n13962) );
  NAND2_X1 U15766 ( .A1(n13936), .A2(n13959), .ZN(n13960) );
  OAI211_X1 U15767 ( .C1(P1_EBX_REG_14__SCAN_IN), .C2(n15972), .A(n13960), .B(
        n14002), .ZN(n13961) );
  MUX2_X1 U15768 ( .A(n13997), .B(n14002), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n13963) );
  OAI21_X1 U15769 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15973), .A(
        n13963), .ZN(n13964) );
  INV_X1 U15770 ( .A(n13964), .ZN(n20506) );
  OR2_X1 U15771 ( .A1(n13925), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n13968) );
  INV_X1 U15772 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n22034) );
  NAND2_X1 U15773 ( .A1(n13936), .A2(n22034), .ZN(n13966) );
  INV_X1 U15774 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n22171) );
  NAND2_X1 U15775 ( .A1(n13918), .A2(n22171), .ZN(n13965) );
  NAND3_X1 U15776 ( .A1(n13966), .A2(n14002), .A3(n13965), .ZN(n13967) );
  NAND2_X1 U15777 ( .A1(n13968), .A2(n13967), .ZN(n16176) );
  MUX2_X1 U15778 ( .A(n13997), .B(n14002), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n13969) );
  OAI21_X1 U15779 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n15973), .A(
        n13969), .ZN(n16127) );
  OR2_X1 U15780 ( .A1(n13925), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n13972) );
  NAND2_X1 U15781 ( .A1(n13936), .A2(n22022), .ZN(n13970) );
  OAI211_X1 U15782 ( .C1(P1_EBX_REG_18__SCAN_IN), .C2(n15972), .A(n13970), .B(
        n14002), .ZN(n13971) );
  MUX2_X1 U15783 ( .A(n13997), .B(n14002), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n13973) );
  OAI21_X1 U15784 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n15973), .A(
        n13973), .ZN(n20519) );
  OR2_X1 U15785 ( .A1(n13925), .A2(P1_EBX_REG_20__SCAN_IN), .ZN(n13978) );
  INV_X1 U15786 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16569) );
  NAND2_X1 U15787 ( .A1(n13936), .A2(n16569), .ZN(n13976) );
  INV_X1 U15788 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n13974) );
  NAND2_X1 U15789 ( .A1(n13918), .A2(n13974), .ZN(n13975) );
  NAND3_X1 U15790 ( .A1(n13976), .A2(n14002), .A3(n13975), .ZN(n13977) );
  NAND2_X1 U15791 ( .A1(n13978), .A2(n13977), .ZN(n16117) );
  INV_X1 U15792 ( .A(n13997), .ZN(n13979) );
  INV_X1 U15793 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n20518) );
  NAND2_X1 U15794 ( .A1(n13979), .A2(n20518), .ZN(n13982) );
  NAND2_X1 U15795 ( .A1(n14002), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13980) );
  OAI211_X1 U15796 ( .C1(P1_EBX_REG_21__SCAN_IN), .C2(n15972), .A(n13936), .B(
        n13980), .ZN(n13981) );
  OR2_X1 U15797 ( .A1(n13925), .A2(P1_EBX_REG_22__SCAN_IN), .ZN(n13985) );
  NAND2_X1 U15798 ( .A1(n13936), .A2(n16432), .ZN(n13983) );
  OAI211_X1 U15799 ( .C1(P1_EBX_REG_22__SCAN_IN), .C2(n15972), .A(n13983), .B(
        n14002), .ZN(n13984) );
  NAND2_X1 U15800 ( .A1(n13985), .A2(n13984), .ZN(n16161) );
  MUX2_X1 U15801 ( .A(n13997), .B(n14002), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n13986) );
  OAI21_X1 U15802 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15973), .A(
        n13986), .ZN(n16524) );
  OR2_X1 U15803 ( .A1(n13925), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n13989) );
  INV_X1 U15804 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16325) );
  NAND2_X1 U15805 ( .A1(n13936), .A2(n16325), .ZN(n13987) );
  OAI211_X1 U15806 ( .C1(P1_EBX_REG_24__SCAN_IN), .C2(n15972), .A(n13987), .B(
        n14002), .ZN(n13988) );
  MUX2_X1 U15807 ( .A(n13997), .B(n14002), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n13992) );
  INV_X1 U15808 ( .A(n15973), .ZN(n14001) );
  INV_X1 U15809 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n13990) );
  NAND2_X1 U15810 ( .A1(n14001), .A2(n13990), .ZN(n13991) );
  OR2_X1 U15811 ( .A1(n13925), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n13996) );
  NAND2_X1 U15812 ( .A1(n14002), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13993) );
  NAND2_X1 U15813 ( .A1(n13936), .A2(n13993), .ZN(n13994) );
  OAI21_X1 U15814 ( .B1(P1_EBX_REG_26__SCAN_IN), .B2(n15972), .A(n13994), .ZN(
        n13995) );
  NAND2_X1 U15815 ( .A1(n13996), .A2(n13995), .ZN(n16082) );
  MUX2_X1 U15816 ( .A(n13997), .B(n14002), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n13998) );
  OAI21_X1 U15817 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n15973), .A(
        n13998), .ZN(n16073) );
  INV_X1 U15818 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n17494) );
  OAI21_X1 U15819 ( .B1(n15972), .B2(P1_EBX_REG_28__SCAN_IN), .A(n14002), .ZN(
        n13999) );
  AOI21_X1 U15820 ( .B1(n16291), .B2(n13936), .A(n13999), .ZN(n14000) );
  AOI21_X1 U15821 ( .B1(n11477), .B2(n17494), .A(n14000), .ZN(n16062) );
  NOR2_X1 U15822 ( .A1(n15972), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n14003) );
  AOI21_X1 U15823 ( .B1(n14001), .B2(n13246), .A(n14003), .ZN(n14004) );
  MUX2_X1 U15824 ( .A(n14003), .B(n14004), .S(n14002), .Z(n16053) );
  AOI22_X1 U15825 ( .A1(n16052), .A2(n14838), .B1(n14004), .B2(n11210), .ZN(
        n14005) );
  XOR2_X1 U15826 ( .A(n15971), .B(n14005), .Z(n16465) );
  INV_X1 U15827 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n16043) );
  NAND2_X1 U15828 ( .A1(n14009), .A2(n14008), .ZN(P1_U2842) );
  INV_X1 U15829 ( .A(n19259), .ZN(n14010) );
  NAND2_X1 U15830 ( .A1(n15441), .A2(n14010), .ZN(n14015) );
  NAND2_X1 U15831 ( .A1(n11772), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14011) );
  NAND2_X1 U15832 ( .A1(n19897), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n14020) );
  AOI21_X1 U15833 ( .B1(n19809), .B2(n14020), .A(n19942), .ZN(n14013) );
  INV_X1 U15834 ( .A(n14020), .ZN(n14012) );
  NAND2_X1 U15835 ( .A1(n14012), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19755) );
  AOI21_X1 U15836 ( .B1(n14027), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19786), .ZN(n14014) );
  INV_X1 U15837 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n20152) );
  NOR2_X1 U15838 ( .A1(n14210), .A2(n20152), .ZN(n14017) );
  INV_X1 U15839 ( .A(n19897), .ZN(n14025) );
  NAND2_X1 U15840 ( .A1(n14025), .A2(n19832), .ZN(n14019) );
  NAND2_X1 U15841 ( .A1(n14020), .A2(n14019), .ZN(n19787) );
  NOR2_X1 U15842 ( .A1(n19787), .A2(n19942), .ZN(n14021) );
  AOI21_X1 U15843 ( .B1(n14027), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n14021), .ZN(n14022) );
  INV_X1 U15844 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n20194) );
  OAI21_X1 U15845 ( .B1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n14025), .ZN(n19858) );
  NOR2_X1 U15846 ( .A1(n19858), .A2(n19942), .ZN(n19911) );
  AOI21_X1 U15847 ( .B1(n14027), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n19911), .ZN(n14026) );
  NAND2_X1 U15848 ( .A1(n11772), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n14032) );
  AND2_X1 U15849 ( .A1(n14033), .A2(n14032), .ZN(n14034) );
  INV_X1 U15850 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n20112) );
  NOR2_X1 U15851 ( .A1(n14210), .A2(n20112), .ZN(n14975) );
  INV_X1 U15852 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n20009) );
  INV_X1 U15853 ( .A(n15077), .ZN(n14035) );
  AND2_X1 U15854 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n14035), .ZN(
        n14036) );
  AOI22_X1 U15855 ( .A1(n14068), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14069), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14041) );
  AOI22_X1 U15856 ( .A1(n14071), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14072), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14040) );
  AOI22_X1 U15857 ( .A1(n14126), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11942), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14039) );
  AOI22_X1 U15858 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17363), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14038) );
  NAND4_X1 U15859 ( .A1(n14041), .A2(n14040), .A3(n14039), .A4(n14038), .ZN(
        n14047) );
  AOI22_X1 U15860 ( .A1(n11909), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11901), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14045) );
  AOI22_X1 U15861 ( .A1(n14104), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11921), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14044) );
  AOI22_X1 U15862 ( .A1(n11962), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11906), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14043) );
  AOI22_X1 U15863 ( .A1(n11907), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11908), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14042) );
  NAND4_X1 U15864 ( .A1(n14045), .A2(n14044), .A3(n14043), .A4(n14042), .ZN(
        n14046) );
  AOI22_X1 U15865 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n14068), .B1(
        n14069), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14051) );
  AOI22_X1 U15866 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n14072), .B1(
        n14071), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14050) );
  AOI22_X1 U15867 ( .A1(n14126), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11942), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14049) );
  AOI22_X1 U15868 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12556), .B1(
        n17363), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14048) );
  NAND4_X1 U15869 ( .A1(n14051), .A2(n14050), .A3(n14049), .A4(n14048), .ZN(
        n14057) );
  AOI22_X1 U15870 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11901), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14055) );
  AOI22_X1 U15871 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n11921), .B1(
        n14104), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14054) );
  AOI22_X1 U15872 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n11906), .B1(
        n11962), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14053) );
  AOI22_X1 U15873 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n11907), .B1(
        n11908), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14052) );
  NAND4_X1 U15874 ( .A1(n14055), .A2(n14054), .A3(n14053), .A4(n14052), .ZN(
        n14056) );
  NOR2_X1 U15875 ( .A1(n14057), .A2(n14056), .ZN(n15834) );
  AOI22_X1 U15876 ( .A1(n14068), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14069), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14061) );
  AOI22_X1 U15877 ( .A1(n14071), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14072), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14060) );
  AOI22_X1 U15878 ( .A1(n14126), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11942), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14059) );
  AOI22_X1 U15879 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17363), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14058) );
  NAND4_X1 U15880 ( .A1(n14061), .A2(n14060), .A3(n14059), .A4(n14058), .ZN(
        n14067) );
  AOI22_X1 U15881 ( .A1(n11909), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11901), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14065) );
  AOI22_X1 U15882 ( .A1(n14104), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11921), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14064) );
  AOI22_X1 U15883 ( .A1(n11962), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11906), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14063) );
  AOI22_X1 U15884 ( .A1(n11907), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11908), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14062) );
  NAND4_X1 U15885 ( .A1(n14065), .A2(n14064), .A3(n14063), .A4(n14062), .ZN(
        n14066) );
  INV_X1 U15886 ( .A(n14068), .ZN(n14099) );
  INV_X1 U15887 ( .A(n14069), .ZN(n14098) );
  OAI22_X1 U15888 ( .A1(n14099), .A2(n20152), .B1(n14098), .B2(n14070), .ZN(
        n14086) );
  INV_X1 U15889 ( .A(n14071), .ZN(n14103) );
  INV_X1 U15890 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14074) );
  INV_X1 U15891 ( .A(n14072), .ZN(n14101) );
  INV_X1 U15892 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14073) );
  OAI22_X1 U15893 ( .A1(n14103), .A2(n14074), .B1(n14101), .B2(n14073), .ZN(
        n14085) );
  INV_X1 U15894 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14078) );
  AOI22_X1 U15895 ( .A1(n14126), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11942), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14076) );
  NAND2_X1 U15896 ( .A1(n17363), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n14075) );
  OAI211_X1 U15897 ( .C1(n14078), .C2(n14077), .A(n14076), .B(n14075), .ZN(
        n14084) );
  AOI22_X1 U15898 ( .A1(n11909), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11901), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14082) );
  AOI22_X1 U15899 ( .A1(n14104), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11921), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14081) );
  AOI22_X1 U15900 ( .A1(n11962), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11906), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14080) );
  AOI22_X1 U15901 ( .A1(n11907), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11908), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14079) );
  NAND4_X1 U15902 ( .A1(n14082), .A2(n14081), .A3(n14080), .A4(n14079), .ZN(
        n14083) );
  NOR4_X1 U15903 ( .A1(n14086), .A2(n14085), .A3(n14084), .A4(n14083), .ZN(
        n15911) );
  AOI22_X1 U15904 ( .A1(n14068), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n14069), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14090) );
  AOI22_X1 U15905 ( .A1(n14071), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n14072), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14089) );
  AOI22_X1 U15906 ( .A1(n14126), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11942), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14088) );
  AOI22_X1 U15907 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17363), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14087) );
  NAND4_X1 U15908 ( .A1(n14090), .A2(n14089), .A3(n14088), .A4(n14087), .ZN(
        n14096) );
  AOI22_X1 U15909 ( .A1(n11909), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11901), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14094) );
  AOI22_X1 U15910 ( .A1(n14104), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11921), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14093) );
  AOI22_X1 U15911 ( .A1(n11962), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11906), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14092) );
  AOI22_X1 U15912 ( .A1(n11907), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11908), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14091) );
  NAND4_X1 U15913 ( .A1(n14094), .A2(n14093), .A3(n14092), .A4(n14091), .ZN(
        n14095) );
  OR2_X1 U15914 ( .A1(n14096), .A2(n14095), .ZN(n16735) );
  INV_X1 U15915 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n20059) );
  OAI22_X1 U15916 ( .A1(n20059), .A2(n14099), .B1(n14098), .B2(n14097), .ZN(
        n14114) );
  INV_X1 U15917 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14102) );
  INV_X1 U15918 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14100) );
  OAI22_X1 U15919 ( .A1(n14103), .A2(n14102), .B1(n14101), .B2(n14100), .ZN(
        n14113) );
  AOI22_X1 U15920 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n11901), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14108) );
  AOI22_X1 U15921 ( .A1(n14104), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11921), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14107) );
  AOI22_X1 U15922 ( .A1(n11962), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11906), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14106) );
  AOI22_X1 U15923 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n11908), .B1(
        n11907), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14105) );
  NAND4_X1 U15924 ( .A1(n14108), .A2(n14107), .A3(n14106), .A4(n14105), .ZN(
        n14112) );
  AOI22_X1 U15925 ( .A1(n14126), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11942), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14110) );
  AOI22_X1 U15926 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17363), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14109) );
  NAND2_X1 U15927 ( .A1(n14110), .A2(n14109), .ZN(n14111) );
  NOR4_X1 U15928 ( .A1(n14114), .A2(n14113), .A3(n14112), .A4(n14111), .ZN(
        n16731) );
  AOI22_X1 U15929 ( .A1(n14068), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14069), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14118) );
  AOI22_X1 U15930 ( .A1(n14071), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n14072), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14117) );
  AOI22_X1 U15931 ( .A1(n14126), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11942), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14116) );
  AOI22_X1 U15932 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17363), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14115) );
  NAND4_X1 U15933 ( .A1(n14118), .A2(n14117), .A3(n14116), .A4(n14115), .ZN(
        n14125) );
  AOI22_X1 U15934 ( .A1(n11909), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11901), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14123) );
  AOI22_X1 U15935 ( .A1(n14104), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11921), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14122) );
  AOI22_X1 U15936 ( .A1(n11962), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11906), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14121) );
  AOI22_X1 U15937 ( .A1(n11907), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11908), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14120) );
  NAND4_X1 U15938 ( .A1(n14123), .A2(n14122), .A3(n14121), .A4(n14120), .ZN(
        n14124) );
  AOI22_X1 U15939 ( .A1(n14068), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n14069), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14130) );
  AOI22_X1 U15940 ( .A1(n14071), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14072), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14129) );
  AOI22_X1 U15941 ( .A1(n14126), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11942), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14128) );
  AOI22_X1 U15942 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17363), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14127) );
  NAND4_X1 U15943 ( .A1(n14130), .A2(n14129), .A3(n14128), .A4(n14127), .ZN(
        n14136) );
  AOI22_X1 U15944 ( .A1(n11909), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11901), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14134) );
  AOI22_X1 U15945 ( .A1(n14104), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11921), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14133) );
  AOI22_X1 U15946 ( .A1(n11962), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11906), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14132) );
  AOI22_X1 U15947 ( .A1(n11907), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11908), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14131) );
  NAND4_X1 U15948 ( .A1(n14134), .A2(n14133), .A3(n14132), .A4(n14131), .ZN(
        n14135) );
  AOI22_X1 U15949 ( .A1(n14277), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11183), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14145) );
  AND2_X1 U15950 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14138) );
  OR2_X1 U15951 ( .A1(n14138), .A2(n14137), .ZN(n14276) );
  INV_X1 U15952 ( .A(n14276), .ZN(n14255) );
  INV_X1 U15953 ( .A(n14139), .ZN(n14274) );
  NAND2_X1 U15954 ( .A1(n14139), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n14141) );
  NAND2_X1 U15955 ( .A1(n14156), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n14140) );
  AND3_X1 U15956 ( .A1(n14255), .A2(n14141), .A3(n14140), .ZN(n14144) );
  AOI22_X1 U15957 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14142) );
  NAND4_X1 U15958 ( .A1(n14145), .A2(n14144), .A3(n14143), .A4(n14142), .ZN(
        n14153) );
  AOI22_X1 U15959 ( .A1(n11186), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11183), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14151) );
  NAND2_X1 U15960 ( .A1(n14139), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n14147) );
  NAND2_X1 U15961 ( .A1(n14156), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n14146) );
  AND3_X1 U15962 ( .A1(n14147), .A2(n14276), .A3(n14146), .ZN(n14150) );
  AOI22_X1 U15963 ( .A1(n14277), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11883), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14148) );
  NAND4_X1 U15964 ( .A1(n14151), .A2(n14150), .A3(n14149), .A4(n14148), .ZN(
        n14152) );
  AND2_X1 U15965 ( .A1(n14153), .A2(n14152), .ZN(n14154) );
  XNOR2_X1 U15966 ( .A(n14155), .B(n14154), .ZN(n16718) );
  NAND2_X1 U15967 ( .A1(n14155), .A2(n14154), .ZN(n14171) );
  NAND2_X1 U15968 ( .A1(n14139), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n14158) );
  NAND2_X1 U15969 ( .A1(n14156), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n14157) );
  AND3_X1 U15970 ( .A1(n14255), .A2(n14158), .A3(n14157), .ZN(n14161) );
  AOI22_X1 U15971 ( .A1(n14277), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11185), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14160) );
  AOI22_X1 U15972 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11170), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14159) );
  NAND4_X1 U15973 ( .A1(n14162), .A2(n14161), .A3(n14160), .A4(n14159), .ZN(
        n14170) );
  AOI22_X1 U15974 ( .A1(n14277), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11185), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14167) );
  AOI22_X1 U15975 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n11883), .B1(
        n11170), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14166) );
  NAND2_X1 U15976 ( .A1(n14139), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n14164) );
  NAND2_X1 U15977 ( .A1(n14156), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n14163) );
  AND3_X1 U15978 ( .A1(n14164), .A2(n14276), .A3(n14163), .ZN(n14165) );
  NAND4_X1 U15979 ( .A1(n14168), .A2(n14167), .A3(n14166), .A4(n14165), .ZN(
        n14169) );
  NAND2_X1 U15980 ( .A1(n14170), .A2(n14169), .ZN(n14173) );
  NOR2_X1 U15981 ( .A1(n14171), .A2(n14173), .ZN(n14195) );
  INV_X1 U15982 ( .A(n14210), .ZN(n14231) );
  INV_X1 U15983 ( .A(n14171), .ZN(n14172) );
  NAND2_X1 U15984 ( .A1(n14231), .A2(n14172), .ZN(n14174) );
  AOI22_X1 U15985 ( .A1(n14195), .A2(n13896), .B1(n14174), .B2(n14173), .ZN(
        n16711) );
  INV_X1 U15986 ( .A(n14195), .ZN(n14189) );
  AOI22_X1 U15987 ( .A1(n14277), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11184), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14179) );
  NAND2_X1 U15988 ( .A1(n14139), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n14176) );
  NAND2_X1 U15989 ( .A1(n14156), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n14175) );
  AND3_X1 U15990 ( .A1(n14255), .A2(n14176), .A3(n14175), .ZN(n14178) );
  AOI22_X1 U15991 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11170), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14177) );
  NAND4_X1 U15992 ( .A1(n14180), .A2(n14179), .A3(n14178), .A4(n14177), .ZN(
        n14188) );
  AOI22_X1 U15993 ( .A1(n14277), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11185), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14185) );
  AOI22_X1 U15994 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14184) );
  NAND2_X1 U15995 ( .A1(n14139), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n14182) );
  NAND2_X1 U15996 ( .A1(n14156), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n14181) );
  AND3_X1 U15997 ( .A1(n14182), .A2(n14276), .A3(n14181), .ZN(n14183) );
  NAND4_X1 U15998 ( .A1(n14186), .A2(n14185), .A3(n14184), .A4(n14183), .ZN(
        n14187) );
  AND2_X1 U15999 ( .A1(n14188), .A2(n14187), .ZN(n14194) );
  XNOR2_X1 U16000 ( .A(n14189), .B(n14194), .ZN(n14190) );
  NAND2_X1 U16001 ( .A1(n14190), .A2(n14231), .ZN(n14193) );
  INV_X1 U16002 ( .A(n14193), .ZN(n14191) );
  INV_X1 U16003 ( .A(n14194), .ZN(n14192) );
  NOR2_X1 U16004 ( .A1(n13896), .A2(n14192), .ZN(n16705) );
  NAND2_X1 U16005 ( .A1(n14195), .A2(n14194), .ZN(n14211) );
  NAND2_X1 U16006 ( .A1(n14139), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n14197) );
  NAND2_X1 U16007 ( .A1(n14156), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n14196) );
  AND3_X1 U16008 ( .A1(n14255), .A2(n14197), .A3(n14196), .ZN(n14200) );
  AOI22_X1 U16009 ( .A1(n14277), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11184), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14199) );
  AOI22_X1 U16010 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14198) );
  NAND4_X1 U16011 ( .A1(n14201), .A2(n14200), .A3(n14199), .A4(n14198), .ZN(
        n14209) );
  AOI22_X1 U16012 ( .A1(n14277), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11184), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14206) );
  AOI22_X1 U16013 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11170), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14205) );
  NAND2_X1 U16014 ( .A1(n14139), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n14203) );
  NAND2_X1 U16015 ( .A1(n14156), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n14202) );
  AND3_X1 U16016 ( .A1(n14203), .A2(n14276), .A3(n14202), .ZN(n14204) );
  NAND4_X1 U16017 ( .A1(n14207), .A2(n14206), .A3(n14205), .A4(n14204), .ZN(
        n14208) );
  NAND2_X1 U16018 ( .A1(n14209), .A2(n14208), .ZN(n14213) );
  AOI21_X1 U16019 ( .B1(n14211), .B2(n14213), .A(n14210), .ZN(n14212) );
  INV_X1 U16020 ( .A(n14213), .ZN(n14214) );
  NAND2_X1 U16021 ( .A1(n14673), .A2(n14214), .ZN(n16698) );
  INV_X1 U16022 ( .A(n14230), .ZN(n14233) );
  NAND2_X1 U16023 ( .A1(n14139), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n14217) );
  NAND2_X1 U16024 ( .A1(n14156), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n14216) );
  AND3_X1 U16025 ( .A1(n14255), .A2(n14217), .A3(n14216), .ZN(n14220) );
  AOI22_X1 U16026 ( .A1(n14277), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11184), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14219) );
  AOI22_X1 U16027 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14218) );
  NAND4_X1 U16028 ( .A1(n14221), .A2(n14220), .A3(n14219), .A4(n14218), .ZN(
        n14229) );
  AOI22_X1 U16029 ( .A1(n14277), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11184), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14226) );
  AOI22_X1 U16030 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11170), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14225) );
  NAND2_X1 U16031 ( .A1(n14139), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n14223) );
  NAND2_X1 U16032 ( .A1(n14156), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n14222) );
  AND3_X1 U16033 ( .A1(n14223), .A2(n14276), .A3(n14222), .ZN(n14224) );
  NAND4_X1 U16034 ( .A1(n14227), .A2(n14226), .A3(n14225), .A4(n14224), .ZN(
        n14228) );
  NAND2_X1 U16035 ( .A1(n14229), .A2(n14228), .ZN(n14234) );
  INV_X1 U16036 ( .A(n14234), .ZN(n14232) );
  OR2_X1 U16037 ( .A1(n14230), .A2(n14234), .ZN(n16684) );
  OAI211_X1 U16038 ( .C1(n14233), .C2(n14232), .A(n14231), .B(n16684), .ZN(
        n14250) );
  NOR2_X1 U16039 ( .A1(n13896), .A2(n14234), .ZN(n16692) );
  AOI22_X1 U16040 ( .A1(n14277), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11184), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14240) );
  NAND2_X1 U16041 ( .A1(n14139), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n14237) );
  NAND2_X1 U16042 ( .A1(n14156), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n14236) );
  AND3_X1 U16043 ( .A1(n14255), .A2(n14237), .A3(n14236), .ZN(n14239) );
  AOI22_X1 U16044 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14238) );
  NAND4_X1 U16045 ( .A1(n14241), .A2(n14240), .A3(n14239), .A4(n14238), .ZN(
        n14249) );
  AOI22_X1 U16046 ( .A1(n14277), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11184), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14246) );
  AOI22_X1 U16047 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11170), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14245) );
  NAND2_X1 U16048 ( .A1(n14139), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n14243) );
  NAND2_X1 U16049 ( .A1(n14156), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n14242) );
  AND3_X1 U16050 ( .A1(n14243), .A2(n14276), .A3(n14242), .ZN(n14244) );
  NAND4_X1 U16051 ( .A1(n14247), .A2(n14246), .A3(n14245), .A4(n14244), .ZN(
        n14248) );
  AND2_X1 U16052 ( .A1(n14249), .A2(n14248), .ZN(n16685) );
  NAND2_X1 U16053 ( .A1(n14251), .A2(n14250), .ZN(n16689) );
  INV_X1 U16054 ( .A(n16684), .ZN(n14252) );
  NAND3_X1 U16055 ( .A1(n14252), .A2(n16685), .A3(n13896), .ZN(n16676) );
  AOI22_X1 U16056 ( .A1(n11188), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11184), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14258) );
  NAND2_X1 U16057 ( .A1(n14139), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n14254) );
  NAND2_X1 U16058 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n14253) );
  AND3_X1 U16059 ( .A1(n14255), .A2(n14254), .A3(n14253), .ZN(n14257) );
  AOI22_X1 U16060 ( .A1(n14156), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14256) );
  NAND4_X1 U16061 ( .A1(n14259), .A2(n14258), .A3(n14257), .A4(n14256), .ZN(
        n14267) );
  AOI22_X1 U16062 ( .A1(n14277), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11184), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14264) );
  AOI22_X1 U16063 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11170), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14263) );
  NAND2_X1 U16064 ( .A1(n14139), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n14261) );
  NAND2_X1 U16065 ( .A1(n14156), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n14260) );
  AND3_X1 U16066 ( .A1(n14261), .A2(n14276), .A3(n14260), .ZN(n14262) );
  NAND4_X1 U16067 ( .A1(n14265), .A2(n14264), .A3(n14263), .A4(n14262), .ZN(
        n14266) );
  NAND2_X1 U16068 ( .A1(n14267), .A2(n14266), .ZN(n16675) );
  AOI22_X1 U16069 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11170), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14270) );
  NAND2_X1 U16070 ( .A1(n14139), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n14269) );
  NAND2_X1 U16071 ( .A1(n14156), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n14268) );
  NAND4_X1 U16072 ( .A1(n14270), .A2(n14269), .A3(n14268), .A4(n14276), .ZN(
        n14285) );
  AOI22_X1 U16073 ( .A1(n11188), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11184), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14271) );
  NAND2_X1 U16074 ( .A1(n14272), .A2(n14271), .ZN(n14284) );
  NOR2_X1 U16075 ( .A1(n14274), .A2(n14273), .ZN(n14275) );
  AOI211_X1 U16076 ( .C1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .C2(n14156), .A(
        n14276), .B(n14275), .ZN(n14282) );
  AOI22_X1 U16077 ( .A1(n11187), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11184), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14281) );
  AOI22_X1 U16078 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14279) );
  NAND4_X1 U16079 ( .A1(n14282), .A2(n14281), .A3(n14280), .A4(n14279), .ZN(
        n14283) );
  OAI21_X1 U16080 ( .B1(n14285), .B2(n14284), .A(n14283), .ZN(n14286) );
  INV_X1 U16081 ( .A(n14286), .ZN(n14287) );
  XNOR2_X1 U16082 ( .A(n14288), .B(n14287), .ZN(n16020) );
  INV_X1 U16083 ( .A(n19242), .ZN(n14289) );
  NAND2_X1 U16084 ( .A1(n14289), .A2(n19239), .ZN(n15760) );
  INV_X1 U16085 ( .A(n12732), .ZN(n17344) );
  NAND2_X1 U16086 ( .A1(n15760), .A2(n17344), .ZN(n14290) );
  NOR2_X1 U16087 ( .A1(n16829), .A2(n11141), .ZN(n14291) );
  AOI21_X1 U16088 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n11141), .A(n14291), .ZN(
        n14292) );
  OAI21_X1 U16089 ( .B1(n16020), .B2(n16740), .A(n14292), .ZN(P2_U2857) );
  AOI21_X1 U16090 ( .B1(n17866), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14294), .ZN(n14295) );
  OAI21_X1 U16091 ( .B1(n17883), .B2(n14296), .A(n14295), .ZN(n14297) );
  INV_X1 U16092 ( .A(n14297), .ZN(n14298) );
  OAI211_X1 U16093 ( .C1(n14302), .C2(n17860), .A(n14301), .B(n14300), .ZN(
        P2_U2983) );
  INV_X1 U16094 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n21353) );
  INV_X1 U16095 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18473) );
  INV_X1 U16096 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21714) );
  NOR2_X1 U16097 ( .A1(n18473), .A2(n21714), .ZN(n21411) );
  NAND2_X1 U16098 ( .A1(n21411), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n18447) );
  AOI22_X1 U16099 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14306) );
  AOI22_X1 U16100 ( .A1(n11145), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18331), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14305) );
  NOR2_X2 U16101 ( .A1(n14308), .A2(n14307), .ZN(n14342) );
  AOI22_X1 U16102 ( .A1(n18347), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11147), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14304) );
  AOI22_X1 U16103 ( .A1(n18326), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18055), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14303) );
  NAND4_X1 U16104 ( .A1(n14306), .A2(n14305), .A3(n14304), .A4(n14303), .ZN(
        n14316) );
  AOI22_X1 U16105 ( .A1(n18341), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18130), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14314) );
  AOI22_X1 U16106 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18332), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14313) );
  AOI22_X1 U16108 ( .A1(n18348), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14312) );
  NOR2_X2 U16109 ( .A1(n14310), .A2(n21383), .ZN(n14341) );
  AOI22_X1 U16110 ( .A1(n11144), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14311) );
  NAND4_X1 U16111 ( .A1(n14314), .A2(n14313), .A3(n14312), .A4(n14311), .ZN(
        n14315) );
  AOI22_X1 U16112 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18332), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14320) );
  AOI22_X1 U16113 ( .A1(n18348), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n18331), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14319) );
  AOI22_X1 U16114 ( .A1(n18055), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14318) );
  AOI22_X1 U16115 ( .A1(n11147), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n18326), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14317) );
  NAND4_X1 U16116 ( .A1(n14320), .A2(n14319), .A3(n14318), .A4(n14317), .ZN(
        n14326) );
  AOI22_X1 U16117 ( .A1(n11144), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14324) );
  AOI22_X1 U16118 ( .A1(n18341), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14323) );
  AOI22_X1 U16119 ( .A1(n18130), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18347), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14322) );
  AOI22_X1 U16120 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14321) );
  NAND4_X1 U16121 ( .A1(n14324), .A2(n14323), .A3(n14322), .A4(n14321), .ZN(
        n14325) );
  AOI22_X1 U16122 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14349), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14330) );
  AOI22_X1 U16123 ( .A1(n18101), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18130), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14329) );
  AOI22_X1 U16124 ( .A1(n18348), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11147), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14328) );
  AOI22_X1 U16125 ( .A1(n18326), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18055), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14327) );
  NAND4_X1 U16126 ( .A1(n14330), .A2(n14329), .A3(n14328), .A4(n14327), .ZN(
        n14336) );
  AOI22_X1 U16127 ( .A1(n14342), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14334) );
  AOI22_X1 U16128 ( .A1(n18341), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18331), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14333) );
  AOI22_X1 U16129 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14332) );
  AOI22_X1 U16130 ( .A1(n11144), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14341), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14331) );
  NAND4_X1 U16131 ( .A1(n14334), .A2(n14333), .A3(n14332), .A4(n14331), .ZN(
        n14335) );
  AOI22_X1 U16132 ( .A1(n11147), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14340) );
  AOI22_X1 U16133 ( .A1(n11145), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n14349), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14339) );
  AOI22_X1 U16134 ( .A1(n18348), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n18130), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14338) );
  AOI22_X1 U16135 ( .A1(n18326), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11175), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14337) );
  NAND4_X1 U16136 ( .A1(n14340), .A2(n14339), .A3(n14338), .A4(n14337), .ZN(
        n14348) );
  AOI22_X1 U16137 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n18101), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14346) );
  AOI22_X1 U16138 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14389), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14345) );
  AOI22_X1 U16139 ( .A1(n14341), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14342), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14344) );
  AOI22_X1 U16140 ( .A1(n11144), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14447), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14343) );
  NAND4_X1 U16141 ( .A1(n14346), .A2(n14345), .A3(n14344), .A4(n14343), .ZN(
        n14347) );
  AOI22_X1 U16142 ( .A1(n18332), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n14341), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14361) );
  AOI22_X1 U16143 ( .A1(n11144), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14360) );
  INV_X1 U16144 ( .A(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14351) );
  AOI22_X1 U16145 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18165), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14350) );
  OAI21_X1 U16146 ( .B1(n11209), .B2(n14351), .A(n14350), .ZN(n14358) );
  AOI22_X1 U16147 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14356) );
  AOI22_X1 U16148 ( .A1(n18341), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18130), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14355) );
  AOI22_X1 U16149 ( .A1(n18347), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18326), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14354) );
  AOI22_X1 U16150 ( .A1(n11147), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n18055), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14353) );
  NAND4_X1 U16151 ( .A1(n14356), .A2(n14355), .A3(n14354), .A4(n14353), .ZN(
        n14357) );
  AOI211_X1 U16152 ( .C1(n18288), .C2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n14358), .B(n14357), .ZN(n14359) );
  NAND3_X1 U16153 ( .A1(n14361), .A2(n14360), .A3(n14359), .ZN(n14571) );
  NAND2_X1 U16154 ( .A1(n14574), .A2(n14571), .ZN(n14388) );
  NOR2_X1 U16155 ( .A1(n21213), .A2(n14388), .ZN(n14387) );
  AOI22_X1 U16156 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n11144), .B1(
        P3_INSTQUEUE_REG_1__5__SCAN_IN), .B2(n18349), .ZN(n14371) );
  AOI22_X1 U16157 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18341), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14370) );
  AOI22_X1 U16158 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18165), .B1(
        P3_INSTQUEUE_REG_15__5__SCAN_IN), .B2(n18326), .ZN(n14362) );
  OAI21_X1 U16159 ( .B1(n14374), .B2(n18048), .A(n14362), .ZN(n14368) );
  AOI22_X1 U16160 ( .A1(n18332), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14366) );
  AOI22_X1 U16161 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18342), .B1(
        P3_INSTQUEUE_REG_3__5__SCAN_IN), .B2(n18347), .ZN(n14365) );
  AOI22_X1 U16162 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__5__SCAN_IN), .B2(n18350), .ZN(n14364) );
  INV_X4 U16163 ( .A(n18216), .ZN(n18130) );
  AOI22_X1 U16164 ( .A1(n18348), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__5__SCAN_IN), .B2(n18130), .ZN(n14363) );
  NAND4_X1 U16165 ( .A1(n14366), .A2(n14365), .A3(n14364), .A4(n14363), .ZN(
        n14367) );
  AOI211_X1 U16166 ( .C1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .C2(n11175), .A(
        n14368), .B(n14367), .ZN(n14369) );
  NAND3_X1 U16167 ( .A1(n14371), .A2(n14370), .A3(n14369), .ZN(n14570) );
  NAND2_X1 U16168 ( .A1(n14387), .A2(n14570), .ZN(n14385) );
  AOI22_X1 U16169 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18288), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14383) );
  AOI22_X1 U16170 ( .A1(n18130), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n18347), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14382) );
  AOI22_X1 U16171 ( .A1(n18326), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n18055), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14373) );
  OAI21_X1 U16172 ( .B1(n14374), .B2(n18184), .A(n14373), .ZN(n14380) );
  AOI22_X1 U16173 ( .A1(n11144), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14378) );
  AOI22_X1 U16174 ( .A1(n18332), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18331), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14377) );
  AOI22_X1 U16175 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14376) );
  AOI22_X1 U16176 ( .A1(n18341), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14375) );
  NAND4_X1 U16177 ( .A1(n14378), .A2(n14377), .A3(n14376), .A4(n14375), .ZN(
        n14379) );
  AOI211_X1 U16178 ( .C1(n14341), .C2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A(
        n14380), .B(n14379), .ZN(n14381) );
  INV_X1 U16179 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21752) );
  INV_X1 U16180 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18405) );
  NAND2_X1 U16181 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n21513) );
  INV_X1 U16182 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21762) );
  NOR3_X1 U16183 ( .A1(n21513), .A2(n21763), .A3(n21762), .ZN(n21522) );
  NAND2_X1 U16184 ( .A1(n21522), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n21538) );
  INV_X1 U16185 ( .A(n21538), .ZN(n21541) );
  NAND2_X1 U16186 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n21541), .ZN(
        n21561) );
  NOR2_X1 U16187 ( .A1(n18405), .A2(n21561), .ZN(n21725) );
  AOI21_X1 U16188 ( .B1(n21653), .B2(n14384), .A(n18548), .ZN(n14415) );
  INV_X1 U16189 ( .A(n21204), .ZN(n14568) );
  XNOR2_X1 U16190 ( .A(n14568), .B(n14385), .ZN(n14386) );
  NAND2_X1 U16191 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n14386), .ZN(
        n14414) );
  XOR2_X1 U16192 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n14386), .Z(
        n18690) );
  XOR2_X1 U16193 ( .A(n14570), .B(n14387), .Z(n14410) );
  INV_X1 U16194 ( .A(n21213), .ZN(n14584) );
  XNOR2_X1 U16195 ( .A(n14584), .B(n14388), .ZN(n14408) );
  XOR2_X1 U16196 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n14408), .Z(
        n18709) );
  NAND2_X1 U16197 ( .A1(n14577), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14402) );
  XNOR2_X1 U16198 ( .A(n21337), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18746) );
  AOI22_X1 U16199 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18313), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14394) );
  AOI22_X1 U16200 ( .A1(n18101), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18331), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14393) );
  AOI22_X1 U16201 ( .A1(n18130), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n18326), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14392) );
  AOI22_X1 U16202 ( .A1(n11147), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n18055), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14391) );
  NAND4_X1 U16203 ( .A1(n14394), .A2(n14393), .A3(n14392), .A4(n14391), .ZN(
        n14401) );
  AOI22_X1 U16204 ( .A1(n14341), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14342), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14399) );
  AOI22_X1 U16205 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14349), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14398) );
  AOI22_X1 U16206 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18288), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14397) );
  AOI22_X1 U16207 ( .A1(n11144), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14396) );
  NAND4_X1 U16208 ( .A1(n14399), .A2(n14398), .A3(n14397), .A4(n14396), .ZN(
        n14400) );
  NOR2_X1 U16209 ( .A1(n21350), .A2(n21508), .ZN(n18752) );
  NAND2_X1 U16210 ( .A1(n18746), .A2(n18752), .ZN(n18745) );
  NAND2_X1 U16211 ( .A1(n14402), .A2(n18745), .ZN(n18738) );
  NAND2_X1 U16212 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n14404), .ZN(
        n14405) );
  NAND2_X1 U16213 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n14406), .ZN(
        n14407) );
  INV_X1 U16214 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21447) );
  XNOR2_X1 U16215 ( .A(n21447), .B(n14406), .ZN(n18728) );
  XOR2_X1 U16216 ( .A(n14571), .B(n14574), .Z(n18727) );
  NAND2_X1 U16217 ( .A1(n18728), .A2(n18727), .ZN(n18726) );
  NAND2_X1 U16218 ( .A1(n14407), .A2(n18726), .ZN(n18708) );
  NAND2_X1 U16219 ( .A1(n18709), .A2(n18708), .ZN(n18707) );
  NAND2_X1 U16220 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n14408), .ZN(
        n14409) );
  NAND2_X1 U16221 ( .A1(n14410), .A2(n14412), .ZN(n14413) );
  NAND2_X1 U16222 ( .A1(n14413), .A2(n18698), .ZN(n18689) );
  NAND2_X1 U16223 ( .A1(n18690), .A2(n18689), .ZN(n18688) );
  NAND2_X1 U16224 ( .A1(n14415), .A2(n18401), .ZN(n14417) );
  AOI22_X1 U16225 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21668), .B1(
        n18548), .B2(n21495), .ZN(n18666) );
  NAND2_X1 U16226 ( .A1(n21725), .A2(n18639), .ZN(n14420) );
  INV_X1 U16227 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21798) );
  INV_X1 U16228 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n21772) );
  NAND2_X1 U16229 ( .A1(n21798), .A2(n21772), .ZN(n18646) );
  NOR3_X1 U16230 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(n18646), .ZN(n18437) );
  INV_X1 U16231 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n21543) );
  NAND2_X1 U16232 ( .A1(n18437), .A2(n21543), .ZN(n18403) );
  OR3_X1 U16233 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(n18403), .ZN(n14419) );
  INV_X1 U16234 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21750) );
  NAND2_X1 U16235 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21398) );
  INV_X1 U16236 ( .A(n21398), .ZN(n21730) );
  NAND2_X1 U16237 ( .A1(n14421), .A2(n14420), .ZN(n18415) );
  NAND2_X1 U16238 ( .A1(n21730), .A2(n18415), .ZN(n18392) );
  NAND2_X1 U16239 ( .A1(n14422), .A2(n18392), .ZN(n18376) );
  NAND2_X1 U16240 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18376), .ZN(
        n18471) );
  INV_X1 U16241 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18393) );
  NOR2_X1 U16242 ( .A1(n21398), .A2(n18393), .ZN(n21403) );
  INV_X1 U16243 ( .A(n18447), .ZN(n14423) );
  NAND2_X1 U16244 ( .A1(n21403), .A2(n14423), .ZN(n21573) );
  NAND2_X1 U16245 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21692) );
  NOR2_X1 U16246 ( .A1(n21573), .A2(n21692), .ZN(n18534) );
  NAND2_X1 U16247 ( .A1(n21668), .A2(n18393), .ZN(n18394) );
  NOR2_X1 U16248 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18446), .ZN(
        n18494) );
  INV_X1 U16249 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18496) );
  AOI22_X1 U16250 ( .A1(n18534), .A2(n18415), .B1(n18494), .B2(n18496), .ZN(
        n14424) );
  NOR2_X2 U16251 ( .A1(n18445), .A2(n14424), .ZN(n18522) );
  INV_X1 U16252 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n21696) );
  INV_X1 U16253 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21598) );
  OR2_X1 U16254 ( .A1(n18548), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14425) );
  INV_X1 U16255 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n21599) );
  INV_X1 U16256 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21665) );
  NAND2_X1 U16257 ( .A1(n14430), .A2(n21665), .ZN(n21674) );
  INV_X1 U16258 ( .A(n21674), .ZN(n18538) );
  NOR2_X1 U16259 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18548), .ZN(
        n18536) );
  INV_X1 U16260 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n21641) );
  NOR2_X1 U16261 ( .A1(n14430), .A2(n21665), .ZN(n18537) );
  NOR2_X1 U16262 ( .A1(n21654), .A2(n21641), .ZN(n14429) );
  NOR2_X1 U16263 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18569), .ZN(
        n18568) );
  AOI22_X1 U16264 ( .A1(n14430), .A2(n18568), .B1(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n14429), .ZN(n14431) );
  XOR2_X1 U16265 ( .A(n21353), .B(n14431), .Z(n14612) );
  INV_X1 U16266 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21834) );
  OAI22_X1 U16267 ( .A1(n21371), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n21834), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14437) );
  AOI22_X1 U16268 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n21827), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n21382), .ZN(n14467) );
  AND2_X1 U16269 ( .A1(n14468), .A2(n14467), .ZN(n14432) );
  OAI22_X1 U16270 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21838), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n14434), .ZN(n14439) );
  NOR2_X1 U16271 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21838), .ZN(
        n14435) );
  NAND2_X1 U16272 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n14434), .ZN(
        n14440) );
  AOI22_X1 U16273 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n14439), .B1(
        n14435), .B2(n14440), .ZN(n14444) );
  AOI21_X1 U16274 ( .B1(n17368), .B2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n14468), .ZN(n14538) );
  AND2_X1 U16275 ( .A1(n14467), .A2(n14538), .ZN(n14443) );
  NAND2_X1 U16276 ( .A1(n14438), .A2(n14437), .ZN(n14436) );
  OAI211_X1 U16277 ( .C1(n14438), .C2(n14437), .A(n14444), .B(n14436), .ZN(
        n14470) );
  INV_X1 U16278 ( .A(n14470), .ZN(n14539) );
  AOI21_X1 U16279 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n14440), .A(
        n14439), .ZN(n14441) );
  INV_X1 U16280 ( .A(n14469), .ZN(n14442) );
  AOI22_X1 U16281 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n18332), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14456) );
  AOI22_X1 U16282 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18288), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14455) );
  AOI22_X1 U16283 ( .A1(n18326), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11175), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14446) );
  OAI21_X1 U16284 ( .B1(n11209), .B2(n18048), .A(n14446), .ZN(n14453) );
  AOI22_X1 U16285 ( .A1(n11144), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14451) );
  AOI22_X1 U16286 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n18130), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14450) );
  AOI22_X1 U16287 ( .A1(n18347), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n18165), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14449) );
  AOI22_X1 U16288 ( .A1(n11145), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14448) );
  NAND4_X1 U16289 ( .A1(n14451), .A2(n14450), .A3(n14449), .A4(n14448), .ZN(
        n14452) );
  AOI211_X1 U16290 ( .C1(n11147), .C2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n14453), .B(n14452), .ZN(n14454) );
  NAND3_X1 U16291 ( .A1(n14456), .A2(n14455), .A3(n14454), .ZN(n21231) );
  AOI22_X1 U16292 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14466) );
  AOI22_X1 U16293 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11144), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14465) );
  AOI22_X1 U16294 ( .A1(n18350), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18347), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14457) );
  OAI21_X1 U16295 ( .B1(n11209), .B2(n18195), .A(n14457), .ZN(n14463) );
  AOI22_X1 U16296 ( .A1(n18288), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n18130), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14461) );
  AOI22_X1 U16297 ( .A1(n18342), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n18165), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14460) );
  AOI22_X1 U16298 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18326), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14459) );
  AOI22_X1 U16299 ( .A1(n11147), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n14390), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14458) );
  NAND4_X1 U16300 ( .A1(n14461), .A2(n14460), .A3(n14459), .A4(n14458), .ZN(
        n14462) );
  AOI211_X1 U16301 ( .C1(n18332), .C2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A(
        n14463), .B(n14462), .ZN(n14464) );
  XNOR2_X1 U16302 ( .A(n14468), .B(n14467), .ZN(n14471) );
  AOI22_X1 U16303 ( .A1(n11144), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n18347), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14475) );
  AOI22_X1 U16304 ( .A1(n18342), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n18165), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14474) );
  AOI22_X1 U16305 ( .A1(n11145), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11147), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14473) );
  AOI22_X1 U16306 ( .A1(n18326), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n18055), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14472) );
  NAND4_X1 U16307 ( .A1(n14475), .A2(n14474), .A3(n14473), .A4(n14472), .ZN(
        n14481) );
  AOI22_X1 U16308 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n18130), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14479) );
  AOI22_X1 U16309 ( .A1(n18332), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14478) );
  AOI22_X1 U16310 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n18288), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14477) );
  AOI22_X1 U16311 ( .A1(n18341), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14476) );
  NAND4_X1 U16312 ( .A1(n14479), .A2(n14478), .A3(n14477), .A4(n14476), .ZN(
        n14480) );
  INV_X2 U16313 ( .A(n18837), .ZN(n18840) );
  OAI211_X1 U16314 ( .C1(P3_STATE_REG_2__SCAN_IN), .C2(P3_STATE_REG_1__SCAN_IN), .A(n18840), .B(n22345), .ZN(n20735) );
  OAI211_X1 U16315 ( .C1(n19553), .C2(n20741), .A(n14565), .B(n20735), .ZN(
        n14482) );
  NAND2_X1 U16316 ( .A1(n22352), .A2(n14482), .ZN(n21814) );
  NOR3_X1 U16317 ( .A1(n14544), .A2(n21817), .A3(n21814), .ZN(n14537) );
  AOI22_X1 U16318 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11144), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14492) );
  AOI22_X1 U16319 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14342), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14491) );
  INV_X1 U16320 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18296) );
  AOI22_X1 U16321 ( .A1(n18332), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14483) );
  OAI21_X1 U16322 ( .B1(n11209), .B2(n18296), .A(n14483), .ZN(n14489) );
  AOI22_X1 U16323 ( .A1(n18288), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n18165), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14487) );
  AOI22_X1 U16324 ( .A1(n18130), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14486) );
  AOI22_X1 U16325 ( .A1(n18342), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11147), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14485) );
  AOI22_X1 U16326 ( .A1(n18326), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14390), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14484) );
  NAND4_X1 U16327 ( .A1(n14487), .A2(n14486), .A3(n14485), .A4(n14484), .ZN(
        n14488) );
  AOI211_X1 U16328 ( .C1(n11164), .C2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n14489), .B(n14488), .ZN(n14490) );
  NAND3_X1 U16329 ( .A1(n14492), .A2(n14491), .A3(n14490), .ZN(n14555) );
  AOI22_X1 U16330 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14496) );
  AOI22_X1 U16331 ( .A1(n18288), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n14342), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14495) );
  AOI22_X1 U16332 ( .A1(n18165), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18326), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14494) );
  AOI22_X1 U16333 ( .A1(n11147), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11175), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14493) );
  NAND4_X1 U16334 ( .A1(n14496), .A2(n14495), .A3(n14494), .A4(n14493), .ZN(
        n14502) );
  AOI22_X1 U16335 ( .A1(n18332), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14500) );
  AOI22_X1 U16336 ( .A1(n18130), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11144), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14499) );
  AOI22_X1 U16337 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n18341), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14498) );
  AOI22_X1 U16338 ( .A1(n18342), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14497) );
  NAND4_X1 U16339 ( .A1(n14500), .A2(n14499), .A3(n14498), .A4(n14497), .ZN(
        n14501) );
  AOI22_X1 U16340 ( .A1(n18130), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14512) );
  AOI22_X1 U16341 ( .A1(n18288), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18165), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14511) );
  AOI22_X1 U16342 ( .A1(n18332), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14503) );
  OAI21_X1 U16343 ( .B1(n11209), .B2(n18281), .A(n14503), .ZN(n14509) );
  AOI22_X1 U16344 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n18347), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14507) );
  AOI22_X1 U16345 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11144), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14506) );
  AOI22_X1 U16346 ( .A1(n11145), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n18326), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14505) );
  AOI22_X1 U16347 ( .A1(n11147), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11175), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14504) );
  NAND4_X1 U16348 ( .A1(n14507), .A2(n14506), .A3(n14505), .A4(n14504), .ZN(
        n14508) );
  NAND2_X1 U16349 ( .A1(n20736), .A2(n20741), .ZN(n14513) );
  NAND2_X1 U16350 ( .A1(n19553), .A2(n14513), .ZN(n14558) );
  AOI22_X1 U16351 ( .A1(n18130), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14517) );
  AOI22_X1 U16352 ( .A1(n11145), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18165), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14516) );
  AOI22_X1 U16353 ( .A1(n18332), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11147), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14515) );
  AOI22_X1 U16354 ( .A1(n18326), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18055), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14514) );
  NAND4_X1 U16355 ( .A1(n14517), .A2(n14516), .A3(n14515), .A4(n14514), .ZN(
        n14523) );
  AOI22_X1 U16356 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18234), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14521) );
  AOI22_X1 U16357 ( .A1(n18288), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11164), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14520) );
  AOI22_X1 U16358 ( .A1(n11144), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14519) );
  AOI22_X1 U16359 ( .A1(n18342), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14342), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14518) );
  NAND4_X1 U16360 ( .A1(n14521), .A2(n14520), .A3(n14519), .A4(n14518), .ZN(
        n14522) );
  AOI22_X1 U16361 ( .A1(n18342), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18165), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14524) );
  OAI21_X1 U16362 ( .B1(n11209), .B2(n18184), .A(n14524), .ZN(n14529) );
  AOI22_X1 U16363 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11144), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14528) );
  AOI22_X1 U16364 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n18332), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14527) );
  AOI22_X1 U16365 ( .A1(n18347), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11147), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14526) );
  AOI22_X1 U16366 ( .A1(n18326), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18055), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14525) );
  NAND3_X1 U16367 ( .A1(n19511), .A2(n20736), .A3(n21267), .ZN(n14551) );
  NAND2_X1 U16368 ( .A1(n21231), .A2(n21232), .ZN(n14559) );
  NAND2_X1 U16369 ( .A1(n21374), .A2(n14532), .ZN(n14546) );
  NAND2_X1 U16370 ( .A1(n19430), .A2(n21232), .ZN(n14549) );
  OAI211_X1 U16371 ( .C1(n19470), .C2(n17367), .A(n14545), .B(n14549), .ZN(
        n14535) );
  NOR2_X1 U16372 ( .A1(n20736), .A2(n20741), .ZN(n14533) );
  NAND2_X1 U16373 ( .A1(n21267), .A2(n21171), .ZN(n21170) );
  NAND2_X1 U16374 ( .A1(n14533), .A2(n21170), .ZN(n14554) );
  INV_X1 U16375 ( .A(n14554), .ZN(n14534) );
  AOI221_X1 U16376 ( .B1(n14558), .B2(n14546), .C1(n14535), .C2(n14546), .A(
        n14534), .ZN(n14536) );
  OAI221_X1 U16377 ( .B1(n14543), .B2(n18807), .C1(n14543), .C2(n21171), .A(
        n14536), .ZN(n15966) );
  AOI211_X1 U16378 ( .C1(n21813), .C2(n14544), .A(n14537), .B(n15966), .ZN(
        n14542) );
  AOI21_X1 U16379 ( .B1(n14539), .B2(n14538), .A(n21817), .ZN(n14540) );
  INV_X1 U16380 ( .A(n14540), .ZN(n21808) );
  INV_X1 U16381 ( .A(n21374), .ZN(n14560) );
  NAND2_X1 U16382 ( .A1(n19553), .A2(n19511), .ZN(n21358) );
  NOR2_X1 U16383 ( .A1(n20741), .A2(n18807), .ZN(n21166) );
  AND2_X1 U16384 ( .A1(n21267), .A2(n21166), .ZN(n14547) );
  INV_X1 U16385 ( .A(n14545), .ZN(n14563) );
  NAND2_X1 U16386 ( .A1(n14548), .A2(n14555), .ZN(n21359) );
  NAND4_X1 U16387 ( .A1(n19553), .A2(n20736), .A3(n21359), .A4(n14549), .ZN(
        n14550) );
  OAI221_X1 U16388 ( .B1(n19470), .B2(n21267), .C1(n19470), .C2(n14559), .A(
        n14550), .ZN(n14557) );
  OAI21_X1 U16389 ( .B1(n14552), .B2(n19511), .A(n14551), .ZN(n14553) );
  OAI211_X1 U16390 ( .C1(n21171), .C2(n14555), .A(n14554), .B(n14553), .ZN(
        n14556) );
  NOR2_X4 U16391 ( .A1(n15964), .A2(n14564), .ZN(n21795) );
  NAND2_X1 U16392 ( .A1(n14563), .A2(n20741), .ZN(n21357) );
  NAND2_X1 U16393 ( .A1(n14612), .A2(n21801), .ZN(n14610) );
  INV_X1 U16394 ( .A(n18534), .ZN(n14600) );
  INV_X1 U16395 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21544) );
  NAND2_X1 U16396 ( .A1(n21732), .A2(n21541), .ZN(n18612) );
  NAND2_X1 U16397 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n21682), .ZN(
        n18510) );
  NOR2_X1 U16398 ( .A1(n21598), .A2(n18510), .ZN(n18509) );
  NAND2_X1 U16399 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18509), .ZN(
        n21631) );
  NAND2_X1 U16400 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21636) );
  NOR2_X1 U16401 ( .A1(n21636), .A2(n21641), .ZN(n18579) );
  INV_X1 U16402 ( .A(n18579), .ZN(n21644) );
  NOR2_X1 U16403 ( .A1(n21631), .A2(n21644), .ZN(n21627) );
  NAND2_X1 U16404 ( .A1(n21627), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14566) );
  XNOR2_X1 U16405 ( .A(n21353), .B(n14566), .ZN(n14614) );
  NAND2_X1 U16406 ( .A1(n21809), .A2(n21653), .ZN(n21731) );
  INV_X1 U16407 ( .A(n21350), .ZN(n14573) );
  INV_X1 U16408 ( .A(n14571), .ZN(n21217) );
  NOR2_X1 U16409 ( .A1(n14572), .A2(n21217), .ZN(n14583) );
  NAND2_X1 U16410 ( .A1(n14584), .A2(n14583), .ZN(n14569) );
  INV_X1 U16411 ( .A(n14570), .ZN(n21208) );
  NOR2_X1 U16412 ( .A1(n14569), .A2(n21208), .ZN(n14588) );
  NAND2_X1 U16413 ( .A1(n14568), .A2(n14588), .ZN(n14592) );
  NOR2_X1 U16414 ( .A1(n14592), .A2(n21653), .ZN(n14598) );
  INV_X1 U16415 ( .A(n14598), .ZN(n14593) );
  INV_X1 U16416 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21470) );
  XOR2_X1 U16417 ( .A(n14570), .B(n14569), .Z(n14586) );
  NOR2_X1 U16418 ( .A1(n21470), .A2(n14586), .ZN(n14587) );
  XNOR2_X1 U16419 ( .A(n14571), .B(n14572), .ZN(n14580) );
  AND2_X1 U16420 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n14580), .ZN(
        n14581) );
  AOI21_X1 U16421 ( .B1(n14574), .B2(n14573), .A(n14572), .ZN(n14575) );
  INV_X1 U16422 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21444) );
  NOR2_X1 U16423 ( .A1(n14575), .A2(n21444), .ZN(n14579) );
  XOR2_X1 U16424 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n14575), .Z(
        n18736) );
  NOR2_X1 U16425 ( .A1(n14577), .A2(n21508), .ZN(n14578) );
  NAND3_X1 U16426 ( .A1(n21350), .A2(n14577), .A3(n21508), .ZN(n14576) );
  OAI221_X1 U16427 ( .B1(n14578), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n21350), .C2(n14577), .A(n14576), .ZN(n18735) );
  NOR2_X1 U16428 ( .A1(n18736), .A2(n18735), .ZN(n18734) );
  XOR2_X1 U16429 ( .A(n21447), .B(n14580), .Z(n18724) );
  NOR2_X1 U16430 ( .A1(n18725), .A2(n18724), .ZN(n18723) );
  INV_X1 U16431 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n21463) );
  NOR2_X1 U16432 ( .A1(n14582), .A2(n21463), .ZN(n14585) );
  XNOR2_X1 U16433 ( .A(n14584), .B(n14583), .ZN(n18711) );
  XOR2_X1 U16434 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n14586), .Z(
        n18701) );
  NOR2_X1 U16435 ( .A1(n18702), .A2(n18701), .ZN(n18700) );
  XOR2_X1 U16436 ( .A(n21204), .B(n14588), .Z(n14590) );
  NOR2_X1 U16437 ( .A1(n14589), .A2(n14590), .ZN(n14591) );
  INV_X1 U16438 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21787) );
  XNOR2_X1 U16439 ( .A(n21653), .B(n14592), .ZN(n14595) );
  NAND2_X1 U16440 ( .A1(n14594), .A2(n14595), .ZN(n18676) );
  NAND2_X1 U16441 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n18676), .ZN(
        n14597) );
  NOR2_X1 U16442 ( .A1(n14593), .A2(n14597), .ZN(n14599) );
  OR2_X1 U16443 ( .A1(n14595), .A2(n14594), .ZN(n18677) );
  OAI21_X1 U16444 ( .B1(n14598), .B2(n14597), .A(n18677), .ZN(n14596) );
  NAND2_X1 U16445 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18611), .ZN(
        n21555) );
  NOR2_X1 U16446 ( .A1(n21599), .A2(n18501), .ZN(n21635) );
  INV_X1 U16447 ( .A(n21635), .ZN(n21605) );
  INV_X1 U16448 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21786) );
  NOR3_X1 U16449 ( .A1(n21495), .A2(n21787), .A3(n21786), .ZN(n21505) );
  INV_X1 U16450 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21443) );
  OAI21_X1 U16451 ( .B1(n21508), .B2(n21443), .A(n21444), .ZN(n21446) );
  INV_X1 U16452 ( .A(n21446), .ZN(n21448) );
  NAND3_X1 U16453 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21480) );
  NOR2_X1 U16454 ( .A1(n21448), .A2(n21480), .ZN(n21468) );
  NAND2_X1 U16455 ( .A1(n21505), .A2(n21468), .ZN(n21510) );
  NOR2_X1 U16456 ( .A1(n21561), .A2(n21510), .ZN(n21557) );
  NAND3_X1 U16457 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21730), .A3(
        n21557), .ZN(n21735) );
  NOR2_X1 U16458 ( .A1(n21812), .A2(n21735), .ZN(n21401) );
  NOR2_X1 U16459 ( .A1(n18393), .A2(n18447), .ZN(n14601) );
  AOI21_X1 U16460 ( .B1(n21576), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n21776), .ZN(n21399) );
  INV_X1 U16461 ( .A(n21399), .ZN(n21445) );
  NOR3_X1 U16462 ( .A1(n21444), .A2(n21443), .A3(n21480), .ZN(n21466) );
  NAND2_X1 U16463 ( .A1(n21505), .A2(n21466), .ZN(n21775) );
  INV_X1 U16464 ( .A(n21775), .ZN(n21540) );
  NAND2_X1 U16465 ( .A1(n21725), .A2(n21540), .ZN(n21727) );
  NOR2_X1 U16466 ( .A1(n21573), .A2(n21727), .ZN(n21583) );
  AOI22_X1 U16467 ( .A1(n21401), .A2(n14601), .B1(n21445), .B2(n21583), .ZN(
        n21633) );
  NAND3_X1 U16468 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21588) );
  NOR3_X1 U16469 ( .A1(n21588), .A2(n21598), .A3(n21599), .ZN(n21613) );
  INV_X1 U16470 ( .A(n21613), .ZN(n21632) );
  NOR4_X1 U16471 ( .A1(n21633), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n21632), .A4(n21644), .ZN(n14602) );
  NAND2_X1 U16472 ( .A1(n21583), .A2(n21613), .ZN(n21657) );
  INV_X1 U16473 ( .A(n21573), .ZN(n14603) );
  NOR2_X1 U16474 ( .A1(n21508), .A2(n21727), .ZN(n21556) );
  NAND2_X1 U16475 ( .A1(n14603), .A2(n21556), .ZN(n21575) );
  NOR2_X1 U16476 ( .A1(n21632), .A2(n21575), .ZN(n14605) );
  NOR3_X1 U16477 ( .A1(n18393), .A2(n18447), .A3(n21735), .ZN(n21585) );
  AOI21_X1 U16478 ( .B1(n21613), .B2(n21585), .A(n21812), .ZN(n14604) );
  INV_X1 U16479 ( .A(n14604), .ZN(n21615) );
  OAI221_X1 U16480 ( .B1(n21790), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), 
        .C1(n21790), .C2(n14605), .A(n21615), .ZN(n21660) );
  AOI221_X1 U16481 ( .B1(n21636), .B2(n21776), .C1(n21657), .C2(n21776), .A(
        n21660), .ZN(n21629) );
  OAI211_X1 U16482 ( .C1(n21756), .C2(n18579), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n21629), .ZN(n21648) );
  INV_X1 U16483 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n21855) );
  NAND2_X1 U16484 ( .A1(n21855), .A2(n20744), .ZN(n18370) );
  OR2_X1 U16485 ( .A1(n18370), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n17758) );
  NAND2_X1 U16486 ( .A1(n21774), .A2(P3_REIP_REG_31__SCAN_IN), .ZN(n14618) );
  NAND2_X1 U16487 ( .A1(n14610), .A2(n14609), .ZN(P3_U2831) );
  INV_X1 U16488 ( .A(n21813), .ZN(n14611) );
  NAND2_X1 U16489 ( .A1(n14612), .A2(n18661), .ZN(n14631) );
  NAND2_X1 U16490 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18667) );
  INV_X1 U16491 ( .A(n18667), .ZN(n18656) );
  NAND4_X1 U16492 ( .A1(n18656), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n18619) );
  NAND2_X1 U16493 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18386) );
  INV_X1 U16494 ( .A(n18386), .ZN(n14615) );
  INV_X1 U16495 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14617) );
  NAND2_X1 U16496 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n18591), .ZN(
        n18570) );
  INV_X1 U16497 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n21147) );
  NAND2_X1 U16498 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18371) );
  NAND2_X1 U16499 ( .A1(n21855), .A2(n18371), .ZN(n20674) );
  INV_X1 U16500 ( .A(n14618), .ZN(n14625) );
  NAND3_X1 U16501 ( .A1(n18451), .A2(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18488) );
  NOR2_X1 U16502 ( .A1(n21041), .A2(n18488), .ZN(n18504) );
  NAND3_X1 U16503 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A3(n18504), .ZN(n18559) );
  NOR2_X1 U16504 ( .A1(n11362), .A2(n18559), .ZN(n18550) );
  NAND3_X1 U16505 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(n18550), .ZN(n18582) );
  NOR2_X1 U16506 ( .A1(n18592), .A2(n18582), .ZN(n14620) );
  INV_X1 U16507 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20757) );
  INV_X1 U16508 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n21862) );
  NAND2_X1 U16509 ( .A1(n21862), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18754) );
  NAND2_X1 U16510 ( .A1(n21354), .A2(n20744), .ZN(n21863) );
  AOI21_X1 U16511 ( .B1(n18371), .B2(n21863), .A(n21367), .ZN(n19317) );
  NAND2_X1 U16512 ( .A1(n14620), .A2(n18549), .ZN(n18574) );
  XNOR2_X1 U16513 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14623) );
  NOR2_X1 U16514 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18529), .ZN(
        n18594) );
  OAI21_X1 U16515 ( .B1(n19551), .B2(n14620), .A(n18753), .ZN(n14621) );
  AOI21_X1 U16516 ( .B1(n14619), .B2(n11315), .A(n14621), .ZN(n14622) );
  INV_X1 U16517 ( .A(n14622), .ZN(n18584) );
  NOR2_X1 U16518 ( .A1(n18594), .A2(n18584), .ZN(n18573) );
  OAI22_X1 U16519 ( .A1(n18574), .A2(n14623), .B1(n18573), .B2(n21147), .ZN(
        n14624) );
  AOI211_X1 U16520 ( .C1(n20817), .C2(n18593), .A(n14625), .B(n14624), .ZN(
        n14626) );
  INV_X1 U16521 ( .A(n14626), .ZN(n14627) );
  NAND2_X1 U16522 ( .A1(n14631), .A2(n14630), .ZN(P3_U2799) );
  NOR2_X1 U16523 ( .A1(P2_BE_N_REG_3__SCAN_IN), .A2(P2_BE_N_REG_2__SCAN_IN), 
        .ZN(n14633) );
  NOR4_X1 U16524 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_0__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n14632) );
  NAND4_X1 U16525 ( .A1(n14633), .A2(P2_M_IO_N_REG_SCAN_IN), .A3(
        P2_W_R_N_REG_SCAN_IN), .A4(n14632), .ZN(n14656) );
  NOR4_X1 U16526 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n14637) );
  NOR4_X1 U16527 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n14636) );
  NOR4_X1 U16528 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n14635) );
  NOR4_X1 U16529 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n14634) );
  AND4_X1 U16530 ( .A1(n14637), .A2(n14636), .A3(n14635), .A4(n14634), .ZN(
        n14643) );
  NOR4_X1 U16531 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n14641) );
  NOR4_X1 U16532 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n14640) );
  NOR4_X1 U16533 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n14639) );
  INV_X1 U16534 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n14638) );
  AND4_X1 U16535 ( .A1(n14641), .A2(n14640), .A3(n14639), .A4(n14638), .ZN(
        n14642) );
  NAND2_X1 U16536 ( .A1(n14643), .A2(n14642), .ZN(n14644) );
  INV_X1 U16537 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20669) );
  NOR3_X1 U16538 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n20669), .ZN(n14646) );
  NOR4_X1 U16539 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(P1_ADS_N_REG_SCAN_IN), .A3(
        P1_BE_N_REG_1__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n14645) );
  NAND4_X1 U16540 ( .A1(P1_M_IO_N_REG_SCAN_IN), .A2(n15987), .A3(n14646), .A4(
        n14645), .ZN(U214) );
  NOR4_X1 U16541 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n14650) );
  NOR4_X1 U16542 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n14649) );
  NOR4_X1 U16543 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n14648) );
  NOR4_X1 U16544 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n14647) );
  NAND4_X1 U16545 ( .A1(n14650), .A2(n14649), .A3(n14648), .A4(n14647), .ZN(
        n14655) );
  NOR4_X1 U16546 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n14653) );
  NOR4_X1 U16547 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n14652) );
  NOR4_X1 U16548 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n14651) );
  NAND4_X1 U16549 ( .A1(n14653), .A2(n14652), .A3(n14651), .A4(n20360), .ZN(
        n14654) );
  OAI21_X4 U16550 ( .B1(n14655), .B2(n14654), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n15700) );
  NOR2_X1 U16551 ( .A1(n15700), .A2(n14656), .ZN(n20601) );
  NAND2_X1 U16552 ( .A1(n20601), .A2(U214), .ZN(U212) );
  INV_X1 U16553 ( .A(n18852), .ZN(n14658) );
  INV_X1 U16554 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n14657) );
  OAI22_X1 U16555 ( .A1(n14658), .A2(n14657), .B1(n14661), .B2(n19270), .ZN(
        P2_U2816) );
  NOR2_X1 U16556 ( .A1(n14659), .A2(n12471), .ZN(n18880) );
  INV_X1 U16557 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n14660) );
  INV_X1 U16558 ( .A(n14675), .ZN(n14674) );
  OAI211_X1 U16559 ( .C1(n18880), .C2(n14660), .A(n14674), .B(n14661), .ZN(
        P2_U2814) );
  INV_X1 U16560 ( .A(n14661), .ZN(n14662) );
  OAI21_X1 U16561 ( .B1(P2_READREQUEST_REG_SCAN_IN), .B2(n14662), .A(n18852), 
        .ZN(n14663) );
  OAI21_X1 U16562 ( .B1(n14664), .B2(n18852), .A(n14663), .ZN(P2_U3612) );
  OAI21_X1 U16563 ( .B1(n18859), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n14665), .ZN(n19177) );
  INV_X1 U16564 ( .A(n19177), .ZN(n14669) );
  OAI21_X1 U16565 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n14667), .A(
        n14666), .ZN(n19188) );
  NAND2_X1 U16566 ( .A1(n19213), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n19185) );
  OAI21_X1 U16567 ( .B1(n17860), .B2(n19188), .A(n19185), .ZN(n14668) );
  AOI21_X1 U16568 ( .B1(n17879), .B2(n14669), .A(n14668), .ZN(n14672) );
  OAI21_X1 U16569 ( .B1(n17866), .B2(n14670), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14671) );
  OAI211_X1 U16570 ( .C1(n17865), .C2(n18858), .A(n14672), .B(n14671), .ZN(
        P2_U3014) );
  INV_X1 U16571 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n14677) );
  NAND3_X1 U16572 ( .A1(n14675), .A2(n13896), .A3(n19281), .ZN(n14781) );
  AOI22_X1 U16573 ( .A1(n19752), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n15700), .ZN(n20195) );
  NOR2_X1 U16574 ( .A1(n14781), .A2(n20195), .ZN(n14760) );
  AOI21_X1 U16575 ( .B1(n14775), .B2(P2_EAX_REG_17__SCAN_IN), .A(n14760), .ZN(
        n14676) );
  OAI21_X1 U16576 ( .B1(n14749), .B2(n14677), .A(n14676), .ZN(P2_U2953) );
  INV_X1 U16577 ( .A(P2_LWORD_REG_6__SCAN_IN), .ZN(n14679) );
  INV_X1 U16578 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n20615) );
  INV_X1 U16579 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n21207) );
  AOI22_X1 U16580 ( .A1(n19752), .A2(n20615), .B1(n21207), .B2(n15700), .ZN(
        n19961) );
  INV_X1 U16581 ( .A(n19961), .ZN(n19969) );
  NOR2_X1 U16582 ( .A1(n14781), .A2(n19969), .ZN(n14697) );
  AOI21_X1 U16583 ( .B1(n14775), .B2(P2_EAX_REG_6__SCAN_IN), .A(n14697), .ZN(
        n14678) );
  OAI21_X1 U16584 ( .B1(n14749), .B2(n14679), .A(n14678), .ZN(P2_U2973) );
  INV_X1 U16585 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n14681) );
  AOI22_X1 U16586 ( .A1(n19752), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n15700), .ZN(n20019) );
  NOR2_X1 U16587 ( .A1(n14781), .A2(n20019), .ZN(n14705) );
  AOI21_X1 U16588 ( .B1(n14775), .B2(P2_EAX_REG_5__SCAN_IN), .A(n14705), .ZN(
        n14680) );
  OAI21_X1 U16589 ( .B1(n14749), .B2(n14681), .A(n14680), .ZN(P2_U2972) );
  INV_X1 U16590 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n14683) );
  AOI22_X1 U16591 ( .A1(n19752), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n15700), .ZN(n20153) );
  NOR2_X1 U16592 ( .A1(n14781), .A2(n20153), .ZN(n14750) );
  AOI21_X1 U16593 ( .B1(n14775), .B2(P2_EAX_REG_18__SCAN_IN), .A(n14750), .ZN(
        n14682) );
  OAI21_X1 U16594 ( .B1(n14749), .B2(n14683), .A(n14682), .ZN(P2_U2954) );
  INV_X1 U16595 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n14685) );
  AOI22_X1 U16596 ( .A1(n19752), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n15700), .ZN(n19757) );
  NOR2_X1 U16597 ( .A1(n14781), .A2(n19757), .ZN(n14702) );
  AOI21_X1 U16598 ( .B1(n14775), .B2(P2_EAX_REG_7__SCAN_IN), .A(n14702), .ZN(
        n14684) );
  OAI21_X1 U16599 ( .B1(n14749), .B2(n14685), .A(n14684), .ZN(P2_U2974) );
  NAND2_X1 U16600 ( .A1(n14688), .A2(n14687), .ZN(n14689) );
  OR2_X1 U16601 ( .A1(n14690), .A2(n14689), .ZN(n14692) );
  NAND2_X1 U16602 ( .A1(n16032), .A2(n16028), .ZN(n16039) );
  INV_X1 U16603 ( .A(n14782), .ZN(n14696) );
  INV_X1 U16604 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n14695) );
  AND2_X1 U16605 ( .A1(n15786), .A2(n17825), .ZN(n15867) );
  INV_X1 U16606 ( .A(n15867), .ZN(n14694) );
  OAI211_X1 U16607 ( .C1(n14696), .C2(n14695), .A(n14783), .B(n14694), .ZN(
        P1_U2801) );
  INV_X1 U16608 ( .A(P2_UWORD_REG_6__SCAN_IN), .ZN(n14699) );
  AOI21_X1 U16609 ( .B1(n14775), .B2(P2_EAX_REG_22__SCAN_IN), .A(n14697), .ZN(
        n14698) );
  OAI21_X1 U16610 ( .B1(n14780), .B2(n14699), .A(n14698), .ZN(P2_U2958) );
  INV_X1 U16611 ( .A(P2_UWORD_REG_8__SCAN_IN), .ZN(n14701) );
  AOI22_X1 U16612 ( .A1(n19752), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n15700), .ZN(n16788) );
  NOR2_X1 U16613 ( .A1(n14781), .A2(n16788), .ZN(n14766) );
  AOI21_X1 U16614 ( .B1(n14775), .B2(P2_EAX_REG_24__SCAN_IN), .A(n14766), .ZN(
        n14700) );
  OAI21_X1 U16615 ( .B1(n14780), .B2(n14701), .A(n14700), .ZN(P2_U2960) );
  INV_X1 U16616 ( .A(P2_UWORD_REG_7__SCAN_IN), .ZN(n14704) );
  AOI21_X1 U16617 ( .B1(n14775), .B2(P2_EAX_REG_23__SCAN_IN), .A(n14702), .ZN(
        n14703) );
  OAI21_X1 U16618 ( .B1(n14780), .B2(n14704), .A(n14703), .ZN(P2_U2959) );
  INV_X1 U16619 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n14707) );
  AOI21_X1 U16620 ( .B1(n14775), .B2(P2_EAX_REG_21__SCAN_IN), .A(n14705), .ZN(
        n14706) );
  OAI21_X1 U16621 ( .B1(n14780), .B2(n14707), .A(n14706), .ZN(P2_U2957) );
  INV_X1 U16622 ( .A(P2_LWORD_REG_4__SCAN_IN), .ZN(n14709) );
  INV_X1 U16623 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n20611) );
  INV_X1 U16624 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n21216) );
  AOI22_X1 U16625 ( .A1(n19752), .A2(n20611), .B1(n21216), .B2(n15700), .ZN(
        n20061) );
  INV_X1 U16626 ( .A(n20061), .ZN(n20073) );
  NOR2_X1 U16627 ( .A1(n14781), .A2(n20073), .ZN(n14763) );
  AOI21_X1 U16628 ( .B1(n14775), .B2(P2_EAX_REG_4__SCAN_IN), .A(n14763), .ZN(
        n14708) );
  OAI21_X1 U16629 ( .B1(n14780), .B2(n14709), .A(n14708), .ZN(P2_U2971) );
  INV_X1 U16630 ( .A(P2_LWORD_REG_11__SCAN_IN), .ZN(n14711) );
  INV_X1 U16631 ( .A(n14781), .ZN(n14731) );
  AOI22_X1 U16632 ( .A1(n19752), .A2(BUF1_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n15700), .ZN(n14998) );
  INV_X1 U16633 ( .A(n14998), .ZN(n16756) );
  NAND2_X1 U16634 ( .A1(n14731), .A2(n16756), .ZN(n14712) );
  NAND2_X1 U16635 ( .A1(n14775), .A2(P2_EAX_REG_11__SCAN_IN), .ZN(n14710) );
  OAI211_X1 U16636 ( .C1(n14780), .C2(n14711), .A(n14712), .B(n14710), .ZN(
        P2_U2978) );
  INV_X1 U16637 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n16760) );
  INV_X1 U16638 ( .A(n14749), .ZN(n14735) );
  NAND2_X1 U16639 ( .A1(n14735), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n14713) );
  OAI211_X1 U16640 ( .C1(n14788), .C2(n16760), .A(n14713), .B(n14712), .ZN(
        P2_U2963) );
  INV_X1 U16641 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n14956) );
  NAND2_X1 U16642 ( .A1(n14735), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n14716) );
  INV_X1 U16643 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n20630) );
  OR2_X1 U16644 ( .A1(n15700), .A2(n20630), .ZN(n14715) );
  NAND2_X1 U16645 ( .A1(n15700), .A2(BUF2_REG_14__SCAN_IN), .ZN(n14714) );
  NAND2_X1 U16646 ( .A1(n14715), .A2(n14714), .ZN(n19742) );
  NAND2_X1 U16647 ( .A1(n14731), .A2(n19742), .ZN(n14725) );
  OAI211_X1 U16648 ( .C1(n14956), .C2(n14788), .A(n14716), .B(n14725), .ZN(
        P2_U2966) );
  INV_X1 U16649 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n14951) );
  NAND2_X1 U16650 ( .A1(n14735), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n14719) );
  INV_X1 U16651 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n20626) );
  OR2_X1 U16652 ( .A1(n15700), .A2(n20626), .ZN(n14718) );
  NAND2_X1 U16653 ( .A1(n15700), .A2(BUF2_REG_12__SCAN_IN), .ZN(n14717) );
  NAND2_X1 U16654 ( .A1(n14718), .A2(n14717), .ZN(n19745) );
  NAND2_X1 U16655 ( .A1(n14731), .A2(n19745), .ZN(n14733) );
  OAI211_X1 U16656 ( .C1(n14951), .C2(n14788), .A(n14719), .B(n14733), .ZN(
        P2_U2964) );
  INV_X1 U16657 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n16780) );
  NAND2_X1 U16658 ( .A1(n14735), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n14724) );
  INV_X1 U16659 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n14720) );
  OR2_X1 U16660 ( .A1(n15700), .A2(n14720), .ZN(n14722) );
  NAND2_X1 U16661 ( .A1(n15700), .A2(BUF2_REG_9__SCAN_IN), .ZN(n14721) );
  AND2_X1 U16662 ( .A1(n14722), .A2(n14721), .ZN(n16775) );
  INV_X1 U16663 ( .A(n16775), .ZN(n14723) );
  NAND2_X1 U16664 ( .A1(n14731), .A2(n14723), .ZN(n14773) );
  OAI211_X1 U16665 ( .C1(n14788), .C2(n16780), .A(n14724), .B(n14773), .ZN(
        P2_U2961) );
  INV_X1 U16666 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n17947) );
  NAND2_X1 U16667 ( .A1(n14735), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n14726) );
  OAI211_X1 U16668 ( .C1(n17947), .C2(n14788), .A(n14726), .B(n14725), .ZN(
        P2_U2981) );
  INV_X1 U16669 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n16745) );
  NAND2_X1 U16670 ( .A1(n14735), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n14728) );
  AOI22_X1 U16671 ( .A1(n19752), .A2(BUF1_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n15700), .ZN(n16741) );
  INV_X1 U16672 ( .A(n16741), .ZN(n14727) );
  NAND2_X1 U16673 ( .A1(n14731), .A2(n14727), .ZN(n14777) );
  OAI211_X1 U16674 ( .C1(n14788), .C2(n16745), .A(n14728), .B(n14777), .ZN(
        P2_U2965) );
  INV_X1 U16675 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n17939) );
  NAND2_X1 U16676 ( .A1(n14735), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n14732) );
  INV_X1 U16677 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n20622) );
  OR2_X1 U16678 ( .A1(n15700), .A2(n20622), .ZN(n14730) );
  NAND2_X1 U16679 ( .A1(n15700), .A2(BUF2_REG_10__SCAN_IN), .ZN(n14729) );
  AND2_X1 U16680 ( .A1(n14730), .A2(n14729), .ZN(n16770) );
  INV_X1 U16681 ( .A(n16770), .ZN(n19748) );
  NAND2_X1 U16682 ( .A1(n14731), .A2(n19748), .ZN(n14736) );
  OAI211_X1 U16683 ( .C1(n17939), .C2(n14788), .A(n14732), .B(n14736), .ZN(
        P2_U2977) );
  INV_X1 U16684 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n17943) );
  NAND2_X1 U16685 ( .A1(n14735), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n14734) );
  OAI211_X1 U16686 ( .C1(n17943), .C2(n14788), .A(n14734), .B(n14733), .ZN(
        P2_U2979) );
  INV_X1 U16687 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n14799) );
  NAND2_X1 U16688 ( .A1(n14735), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n14737) );
  OAI211_X1 U16689 ( .C1(n14799), .C2(n14788), .A(n14737), .B(n14736), .ZN(
        P2_U2962) );
  INV_X1 U16690 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18877) );
  AOI21_X1 U16691 ( .B1(n14746), .B2(n14739), .A(n14738), .ZN(n17322) );
  NAND2_X1 U16692 ( .A1(n12415), .A2(n17322), .ZN(n14740) );
  NAND2_X1 U16693 ( .A1(n19213), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n17326) );
  OAI211_X1 U16694 ( .C1(n17029), .C2(n18877), .A(n14740), .B(n17326), .ZN(
        n14741) );
  AOI21_X1 U16695 ( .B1(n17850), .B2(n18877), .A(n14741), .ZN(n14748) );
  INV_X1 U16696 ( .A(n14744), .ZN(n14743) );
  OAI222_X1 U16697 ( .A1(n14746), .A2(n14745), .B1(n14746), .B2(n14744), .C1(
        n14743), .C2(n14742), .ZN(n17324) );
  NAND2_X1 U16698 ( .A1(n17324), .A2(n17879), .ZN(n14747) );
  OAI211_X1 U16699 ( .C1(n17336), .C2(n17865), .A(n14748), .B(n14747), .ZN(
        P2_U3013) );
  INV_X1 U16700 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n14752) );
  AOI21_X1 U16701 ( .B1(n14775), .B2(P2_EAX_REG_2__SCAN_IN), .A(n14750), .ZN(
        n14751) );
  OAI21_X1 U16702 ( .B1(n14780), .B2(n14752), .A(n14751), .ZN(P2_U2969) );
  INV_X1 U16703 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n14754) );
  AOI22_X1 U16704 ( .A1(n19752), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n15700), .ZN(n20245) );
  NOR2_X1 U16705 ( .A1(n14781), .A2(n20245), .ZN(n14757) );
  AOI21_X1 U16706 ( .B1(n14775), .B2(P2_EAX_REG_0__SCAN_IN), .A(n14757), .ZN(
        n14753) );
  OAI21_X1 U16707 ( .B1(n14780), .B2(n14754), .A(n14753), .ZN(P2_U2967) );
  INV_X1 U16708 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n14756) );
  AOI22_X1 U16709 ( .A1(n19752), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n15700), .ZN(n20113) );
  NOR2_X1 U16710 ( .A1(n14781), .A2(n20113), .ZN(n14769) );
  AOI21_X1 U16711 ( .B1(n14775), .B2(P2_EAX_REG_19__SCAN_IN), .A(n14769), .ZN(
        n14755) );
  OAI21_X1 U16712 ( .B1(n14780), .B2(n14756), .A(n14755), .ZN(P2_U2955) );
  INV_X1 U16713 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n14759) );
  AOI21_X1 U16714 ( .B1(n14775), .B2(P2_EAX_REG_16__SCAN_IN), .A(n14757), .ZN(
        n14758) );
  OAI21_X1 U16715 ( .B1(n14780), .B2(n14759), .A(n14758), .ZN(P2_U2952) );
  INV_X1 U16716 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n14762) );
  AOI21_X1 U16717 ( .B1(n14775), .B2(P2_EAX_REG_1__SCAN_IN), .A(n14760), .ZN(
        n14761) );
  OAI21_X1 U16718 ( .B1(n14749), .B2(n14762), .A(n14761), .ZN(P2_U2968) );
  INV_X1 U16719 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n14765) );
  AOI21_X1 U16720 ( .B1(n14775), .B2(P2_EAX_REG_20__SCAN_IN), .A(n14763), .ZN(
        n14764) );
  OAI21_X1 U16721 ( .B1(n14749), .B2(n14765), .A(n14764), .ZN(P2_U2956) );
  INV_X1 U16722 ( .A(P2_LWORD_REG_8__SCAN_IN), .ZN(n14768) );
  AOI21_X1 U16723 ( .B1(n14775), .B2(P2_EAX_REG_8__SCAN_IN), .A(n14766), .ZN(
        n14767) );
  OAI21_X1 U16724 ( .B1(n14749), .B2(n14768), .A(n14767), .ZN(P2_U2975) );
  INV_X1 U16725 ( .A(P2_LWORD_REG_3__SCAN_IN), .ZN(n14771) );
  AOI21_X1 U16726 ( .B1(n14775), .B2(P2_EAX_REG_3__SCAN_IN), .A(n14769), .ZN(
        n14770) );
  OAI21_X1 U16727 ( .B1(n14749), .B2(n14771), .A(n14770), .ZN(P2_U2970) );
  INV_X1 U16728 ( .A(P2_LWORD_REG_9__SCAN_IN), .ZN(n14774) );
  NAND2_X1 U16729 ( .A1(n14775), .A2(P2_EAX_REG_9__SCAN_IN), .ZN(n14772) );
  OAI211_X1 U16730 ( .C1(n14749), .C2(n14774), .A(n14773), .B(n14772), .ZN(
        P2_U2976) );
  INV_X1 U16731 ( .A(P2_LWORD_REG_13__SCAN_IN), .ZN(n14778) );
  NAND2_X1 U16732 ( .A1(n14775), .A2(P2_EAX_REG_13__SCAN_IN), .ZN(n14776) );
  OAI211_X1 U16733 ( .C1(n14780), .C2(n14778), .A(n14777), .B(n14776), .ZN(
        P2_U2980) );
  AOI22_X1 U16734 ( .A1(n19752), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n15700), .ZN(n15111) );
  INV_X1 U16735 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n17952) );
  INV_X1 U16736 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n14779) );
  OAI222_X1 U16737 ( .A1(n14781), .A2(n15111), .B1(n14788), .B2(n17952), .C1(
        n14780), .C2(n14779), .ZN(P2_U2982) );
  INV_X1 U16738 ( .A(n21874), .ZN(n14785) );
  OAI21_X1 U16739 ( .B1(n15867), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n14785), 
        .ZN(n14784) );
  OAI21_X1 U16740 ( .B1(n14786), .B2(n14785), .A(n14784), .ZN(P1_U3487) );
  INV_X1 U16741 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n14792) );
  NOR2_X1 U16742 ( .A1(n12471), .A2(n14673), .ZN(n14787) );
  NAND2_X1 U16743 ( .A1(n19242), .A2(n14787), .ZN(n15758) );
  OAI21_X1 U16744 ( .B1(n15758), .B2(n19287), .A(n14788), .ZN(n14790) );
  INV_X1 U16745 ( .A(n22332), .ZN(n14789) );
  NOR2_X1 U16746 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n17768), .ZN(n17937) );
  AOI22_X1 U16747 ( .A1(n17949), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n17928), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n14791) );
  OAI21_X1 U16748 ( .B1(n14792), .B2(n14959), .A(n14791), .ZN(P2_U2929) );
  INV_X1 U16749 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n16799) );
  AOI22_X1 U16750 ( .A1(n17949), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n17928), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n14793) );
  OAI21_X1 U16751 ( .B1(n16799), .B2(n14959), .A(n14793), .ZN(P2_U2928) );
  INV_X1 U16752 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n16806) );
  AOI22_X1 U16753 ( .A1(n17949), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n17928), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n14794) );
  OAI21_X1 U16754 ( .B1(n16806), .B2(n14959), .A(n14794), .ZN(P2_U2930) );
  INV_X1 U16755 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n16787) );
  AOI22_X1 U16756 ( .A1(n17949), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n17928), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n14795) );
  OAI21_X1 U16757 ( .B1(n16787), .B2(n14959), .A(n14795), .ZN(P2_U2927) );
  INV_X1 U16758 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n14797) );
  AOI22_X1 U16759 ( .A1(n17949), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n17928), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n14796) );
  OAI21_X1 U16760 ( .B1(n14797), .B2(n14959), .A(n14796), .ZN(P2_U2931) );
  AOI22_X1 U16761 ( .A1(n17949), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n17928), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n14798) );
  OAI21_X1 U16762 ( .B1(n14799), .B2(n14959), .A(n14798), .ZN(P2_U2925) );
  AOI22_X1 U16763 ( .A1(n17949), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n17928), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n14800) );
  OAI21_X1 U16764 ( .B1(n16780), .B2(n14959), .A(n14800), .ZN(P2_U2926) );
  NAND2_X1 U16765 ( .A1(n13896), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n14801) );
  AND4_X1 U16766 ( .A1(n19970), .A2(n14801), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n19916), .ZN(n14802) );
  NOR2_X1 U16767 ( .A1(n11141), .A2(n18858), .ZN(n14804) );
  AOI21_X1 U16768 ( .B1(P2_EBX_REG_0__SCAN_IN), .B2(n11141), .A(n14804), .ZN(
        n14805) );
  OAI21_X1 U16769 ( .B1(n19925), .B2(n16740), .A(n14805), .ZN(P2_U2887) );
  INV_X1 U16770 ( .A(n19241), .ZN(n14808) );
  AND2_X1 U16771 ( .A1(n12725), .A2(n19281), .ZN(n19246) );
  NAND2_X1 U16772 ( .A1(n19245), .A2(n19246), .ZN(n14806) );
  NOR2_X1 U16773 ( .A1(n19248), .A2(n14806), .ZN(n14807) );
  AOI21_X1 U16774 ( .B1(n19242), .B2(n14808), .A(n14807), .ZN(n15761) );
  NAND2_X1 U16775 ( .A1(n14809), .A2(n12722), .ZN(n14810) );
  NAND2_X1 U16776 ( .A1(n15761), .A2(n14810), .ZN(n14811) );
  NAND2_X1 U16777 ( .A1(n15694), .A2(n12494), .ZN(n15600) );
  INV_X1 U16778 ( .A(n14812), .ZN(n14813) );
  XNOR2_X1 U16779 ( .A(n14814), .B(n14813), .ZN(n17311) );
  INV_X1 U16780 ( .A(n17311), .ZN(n18917) );
  NAND2_X1 U16781 ( .A1(n16817), .A2(n14815), .ZN(n20012) );
  INV_X1 U16782 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n17930) );
  OAI222_X1 U16783 ( .A1(n15600), .A2(n19969), .B1(n18917), .B2(n20018), .C1(
        n17930), .C2(n16817), .ZN(P2_U2913) );
  OAI21_X1 U16784 ( .B1(n14819), .B2(n14818), .A(n14817), .ZN(n18928) );
  OAI222_X1 U16785 ( .A1(n15600), .A2(n19757), .B1(n18928), .B2(n20018), .C1(
        n17932), .C2(n16817), .ZN(P2_U2912) );
  XNOR2_X1 U16786 ( .A(n14820), .B(n14821), .ZN(n19179) );
  XNOR2_X1 U16787 ( .A(n19925), .B(n19179), .ZN(n14826) );
  INV_X1 U16788 ( .A(n15600), .ZN(n20011) );
  INV_X1 U16789 ( .A(n20245), .ZN(n14824) );
  OAI22_X1 U16790 ( .A1(n16818), .A2(n19179), .B1(n16817), .B2(n14822), .ZN(
        n14823) );
  AOI21_X1 U16791 ( .B1(n20011), .B2(n14824), .A(n14823), .ZN(n14825) );
  OAI21_X1 U16792 ( .B1(n14826), .B2(n20012), .A(n14825), .ZN(P2_U2919) );
  INV_X1 U16793 ( .A(n13341), .ZN(n15240) );
  INV_X1 U16794 ( .A(n14828), .ZN(n14830) );
  AND3_X1 U16795 ( .A1(n14919), .A2(n14830), .A3(n14829), .ZN(n14831) );
  NAND2_X1 U16796 ( .A1(n14827), .A2(n14831), .ZN(n14844) );
  INV_X1 U16797 ( .A(n14832), .ZN(n14839) );
  INV_X1 U16798 ( .A(n15239), .ZN(n14870) );
  OAI21_X1 U16799 ( .B1(n12975), .B2(n14833), .A(n14870), .ZN(n14836) );
  AOI21_X1 U16800 ( .B1(n16023), .B2(n12966), .A(n16033), .ZN(n14835) );
  NAND3_X1 U16801 ( .A1(n14836), .A2(n14835), .A3(n14834), .ZN(n14837) );
  AOI21_X1 U16802 ( .B1(n14839), .B2(n14838), .A(n14837), .ZN(n14843) );
  AOI21_X1 U16803 ( .B1(n12951), .B2(n15229), .A(n15146), .ZN(n14841) );
  NAND2_X1 U16804 ( .A1(n14842), .A2(n14841), .ZN(n14850) );
  NAND3_X1 U16805 ( .A1(n14843), .A2(n14840), .A3(n14850), .ZN(n14921) );
  OR2_X1 U16806 ( .A1(n14844), .A2(n14921), .ZN(n16620) );
  OAI22_X1 U16807 ( .A1(n15240), .A2(n16607), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n16592), .ZN(n17788) );
  INV_X1 U16808 ( .A(n22277), .ZN(n16623) );
  OAI22_X1 U16809 ( .A1(n17825), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n16623), .ZN(n14845) );
  AOI21_X1 U16810 ( .B1(n17788), .B2(n16596), .A(n14845), .ZN(n14869) );
  INV_X1 U16811 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n14846) );
  NAND2_X1 U16812 ( .A1(n14847), .A2(n14846), .ZN(n22314) );
  INV_X1 U16813 ( .A(n22314), .ZN(n16040) );
  OAI21_X1 U16814 ( .B1(n15229), .B2(n16040), .A(n21876), .ZN(n15228) );
  AOI211_X1 U16815 ( .C1(n16038), .C2(n22314), .A(n15228), .B(n16036), .ZN(
        n14848) );
  OAI21_X1 U16816 ( .B1(n16613), .B2(n14828), .A(n14848), .ZN(n14856) );
  INV_X1 U16817 ( .A(n16032), .ZN(n14853) );
  INV_X1 U16818 ( .A(n14849), .ZN(n14851) );
  NAND2_X1 U16819 ( .A1(n14851), .A2(n14850), .ZN(n14852) );
  NAND2_X1 U16820 ( .A1(n14853), .A2(n14852), .ZN(n14905) );
  NAND2_X1 U16821 ( .A1(n16030), .A2(n16036), .ZN(n14855) );
  OR2_X1 U16822 ( .A1(n15239), .A2(n12966), .ZN(n14854) );
  NAND4_X1 U16823 ( .A1(n14856), .A2(n14905), .A3(n14855), .A4(n14854), .ZN(
        n14862) );
  NAND2_X1 U16824 ( .A1(n16028), .A2(n21876), .ZN(n14857) );
  OR2_X1 U16825 ( .A1(n11162), .A2(n14857), .ZN(n14861) );
  NAND2_X1 U16826 ( .A1(n14858), .A2(n12946), .ZN(n14859) );
  NOR2_X1 U16827 ( .A1(n16592), .A2(n14859), .ZN(n14907) );
  NAND2_X1 U16828 ( .A1(n14907), .A2(n16029), .ZN(n14860) );
  INV_X1 U16829 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n22269) );
  NOR3_X1 U16830 ( .A1(n22269), .A2(n22274), .A3(n22273), .ZN(n14864) );
  NOR2_X1 U16831 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n22435), .ZN(n14863) );
  OR2_X1 U16832 ( .A1(n14864), .A2(n14863), .ZN(n14865) );
  AOI21_X1 U16833 ( .B1(n17803), .B2(n16042), .A(n14865), .ZN(n16626) );
  INV_X1 U16834 ( .A(n16613), .ZN(n14867) );
  NOR2_X1 U16835 ( .A1(n14867), .A2(n14866), .ZN(n17787) );
  AOI22_X1 U16836 ( .A1(n16626), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n16596), .B2(n17787), .ZN(n14868) );
  OAI21_X1 U16837 ( .B1(n14869), .B2(n16626), .A(n14868), .ZN(P1_U3474) );
  XNOR2_X1 U16838 ( .A(n16595), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14874) );
  NOR2_X1 U16839 ( .A1(n14870), .A2(n21878), .ZN(n16041) );
  AND2_X1 U16840 ( .A1(n14871), .A2(n16041), .ZN(n16611) );
  XNOR2_X1 U16841 ( .A(n14872), .B(n12838), .ZN(n14877) );
  INV_X1 U16842 ( .A(n14877), .ZN(n14873) );
  AOI22_X1 U16843 ( .A1(n16613), .A2(n14874), .B1(n16611), .B2(n14873), .ZN(
        n14876) );
  NAND3_X1 U16844 ( .A1(n16607), .A2(n12975), .A3(n14877), .ZN(n14875) );
  OAI211_X1 U16845 ( .C1(n15337), .C2(n16607), .A(n14876), .B(n14875), .ZN(
        n17784) );
  OAI22_X1 U16846 ( .A1(n22064), .A2(n16449), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n16599) );
  INV_X1 U16847 ( .A(n16599), .ZN(n14878) );
  INV_X1 U16848 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21908) );
  NOR2_X1 U16849 ( .A1(n17825), .A2(n21908), .ZN(n16598) );
  AOI222_X1 U16850 ( .A1(n17784), .A2(n16596), .B1(n14878), .B2(n16598), .C1(
        n22277), .C2(n14877), .ZN(n14879) );
  MUX2_X1 U16851 ( .A(n14879), .B(n12838), .S(n16626), .Z(n14880) );
  INV_X1 U16852 ( .A(n14880), .ZN(P1_U3472) );
  XNOR2_X2 U16853 ( .A(n14883), .B(n14882), .ZN(n19820) );
  MUX2_X1 U16854 ( .A(n17336), .B(n18871), .S(n11141), .Z(n14884) );
  OAI21_X1 U16855 ( .B1(n19820), .B2(n16740), .A(n14884), .ZN(P2_U2886) );
  INV_X1 U16856 ( .A(n16626), .ZN(n16601) );
  INV_X1 U16857 ( .A(n15092), .ZN(n15248) );
  NOR2_X1 U16858 ( .A1(n14885), .A2(n15248), .ZN(n14886) );
  XNOR2_X1 U16859 ( .A(n14886), .B(n17802), .ZN(n22075) );
  INV_X1 U16860 ( .A(n14827), .ZN(n17799) );
  NAND4_X1 U16861 ( .A1(n22075), .A2(n16596), .A3(n17799), .A4(n16601), .ZN(
        n14887) );
  OAI21_X1 U16862 ( .B1(n17802), .B2(n16601), .A(n14887), .ZN(P1_U3468) );
  MUX2_X1 U16863 ( .A(n16014), .B(n15746), .S(n11141), .Z(n14890) );
  OAI21_X1 U16864 ( .B1(n19879), .B2(n16740), .A(n14890), .ZN(P2_U2885) );
  AOI21_X1 U16865 ( .B1(n14891), .B2(n14817), .A(n14926), .ZN(n19190) );
  INV_X1 U16866 ( .A(n19190), .ZN(n14892) );
  INV_X1 U16867 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n17934) );
  OAI222_X1 U16868 ( .A1(n15600), .A2(n16788), .B1(n14892), .B2(n20018), .C1(
        n17934), .C2(n16817), .ZN(P2_U2911) );
  OAI21_X1 U16869 ( .B1(n14894), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n14893), .ZN(n14942) );
  INV_X1 U16870 ( .A(n21876), .ZN(n22305) );
  AOI21_X1 U16871 ( .B1(n15229), .B2(n22314), .A(n22305), .ZN(n14895) );
  NAND2_X1 U16872 ( .A1(n16028), .A2(n14895), .ZN(n14901) );
  INV_X1 U16873 ( .A(n15228), .ZN(n14896) );
  NAND2_X1 U16874 ( .A1(n14828), .A2(n14896), .ZN(n14897) );
  NAND3_X1 U16875 ( .A1(n14897), .A2(n16021), .A3(n15992), .ZN(n14898) );
  NAND2_X1 U16876 ( .A1(n14898), .A2(n16029), .ZN(n14900) );
  MUX2_X1 U16877 ( .A(n14901), .B(n14900), .S(n14899), .Z(n14904) );
  NAND3_X1 U16878 ( .A1(n16036), .A2(n14902), .A3(n15229), .ZN(n14903) );
  NAND3_X1 U16879 ( .A1(n14905), .A2(n14904), .A3(n14903), .ZN(n14906) );
  NOR2_X1 U16880 ( .A1(n17804), .A2(n14907), .ZN(n16024) );
  OAI22_X1 U16881 ( .A1(n12961), .A2(n14908), .B1(n16038), .B2(n15379), .ZN(
        n14909) );
  INV_X1 U16882 ( .A(n14909), .ZN(n14910) );
  NAND3_X1 U16883 ( .A1(n16024), .A2(n14910), .A3(n11162), .ZN(n14911) );
  OAI22_X1 U16884 ( .A1(n12955), .A2(n14908), .B1(n16038), .B2(n15229), .ZN(
        n14912) );
  NOR2_X1 U16885 ( .A1(n15973), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14913) );
  OR2_X1 U16886 ( .A1(n14914), .A2(n14913), .ZN(n15236) );
  INV_X1 U16887 ( .A(n15236), .ZN(n14917) );
  INV_X1 U16888 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n15237) );
  NOR2_X1 U16889 ( .A1(n22049), .A2(n15237), .ZN(n14946) );
  INV_X1 U16890 ( .A(n14923), .ZN(n14915) );
  NAND2_X1 U16891 ( .A1(n14915), .A2(n22049), .ZN(n22062) );
  AOI21_X1 U16892 ( .B1(n21892), .B2(n22062), .A(n21908), .ZN(n14916) );
  AOI211_X1 U16893 ( .C1(n22056), .C2(n14917), .A(n14946), .B(n14916), .ZN(
        n14924) );
  OAI21_X1 U16894 ( .B1(n14919), .B2(n16021), .A(n14918), .ZN(n14920) );
  OR2_X1 U16895 ( .A1(n14921), .A2(n14920), .ZN(n14922) );
  NAND2_X1 U16896 ( .A1(n14923), .A2(n14922), .ZN(n21888) );
  INV_X1 U16897 ( .A(n21888), .ZN(n16536) );
  OAI21_X1 U16898 ( .B1(n16536), .B2(n22007), .A(n21908), .ZN(n22063) );
  OAI211_X1 U16899 ( .C1(n14942), .C2(n22031), .A(n14924), .B(n22063), .ZN(
        P1_U3031) );
  OAI21_X1 U16900 ( .B1(n14926), .B2(n14925), .A(n15767), .ZN(n18946) );
  INV_X1 U16901 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n17936) );
  OAI222_X1 U16902 ( .A1(n15600), .A2(n16775), .B1(n18946), .B2(n20018), .C1(
        n17936), .C2(n16817), .ZN(P2_U2910) );
  INV_X1 U16903 ( .A(n14927), .ZN(n14930) );
  OAI21_X1 U16904 ( .B1(n14930), .B2(n14929), .A(n14928), .ZN(n15247) );
  AND2_X1 U16905 ( .A1(n15229), .A2(n21876), .ZN(n14934) );
  NOR2_X1 U16906 ( .A1(n14829), .A2(n14932), .ZN(n14933) );
  INV_X1 U16907 ( .A(n15987), .ZN(n15991) );
  NAND2_X1 U16908 ( .A1(n15991), .A2(DATAI_0_), .ZN(n14940) );
  NAND2_X1 U16909 ( .A1(n15987), .A2(BUF1_REG_0__SCAN_IN), .ZN(n14939) );
  AND2_X1 U16910 ( .A1(n14940), .A2(n14939), .ZN(n15481) );
  INV_X1 U16911 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20416) );
  OAI222_X1 U16912 ( .A1(n15247), .A2(n16238), .B1(n16268), .B2(n15481), .C1(
        n16265), .C2(n20416), .ZN(P1_U2904) );
  INV_X1 U16913 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n15696) );
  AOI22_X1 U16914 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n17948), .B1(n17949), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n14941) );
  OAI21_X1 U16915 ( .B1(n15696), .B2(n14959), .A(n14941), .ZN(P2_U2935) );
  INV_X1 U16916 ( .A(n14942), .ZN(n14947) );
  INV_X1 U16917 ( .A(n20588), .ZN(n16405) );
  INV_X1 U16918 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14943) );
  AOI21_X1 U16919 ( .B1(n16405), .B2(n14944), .A(n14943), .ZN(n14945) );
  AOI211_X1 U16920 ( .C1(n14947), .C2(n20591), .A(n14946), .B(n14945), .ZN(
        n14948) );
  OAI21_X1 U16921 ( .B1(n16428), .B2(n15247), .A(n14948), .ZN(P1_U2999) );
  AOI22_X1 U16922 ( .A1(n17949), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n17948), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n14949) );
  OAI21_X1 U16923 ( .B1(n16745), .B2(n14959), .A(n14949), .ZN(P2_U2922) );
  AOI22_X1 U16924 ( .A1(n17949), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n17948), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n14950) );
  OAI21_X1 U16925 ( .B1(n14951), .B2(n14959), .A(n14950), .ZN(P2_U2923) );
  AOI22_X1 U16926 ( .A1(n17949), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n17948), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n14952) );
  OAI21_X1 U16927 ( .B1(n16760), .B2(n14959), .A(n14952), .ZN(P2_U2924) );
  INV_X1 U16928 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n14954) );
  AOI22_X1 U16929 ( .A1(n17937), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n17948), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n14953) );
  OAI21_X1 U16930 ( .B1(n14954), .B2(n14959), .A(n14953), .ZN(P2_U2934) );
  AOI22_X1 U16931 ( .A1(n17937), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n17948), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n14955) );
  OAI21_X1 U16932 ( .B1(n14956), .B2(n14959), .A(n14955), .ZN(P2_U2921) );
  INV_X1 U16933 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n15879) );
  AOI22_X1 U16934 ( .A1(n17937), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n17948), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n14957) );
  OAI21_X1 U16935 ( .B1(n15879), .B2(n14959), .A(n14957), .ZN(P2_U2933) );
  INV_X1 U16936 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n16816) );
  AOI22_X1 U16937 ( .A1(n17937), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n17948), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n14958) );
  OAI21_X1 U16938 ( .B1(n16816), .B2(n14959), .A(n14958), .ZN(P2_U2932) );
  NOR2_X1 U16939 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n22278) );
  INV_X1 U16940 ( .A(n22278), .ZN(n14960) );
  INV_X1 U16941 ( .A(n12849), .ZN(n14962) );
  OAI21_X1 U16942 ( .B1(n14962), .B2(n14961), .A(n17802), .ZN(n14963) );
  NAND2_X1 U16943 ( .A1(n14963), .A2(n22269), .ZN(n16587) );
  OR2_X1 U16944 ( .A1(n22274), .A2(n22273), .ZN(n14964) );
  AOI21_X1 U16945 ( .B1(n16587), .B2(n22269), .A(n14964), .ZN(n14965) );
  OR2_X1 U16946 ( .A1(n15124), .A2(n14965), .ZN(n17826) );
  NAND2_X1 U16947 ( .A1(n17826), .A2(n15786), .ZN(n15034) );
  INV_X1 U16948 ( .A(n15335), .ZN(n14967) );
  INV_X1 U16949 ( .A(n14966), .ZN(n15451) );
  NAND2_X1 U16950 ( .A1(n15451), .A2(n22286), .ZN(n15288) );
  NAND2_X1 U16951 ( .A1(n14967), .A2(n15288), .ZN(n14973) );
  NAND2_X1 U16952 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n22435), .ZN(n16589) );
  NAND2_X1 U16953 ( .A1(n17826), .A2(n16589), .ZN(n15036) );
  INV_X1 U16954 ( .A(n15036), .ZN(n14971) );
  INV_X1 U16955 ( .A(n14969), .ZN(n22427) );
  INV_X1 U16956 ( .A(n17826), .ZN(n14970) );
  AOI22_X1 U16957 ( .A1(n14971), .A2(n22427), .B1(n14970), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n14972) );
  OAI21_X1 U16958 ( .B1(n15034), .B2(n14973), .A(n14972), .ZN(P1_U3477) );
  OR2_X1 U16959 ( .A1(n14976), .A2(n14975), .ZN(n14977) );
  NAND2_X1 U16960 ( .A1(n14974), .A2(n14977), .ZN(n20013) );
  OR2_X1 U16961 ( .A1(n14979), .A2(n14978), .ZN(n14981) );
  NAND2_X1 U16962 ( .A1(n14981), .A2(n14980), .ZN(n19201) );
  MUX2_X1 U16963 ( .A(n12275), .B(n19201), .S(n16727), .Z(n14982) );
  OAI21_X1 U16964 ( .B1(n20013), .B2(n16740), .A(n14982), .ZN(P2_U2883) );
  INV_X1 U16965 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n15635) );
  MUX2_X1 U16966 ( .A(n15635), .B(n15437), .S(n16727), .Z(n14987) );
  OAI21_X1 U16967 ( .B1(n19880), .B2(n16740), .A(n14987), .ZN(P2_U2884) );
  OAI222_X1 U16968 ( .A1(n15236), .A2(n20510), .B1(n20524), .B2(n14988), .C1(
        n15247), .C2(n16189), .ZN(P1_U2872) );
  XOR2_X1 U16969 ( .A(n14974), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n14992)
         );
  AOI21_X1 U16970 ( .B1(n14989), .B2(n14980), .A(n11263), .ZN(n18903) );
  NOR2_X1 U16971 ( .A1(n16727), .A2(n12046), .ZN(n14990) );
  AOI21_X1 U16972 ( .B1(n18903), .B2(n16727), .A(n14990), .ZN(n14991) );
  OAI21_X1 U16973 ( .B1(n14992), .B2(n16740), .A(n14991), .ZN(P2_U2882) );
  OR2_X1 U16974 ( .A1(n14994), .A2(n14995), .ZN(n14996) );
  AND2_X1 U16975 ( .A1(n14993), .A2(n14996), .ZN(n18955) );
  INV_X1 U16976 ( .A(n18955), .ZN(n14997) );
  INV_X1 U16977 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n17941) );
  OAI222_X1 U16978 ( .A1(n15600), .A2(n14998), .B1(n14997), .B2(n20018), .C1(
        n17941), .C2(n16817), .ZN(P2_U2908) );
  XNOR2_X1 U16979 ( .A(n15333), .B(n15335), .ZN(n15000) );
  OAI222_X1 U16980 ( .A1(n15036), .A2(n15337), .B1(n17826), .B2(n17795), .C1(
        n15000), .C2(n15034), .ZN(P1_U3476) );
  OR2_X1 U16981 ( .A1(n15002), .A2(n15001), .ZN(n15003) );
  NAND2_X1 U16982 ( .A1(n15049), .A2(n15003), .ZN(n22069) );
  NAND2_X1 U16983 ( .A1(n15991), .A2(DATAI_1_), .ZN(n15005) );
  NAND2_X1 U16984 ( .A1(n15987), .A2(BUF1_REG_1__SCAN_IN), .ZN(n15004) );
  AND2_X1 U16985 ( .A1(n15005), .A2(n15004), .ZN(n15494) );
  OAI222_X1 U16986 ( .A1(n22069), .A2(n16238), .B1(n16268), .B2(n15494), .C1(
        n16265), .C2(n13333), .ZN(P1_U2903) );
  XNOR2_X1 U16987 ( .A(n15006), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n15012) );
  NAND2_X1 U16988 ( .A1(n15008), .A2(n15009), .ZN(n15010) );
  NAND2_X1 U16989 ( .A1(n15007), .A2(n15010), .ZN(n18927) );
  MUX2_X1 U16990 ( .A(n18927), .B(n12285), .S(n11141), .Z(n15011) );
  OAI21_X1 U16991 ( .B1(n15012), .B2(n16740), .A(n15011), .ZN(P2_U2880) );
  INV_X1 U16992 ( .A(n19820), .ZN(n19913) );
  OAI21_X1 U16993 ( .B1(n15015), .B2(n15014), .A(n15013), .ZN(n17323) );
  XNOR2_X1 U16994 ( .A(n19913), .B(n17323), .ZN(n15017) );
  NOR2_X1 U16995 ( .A1(n19925), .A2(n19179), .ZN(n15016) );
  NOR2_X1 U16996 ( .A1(n15017), .A2(n15016), .ZN(n15201) );
  AOI21_X1 U16997 ( .B1(n15017), .B2(n15016), .A(n15201), .ZN(n15021) );
  AOI22_X1 U16998 ( .A1(n20067), .A2(n17323), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n20060), .ZN(n15020) );
  INV_X1 U16999 ( .A(n20195), .ZN(n15018) );
  NAND2_X1 U17000 ( .A1(n20011), .A2(n15018), .ZN(n15019) );
  OAI211_X1 U17001 ( .C1(n15021), .C2(n20012), .A(n15020), .B(n15019), .ZN(
        P2_U2918) );
  OR2_X1 U17002 ( .A1(n15022), .A2(n11263), .ZN(n15023) );
  NAND2_X1 U17003 ( .A1(n15008), .A2(n15023), .ZN(n18916) );
  NOR2_X1 U17004 ( .A1(n14974), .A2(n20059), .ZN(n15025) );
  INV_X1 U17005 ( .A(n15006), .ZN(n15024) );
  OAI211_X1 U17006 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n15025), .A(
        n15024), .B(n16732), .ZN(n15027) );
  NAND2_X1 U17007 ( .A1(n11141), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n15026) );
  OAI211_X1 U17008 ( .C1(n18916), .C2(n11141), .A(n15027), .B(n15026), .ZN(
        P2_U2881) );
  XNOR2_X1 U17009 ( .A(n15028), .B(n15972), .ZN(n22055) );
  INV_X1 U17010 ( .A(n20524), .ZN(n16183) );
  AOI22_X1 U17011 ( .A1(n20528), .A2(n22055), .B1(n16183), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n15029) );
  OAI21_X1 U17012 ( .B1(n22069), .B2(n16189), .A(n15029), .ZN(P1_U2871) );
  INV_X1 U17013 ( .A(n16621), .ZN(n15035) );
  NAND2_X1 U17014 ( .A1(n15333), .A2(n15031), .ZN(n15458) );
  INV_X1 U17015 ( .A(n15458), .ZN(n15452) );
  NAND2_X1 U17016 ( .A1(n15452), .A2(n15335), .ZN(n15250) );
  NOR2_X1 U17017 ( .A1(n14999), .A2(n15031), .ZN(n15287) );
  NAND2_X1 U17018 ( .A1(n15087), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n15103) );
  INV_X1 U17019 ( .A(n15103), .ZN(n15032) );
  AOI21_X1 U17020 ( .B1(n13319), .B2(n15250), .A(n15032), .ZN(n15033) );
  OAI222_X1 U17021 ( .A1(n17826), .A2(n15570), .B1(n15036), .B2(n15035), .C1(
        n15034), .C2(n15033), .ZN(P1_U3475) );
  INV_X1 U17022 ( .A(n15037), .ZN(n15846) );
  AOI21_X1 U17023 ( .B1(n15039), .B2(n15846), .A(n15038), .ZN(n17226) );
  INV_X1 U17024 ( .A(n17226), .ZN(n18970) );
  INV_X1 U17025 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n17945) );
  OAI222_X1 U17026 ( .A1(n15600), .A2(n16741), .B1(n18970), .B2(n20018), .C1(
        n17945), .C2(n16817), .ZN(P2_U2906) );
  XNOR2_X1 U17027 ( .A(n15040), .B(n15056), .ZN(n15046) );
  OR2_X1 U17028 ( .A1(n15042), .A2(n15043), .ZN(n15044) );
  NAND2_X1 U17029 ( .A1(n15041), .A2(n15044), .ZN(n18941) );
  MUX2_X1 U17030 ( .A(n18941), .B(n12132), .S(n11141), .Z(n15045) );
  OAI21_X1 U17031 ( .B1(n15046), .B2(n16740), .A(n15045), .ZN(P2_U2878) );
  INV_X1 U17032 ( .A(n15047), .ZN(n15048) );
  AOI21_X1 U17033 ( .B1(n15050), .B2(n15049), .A(n15048), .ZN(n15276) );
  INV_X1 U17034 ( .A(n15276), .ZN(n15084) );
  NAND2_X1 U17035 ( .A1(n15991), .A2(DATAI_2_), .ZN(n15052) );
  NAND2_X1 U17036 ( .A1(n15987), .A2(BUF1_REG_2__SCAN_IN), .ZN(n15051) );
  OAI222_X1 U17037 ( .A1(n15084), .A2(n16238), .B1(n16268), .B2(n15496), .C1(
        n16265), .C2(n13327), .ZN(P1_U2902) );
  INV_X1 U17038 ( .A(n15053), .ZN(n15054) );
  AOI21_X1 U17039 ( .B1(n15055), .B2(n15041), .A(n15054), .ZN(n17267) );
  INV_X1 U17040 ( .A(n17267), .ZN(n15062) );
  AND2_X1 U17041 ( .A1(n15040), .A2(n15056), .ZN(n15059) );
  OAI211_X1 U17042 ( .C1(n15059), .C2(n15058), .A(n16732), .B(n15057), .ZN(
        n15061) );
  NAND2_X1 U17043 ( .A1(n11141), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n15060) );
  OAI211_X1 U17044 ( .C1(n15062), .C2(n11141), .A(n15061), .B(n15060), .ZN(
        P2_U2877) );
  NAND2_X1 U17045 ( .A1(n16613), .A2(n15063), .ZN(n15064) );
  NOR2_X4 U17046 ( .A1(n20414), .A2(n21877), .ZN(n20429) );
  AOI22_X1 U17047 ( .A1(n20425), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n20429), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n15066) );
  OAI21_X1 U17048 ( .B1(n13540), .B2(n15623), .A(n15066), .ZN(P1_U2919) );
  INV_X1 U17049 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n15526) );
  AOI22_X1 U17050 ( .A1(n21877), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n20429), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n15067) );
  OAI21_X1 U17051 ( .B1(n15526), .B2(n15623), .A(n15067), .ZN(P1_U2918) );
  AOI22_X1 U17052 ( .A1(n20588), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n22052), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n15068) );
  OAI21_X1 U17053 ( .B1(n20594), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n15068), .ZN(n15069) );
  INV_X1 U17054 ( .A(n15069), .ZN(n15073) );
  OR2_X1 U17055 ( .A1(n15070), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n22054) );
  NAND3_X1 U17056 ( .A1(n22054), .A2(n15071), .A3(n20591), .ZN(n15072) );
  OAI211_X1 U17057 ( .C1(n22069), .C2(n16428), .A(n15073), .B(n15072), .ZN(
        P1_U2998) );
  AOI21_X1 U17058 ( .B1(n15074), .B2(n15007), .A(n15042), .ZN(n19192) );
  INV_X1 U17059 ( .A(n19192), .ZN(n15075) );
  NOR2_X1 U17060 ( .A1(n15075), .A2(n11141), .ZN(n15079) );
  NAND2_X1 U17061 ( .A1(n15006), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n15076) );
  AOI211_X1 U17062 ( .C1(n15077), .C2(n15076), .A(n16740), .B(n15040), .ZN(
        n15078) );
  AOI211_X1 U17063 ( .C1(P2_EBX_REG_8__SCAN_IN), .C2(n11141), .A(n15079), .B(
        n15078), .ZN(n15080) );
  INV_X1 U17064 ( .A(n15080), .ZN(P2_U2879) );
  NAND2_X1 U17065 ( .A1(n15082), .A2(n15081), .ZN(n15083) );
  NAND2_X1 U17066 ( .A1(n15374), .A2(n15083), .ZN(n21919) );
  INV_X1 U17067 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n15085) );
  OAI222_X1 U17068 ( .A1(n21919), .A2(n20510), .B1(n15085), .B2(n20524), .C1(
        n16189), .C2(n15084), .ZN(P1_U2870) );
  INV_X1 U17069 ( .A(DATAI_31_), .ZN(n15086) );
  INV_X1 U17070 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n20667) );
  OAI22_X1 U17071 ( .A1(n15086), .A2(n15164), .B1(n20667), .B2(n15161), .ZN(
        n22662) );
  INV_X1 U17072 ( .A(n22662), .ZN(n22681) );
  INV_X1 U17073 ( .A(DATAI_23_), .ZN(n15089) );
  INV_X1 U17074 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n20649) );
  OR2_X1 U17075 ( .A1(n15161), .A2(n20649), .ZN(n15088) );
  NAND2_X1 U17076 ( .A1(n15991), .A2(DATAI_7_), .ZN(n15091) );
  NAND2_X1 U17077 ( .A1(n15987), .A2(BUF1_REG_7__SCAN_IN), .ZN(n15090) );
  NOR2_X1 U17078 ( .A1(n15337), .A2(n15092), .ZN(n22396) );
  INV_X1 U17079 ( .A(n15093), .ZN(n15094) );
  AND2_X1 U17080 ( .A1(n13341), .A2(n15094), .ZN(n15338) );
  NOR2_X1 U17081 ( .A1(n15095), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n15100) );
  AOI21_X1 U17082 ( .B1(n22396), .B2(n15338), .A(n15100), .ZN(n15102) );
  INV_X1 U17083 ( .A(n15102), .ZN(n15096) );
  NAND2_X1 U17084 ( .A1(n15096), .A2(n15786), .ZN(n15098) );
  NOR3_X1 U17085 ( .A1(n17795), .A2(n22374), .A3(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n22398) );
  NAND2_X1 U17086 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n22398), .ZN(n15097) );
  AND2_X1 U17087 ( .A1(n15098), .A2(n15097), .ZN(n15170) );
  INV_X1 U17088 ( .A(n15100), .ZN(n15169) );
  OAI22_X1 U17089 ( .A1(n22667), .A2(n15170), .B1(n22639), .B2(n15169), .ZN(
        n15101) );
  AOI21_X1 U17090 ( .B1(n22531), .B2(n22675), .A(n15101), .ZN(n15106) );
  NAND3_X1 U17091 ( .A1(n15103), .A2(n15786), .A3(n15102), .ZN(n15104) );
  NAND2_X1 U17092 ( .A1(n15172), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n15105) );
  OAI211_X1 U17093 ( .C1(n15175), .C2(n22681), .A(n15106), .B(n15105), .ZN(
        P1_U3096) );
  INV_X1 U17094 ( .A(n15108), .ZN(n15109) );
  OAI21_X1 U17095 ( .B1(n15107), .B2(n15110), .A(n15109), .ZN(n18986) );
  OAI222_X1 U17096 ( .A1(n15600), .A2(n15111), .B1(n18986), .B2(n20018), .C1(
        n17952), .C2(n16817), .ZN(P2_U2904) );
  INV_X1 U17097 ( .A(DATAI_28_), .ZN(n15113) );
  INV_X1 U17098 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n20659) );
  OR2_X1 U17099 ( .A1(n15161), .A2(n20659), .ZN(n15112) );
  OAI21_X1 U17100 ( .B1(n15164), .B2(n15113), .A(n15112), .ZN(n22555) );
  INV_X1 U17101 ( .A(n22555), .ZN(n22536) );
  NAND2_X1 U17102 ( .A1(n15172), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n15118) );
  INV_X1 U17103 ( .A(DATAI_20_), .ZN(n15114) );
  INV_X1 U17104 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n20642) );
  OAI22_X1 U17105 ( .A1(n15114), .A2(n15164), .B1(n20642), .B2(n15161), .ZN(
        n22547) );
  NOR2_X1 U17106 ( .A1(n15987), .A2(DATAI_4_), .ZN(n15115) );
  AOI21_X1 U17107 ( .B1(n15987), .B2(n20611), .A(n15115), .ZN(n16235) );
  NAND2_X1 U17108 ( .A1(n15124), .A2(n16235), .ZN(n22550) );
  OAI22_X1 U17109 ( .A1(n22535), .A2(n15169), .B1(n22550), .B2(n15170), .ZN(
        n15116) );
  AOI21_X1 U17110 ( .B1(n22531), .B2(n22547), .A(n15116), .ZN(n15117) );
  OAI211_X1 U17111 ( .C1(n22536), .C2(n15175), .A(n15118), .B(n15117), .ZN(
        P1_U3093) );
  INV_X1 U17112 ( .A(DATAI_29_), .ZN(n15120) );
  INV_X1 U17113 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20661) );
  OR2_X1 U17114 ( .A1(n15161), .A2(n20661), .ZN(n15119) );
  OAI21_X1 U17115 ( .B1(n15164), .B2(n15120), .A(n15119), .ZN(n22580) );
  INV_X1 U17116 ( .A(n22580), .ZN(n22574) );
  NAND2_X1 U17117 ( .A1(n15172), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n15127) );
  INV_X1 U17118 ( .A(DATAI_21_), .ZN(n15122) );
  INV_X1 U17119 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20644) );
  OR2_X1 U17120 ( .A1(n15161), .A2(n20644), .ZN(n15121) );
  OAI21_X1 U17121 ( .B1(n15164), .B2(n15122), .A(n15121), .ZN(n22579) );
  NOR2_X1 U17122 ( .A1(n15168), .A2(n16022), .ZN(n22578) );
  INV_X1 U17123 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n20613) );
  NOR2_X1 U17124 ( .A1(n15987), .A2(DATAI_5_), .ZN(n15123) );
  AOI21_X1 U17125 ( .B1(n15987), .B2(n20613), .A(n15123), .ZN(n16231) );
  NAND2_X1 U17126 ( .A1(n15124), .A2(n16231), .ZN(n22583) );
  OAI22_X1 U17127 ( .A1(n22573), .A2(n15169), .B1(n22583), .B2(n15170), .ZN(
        n15125) );
  AOI21_X1 U17128 ( .B1(n22531), .B2(n22579), .A(n15125), .ZN(n15126) );
  OAI211_X1 U17129 ( .C1(n22574), .C2(n15175), .A(n15127), .B(n15126), .ZN(
        P1_U3094) );
  INV_X1 U17130 ( .A(DATAI_26_), .ZN(n15129) );
  INV_X1 U17131 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n20655) );
  OR2_X1 U17132 ( .A1(n15161), .A2(n20655), .ZN(n15128) );
  OAI21_X1 U17133 ( .B1(n15164), .B2(n15129), .A(n15128), .ZN(n22489) );
  INV_X1 U17134 ( .A(n22489), .ZN(n22483) );
  INV_X1 U17135 ( .A(DATAI_18_), .ZN(n15131) );
  INV_X1 U17136 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n20638) );
  OR2_X1 U17137 ( .A1(n15161), .A2(n20638), .ZN(n15130) );
  OAI21_X1 U17138 ( .B1(n15164), .B2(n15131), .A(n15130), .ZN(n22488) );
  NOR2_X1 U17139 ( .A1(n15168), .A2(n14899), .ZN(n22487) );
  OAI22_X1 U17140 ( .A1(n22492), .A2(n15170), .B1(n22482), .B2(n15169), .ZN(
        n15132) );
  AOI21_X1 U17141 ( .B1(n22531), .B2(n22488), .A(n15132), .ZN(n15134) );
  NAND2_X1 U17142 ( .A1(n15172), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n15133) );
  OAI211_X1 U17143 ( .C1(n22483), .C2(n15175), .A(n15134), .B(n15133), .ZN(
        P1_U3091) );
  INV_X1 U17144 ( .A(DATAI_25_), .ZN(n15136) );
  INV_X1 U17145 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n20653) );
  OR2_X1 U17146 ( .A1(n15161), .A2(n20653), .ZN(n15135) );
  OAI21_X1 U17147 ( .B1(n15164), .B2(n15136), .A(n15135), .ZN(n22466) );
  INV_X1 U17148 ( .A(n22466), .ZN(n22460) );
  INV_X1 U17149 ( .A(DATAI_17_), .ZN(n15138) );
  INV_X1 U17150 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n20636) );
  OR2_X1 U17151 ( .A1(n15161), .A2(n20636), .ZN(n15137) );
  OAI21_X1 U17152 ( .B1(n15164), .B2(n15138), .A(n15137), .ZN(n22465) );
  NOR2_X1 U17153 ( .A1(n15168), .A2(n15379), .ZN(n22464) );
  OAI22_X1 U17154 ( .A1(n22469), .A2(n15170), .B1(n22459), .B2(n15169), .ZN(
        n15139) );
  AOI21_X1 U17155 ( .B1(n22531), .B2(n22465), .A(n15139), .ZN(n15141) );
  NAND2_X1 U17156 ( .A1(n15172), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n15140) );
  OAI211_X1 U17157 ( .C1(n22460), .C2(n15175), .A(n15141), .B(n15140), .ZN(
        P1_U3090) );
  INV_X1 U17158 ( .A(DATAI_24_), .ZN(n15143) );
  INV_X1 U17159 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n20651) );
  OR2_X1 U17160 ( .A1(n15161), .A2(n20651), .ZN(n15142) );
  OAI21_X1 U17161 ( .B1(n15164), .B2(n15143), .A(n15142), .ZN(n22442) );
  INV_X1 U17162 ( .A(n22442), .ZN(n22401) );
  INV_X1 U17163 ( .A(DATAI_16_), .ZN(n15145) );
  INV_X1 U17164 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n20634) );
  OR2_X1 U17165 ( .A1(n15161), .A2(n20634), .ZN(n15144) );
  OAI21_X1 U17166 ( .B1(n15164), .B2(n15145), .A(n15144), .ZN(n22434) );
  NOR2_X1 U17167 ( .A1(n15168), .A2(n15146), .ZN(n22433) );
  OAI22_X1 U17168 ( .A1(n22445), .A2(n15170), .B1(n22400), .B2(n15169), .ZN(
        n15147) );
  AOI21_X1 U17169 ( .B1(n22531), .B2(n22434), .A(n15147), .ZN(n15149) );
  NAND2_X1 U17170 ( .A1(n15172), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n15148) );
  OAI211_X1 U17171 ( .C1(n22401), .C2(n15175), .A(n15149), .B(n15148), .ZN(
        P1_U3089) );
  INV_X1 U17172 ( .A(DATAI_30_), .ZN(n15151) );
  INV_X1 U17173 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20665) );
  OR2_X1 U17174 ( .A1(n15161), .A2(n20665), .ZN(n15150) );
  OAI21_X1 U17175 ( .B1(n15164), .B2(n15151), .A(n15150), .ZN(n22610) );
  INV_X1 U17176 ( .A(n22610), .ZN(n22603) );
  INV_X1 U17177 ( .A(DATAI_22_), .ZN(n15153) );
  INV_X1 U17178 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n20646) );
  OR2_X1 U17179 ( .A1(n15161), .A2(n20646), .ZN(n15152) );
  OAI21_X1 U17180 ( .B1(n15164), .B2(n15153), .A(n15152), .ZN(n22609) );
  NAND2_X1 U17181 ( .A1(n15991), .A2(DATAI_6_), .ZN(n15155) );
  NAND2_X1 U17182 ( .A1(n15987), .A2(BUF1_REG_6__SCAN_IN), .ZN(n15154) );
  AND2_X1 U17183 ( .A1(n15155), .A2(n15154), .ZN(n15559) );
  NOR2_X1 U17184 ( .A1(n15168), .A2(n16023), .ZN(n22608) );
  OAI22_X1 U17185 ( .A1(n22613), .A2(n15170), .B1(n22601), .B2(n15169), .ZN(
        n15156) );
  AOI21_X1 U17186 ( .B1(n22531), .B2(n22609), .A(n15156), .ZN(n15158) );
  NAND2_X1 U17187 ( .A1(n15172), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n15157) );
  OAI211_X1 U17188 ( .C1(n22603), .C2(n15175), .A(n15158), .B(n15157), .ZN(
        P1_U3095) );
  INV_X1 U17189 ( .A(DATAI_27_), .ZN(n15160) );
  INV_X1 U17190 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n20657) );
  OR2_X1 U17191 ( .A1(n15161), .A2(n20657), .ZN(n15159) );
  OAI21_X1 U17192 ( .B1(n15164), .B2(n15160), .A(n15159), .ZN(n22513) );
  INV_X1 U17193 ( .A(n22513), .ZN(n22507) );
  INV_X1 U17194 ( .A(DATAI_19_), .ZN(n15163) );
  INV_X1 U17195 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n20640) );
  OR2_X1 U17196 ( .A1(n15161), .A2(n20640), .ZN(n15162) );
  OAI21_X1 U17197 ( .B1(n15164), .B2(n15163), .A(n15162), .ZN(n22512) );
  NAND2_X1 U17198 ( .A1(n15991), .A2(DATAI_3_), .ZN(n15166) );
  NAND2_X1 U17199 ( .A1(n15987), .A2(BUF1_REG_3__SCAN_IN), .ZN(n15165) );
  AND2_X1 U17200 ( .A1(n15166), .A2(n15165), .ZN(n15492) );
  NOR2_X1 U17201 ( .A1(n15168), .A2(n15167), .ZN(n22511) );
  OAI22_X1 U17202 ( .A1(n22516), .A2(n15170), .B1(n22506), .B2(n15169), .ZN(
        n15171) );
  AOI21_X1 U17203 ( .B1(n22531), .B2(n22512), .A(n15171), .ZN(n15174) );
  NAND2_X1 U17204 ( .A1(n15172), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n15173) );
  OAI211_X1 U17205 ( .C1(n22507), .C2(n15175), .A(n15174), .B(n15173), .ZN(
        P1_U3092) );
  NOR2_X1 U17206 ( .A1(n22370), .A2(n14966), .ZN(n15176) );
  NAND2_X1 U17207 ( .A1(n15176), .A2(n13338), .ZN(n22366) );
  NAND2_X1 U17208 ( .A1(n15176), .A2(n15568), .ZN(n22623) );
  NOR3_X1 U17209 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n22360) );
  INV_X1 U17210 ( .A(n15337), .ZN(n15177) );
  INV_X1 U17211 ( .A(n22382), .ZN(n15178) );
  INV_X1 U17212 ( .A(n15454), .ZN(n15571) );
  INV_X1 U17213 ( .A(n22360), .ZN(n15180) );
  NOR2_X1 U17214 ( .A1(n22415), .A2(n15180), .ZN(n15197) );
  AOI21_X1 U17215 ( .B1(n15178), .B2(n15571), .A(n15197), .ZN(n15181) );
  OAI211_X1 U17216 ( .C1(n22370), .C2(n22286), .A(n15786), .B(n15181), .ZN(
        n15179) );
  OAI211_X1 U17217 ( .C1(n15786), .C2(n22360), .A(n22387), .B(n15179), .ZN(
        n15196) );
  AOI22_X1 U17218 ( .A1(n22589), .A2(n22579), .B1(n15196), .B2(
        P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15183) );
  OAI22_X1 U17219 ( .A1(n15181), .A2(n22424), .B1(n15180), .B2(n15575), .ZN(
        n15198) );
  INV_X1 U17220 ( .A(n22583), .ZN(n15587) );
  AOI22_X1 U17221 ( .A1(n15198), .A2(n15587), .B1(n22578), .B2(n15197), .ZN(
        n15182) );
  OAI211_X1 U17222 ( .C1(n22574), .C2(n22366), .A(n15183), .B(n15182), .ZN(
        P1_U3046) );
  AOI22_X1 U17223 ( .A1(n22589), .A2(n22512), .B1(n15196), .B2(
        P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15185) );
  AOI22_X1 U17224 ( .A1(n16643), .A2(n15198), .B1(n22511), .B2(n15197), .ZN(
        n15184) );
  OAI211_X1 U17225 ( .C1(n22507), .C2(n22366), .A(n15185), .B(n15184), .ZN(
        P1_U3044) );
  AOI22_X1 U17226 ( .A1(n22589), .A2(n22609), .B1(n15196), .B2(
        P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n15187) );
  AOI22_X1 U17227 ( .A1(n16648), .A2(n15198), .B1(n22608), .B2(n15197), .ZN(
        n15186) );
  OAI211_X1 U17228 ( .C1(n22603), .C2(n22366), .A(n15187), .B(n15186), .ZN(
        P1_U3047) );
  AOI22_X1 U17229 ( .A1(n22589), .A2(n22488), .B1(n15196), .B2(
        P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15189) );
  AOI22_X1 U17230 ( .A1(n16638), .A2(n15198), .B1(n22487), .B2(n15197), .ZN(
        n15188) );
  OAI211_X1 U17231 ( .C1(n22483), .C2(n22366), .A(n15189), .B(n15188), .ZN(
        P1_U3043) );
  AOI22_X1 U17232 ( .A1(n22589), .A2(n22465), .B1(n15196), .B2(
        P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15191) );
  AOI22_X1 U17233 ( .A1(n16633), .A2(n15198), .B1(n22464), .B2(n15197), .ZN(
        n15190) );
  OAI211_X1 U17234 ( .C1(n22460), .C2(n22366), .A(n15191), .B(n15190), .ZN(
        P1_U3042) );
  AOI22_X1 U17235 ( .A1(n22589), .A2(n22434), .B1(n15196), .B2(
        P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15193) );
  AOI22_X1 U17236 ( .A1(n16628), .A2(n15198), .B1(n22433), .B2(n15197), .ZN(
        n15192) );
  OAI211_X1 U17237 ( .C1(n22401), .C2(n22366), .A(n15193), .B(n15192), .ZN(
        P1_U3041) );
  AOI22_X1 U17238 ( .A1(n22589), .A2(n22675), .B1(n15196), .B2(
        P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15195) );
  AOI22_X1 U17239 ( .A1(n22674), .A2(n15198), .B1(n22671), .B2(n15197), .ZN(
        n15194) );
  OAI211_X1 U17240 ( .C1(n22681), .C2(n22366), .A(n15195), .B(n15194), .ZN(
        P1_U3048) );
  AOI22_X1 U17241 ( .A1(n22589), .A2(n22547), .B1(n15196), .B2(
        P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15200) );
  INV_X1 U17242 ( .A(n22550), .ZN(n22552) );
  AOI22_X1 U17243 ( .A1(n15198), .A2(n22552), .B1(n22554), .B2(n15197), .ZN(
        n15199) );
  OAI211_X1 U17244 ( .C1(n22536), .C2(n22366), .A(n15200), .B(n15199), .ZN(
        P1_U3045) );
  INV_X1 U17245 ( .A(n17323), .ZN(n18873) );
  AOI21_X1 U17246 ( .B1(n18873), .B2(n19820), .A(n15201), .ZN(n15413) );
  XNOR2_X1 U17247 ( .A(n15202), .B(n15203), .ZN(n17889) );
  INV_X1 U17248 ( .A(n17889), .ZN(n15751) );
  XNOR2_X1 U17249 ( .A(n15413), .B(n15751), .ZN(n15412) );
  XNOR2_X1 U17250 ( .A(n15412), .B(n19879), .ZN(n15204) );
  NAND2_X1 U17251 ( .A1(n15204), .A2(n20068), .ZN(n15206) );
  AOI22_X1 U17252 ( .A1(n20067), .A2(n17889), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n20060), .ZN(n15205) );
  OAI211_X1 U17253 ( .C1(n20153), .C2(n15600), .A(n15206), .B(n15205), .ZN(
        P2_U2917) );
  XOR2_X1 U17254 ( .A(n15207), .B(n15208), .Z(n15384) );
  INV_X1 U17255 ( .A(n15384), .ZN(n15375) );
  OAI222_X1 U17256 ( .A1(n15375), .A2(n16238), .B1(n16268), .B2(n15492), .C1(
        n16265), .C2(n13322), .ZN(P1_U2901) );
  OR2_X1 U17257 ( .A1(n15210), .A2(n15209), .ZN(n15211) );
  NAND2_X1 U17258 ( .A1(n15212), .A2(n15211), .ZN(n21915) );
  AOI22_X1 U17259 ( .A1(n20588), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n22052), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n15213) );
  OAI21_X1 U17260 ( .B1(n20594), .B2(n15286), .A(n15213), .ZN(n15214) );
  AOI21_X1 U17261 ( .B1(n15276), .B2(n20555), .A(n15214), .ZN(n15215) );
  OAI21_X1 U17262 ( .B1(n22268), .B2(n21915), .A(n15215), .ZN(P1_U2997) );
  OAI21_X1 U17263 ( .B1(n15218), .B2(n15217), .A(n15216), .ZN(n21932) );
  AOI22_X1 U17264 ( .A1(n20588), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n22052), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n15219) );
  OAI21_X1 U17265 ( .B1(n20594), .B2(n15395), .A(n15219), .ZN(n15220) );
  AOI21_X1 U17266 ( .B1(n15384), .B2(n20555), .A(n15220), .ZN(n15221) );
  OAI21_X1 U17267 ( .B1(n21932), .B2(n22268), .A(n15221), .ZN(P1_U2996) );
  NAND2_X1 U17268 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n22278), .ZN(n17819) );
  INV_X1 U17269 ( .A(n17819), .ZN(n15222) );
  AND2_X1 U17270 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n22274), .ZN(n15223) );
  NAND2_X1 U17271 ( .A1(n13791), .A2(n15223), .ZN(n15224) );
  NOR2_X1 U17272 ( .A1(n15243), .A2(n17825), .ZN(n15226) );
  NAND2_X1 U17273 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n22104), .ZN(n15238) );
  NOR2_X1 U17274 ( .A1(n16037), .A2(n15238), .ZN(n15227) );
  OR2_X1 U17275 ( .A1(n22262), .A2(n15227), .ZN(n22099) );
  INV_X1 U17276 ( .A(n22099), .ZN(n22085) );
  AND2_X1 U17277 ( .A1(n15229), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n15230) );
  NAND2_X1 U17278 ( .A1(n16021), .A2(n15233), .ZN(n15232) );
  NOR2_X1 U17279 ( .A1(n15230), .A2(n15232), .ZN(n15231) );
  NAND2_X1 U17280 ( .A1(n22104), .A2(n22220), .ZN(n22166) );
  NAND2_X1 U17281 ( .A1(P1_EBX_REG_31__SCAN_IN), .A2(n15233), .ZN(n15234) );
  AOI21_X1 U17282 ( .B1(n21876), .B2(n22286), .A(n15234), .ZN(n15235) );
  OAI22_X1 U17283 ( .A1(n22177), .A2(n15237), .B1(n22267), .B2(n15236), .ZN(
        n15242) );
  NOR2_X1 U17284 ( .A1(n15239), .A2(n15238), .ZN(n22074) );
  INV_X1 U17285 ( .A(n22074), .ZN(n15277) );
  NOR2_X1 U17286 ( .A1(n15240), .A2(n15277), .ZN(n15241) );
  AOI211_X1 U17287 ( .C1(n22235), .C2(P1_EBX_REG_0__SCAN_IN), .A(n15242), .B(
        n15241), .ZN(n15246) );
  OAI21_X1 U17288 ( .B1(n22244), .B2(n22260), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15245) );
  OAI211_X1 U17289 ( .C1(n22085), .C2(n15247), .A(n15246), .B(n15245), .ZN(
        P1_U2840) );
  NOR3_X1 U17290 ( .A1(n15570), .A2(n17795), .A3(n22374), .ZN(n15544) );
  INV_X1 U17291 ( .A(n15338), .ZN(n22381) );
  OR2_X1 U17292 ( .A1(n22428), .A2(n22381), .ZN(n15249) );
  NAND2_X1 U17293 ( .A1(n15249), .A2(n22670), .ZN(n15254) );
  INV_X1 U17294 ( .A(n15254), .ZN(n15251) );
  NAND2_X1 U17295 ( .A1(n15251), .A2(n15250), .ZN(n15252) );
  OR2_X1 U17296 ( .A1(n22424), .A2(n15252), .ZN(n15253) );
  OAI211_X1 U17297 ( .C1(n15786), .C2(n15544), .A(n22387), .B(n15253), .ZN(
        n22677) );
  NAND2_X1 U17298 ( .A1(n14966), .A2(n13338), .ZN(n22369) );
  NAND2_X1 U17299 ( .A1(n14966), .A2(n15568), .ZN(n15655) );
  INV_X1 U17300 ( .A(n22465), .ZN(n22452) );
  OAI22_X1 U17301 ( .A1(n22460), .A2(n22680), .B1(n22615), .B2(n22452), .ZN(
        n15256) );
  AOI22_X1 U17302 ( .A1(n15254), .A2(n15786), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15544), .ZN(n22669) );
  OAI22_X1 U17303 ( .A1(n22469), .A2(n22669), .B1(n22670), .B2(n22459), .ZN(
        n15255) );
  AOI211_X1 U17304 ( .C1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .C2(n22677), .A(
        n15256), .B(n15255), .ZN(n15257) );
  INV_X1 U17305 ( .A(n15257), .ZN(P1_U3154) );
  OAI22_X1 U17306 ( .A1(n22573), .A2(n22670), .B1(n22583), .B2(n22669), .ZN(
        n15259) );
  INV_X1 U17307 ( .A(n22579), .ZN(n22567) );
  OAI22_X1 U17308 ( .A1(n22574), .A2(n22680), .B1(n22615), .B2(n22567), .ZN(
        n15258) );
  AOI211_X1 U17309 ( .C1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .C2(n22677), .A(
        n15259), .B(n15258), .ZN(n15260) );
  INV_X1 U17310 ( .A(n15260), .ZN(P1_U3158) );
  INV_X1 U17311 ( .A(n22488), .ZN(n22476) );
  OAI22_X1 U17312 ( .A1(n22483), .A2(n22680), .B1(n22615), .B2(n22476), .ZN(
        n15262) );
  OAI22_X1 U17313 ( .A1(n22492), .A2(n22669), .B1(n22670), .B2(n22482), .ZN(
        n15261) );
  AOI211_X1 U17314 ( .C1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .C2(n22677), .A(
        n15262), .B(n15261), .ZN(n15263) );
  INV_X1 U17315 ( .A(n15263), .ZN(P1_U3155) );
  INV_X1 U17316 ( .A(n22609), .ZN(n22587) );
  OAI22_X1 U17317 ( .A1(n22603), .A2(n22680), .B1(n22615), .B2(n22587), .ZN(
        n15265) );
  OAI22_X1 U17318 ( .A1(n22613), .A2(n22669), .B1(n22670), .B2(n22601), .ZN(
        n15264) );
  AOI211_X1 U17319 ( .C1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .C2(n22677), .A(
        n15265), .B(n15264), .ZN(n15266) );
  INV_X1 U17320 ( .A(n15266), .ZN(P1_U3159) );
  INV_X1 U17321 ( .A(n22512), .ZN(n22499) );
  OAI22_X1 U17322 ( .A1(n22507), .A2(n22680), .B1(n22615), .B2(n22499), .ZN(
        n15268) );
  OAI22_X1 U17323 ( .A1(n22516), .A2(n22669), .B1(n22670), .B2(n22506), .ZN(
        n15267) );
  AOI211_X1 U17324 ( .C1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .C2(n22677), .A(
        n15268), .B(n15267), .ZN(n15269) );
  INV_X1 U17325 ( .A(n15269), .ZN(P1_U3156) );
  OAI22_X1 U17326 ( .A1(n22535), .A2(n22670), .B1(n22550), .B2(n22669), .ZN(
        n15271) );
  OAI22_X1 U17327 ( .A1(n22536), .A2(n22680), .B1(n22615), .B2(n22560), .ZN(
        n15270) );
  AOI211_X1 U17328 ( .C1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .C2(n22677), .A(
        n15271), .B(n15270), .ZN(n15272) );
  INV_X1 U17329 ( .A(n15272), .ZN(P1_U3157) );
  INV_X1 U17330 ( .A(n22434), .ZN(n15810) );
  OAI22_X1 U17331 ( .A1(n22401), .A2(n22680), .B1(n22615), .B2(n15810), .ZN(
        n15274) );
  OAI22_X1 U17332 ( .A1(n22445), .A2(n22669), .B1(n22670), .B2(n22400), .ZN(
        n15273) );
  AOI211_X1 U17333 ( .C1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .C2(n22677), .A(
        n15274), .B(n15273), .ZN(n15275) );
  INV_X1 U17334 ( .A(n15275), .ZN(P1_U3153) );
  NAND2_X1 U17335 ( .A1(n15276), .A2(n22099), .ZN(n15285) );
  NOR2_X1 U17336 ( .A1(n15337), .A2(n15277), .ZN(n15283) );
  OAI21_X1 U17337 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n22220), .A(n22104), .ZN(
        n15278) );
  AOI22_X1 U17338 ( .A1(n22235), .A2(P1_EBX_REG_2__SCAN_IN), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n15278), .ZN(n15281) );
  INV_X1 U17339 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n15279) );
  NAND3_X1 U17340 ( .A1(n22236), .A2(P1_REIP_REG_1__SCAN_IN), .A3(n15279), 
        .ZN(n15280) );
  OAI211_X1 U17341 ( .C1(n21919), .C2(n22267), .A(n15281), .B(n15280), .ZN(
        n15282) );
  AOI211_X1 U17342 ( .C1(n22244), .C2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n15283), .B(n15282), .ZN(n15284) );
  OAI211_X1 U17343 ( .C1(n22251), .C2(n15286), .A(n15285), .B(n15284), .ZN(
        P1_U2838) );
  OR3_X1 U17344 ( .A1(n17795), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n15657) );
  NAND3_X1 U17345 ( .A1(n15291), .A2(n15786), .A3(n15288), .ZN(n15290) );
  INV_X1 U17346 ( .A(n22387), .ZN(n15289) );
  INV_X1 U17347 ( .A(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15296) );
  NOR2_X1 U17348 ( .A1(n22415), .A2(n15657), .ZN(n15321) );
  AOI21_X1 U17349 ( .B1(n22396), .B2(n15571), .A(n15321), .ZN(n15292) );
  OAI22_X1 U17350 ( .A1(n15292), .A2(n22424), .B1(n15657), .B2(n15575), .ZN(
        n15322) );
  AOI22_X1 U17351 ( .A1(n22578), .A2(n15321), .B1(n15587), .B2(n15322), .ZN(
        n15293) );
  OAI21_X1 U17352 ( .B1(n22640), .B2(n22567), .A(n15293), .ZN(n15294) );
  AOI21_X1 U17353 ( .B1(n15688), .B2(n22580), .A(n15294), .ZN(n15295) );
  OAI21_X1 U17354 ( .B1(n15327), .B2(n15296), .A(n15295), .ZN(P1_U3078) );
  INV_X1 U17355 ( .A(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15300) );
  AOI22_X1 U17356 ( .A1(n22554), .A2(n15321), .B1(n22552), .B2(n15322), .ZN(
        n15297) );
  OAI21_X1 U17357 ( .B1(n22640), .B2(n22560), .A(n15297), .ZN(n15298) );
  AOI21_X1 U17358 ( .B1(n15688), .B2(n22555), .A(n15298), .ZN(n15299) );
  OAI21_X1 U17359 ( .B1(n15327), .B2(n15300), .A(n15299), .ZN(P1_U3077) );
  INV_X1 U17360 ( .A(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15304) );
  AOI22_X1 U17361 ( .A1(n16643), .A2(n15322), .B1(n22511), .B2(n15321), .ZN(
        n15301) );
  OAI21_X1 U17362 ( .B1(n22640), .B2(n22499), .A(n15301), .ZN(n15302) );
  AOI21_X1 U17363 ( .B1(n15688), .B2(n22513), .A(n15302), .ZN(n15303) );
  OAI21_X1 U17364 ( .B1(n15327), .B2(n15304), .A(n15303), .ZN(P1_U3076) );
  INV_X1 U17365 ( .A(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15308) );
  AOI22_X1 U17366 ( .A1(n16638), .A2(n15322), .B1(n22487), .B2(n15321), .ZN(
        n15305) );
  OAI21_X1 U17367 ( .B1(n22640), .B2(n22476), .A(n15305), .ZN(n15306) );
  AOI21_X1 U17368 ( .B1(n15688), .B2(n22489), .A(n15306), .ZN(n15307) );
  OAI21_X1 U17369 ( .B1(n15327), .B2(n15308), .A(n15307), .ZN(P1_U3075) );
  INV_X1 U17370 ( .A(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15312) );
  INV_X1 U17371 ( .A(n22675), .ZN(n22630) );
  AOI22_X1 U17372 ( .A1(n22674), .A2(n15322), .B1(n22671), .B2(n15321), .ZN(
        n15309) );
  OAI21_X1 U17373 ( .B1(n22640), .B2(n22630), .A(n15309), .ZN(n15310) );
  AOI21_X1 U17374 ( .B1(n15688), .B2(n22662), .A(n15310), .ZN(n15311) );
  OAI21_X1 U17375 ( .B1(n15327), .B2(n15312), .A(n15311), .ZN(P1_U3080) );
  INV_X1 U17376 ( .A(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n15316) );
  AOI22_X1 U17377 ( .A1(n16633), .A2(n15322), .B1(n22464), .B2(n15321), .ZN(
        n15313) );
  OAI21_X1 U17378 ( .B1(n22640), .B2(n22452), .A(n15313), .ZN(n15314) );
  AOI21_X1 U17379 ( .B1(n15688), .B2(n22466), .A(n15314), .ZN(n15315) );
  OAI21_X1 U17380 ( .B1(n15327), .B2(n15316), .A(n15315), .ZN(P1_U3074) );
  INV_X1 U17381 ( .A(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15320) );
  AOI22_X1 U17382 ( .A1(n16628), .A2(n15322), .B1(n22433), .B2(n15321), .ZN(
        n15317) );
  OAI21_X1 U17383 ( .B1(n22640), .B2(n15810), .A(n15317), .ZN(n15318) );
  AOI21_X1 U17384 ( .B1(n15688), .B2(n22442), .A(n15318), .ZN(n15319) );
  OAI21_X1 U17385 ( .B1(n15327), .B2(n15320), .A(n15319), .ZN(P1_U3073) );
  INV_X1 U17386 ( .A(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n15326) );
  AOI22_X1 U17387 ( .A1(n16648), .A2(n15322), .B1(n22608), .B2(n15321), .ZN(
        n15323) );
  OAI21_X1 U17388 ( .B1(n22640), .B2(n22587), .A(n15323), .ZN(n15324) );
  AOI21_X1 U17389 ( .B1(n15688), .B2(n22610), .A(n15324), .ZN(n15325) );
  OAI21_X1 U17390 ( .B1(n15327), .B2(n15326), .A(n15325), .ZN(P1_U3079) );
  INV_X1 U17391 ( .A(n16235), .ZN(n15332) );
  INV_X1 U17392 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20421) );
  AND2_X1 U17393 ( .A1(n15330), .A2(n15329), .ZN(n15331) );
  OR2_X1 U17394 ( .A1(n15328), .A2(n15331), .ZN(n22086) );
  OAI222_X1 U17395 ( .A1(n16268), .A2(n15332), .B1(n16265), .B2(n20421), .C1(
        n16238), .C2(n22086), .ZN(P1_U2900) );
  INV_X1 U17396 ( .A(n22370), .ZN(n15334) );
  AOI21_X1 U17397 ( .B1(n15334), .B2(n15335), .A(n22424), .ZN(n22386) );
  AND3_X1 U17398 ( .A1(n22386), .A2(n15335), .A3(n14999), .ZN(n15336) );
  NOR3_X1 U17399 ( .A1(n15570), .A2(n22374), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n22414) );
  NAND2_X1 U17400 ( .A1(n22543), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n15346) );
  AND2_X1 U17401 ( .A1(n16621), .A2(n15337), .ZN(n22410) );
  NAND2_X1 U17402 ( .A1(n22410), .A2(n15338), .ZN(n15340) );
  INV_X1 U17403 ( .A(n22414), .ZN(n15339) );
  NOR2_X1 U17404 ( .A1(n22415), .A2(n15339), .ZN(n22541) );
  INV_X1 U17405 ( .A(n22541), .ZN(n15369) );
  NAND2_X1 U17406 ( .A1(n15340), .A2(n15369), .ZN(n15341) );
  NAND2_X1 U17407 ( .A1(n15341), .A2(n15786), .ZN(n15343) );
  NAND2_X1 U17408 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n22414), .ZN(n15342) );
  AND2_X1 U17409 ( .A1(n15343), .A2(n15342), .ZN(n22540) );
  OAI22_X1 U17410 ( .A1(n22445), .A2(n22540), .B1(n22400), .B2(n15369), .ZN(
        n15344) );
  AOI21_X1 U17411 ( .B1(n22654), .B2(n22442), .A(n15344), .ZN(n15345) );
  OAI211_X1 U17412 ( .C1(n15810), .C2(n22546), .A(n15346), .B(n15345), .ZN(
        P1_U3121) );
  NAND2_X1 U17413 ( .A1(n22543), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n15349) );
  OAI22_X1 U17414 ( .A1(n22573), .A2(n15369), .B1(n22583), .B2(n22540), .ZN(
        n15347) );
  AOI21_X1 U17415 ( .B1(n22654), .B2(n22580), .A(n15347), .ZN(n15348) );
  OAI211_X1 U17416 ( .C1(n22567), .C2(n22546), .A(n15349), .B(n15348), .ZN(
        P1_U3126) );
  NAND2_X1 U17417 ( .A1(n22543), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n15352) );
  OAI22_X1 U17418 ( .A1(n22469), .A2(n22540), .B1(n22459), .B2(n15369), .ZN(
        n15350) );
  AOI21_X1 U17419 ( .B1(n22654), .B2(n22466), .A(n15350), .ZN(n15351) );
  OAI211_X1 U17420 ( .C1(n22452), .C2(n22546), .A(n15352), .B(n15351), .ZN(
        P1_U3122) );
  NAND2_X1 U17421 ( .A1(n22543), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n15355) );
  OAI22_X1 U17422 ( .A1(n22667), .A2(n22540), .B1(n22639), .B2(n15369), .ZN(
        n15353) );
  AOI21_X1 U17423 ( .B1(n22662), .B2(n22654), .A(n15353), .ZN(n15354) );
  OAI211_X1 U17424 ( .C1(n22630), .C2(n22546), .A(n15355), .B(n15354), .ZN(
        P1_U3128) );
  AND2_X1 U17425 ( .A1(n15404), .A2(n15356), .ZN(n15357) );
  OR2_X1 U17426 ( .A1(n15357), .A2(n15626), .ZN(n17246) );
  OAI211_X1 U17427 ( .C1(n15358), .C2(n15360), .A(n15359), .B(n16732), .ZN(
        n15362) );
  NAND2_X1 U17428 ( .A1(n11141), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n15361) );
  OAI211_X1 U17429 ( .C1(n17246), .C2(n11141), .A(n15362), .B(n15361), .ZN(
        P2_U2875) );
  NAND2_X1 U17430 ( .A1(n22543), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n15365) );
  OAI22_X1 U17431 ( .A1(n22492), .A2(n22540), .B1(n22482), .B2(n15369), .ZN(
        n15363) );
  AOI21_X1 U17432 ( .B1(n22654), .B2(n22489), .A(n15363), .ZN(n15364) );
  OAI211_X1 U17433 ( .C1(n22476), .C2(n22546), .A(n15365), .B(n15364), .ZN(
        P1_U3123) );
  NAND2_X1 U17434 ( .A1(n22543), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n15368) );
  OAI22_X1 U17435 ( .A1(n22516), .A2(n22540), .B1(n22506), .B2(n15369), .ZN(
        n15366) );
  AOI21_X1 U17436 ( .B1(n22654), .B2(n22513), .A(n15366), .ZN(n15367) );
  OAI211_X1 U17437 ( .C1(n22499), .C2(n22546), .A(n15368), .B(n15367), .ZN(
        P1_U3124) );
  NAND2_X1 U17438 ( .A1(n22543), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n15372) );
  OAI22_X1 U17439 ( .A1(n22613), .A2(n22540), .B1(n22601), .B2(n15369), .ZN(
        n15370) );
  AOI21_X1 U17440 ( .B1(n22654), .B2(n22610), .A(n15370), .ZN(n15371) );
  OAI211_X1 U17441 ( .C1(n22587), .C2(n22546), .A(n15372), .B(n15371), .ZN(
        P1_U3127) );
  AOI21_X1 U17442 ( .B1(n15374), .B2(n15373), .A(n15397), .ZN(n21931) );
  INV_X1 U17443 ( .A(n21931), .ZN(n15389) );
  INV_X1 U17444 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n15376) );
  OAI222_X1 U17445 ( .A1(n15389), .A2(n20510), .B1(n15376), .B2(n20524), .C1(
        n16189), .C2(n15375), .ZN(P1_U2869) );
  INV_X1 U17446 ( .A(n15522), .ZN(n15383) );
  INV_X1 U17447 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n20632) );
  NAND2_X1 U17448 ( .A1(n15987), .A2(n20632), .ZN(n15380) );
  OAI21_X1 U17449 ( .B1(n15987), .B2(DATAI_15_), .A(n15380), .ZN(n16262) );
  INV_X1 U17450 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n15382) );
  INV_X1 U17451 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n16263) );
  OAI222_X1 U17452 ( .A1(n15383), .A2(n16262), .B1(n15382), .B2(n15381), .C1(
        n16263), .C2(n15535), .ZN(P1_U2967) );
  NAND2_X1 U17453 ( .A1(n15384), .A2(n22099), .ZN(n15394) );
  OAI221_X1 U17454 ( .B1(n22220), .B2(P1_REIP_REG_2__SCAN_IN), .C1(n22220), 
        .C2(P1_REIP_REG_1__SCAN_IN), .A(n22104), .ZN(n15385) );
  AOI22_X1 U17455 ( .A1(n22235), .A2(P1_EBX_REG_3__SCAN_IN), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n15385), .ZN(n15388) );
  INV_X1 U17456 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n15386) );
  NAND4_X1 U17457 ( .A1(n22236), .A2(P1_REIP_REG_2__SCAN_IN), .A3(
        P1_REIP_REG_1__SCAN_IN), .A4(n15386), .ZN(n15387) );
  OAI211_X1 U17458 ( .C1(n15389), .C2(n22267), .A(n15388), .B(n15387), .ZN(
        n15392) );
  INV_X1 U17459 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n15390) );
  NOR2_X1 U17460 ( .A1(n22256), .A2(n15390), .ZN(n15391) );
  AOI211_X1 U17461 ( .C1(n22074), .C2(n16621), .A(n15392), .B(n15391), .ZN(
        n15393) );
  OAI211_X1 U17462 ( .C1(n22251), .C2(n15395), .A(n15394), .B(n15393), .ZN(
        P1_U2837) );
  INV_X1 U17463 ( .A(n22086), .ZN(n20535) );
  OR2_X1 U17464 ( .A1(n15397), .A2(n15396), .ZN(n15398) );
  NAND2_X1 U17465 ( .A1(n20526), .A2(n15398), .ZN(n22077) );
  OAI22_X1 U17466 ( .A1(n22077), .A2(n20510), .B1(n15399), .B2(n20524), .ZN(
        n15400) );
  AOI21_X1 U17467 ( .B1(n20535), .B2(n13916), .A(n15400), .ZN(n15401) );
  INV_X1 U17468 ( .A(n15401), .ZN(P1_U2868) );
  NAND2_X1 U17469 ( .A1(n15053), .A2(n15402), .ZN(n15403) );
  NAND2_X1 U17470 ( .A1(n15404), .A2(n15403), .ZN(n18947) );
  NOR2_X1 U17471 ( .A1(n18947), .A2(n11141), .ZN(n15407) );
  AOI211_X1 U17472 ( .C1(n15405), .C2(n15057), .A(n16740), .B(n15358), .ZN(
        n15406) );
  AOI211_X1 U17473 ( .C1(P2_EBX_REG_11__SCAN_IN), .C2(n11141), .A(n15407), .B(
        n15406), .ZN(n15408) );
  INV_X1 U17474 ( .A(n15408), .ZN(P2_U2876) );
  OR2_X1 U17475 ( .A1(n11267), .A2(n15409), .ZN(n15411) );
  NAND2_X1 U17476 ( .A1(n15411), .A2(n15410), .ZN(n17898) );
  NAND2_X1 U17477 ( .A1(n15412), .A2(n17899), .ZN(n15416) );
  INV_X1 U17478 ( .A(n17898), .ZN(n15640) );
  XNOR2_X1 U17479 ( .A(n19880), .B(n15640), .ZN(n15414) );
  NAND2_X1 U17480 ( .A1(n15413), .A2(n17889), .ZN(n15415) );
  NAND3_X1 U17481 ( .A1(n15416), .A2(n15414), .A3(n15415), .ZN(n15596) );
  INV_X1 U17482 ( .A(n15596), .ZN(n15418) );
  AOI21_X1 U17483 ( .B1(n15416), .B2(n15415), .A(n15414), .ZN(n15417) );
  OAI21_X1 U17484 ( .B1(n15418), .B2(n15417), .A(n20068), .ZN(n15421) );
  INV_X1 U17485 ( .A(n20113), .ZN(n15419) );
  AOI22_X1 U17486 ( .A1(n20011), .A2(n15419), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n20060), .ZN(n15420) );
  OAI211_X1 U17487 ( .C1(n17898), .C2(n16818), .A(n15421), .B(n15420), .ZN(
        P2_U2916) );
  OR2_X1 U17488 ( .A1(n15328), .A2(n15423), .ZN(n15424) );
  AND2_X1 U17489 ( .A1(n15422), .A2(n15424), .ZN(n22100) );
  INV_X1 U17490 ( .A(n22100), .ZN(n15427) );
  INV_X1 U17491 ( .A(n16231), .ZN(n15425) );
  OAI222_X1 U17492 ( .A1(n15427), .A2(n16238), .B1(n16265), .B2(n15426), .C1(
        n15425), .C2(n16268), .ZN(P1_U2899) );
  XNOR2_X1 U17493 ( .A(n17843), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n15429) );
  NOR2_X1 U17494 ( .A1(n15429), .A2(n15428), .ZN(n17842) );
  AOI21_X1 U17495 ( .B1(n15429), .B2(n15428), .A(n17842), .ZN(n15440) );
  NAND2_X1 U17496 ( .A1(n15431), .A2(n15432), .ZN(n15447) );
  NAND3_X1 U17497 ( .A1(n15430), .A2(n15447), .A3(n12415), .ZN(n15436) );
  OAI22_X1 U17498 ( .A1(n15433), .A2(n17029), .B1(n12520), .B2(n18976), .ZN(
        n15434) );
  AOI21_X1 U17499 ( .B1(n17850), .B2(n15634), .A(n15434), .ZN(n15435) );
  OAI211_X1 U17500 ( .C1(n17865), .C2(n15437), .A(n15436), .B(n15435), .ZN(
        n15438) );
  AOI21_X1 U17501 ( .B1(n15440), .B2(n17879), .A(n15438), .ZN(n15439) );
  INV_X1 U17502 ( .A(n15439), .ZN(P2_U3011) );
  INV_X1 U17503 ( .A(n15440), .ZN(n15450) );
  AND2_X1 U17504 ( .A1(n17174), .A2(n16004), .ZN(n15443) );
  OR2_X1 U17505 ( .A1(n15443), .A2(n15442), .ZN(n17294) );
  INV_X1 U17506 ( .A(n17309), .ZN(n15444) );
  MUX2_X1 U17507 ( .A(n17294), .B(n15444), .S(n15820), .Z(n15446) );
  OAI22_X1 U17508 ( .A1(n17898), .A2(n19180), .B1(n12520), .B2(n18976), .ZN(
        n15445) );
  AOI211_X1 U17509 ( .C1(n19202), .C2(n15441), .A(n15446), .B(n15445), .ZN(
        n15449) );
  NAND3_X1 U17510 ( .A1(n15430), .A2(n15447), .A3(n12758), .ZN(n15448) );
  OAI211_X1 U17511 ( .C1(n15450), .C2(n19178), .A(n15449), .B(n15448), .ZN(
        P2_U3043) );
  NOR3_X1 U17512 ( .A1(n17795), .A2(n15570), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n15460) );
  INV_X1 U17513 ( .A(n15460), .ZN(n22432) );
  OR2_X1 U17514 ( .A1(n22415), .A2(n22432), .ZN(n15536) );
  OAI21_X1 U17515 ( .B1(n22428), .B2(n15454), .A(n15536), .ZN(n15456) );
  AOI22_X1 U17516 ( .A1(n15456), .A2(n15786), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15460), .ZN(n15537) );
  OAI22_X1 U17517 ( .A1(n22535), .A2(n15536), .B1(n22550), .B2(n15537), .ZN(
        n15455) );
  AOI21_X1 U17518 ( .B1(n22661), .B2(n22555), .A(n15455), .ZN(n15462) );
  INV_X1 U17519 ( .A(n15456), .ZN(n15457) );
  OAI211_X1 U17520 ( .C1(n15458), .C2(n22286), .A(n15786), .B(n15457), .ZN(
        n15459) );
  NAND2_X1 U17521 ( .A1(n15539), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n15461) );
  OAI211_X1 U17522 ( .C1(n15542), .C2(n22560), .A(n15462), .B(n15461), .ZN(
        P1_U3141) );
  OAI22_X1 U17523 ( .A1(n22445), .A2(n15537), .B1(n22400), .B2(n15536), .ZN(
        n15463) );
  AOI21_X1 U17524 ( .B1(n22661), .B2(n22442), .A(n15463), .ZN(n15465) );
  NAND2_X1 U17525 ( .A1(n15539), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n15464) );
  OAI211_X1 U17526 ( .C1(n15810), .C2(n15542), .A(n15465), .B(n15464), .ZN(
        P1_U3137) );
  OAI22_X1 U17527 ( .A1(n22469), .A2(n15537), .B1(n22459), .B2(n15536), .ZN(
        n15466) );
  AOI21_X1 U17528 ( .B1(n22661), .B2(n22466), .A(n15466), .ZN(n15468) );
  NAND2_X1 U17529 ( .A1(n15539), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n15467) );
  OAI211_X1 U17530 ( .C1(n22452), .C2(n15542), .A(n15468), .B(n15467), .ZN(
        P1_U3138) );
  OAI22_X1 U17531 ( .A1(n22613), .A2(n15537), .B1(n22601), .B2(n15536), .ZN(
        n15469) );
  AOI21_X1 U17532 ( .B1(n22661), .B2(n22610), .A(n15469), .ZN(n15471) );
  NAND2_X1 U17533 ( .A1(n15539), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n15470) );
  OAI211_X1 U17534 ( .C1(n22587), .C2(n15542), .A(n15471), .B(n15470), .ZN(
        P1_U3143) );
  OAI22_X1 U17535 ( .A1(n22516), .A2(n15537), .B1(n22506), .B2(n15536), .ZN(
        n15472) );
  AOI21_X1 U17536 ( .B1(n22661), .B2(n22513), .A(n15472), .ZN(n15474) );
  NAND2_X1 U17537 ( .A1(n15539), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n15473) );
  OAI211_X1 U17538 ( .C1(n22499), .C2(n15542), .A(n15474), .B(n15473), .ZN(
        P1_U3140) );
  OAI22_X1 U17539 ( .A1(n22492), .A2(n15537), .B1(n22482), .B2(n15536), .ZN(
        n15475) );
  AOI21_X1 U17540 ( .B1(n22661), .B2(n22489), .A(n15475), .ZN(n15477) );
  NAND2_X1 U17541 ( .A1(n15539), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n15476) );
  OAI211_X1 U17542 ( .C1(n22476), .C2(n15542), .A(n15477), .B(n15476), .ZN(
        P1_U3139) );
  OAI22_X1 U17543 ( .A1(n22573), .A2(n15536), .B1(n22583), .B2(n15537), .ZN(
        n15478) );
  AOI21_X1 U17544 ( .B1(n22661), .B2(n22580), .A(n15478), .ZN(n15480) );
  NAND2_X1 U17545 ( .A1(n15539), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n15479) );
  OAI211_X1 U17546 ( .C1(n15542), .C2(n22567), .A(n15480), .B(n15479), .ZN(
        P1_U3142) );
  INV_X1 U17547 ( .A(n15481), .ZN(n16254) );
  NAND2_X1 U17548 ( .A1(n15522), .A2(n16254), .ZN(n15508) );
  NAND2_X1 U17549 ( .A1(n15532), .A2(P1_UWORD_REG_0__SCAN_IN), .ZN(n15482) );
  OAI211_X1 U17550 ( .C1(n13524), .C2(n15529), .A(n15508), .B(n15482), .ZN(
        P1_U2937) );
  INV_X1 U17551 ( .A(n15649), .ZN(n16222) );
  NAND2_X1 U17552 ( .A1(n15522), .A2(n16222), .ZN(n15490) );
  NAND2_X1 U17553 ( .A1(n15532), .A2(P1_LWORD_REG_7__SCAN_IN), .ZN(n15483) );
  OAI211_X1 U17554 ( .C1(n13316), .C2(n15535), .A(n15490), .B(n15483), .ZN(
        P1_U2959) );
  INV_X1 U17555 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n15605) );
  NAND2_X1 U17556 ( .A1(n15522), .A2(n16231), .ZN(n15505) );
  NAND2_X1 U17557 ( .A1(n15532), .A2(P1_UWORD_REG_5__SCAN_IN), .ZN(n15484) );
  OAI211_X1 U17558 ( .C1(n15529), .C2(n15605), .A(n15505), .B(n15484), .ZN(
        P1_U2942) );
  INV_X1 U17559 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n15617) );
  NAND2_X1 U17560 ( .A1(n15522), .A2(n16235), .ZN(n15503) );
  NAND2_X1 U17561 ( .A1(n15532), .A2(P1_UWORD_REG_4__SCAN_IN), .ZN(n15485) );
  OAI211_X1 U17562 ( .C1(n15617), .C2(n15529), .A(n15503), .B(n15485), .ZN(
        P1_U2941) );
  MUX2_X1 U17563 ( .A(DATAI_13_), .B(BUF1_REG_13__SCAN_IN), .S(n15987), .Z(
        n16264) );
  NAND2_X1 U17564 ( .A1(n15522), .A2(n16264), .ZN(n15499) );
  NAND2_X1 U17565 ( .A1(n15532), .A2(P1_LWORD_REG_13__SCAN_IN), .ZN(n15486) );
  OAI211_X1 U17566 ( .C1(n16266), .C2(n15529), .A(n15499), .B(n15486), .ZN(
        P1_U2965) );
  MUX2_X1 U17567 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n15987), .Z(
        n16208) );
  NAND2_X1 U17568 ( .A1(n15522), .A2(n16208), .ZN(n15520) );
  NAND2_X1 U17569 ( .A1(n15532), .A2(P1_LWORD_REG_10__SCAN_IN), .ZN(n15487) );
  OAI211_X1 U17570 ( .C1(n15904), .C2(n15535), .A(n15520), .B(n15487), .ZN(
        P1_U2962) );
  INV_X1 U17571 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20435) );
  MUX2_X1 U17572 ( .A(DATAI_14_), .B(BUF1_REG_14__SCAN_IN), .S(n15987), .Z(
        n16194) );
  NAND2_X1 U17573 ( .A1(n15522), .A2(n16194), .ZN(n15534) );
  NAND2_X1 U17574 ( .A1(n15532), .A2(P1_LWORD_REG_14__SCAN_IN), .ZN(n15488) );
  OAI211_X1 U17575 ( .C1(n20435), .C2(n15529), .A(n15534), .B(n15488), .ZN(
        P1_U2966) );
  INV_X1 U17576 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n15603) );
  NAND2_X1 U17577 ( .A1(n15532), .A2(P1_UWORD_REG_7__SCAN_IN), .ZN(n15489) );
  OAI211_X1 U17578 ( .C1(n15529), .C2(n15603), .A(n15490), .B(n15489), .ZN(
        P1_U2944) );
  MUX2_X1 U17579 ( .A(DATAI_12_), .B(BUF1_REG_12__SCAN_IN), .S(n15987), .Z(
        n16201) );
  NAND2_X1 U17580 ( .A1(n15522), .A2(n16201), .ZN(n15516) );
  NAND2_X1 U17581 ( .A1(n15532), .A2(P1_UWORD_REG_12__SCAN_IN), .ZN(n15491) );
  OAI211_X1 U17582 ( .C1(n15535), .C2(n15621), .A(n15516), .B(n15491), .ZN(
        P1_U2949) );
  INV_X1 U17583 ( .A(n15492), .ZN(n16242) );
  NAND2_X1 U17584 ( .A1(n15522), .A2(n16242), .ZN(n15531) );
  NAND2_X1 U17585 ( .A1(n15532), .A2(P1_UWORD_REG_3__SCAN_IN), .ZN(n15493) );
  OAI211_X1 U17586 ( .C1(n13575), .C2(n15529), .A(n15531), .B(n15493), .ZN(
        P1_U2940) );
  INV_X1 U17587 ( .A(n15494), .ZN(n16249) );
  NAND2_X1 U17588 ( .A1(n15522), .A2(n16249), .ZN(n15501) );
  NAND2_X1 U17589 ( .A1(n15532), .A2(P1_LWORD_REG_1__SCAN_IN), .ZN(n15495) );
  OAI211_X1 U17590 ( .C1(n13333), .C2(n15535), .A(n15501), .B(n15495), .ZN(
        P1_U2953) );
  INV_X1 U17591 ( .A(n15496), .ZN(n16246) );
  NAND2_X1 U17592 ( .A1(n15522), .A2(n16246), .ZN(n15525) );
  NAND2_X1 U17593 ( .A1(n15532), .A2(P1_LWORD_REG_2__SCAN_IN), .ZN(n15497) );
  OAI211_X1 U17594 ( .C1(n13327), .C2(n15535), .A(n15525), .B(n15497), .ZN(
        P1_U2954) );
  INV_X1 U17595 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n15607) );
  NAND2_X1 U17596 ( .A1(n15532), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n15498) );
  OAI211_X1 U17597 ( .C1(n15535), .C2(n15607), .A(n15499), .B(n15498), .ZN(
        P1_U2950) );
  NAND2_X1 U17598 ( .A1(n15532), .A2(P1_UWORD_REG_1__SCAN_IN), .ZN(n15500) );
  OAI211_X1 U17599 ( .C1(n13540), .C2(n15529), .A(n15501), .B(n15500), .ZN(
        P1_U2938) );
  NAND2_X1 U17600 ( .A1(n15532), .A2(P1_LWORD_REG_4__SCAN_IN), .ZN(n15502) );
  OAI211_X1 U17601 ( .C1(n20421), .C2(n15535), .A(n15503), .B(n15502), .ZN(
        P1_U2956) );
  NAND2_X1 U17602 ( .A1(n15532), .A2(P1_LWORD_REG_5__SCAN_IN), .ZN(n15504) );
  OAI211_X1 U17603 ( .C1(n15426), .C2(n15535), .A(n15505), .B(n15504), .ZN(
        P1_U2957) );
  INV_X1 U17604 ( .A(n15559), .ZN(n16225) );
  NAND2_X1 U17605 ( .A1(n15522), .A2(n16225), .ZN(n15513) );
  NAND2_X1 U17606 ( .A1(n15532), .A2(P1_LWORD_REG_6__SCAN_IN), .ZN(n15506) );
  OAI211_X1 U17607 ( .C1(n13370), .C2(n15535), .A(n15513), .B(n15506), .ZN(
        P1_U2958) );
  NAND2_X1 U17608 ( .A1(n15532), .A2(P1_LWORD_REG_0__SCAN_IN), .ZN(n15507) );
  OAI211_X1 U17609 ( .C1(n20416), .C2(n15535), .A(n15508), .B(n15507), .ZN(
        P1_U2952) );
  INV_X1 U17610 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n15609) );
  MUX2_X1 U17611 ( .A(DATAI_9_), .B(BUF1_REG_9__SCAN_IN), .S(n15987), .Z(
        n16212) );
  NAND2_X1 U17612 ( .A1(n15522), .A2(n16212), .ZN(n15511) );
  NAND2_X1 U17613 ( .A1(n15532), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n15509) );
  OAI211_X1 U17614 ( .C1(n15529), .C2(n15609), .A(n15511), .B(n15509), .ZN(
        P1_U2946) );
  NAND2_X1 U17615 ( .A1(n15532), .A2(P1_LWORD_REG_9__SCAN_IN), .ZN(n15510) );
  OAI211_X1 U17616 ( .C1(n15902), .C2(n15535), .A(n15511), .B(n15510), .ZN(
        P1_U2961) );
  INV_X1 U17617 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n15611) );
  NAND2_X1 U17618 ( .A1(n15532), .A2(P1_UWORD_REG_6__SCAN_IN), .ZN(n15512) );
  OAI211_X1 U17619 ( .C1(n15529), .C2(n15611), .A(n15513), .B(n15512), .ZN(
        P1_U2943) );
  MUX2_X1 U17620 ( .A(DATAI_11_), .B(BUF1_REG_11__SCAN_IN), .S(n15987), .Z(
        n16204) );
  NAND2_X1 U17621 ( .A1(n15522), .A2(n16204), .ZN(n15518) );
  NAND2_X1 U17622 ( .A1(n15532), .A2(P1_LWORD_REG_11__SCAN_IN), .ZN(n15514) );
  OAI211_X1 U17623 ( .C1(n15924), .C2(n15529), .A(n15518), .B(n15514), .ZN(
        P1_U2963) );
  NAND2_X1 U17624 ( .A1(n15532), .A2(P1_LWORD_REG_12__SCAN_IN), .ZN(n15515) );
  OAI211_X1 U17625 ( .C1(n15932), .C2(n15529), .A(n15516), .B(n15515), .ZN(
        P1_U2964) );
  NAND2_X1 U17626 ( .A1(n15532), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n15517) );
  OAI211_X1 U17627 ( .C1(n13743), .C2(n15535), .A(n15518), .B(n15517), .ZN(
        P1_U2948) );
  INV_X1 U17628 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n15619) );
  NAND2_X1 U17629 ( .A1(n15532), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n15519) );
  OAI211_X1 U17630 ( .C1(n15535), .C2(n15619), .A(n15520), .B(n15519), .ZN(
        P1_U2947) );
  INV_X1 U17631 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20427) );
  INV_X1 U17632 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n20619) );
  NOR2_X1 U17633 ( .A1(n15987), .A2(DATAI_8_), .ZN(n15521) );
  AOI21_X1 U17634 ( .B1(n15987), .B2(n20619), .A(n15521), .ZN(n16216) );
  NAND2_X1 U17635 ( .A1(n15522), .A2(n16216), .ZN(n15528) );
  NAND2_X1 U17636 ( .A1(n15532), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n15523) );
  OAI211_X1 U17637 ( .C1(n20427), .C2(n15535), .A(n15528), .B(n15523), .ZN(
        P1_U2960) );
  NAND2_X1 U17638 ( .A1(n15532), .A2(P1_UWORD_REG_2__SCAN_IN), .ZN(n15524) );
  OAI211_X1 U17639 ( .C1(n15526), .C2(n15529), .A(n15525), .B(n15524), .ZN(
        P1_U2939) );
  INV_X1 U17640 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n15624) );
  NAND2_X1 U17641 ( .A1(n15532), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n15527) );
  OAI211_X1 U17642 ( .C1(n15529), .C2(n15624), .A(n15528), .B(n15527), .ZN(
        P1_U2945) );
  NAND2_X1 U17643 ( .A1(n15532), .A2(P1_LWORD_REG_3__SCAN_IN), .ZN(n15530) );
  OAI211_X1 U17644 ( .C1(n13322), .C2(n15535), .A(n15531), .B(n15530), .ZN(
        P1_U2955) );
  NAND2_X1 U17645 ( .A1(n15532), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n15533) );
  OAI211_X1 U17646 ( .C1(n15535), .C2(n15614), .A(n15534), .B(n15533), .ZN(
        P1_U2951) );
  OAI22_X1 U17647 ( .A1(n22667), .A2(n15537), .B1(n22639), .B2(n15536), .ZN(
        n15538) );
  AOI21_X1 U17648 ( .B1(n22662), .B2(n22661), .A(n15538), .ZN(n15541) );
  NAND2_X1 U17649 ( .A1(n15539), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n15540) );
  OAI211_X1 U17650 ( .C1(n22630), .C2(n15542), .A(n15541), .B(n15540), .ZN(
        P1_U3144) );
  OAI21_X1 U17651 ( .B1(n22556), .B2(n16653), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n15543) );
  OR2_X1 U17652 ( .A1(n22428), .A2(n14969), .ZN(n15550) );
  AOI21_X1 U17653 ( .B1(n15543), .B2(n15550), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n15546) );
  INV_X1 U17654 ( .A(n15544), .ZN(n15545) );
  NOR2_X1 U17655 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15545), .ZN(
        n22553) );
  OR2_X1 U17656 ( .A1(n22372), .A2(n15570), .ZN(n15548) );
  NAND2_X1 U17657 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n15548), .ZN(n22416) );
  NOR2_X1 U17658 ( .A1(n15547), .A2(n15575), .ZN(n22412) );
  INV_X1 U17659 ( .A(n22557), .ZN(n15555) );
  INV_X1 U17660 ( .A(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15554) );
  AND2_X1 U17661 ( .A1(n15547), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n22430) );
  INV_X1 U17662 ( .A(n15548), .ZN(n22411) );
  NAND2_X1 U17663 ( .A1(n22430), .A2(n22411), .ZN(n15549) );
  OAI21_X1 U17664 ( .B1(n15550), .B2(n22424), .A(n15549), .ZN(n22551) );
  AOI22_X1 U17665 ( .A1(n22578), .A2(n22553), .B1(n15587), .B2(n22551), .ZN(
        n15551) );
  OAI21_X1 U17666 ( .B1(n22680), .B2(n22567), .A(n15551), .ZN(n15552) );
  AOI21_X1 U17667 ( .B1(n22556), .B2(n22580), .A(n15552), .ZN(n15553) );
  OAI21_X1 U17668 ( .B1(n15555), .B2(n15554), .A(n15553), .ZN(P1_U3150) );
  NAND2_X1 U17669 ( .A1(n15422), .A2(n15557), .ZN(n15558) );
  AND2_X1 U17670 ( .A1(n15556), .A2(n15558), .ZN(n22112) );
  INV_X1 U17671 ( .A(n22112), .ZN(n15560) );
  OAI222_X1 U17672 ( .A1(n15560), .A2(n16238), .B1(n16268), .B2(n15559), .C1(
        n16265), .C2(n13370), .ZN(P1_U2898) );
  NAND2_X1 U17673 ( .A1(n11247), .A2(n15561), .ZN(n15562) );
  AND2_X1 U17674 ( .A1(n11241), .A2(n15562), .ZN(n16960) );
  INV_X1 U17675 ( .A(n16960), .ZN(n17219) );
  OAI211_X1 U17676 ( .C1(n15563), .C2(n15565), .A(n15564), .B(n16732), .ZN(
        n15567) );
  NAND2_X1 U17677 ( .A1(n11141), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n15566) );
  OAI211_X1 U17678 ( .C1(n17219), .C2(n11141), .A(n15567), .B(n15566), .ZN(
        P2_U2873) );
  NAND2_X1 U17679 ( .A1(n15569), .A2(n13338), .ZN(n22652) );
  NOR3_X1 U17680 ( .A1(n15570), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n15574) );
  INV_X1 U17681 ( .A(n15574), .ZN(n15779) );
  NOR2_X1 U17682 ( .A1(n22415), .A2(n15779), .ZN(n22647) );
  AOI21_X1 U17683 ( .B1(n22410), .B2(n15571), .A(n22647), .ZN(n15576) );
  OAI211_X1 U17684 ( .C1(n15572), .C2(n22286), .A(n15786), .B(n15576), .ZN(
        n15573) );
  OAI211_X1 U17685 ( .C1(n15786), .C2(n15574), .A(n15573), .B(n22387), .ZN(
        n22649) );
  AOI22_X1 U17686 ( .A1(n15780), .A2(n22466), .B1(n22649), .B2(
        P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n15578) );
  OAI22_X1 U17687 ( .A1(n15576), .A2(n22424), .B1(n15779), .B2(n15575), .ZN(
        n22648) );
  AOI22_X1 U17688 ( .A1(n16633), .A2(n22648), .B1(n22464), .B2(n22647), .ZN(
        n15577) );
  OAI211_X1 U17689 ( .C1(n22452), .C2(n22604), .A(n15578), .B(n15577), .ZN(
        P1_U3106) );
  AOI22_X1 U17690 ( .A1(n15780), .A2(n22442), .B1(n22649), .B2(
        P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15580) );
  AOI22_X1 U17691 ( .A1(n16628), .A2(n22648), .B1(n22433), .B2(n22647), .ZN(
        n15579) );
  OAI211_X1 U17692 ( .C1(n15810), .C2(n22604), .A(n15580), .B(n15579), .ZN(
        P1_U3105) );
  AOI22_X1 U17693 ( .A1(n15780), .A2(n22513), .B1(n22649), .B2(
        P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15582) );
  AOI22_X1 U17694 ( .A1(n16643), .A2(n22648), .B1(n22511), .B2(n22647), .ZN(
        n15581) );
  OAI211_X1 U17695 ( .C1(n22499), .C2(n22604), .A(n15582), .B(n15581), .ZN(
        P1_U3108) );
  AOI22_X1 U17696 ( .A1(n15780), .A2(n22610), .B1(n22649), .B2(
        P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n15584) );
  AOI22_X1 U17697 ( .A1(n16648), .A2(n22648), .B1(n22608), .B2(n22647), .ZN(
        n15583) );
  OAI211_X1 U17698 ( .C1(n22587), .C2(n22604), .A(n15584), .B(n15583), .ZN(
        P1_U3111) );
  AOI22_X1 U17699 ( .A1(n15780), .A2(n22555), .B1(n22649), .B2(
        P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n15586) );
  AOI22_X1 U17700 ( .A1(n22554), .A2(n22647), .B1(n22648), .B2(n22552), .ZN(
        n15585) );
  OAI211_X1 U17701 ( .C1(n22560), .C2(n22604), .A(n15586), .B(n15585), .ZN(
        P1_U3109) );
  AOI22_X1 U17702 ( .A1(n15780), .A2(n22580), .B1(n22649), .B2(
        P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15589) );
  AOI22_X1 U17703 ( .A1(n22578), .A2(n22647), .B1(n22648), .B2(n15587), .ZN(
        n15588) );
  OAI211_X1 U17704 ( .C1(n22567), .C2(n22604), .A(n15589), .B(n15588), .ZN(
        P1_U3110) );
  AOI22_X1 U17705 ( .A1(n15780), .A2(n22489), .B1(n22649), .B2(
        P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15591) );
  AOI22_X1 U17706 ( .A1(n16638), .A2(n22648), .B1(n22487), .B2(n22647), .ZN(
        n15590) );
  OAI211_X1 U17707 ( .C1(n22476), .C2(n22604), .A(n15591), .B(n15590), .ZN(
        P1_U3107) );
  NAND2_X1 U17708 ( .A1(n19880), .A2(n17898), .ZN(n15595) );
  NAND2_X1 U17709 ( .A1(n15592), .A2(n15410), .ZN(n15594) );
  INV_X1 U17710 ( .A(n15817), .ZN(n15593) );
  AOI21_X1 U17711 ( .B1(n15596), .B2(n15595), .A(n19207), .ZN(n20014) );
  XOR2_X1 U17712 ( .A(n20013), .B(n20014), .Z(n15597) );
  NAND2_X1 U17713 ( .A1(n15597), .A2(n20068), .ZN(n15599) );
  AOI22_X1 U17714 ( .A1(n20067), .A2(n19207), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n20060), .ZN(n15598) );
  OAI211_X1 U17715 ( .C1(n20073), .C2(n15600), .A(n15599), .B(n15598), .ZN(
        P2_U2915) );
  AOI22_X1 U17716 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20425), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n20429), .ZN(n15601) );
  OAI21_X1 U17717 ( .B1(n13524), .B2(n15623), .A(n15601), .ZN(P1_U2920) );
  AOI22_X1 U17718 ( .A1(n20425), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n20429), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n15602) );
  OAI21_X1 U17719 ( .B1(n15603), .B2(n15623), .A(n15602), .ZN(P1_U2913) );
  AOI22_X1 U17720 ( .A1(n21877), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n20429), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n15604) );
  OAI21_X1 U17721 ( .B1(n15605), .B2(n15623), .A(n15604), .ZN(P1_U2915) );
  AOI22_X1 U17722 ( .A1(n21877), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n20429), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n15606) );
  OAI21_X1 U17723 ( .B1(n15607), .B2(n15623), .A(n15606), .ZN(P1_U2907) );
  AOI22_X1 U17724 ( .A1(n21877), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n20429), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n15608) );
  OAI21_X1 U17725 ( .B1(n15609), .B2(n15623), .A(n15608), .ZN(P1_U2911) );
  AOI22_X1 U17726 ( .A1(n21877), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n20429), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n15610) );
  OAI21_X1 U17727 ( .B1(n15611), .B2(n15623), .A(n15610), .ZN(P1_U2914) );
  AOI22_X1 U17728 ( .A1(n21877), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n20429), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n15612) );
  OAI21_X1 U17729 ( .B1(n13743), .B2(n15623), .A(n15612), .ZN(P1_U2909) );
  AOI22_X1 U17730 ( .A1(n21877), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(n20429), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n15613) );
  OAI21_X1 U17731 ( .B1(n15614), .B2(n15623), .A(n15613), .ZN(P1_U2906) );
  AOI22_X1 U17732 ( .A1(n21877), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n20429), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n15615) );
  OAI21_X1 U17733 ( .B1(n13575), .B2(n15623), .A(n15615), .ZN(P1_U2917) );
  AOI22_X1 U17734 ( .A1(n21877), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n20429), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n15616) );
  OAI21_X1 U17735 ( .B1(n15617), .B2(n15623), .A(n15616), .ZN(P1_U2916) );
  AOI22_X1 U17736 ( .A1(n21877), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n20429), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n15618) );
  OAI21_X1 U17737 ( .B1(n15619), .B2(n15623), .A(n15618), .ZN(P1_U2910) );
  AOI22_X1 U17738 ( .A1(n21877), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n20429), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n15620) );
  OAI21_X1 U17739 ( .B1(n15621), .B2(n15623), .A(n15620), .ZN(P1_U2908) );
  AOI22_X1 U17740 ( .A1(n21877), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n20429), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n15622) );
  OAI21_X1 U17741 ( .B1(n15624), .B2(n15623), .A(n15622), .ZN(P1_U2912) );
  OR2_X1 U17742 ( .A1(n15626), .A2(n15625), .ZN(n15627) );
  AND2_X1 U17743 ( .A1(n15627), .A2(n11247), .ZN(n18968) );
  INV_X1 U17744 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n18967) );
  NOR2_X1 U17745 ( .A1(n16727), .A2(n18967), .ZN(n15630) );
  AOI211_X1 U17746 ( .C1(n15628), .C2(n15359), .A(n16740), .B(n15563), .ZN(
        n15629) );
  AOI211_X1 U17747 ( .C1(n18968), .C2(n16727), .A(n15630), .B(n15629), .ZN(
        n15631) );
  INV_X1 U17748 ( .A(n15631), .ZN(P2_U2874) );
  NAND2_X1 U17749 ( .A1(n19029), .A2(n15632), .ZN(n15633) );
  XNOR2_X1 U17750 ( .A(n15634), .B(n15633), .ZN(n15644) );
  INV_X1 U17751 ( .A(n18880), .ZN(n18886) );
  AOI22_X1 U17752 ( .A1(n19134), .A2(P2_REIP_REG_3__SCAN_IN), .B1(n19135), 
        .B2(P2_EBX_REG_3__SCAN_IN), .ZN(n15637) );
  NAND2_X1 U17753 ( .A1(n19157), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n15636) );
  OAI211_X1 U17754 ( .C1(n15638), .C2(n19149), .A(n15637), .B(n15636), .ZN(
        n15639) );
  AOI21_X1 U17755 ( .B1(n15640), .B2(n19159), .A(n15639), .ZN(n15642) );
  NAND2_X1 U17756 ( .A1(n15441), .A2(n19160), .ZN(n15641) );
  OAI211_X1 U17757 ( .C1(n19880), .C2(n18886), .A(n15642), .B(n15641), .ZN(
        n15643) );
  AOI21_X1 U17758 ( .B1(n15644), .B2(n19127), .A(n15643), .ZN(n15645) );
  INV_X1 U17759 ( .A(n15645), .ZN(P2_U2852) );
  INV_X1 U17760 ( .A(n15646), .ZN(n15647) );
  AOI21_X1 U17761 ( .B1(n15648), .B2(n15556), .A(n15647), .ZN(n20554) );
  INV_X1 U17762 ( .A(n20554), .ZN(n22122) );
  OAI222_X1 U17763 ( .A1(n22122), .A2(n16238), .B1(n16268), .B2(n15649), .C1(
        n16265), .C2(n13316), .ZN(P1_U2897) );
  AND2_X1 U17764 ( .A1(n15652), .A2(n15651), .ZN(n15653) );
  NOR2_X1 U17765 ( .A1(n15650), .A2(n15653), .ZN(n21960) );
  INV_X1 U17766 ( .A(n21960), .ZN(n22119) );
  INV_X1 U17767 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n15654) );
  OAI222_X1 U17768 ( .A1(n22119), .A2(n20510), .B1(n15654), .B2(n20524), .C1(
        n22122), .C2(n16189), .ZN(P1_U2865) );
  INV_X1 U17769 ( .A(n22631), .ZN(n22594) );
  OAI21_X1 U17770 ( .B1(n15688), .B2(n22594), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n15656) );
  NAND2_X1 U17771 ( .A1(n22396), .A2(n14969), .ZN(n15659) );
  AOI21_X1 U17772 ( .B1(n15656), .B2(n15659), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n15658) );
  NOR2_X1 U17773 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15657), .ZN(
        n15662) );
  NAND2_X1 U17774 ( .A1(n15684), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n15665) );
  INV_X1 U17775 ( .A(n15659), .ZN(n15661) );
  INV_X1 U17776 ( .A(n15785), .ZN(n15660) );
  NAND2_X1 U17777 ( .A1(n15660), .A2(n22372), .ZN(n22362) );
  INV_X1 U17778 ( .A(n22362), .ZN(n22358) );
  AOI22_X1 U17779 ( .A1(n15661), .A2(n15786), .B1(n22430), .B2(n22358), .ZN(
        n15686) );
  INV_X1 U17780 ( .A(n15662), .ZN(n15685) );
  OAI22_X1 U17781 ( .A1(n22613), .A2(n15686), .B1(n15685), .B2(n22601), .ZN(
        n15663) );
  AOI21_X1 U17782 ( .B1(n15688), .B2(n22609), .A(n15663), .ZN(n15664) );
  OAI211_X1 U17783 ( .C1(n22603), .C2(n22631), .A(n15665), .B(n15664), .ZN(
        P1_U3071) );
  NAND2_X1 U17784 ( .A1(n15684), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n15668) );
  OAI22_X1 U17785 ( .A1(n22516), .A2(n15686), .B1(n15685), .B2(n22506), .ZN(
        n15666) );
  AOI21_X1 U17786 ( .B1(n15688), .B2(n22512), .A(n15666), .ZN(n15667) );
  OAI211_X1 U17787 ( .C1(n22507), .C2(n22631), .A(n15668), .B(n15667), .ZN(
        P1_U3068) );
  NAND2_X1 U17788 ( .A1(n15684), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n15671) );
  OAI22_X1 U17789 ( .A1(n22469), .A2(n15686), .B1(n15685), .B2(n22459), .ZN(
        n15669) );
  AOI21_X1 U17790 ( .B1(n15688), .B2(n22465), .A(n15669), .ZN(n15670) );
  OAI211_X1 U17791 ( .C1(n22460), .C2(n22631), .A(n15671), .B(n15670), .ZN(
        P1_U3066) );
  NAND2_X1 U17792 ( .A1(n15684), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n15674) );
  OAI22_X1 U17793 ( .A1(n22492), .A2(n15686), .B1(n15685), .B2(n22482), .ZN(
        n15672) );
  AOI21_X1 U17794 ( .B1(n15688), .B2(n22488), .A(n15672), .ZN(n15673) );
  OAI211_X1 U17795 ( .C1(n22483), .C2(n22631), .A(n15674), .B(n15673), .ZN(
        P1_U3067) );
  NAND2_X1 U17796 ( .A1(n15684), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n15677) );
  OAI22_X1 U17797 ( .A1(n22535), .A2(n15685), .B1(n15686), .B2(n22550), .ZN(
        n15675) );
  AOI21_X1 U17798 ( .B1(n15688), .B2(n22547), .A(n15675), .ZN(n15676) );
  OAI211_X1 U17799 ( .C1(n22536), .C2(n22631), .A(n15677), .B(n15676), .ZN(
        P1_U3069) );
  NAND2_X1 U17800 ( .A1(n15684), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n15680) );
  OAI22_X1 U17801 ( .A1(n22667), .A2(n15686), .B1(n15685), .B2(n22639), .ZN(
        n15678) );
  AOI21_X1 U17802 ( .B1(n15688), .B2(n22675), .A(n15678), .ZN(n15679) );
  OAI211_X1 U17803 ( .C1(n22631), .C2(n22681), .A(n15680), .B(n15679), .ZN(
        P1_U3072) );
  NAND2_X1 U17804 ( .A1(n15684), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n15683) );
  OAI22_X1 U17805 ( .A1(n22573), .A2(n15685), .B1(n15686), .B2(n22583), .ZN(
        n15681) );
  AOI21_X1 U17806 ( .B1(n15688), .B2(n22579), .A(n15681), .ZN(n15682) );
  OAI211_X1 U17807 ( .C1(n22574), .C2(n22631), .A(n15683), .B(n15682), .ZN(
        P1_U3070) );
  NAND2_X1 U17808 ( .A1(n15684), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n15690) );
  OAI22_X1 U17809 ( .A1(n22445), .A2(n15686), .B1(n22400), .B2(n15685), .ZN(
        n15687) );
  AOI21_X1 U17810 ( .B1(n15688), .B2(n22434), .A(n15687), .ZN(n15689) );
  OAI211_X1 U17811 ( .C1(n22401), .C2(n22631), .A(n15690), .B(n15689), .ZN(
        P1_U3065) );
  OAI21_X1 U17812 ( .B1(n15691), .B2(n15693), .A(n15692), .ZN(n15718) );
  AND2_X1 U17813 ( .A1(n15694), .A2(n11772), .ZN(n15701) );
  OAI21_X1 U17814 ( .B1(n15695), .B2(n15108), .A(n15839), .ZN(n18998) );
  OAI22_X1 U17815 ( .A1(n16818), .A2(n18998), .B1(n16817), .B2(n15696), .ZN(
        n15699) );
  AND2_X1 U17816 ( .A1(n16817), .A2(n15697), .ZN(n20062) );
  NOR2_X1 U17817 ( .A1(n16819), .A2(n20245), .ZN(n15698) );
  AOI211_X1 U17818 ( .C1(BUF1_REG_16__SCAN_IN), .C2(n20064), .A(n15699), .B(
        n15698), .ZN(n15703) );
  NAND2_X1 U17819 ( .A1(n20063), .A2(BUF2_REG_16__SCAN_IN), .ZN(n15702) );
  OAI211_X1 U17820 ( .C1(n15718), .C2(n20012), .A(n15703), .B(n15702), .ZN(
        P2_U2903) );
  AOI21_X1 U17821 ( .B1(n15704), .B2(n15646), .A(n11194), .ZN(n22133) );
  INV_X1 U17822 ( .A(n22133), .ZN(n15859) );
  INV_X1 U17823 ( .A(n16268), .ZN(n15946) );
  AOI22_X1 U17824 ( .A1(n15946), .A2(n16216), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n16252), .ZN(n15705) );
  OAI21_X1 U17825 ( .B1(n15859), .B2(n16238), .A(n15705), .ZN(P1_U2896) );
  AND2_X1 U17826 ( .A1(n11241), .A2(n15707), .ZN(n15708) );
  NOR2_X1 U17827 ( .A1(n15706), .A2(n15708), .ZN(n18982) );
  NOR2_X1 U17828 ( .A1(n16727), .A2(n12144), .ZN(n15711) );
  AOI211_X1 U17829 ( .C1(n15709), .C2(n15564), .A(n16740), .B(n15691), .ZN(
        n15710) );
  AOI211_X1 U17830 ( .C1(n18982), .C2(n16727), .A(n15711), .B(n15710), .ZN(
        n15712) );
  INV_X1 U17831 ( .A(n15712), .ZN(P2_U2872) );
  NOR2_X1 U17832 ( .A1(n15706), .A2(n15714), .ZN(n15715) );
  OR2_X1 U17833 ( .A1(n15713), .A2(n15715), .ZN(n16928) );
  NOR2_X1 U17834 ( .A1(n16928), .A2(n11141), .ZN(n15716) );
  AOI21_X1 U17835 ( .B1(P2_EBX_REG_16__SCAN_IN), .B2(n11141), .A(n15716), .ZN(
        n15717) );
  OAI21_X1 U17836 ( .B1(n15718), .B2(n16740), .A(n15717), .ZN(P2_U2871) );
  NOR2_X1 U17837 ( .A1(n19015), .A2(n15719), .ZN(n15720) );
  XNOR2_X1 U17838 ( .A(n15720), .B(n16958), .ZN(n15731) );
  INV_X1 U17839 ( .A(n19135), .ZN(n19153) );
  NAND2_X1 U17840 ( .A1(n16960), .A2(n19160), .ZN(n15725) );
  AOI22_X1 U17841 ( .A1(n19157), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n19136), .B2(n15721), .ZN(n15722) );
  OAI21_X1 U17842 ( .B1(n17966), .B2(n19151), .A(n15722), .ZN(n15723) );
  NOR2_X1 U17843 ( .A1(n17016), .A2(n15723), .ZN(n15724) );
  OAI211_X1 U17844 ( .C1(n19153), .C2(n15726), .A(n15725), .B(n15724), .ZN(
        n15730) );
  NOR2_X1 U17845 ( .A1(n15038), .A2(n15727), .ZN(n15728) );
  OR2_X1 U17846 ( .A1(n15107), .A2(n15728), .ZN(n19744) );
  NOR2_X1 U17847 ( .A1(n19744), .A2(n19133), .ZN(n15729) );
  AOI211_X1 U17848 ( .C1(n15731), .C2(n19127), .A(n15730), .B(n15729), .ZN(
        n15732) );
  INV_X1 U17849 ( .A(n15732), .ZN(P2_U2841) );
  NOR2_X1 U17850 ( .A1(n19015), .A2(n15733), .ZN(n15734) );
  XNOR2_X1 U17851 ( .A(n15734), .B(n17882), .ZN(n15742) );
  AOI22_X1 U17852 ( .A1(n15735), .A2(n19136), .B1(n19157), .B2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n15736) );
  OAI21_X1 U17853 ( .B1(n12542), .B2(n19151), .A(n15736), .ZN(n15741) );
  NAND2_X1 U17854 ( .A1(n19192), .A2(n19160), .ZN(n15738) );
  AOI21_X1 U17855 ( .B1(n19159), .B2(n19190), .A(n17016), .ZN(n15737) );
  OAI211_X1 U17856 ( .C1(n19153), .C2(n15739), .A(n15738), .B(n15737), .ZN(
        n15740) );
  AOI211_X1 U17857 ( .C1(n15742), .C2(n19127), .A(n15741), .B(n15740), .ZN(
        n15743) );
  INV_X1 U17858 ( .A(n15743), .ZN(P2_U2847) );
  NOR2_X1 U17859 ( .A1(n19015), .A2(n17338), .ZN(n15744) );
  XNOR2_X1 U17860 ( .A(n15744), .B(n17836), .ZN(n15745) );
  NAND2_X1 U17861 ( .A1(n15745), .A2(n19127), .ZN(n15754) );
  OAI22_X1 U17862 ( .A1(n15746), .A2(n19153), .B1(n17956), .B2(n19151), .ZN(
        n15749) );
  NOR2_X1 U17863 ( .A1(n19149), .A2(n15747), .ZN(n15748) );
  AOI211_X1 U17864 ( .C1(n19157), .C2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n15749), .B(n15748), .ZN(n15750) );
  OAI21_X1 U17865 ( .B1(n15751), .B2(n19133), .A(n15750), .ZN(n15752) );
  AOI21_X1 U17866 ( .B1(n17838), .B2(n19160), .A(n15752), .ZN(n15753) );
  OAI211_X1 U17867 ( .C1(n18886), .C2(n19879), .A(n15754), .B(n15753), .ZN(
        P2_U2853) );
  INV_X1 U17868 ( .A(n17364), .ZN(n17335) );
  INV_X1 U17869 ( .A(n12690), .ZN(n15756) );
  AND2_X1 U17870 ( .A1(n15756), .A2(n15755), .ZN(n17329) );
  INV_X1 U17871 ( .A(n12709), .ZN(n17357) );
  MUX2_X1 U17872 ( .A(n17329), .B(n17357), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n15757) );
  OAI21_X1 U17873 ( .B1(n18858), .B2(n17335), .A(n15757), .ZN(n19219) );
  AOI22_X1 U17874 ( .A1(n19015), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n18857), .B2(n19029), .ZN(n17337) );
  AOI222_X1 U17875 ( .A1(n19219), .A2(n19170), .B1(n19915), .B2(n19279), .C1(
        P2_STATE2_REG_1__SCAN_IN), .C2(n17337), .ZN(n15766) );
  NOR2_X1 U17876 ( .A1(n19270), .A2(n17768), .ZN(n19269) );
  INV_X1 U17877 ( .A(n15758), .ZN(n15759) );
  NAND2_X1 U17878 ( .A1(n15759), .A2(n19247), .ZN(n15763) );
  AND4_X1 U17879 ( .A1(n15763), .A2(n15762), .A3(n15761), .A4(n15760), .ZN(
        n19255) );
  OAI22_X1 U17880 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19916), .B1(n19255), 
        .B2(n19287), .ZN(n15764) );
  NAND2_X1 U17881 ( .A1(n19166), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15765) );
  OAI21_X1 U17882 ( .B1(n15766), .B2(n19166), .A(n15765), .ZN(P2_U3601) );
  AOI21_X1 U17883 ( .B1(n15768), .B2(n15767), .A(n14994), .ZN(n17273) );
  INV_X1 U17884 ( .A(n17273), .ZN(n19750) );
  NOR2_X1 U17885 ( .A1(n19015), .A2(n15769), .ZN(n15770) );
  XNOR2_X1 U17886 ( .A(n15770), .B(n17005), .ZN(n15771) );
  NAND2_X1 U17887 ( .A1(n15771), .A2(n19127), .ZN(n15778) );
  OAI21_X1 U17888 ( .B1(n19153), .B2(n15772), .A(n18976), .ZN(n15776) );
  AOI22_X1 U17889 ( .A1(n15773), .A2(n19136), .B1(n19157), .B2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n15774) );
  OAI21_X1 U17890 ( .B1(n12571), .B2(n19151), .A(n15774), .ZN(n15775) );
  AOI211_X1 U17891 ( .C1(n19160), .C2(n17267), .A(n15776), .B(n15775), .ZN(
        n15777) );
  OAI211_X1 U17892 ( .C1(n19133), .C2(n19750), .A(n15778), .B(n15777), .ZN(
        P2_U2845) );
  NOR2_X1 U17893 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15779), .ZN(
        n22529) );
  OAI21_X1 U17894 ( .B1(n15780), .B2(n22531), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n15781) );
  AOI21_X1 U17895 ( .B1(n22410), .B2(n14969), .A(n22529), .ZN(n15784) );
  NAND2_X1 U17896 ( .A1(n15781), .A2(n15784), .ZN(n15783) );
  NAND2_X1 U17897 ( .A1(n22532), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n15790) );
  INV_X1 U17898 ( .A(n15784), .ZN(n15787) );
  NAND2_X1 U17899 ( .A1(n15785), .A2(n22372), .ZN(n22437) );
  INV_X1 U17900 ( .A(n22437), .ZN(n22429) );
  AOI22_X1 U17901 ( .A1(n15787), .A2(n15786), .B1(n22412), .B2(n22429), .ZN(
        n22528) );
  INV_X1 U17902 ( .A(n22529), .ZN(n15806) );
  OAI22_X1 U17903 ( .A1(n22516), .A2(n22528), .B1(n22506), .B2(n15806), .ZN(
        n15788) );
  AOI21_X1 U17904 ( .B1(n22531), .B2(n22513), .A(n15788), .ZN(n15789) );
  OAI211_X1 U17905 ( .C1(n22499), .C2(n22652), .A(n15790), .B(n15789), .ZN(
        P1_U3100) );
  NAND2_X1 U17906 ( .A1(n22532), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n15793) );
  OAI22_X1 U17907 ( .A1(n22528), .A2(n22583), .B1(n22573), .B2(n15806), .ZN(
        n15791) );
  AOI21_X1 U17908 ( .B1(n22531), .B2(n22580), .A(n15791), .ZN(n15792) );
  OAI211_X1 U17909 ( .C1(n22567), .C2(n22652), .A(n15793), .B(n15792), .ZN(
        P1_U3102) );
  NAND2_X1 U17910 ( .A1(n22532), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n15796) );
  OAI22_X1 U17911 ( .A1(n22613), .A2(n22528), .B1(n22601), .B2(n15806), .ZN(
        n15794) );
  AOI21_X1 U17912 ( .B1(n22531), .B2(n22610), .A(n15794), .ZN(n15795) );
  OAI211_X1 U17913 ( .C1(n22587), .C2(n22652), .A(n15796), .B(n15795), .ZN(
        P1_U3103) );
  NAND2_X1 U17914 ( .A1(n22532), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n15799) );
  OAI22_X1 U17915 ( .A1(n22667), .A2(n22528), .B1(n22639), .B2(n15806), .ZN(
        n15797) );
  AOI21_X1 U17916 ( .B1(n22662), .B2(n22531), .A(n15797), .ZN(n15798) );
  OAI211_X1 U17917 ( .C1(n22630), .C2(n22652), .A(n15799), .B(n15798), .ZN(
        P1_U3104) );
  NAND2_X1 U17918 ( .A1(n22532), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n15802) );
  OAI22_X1 U17919 ( .A1(n22469), .A2(n22528), .B1(n22459), .B2(n15806), .ZN(
        n15800) );
  AOI21_X1 U17920 ( .B1(n22531), .B2(n22466), .A(n15800), .ZN(n15801) );
  OAI211_X1 U17921 ( .C1(n22452), .C2(n22652), .A(n15802), .B(n15801), .ZN(
        P1_U3098) );
  NAND2_X1 U17922 ( .A1(n22532), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n15805) );
  OAI22_X1 U17923 ( .A1(n22492), .A2(n22528), .B1(n22482), .B2(n15806), .ZN(
        n15803) );
  AOI21_X1 U17924 ( .B1(n22531), .B2(n22489), .A(n15803), .ZN(n15804) );
  OAI211_X1 U17925 ( .C1(n22476), .C2(n22652), .A(n15805), .B(n15804), .ZN(
        P1_U3099) );
  NAND2_X1 U17926 ( .A1(n22532), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n15809) );
  OAI22_X1 U17927 ( .A1(n22445), .A2(n22528), .B1(n22400), .B2(n15806), .ZN(
        n15807) );
  AOI21_X1 U17928 ( .B1(n22531), .B2(n22442), .A(n15807), .ZN(n15808) );
  OAI211_X1 U17929 ( .C1(n15810), .C2(n22652), .A(n15809), .B(n15808), .ZN(
        P1_U3097) );
  INV_X1 U17930 ( .A(n15811), .ZN(n17023) );
  OAI21_X1 U17931 ( .B1(n15813), .B2(n15812), .A(n17023), .ZN(n17852) );
  INV_X1 U17932 ( .A(n15814), .ZN(n15815) );
  AOI21_X1 U17933 ( .B1(n12384), .B2(n15816), .A(n15815), .ZN(n17851) );
  NAND2_X1 U17934 ( .A1(n17851), .A2(n12758), .ZN(n15824) );
  XNOR2_X1 U17935 ( .A(n15818), .B(n15817), .ZN(n20017) );
  NOR2_X1 U17936 ( .A1(n17309), .A2(n15820), .ZN(n19205) );
  OAI221_X1 U17937 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C1(n19204), .C2(n12384), .A(
        n19205), .ZN(n15819) );
  NAND2_X1 U17938 ( .A1(n17016), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n17853) );
  OAI211_X1 U17939 ( .C1(n19180), .C2(n20017), .A(n15819), .B(n17853), .ZN(
        n15822) );
  AOI21_X1 U17940 ( .B1(n15820), .B2(n19183), .A(n17294), .ZN(n19206) );
  NOR2_X1 U17941 ( .A1(n19206), .A2(n12384), .ZN(n15821) );
  AOI211_X1 U17942 ( .C1(n18903), .C2(n19202), .A(n15822), .B(n15821), .ZN(
        n15823) );
  OAI211_X1 U17943 ( .C1(n19178), .C2(n17852), .A(n15824), .B(n15823), .ZN(
        P2_U3041) );
  OAI21_X1 U17944 ( .B1(n15827), .B2(n15826), .A(n11149), .ZN(n21964) );
  AOI22_X1 U17945 ( .A1(n20588), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n22052), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n15828) );
  OAI21_X1 U17946 ( .B1(n20594), .B2(n22131), .A(n15828), .ZN(n15829) );
  AOI21_X1 U17947 ( .B1(n22133), .B2(n20555), .A(n15829), .ZN(n15830) );
  OAI21_X1 U17948 ( .B1(n21964), .B2(n22268), .A(n15830), .ZN(P1_U2991) );
  OAI21_X1 U17949 ( .B1(n15713), .B2(n15832), .A(n15831), .ZN(n19005) );
  AOI21_X1 U17950 ( .B1(n15834), .B2(n15692), .A(n15833), .ZN(n15837) );
  NAND2_X1 U17951 ( .A1(n15837), .A2(n16732), .ZN(n15836) );
  NAND2_X1 U17952 ( .A1(n11141), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n15835) );
  OAI211_X1 U17953 ( .C1(n19005), .C2(n11141), .A(n15836), .B(n15835), .ZN(
        P2_U2870) );
  INV_X1 U17954 ( .A(n20063), .ZN(n16824) );
  INV_X1 U17955 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n15845) );
  NAND2_X1 U17956 ( .A1(n15837), .A2(n20068), .ZN(n15844) );
  INV_X1 U17957 ( .A(n15838), .ZN(n15840) );
  XNOR2_X1 U17958 ( .A(n15840), .B(n15839), .ZN(n19006) );
  AOI22_X1 U17959 ( .A1(n20067), .A2(n19006), .B1(P2_EAX_REG_17__SCAN_IN), 
        .B2(n20060), .ZN(n15841) );
  OAI21_X1 U17960 ( .B1(n20195), .B2(n16819), .A(n15841), .ZN(n15842) );
  AOI21_X1 U17961 ( .B1(n20064), .B2(BUF1_REG_17__SCAN_IN), .A(n15842), .ZN(
        n15843) );
  OAI211_X1 U17962 ( .C1(n16824), .C2(n15845), .A(n15844), .B(n15843), .ZN(
        P2_U2902) );
  AOI21_X1 U17963 ( .B1(n15847), .B2(n14993), .A(n15037), .ZN(n17249) );
  INV_X1 U17964 ( .A(n17249), .ZN(n19747) );
  INV_X1 U17965 ( .A(n17246), .ZN(n16984) );
  NAND2_X1 U17966 ( .A1(n19157), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15849) );
  AOI21_X1 U17967 ( .B1(n19135), .B2(P2_EBX_REG_12__SCAN_IN), .A(n17016), .ZN(
        n15848) );
  OAI211_X1 U17968 ( .C1(n19151), .C2(n17965), .A(n15849), .B(n15848), .ZN(
        n15852) );
  NOR2_X1 U17969 ( .A1(n15850), .A2(n19149), .ZN(n15851) );
  AOI211_X1 U17970 ( .C1(n19160), .C2(n16984), .A(n15852), .B(n15851), .ZN(
        n15856) );
  NOR2_X1 U17971 ( .A1(n19015), .A2(n15853), .ZN(n18957) );
  XNOR2_X1 U17972 ( .A(n18957), .B(n16982), .ZN(n15854) );
  NAND2_X1 U17973 ( .A1(n15854), .A2(n19127), .ZN(n15855) );
  OAI211_X1 U17974 ( .C1(n19747), .C2(n19133), .A(n15856), .B(n15855), .ZN(
        P2_U2843) );
  OR2_X1 U17975 ( .A1(n15650), .A2(n15857), .ZN(n15858) );
  NAND2_X1 U17976 ( .A1(n15866), .A2(n15858), .ZN(n22129) );
  INV_X1 U17977 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n22128) );
  OAI222_X1 U17978 ( .A1(n22129), .A2(n20510), .B1(n22128), .B2(n20524), .C1(
        n16189), .C2(n15859), .ZN(P1_U2864) );
  OAI21_X1 U17979 ( .B1(n11194), .B2(n15861), .A(n11617), .ZN(n15917) );
  INV_X1 U17980 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n17481) );
  INV_X1 U17981 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21922) );
  NAND3_X1 U17982 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n22081) );
  NOR2_X1 U17983 ( .A1(n21922), .A2(n22081), .ZN(n22096) );
  NAND2_X1 U17984 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n22096), .ZN(n22106) );
  NOR2_X1 U17985 ( .A1(n17481), .A2(n22106), .ZN(n22116) );
  NAND2_X1 U17986 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n22116), .ZN(n15862) );
  NOR2_X1 U17987 ( .A1(n15862), .A2(n22220), .ZN(n22127) );
  NAND2_X1 U17988 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n22127), .ZN(n15886) );
  INV_X1 U17989 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n15916) );
  INV_X1 U17990 ( .A(n15862), .ZN(n15863) );
  NAND2_X1 U17991 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n15863), .ZN(n15887) );
  INV_X1 U17992 ( .A(n22104), .ZN(n16098) );
  AOI21_X1 U17993 ( .B1(n22236), .B2(n15887), .A(n16098), .ZN(n22136) );
  INV_X1 U17994 ( .A(n15889), .ZN(n15864) );
  AOI21_X1 U17995 ( .B1(n15866), .B2(n15865), .A(n15864), .ZN(n21977) );
  AOI22_X1 U17996 ( .A1(n21977), .A2(n22199), .B1(n22235), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n15868) );
  NAND2_X1 U17997 ( .A1(n22104), .A2(n15867), .ZN(n22092) );
  OAI211_X1 U17998 ( .C1(n22256), .C2(n15869), .A(n15868), .B(n22092), .ZN(
        n15870) );
  INV_X1 U17999 ( .A(n15870), .ZN(n15871) );
  OAI221_X1 U18000 ( .B1(P1_REIP_REG_9__SCAN_IN), .B2(n15886), .C1(n15916), 
        .C2(n22136), .A(n15871), .ZN(n15872) );
  AOI21_X1 U18001 ( .B1(n15920), .B2(n22260), .A(n15872), .ZN(n15873) );
  OAI21_X1 U18002 ( .B1(n15917), .B2(n22246), .A(n15873), .ZN(P1_U2831) );
  AOI22_X1 U18003 ( .A1(n21977), .A2(n20528), .B1(n16183), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n15874) );
  OAI21_X1 U18004 ( .B1(n15917), .B2(n16189), .A(n15874), .ZN(P1_U2863) );
  OAI21_X1 U18005 ( .B1(n15833), .B2(n15876), .A(n15875), .ZN(n15901) );
  XOR2_X1 U18006 ( .A(n15878), .B(n15877), .Z(n17163) );
  INV_X1 U18007 ( .A(n17163), .ZN(n19018) );
  OAI22_X1 U18008 ( .A1(n16818), .A2(n19018), .B1(n16817), .B2(n15879), .ZN(
        n15881) );
  NOR2_X1 U18009 ( .A1(n16819), .A2(n20153), .ZN(n15880) );
  AOI211_X1 U18010 ( .C1(BUF1_REG_18__SCAN_IN), .C2(n20064), .A(n15881), .B(
        n15880), .ZN(n15883) );
  NAND2_X1 U18011 ( .A1(n20063), .A2(BUF2_REG_18__SCAN_IN), .ZN(n15882) );
  OAI211_X1 U18012 ( .C1(n15901), .C2(n20012), .A(n15883), .B(n15882), .ZN(
        P2_U2901) );
  OAI21_X1 U18013 ( .B1(n15860), .B2(n15885), .A(n15884), .ZN(n16427) );
  INV_X1 U18014 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n16422) );
  OAI21_X1 U18015 ( .B1(n15916), .B2(n15886), .A(n16422), .ZN(n15895) );
  NOR3_X1 U18016 ( .A1(n16422), .A2(n15916), .A3(n15887), .ZN(n15976) );
  OAI21_X1 U18017 ( .B1(n15976), .B2(n22220), .A(n22104), .ZN(n22141) );
  AND2_X1 U18018 ( .A1(n15889), .A2(n15888), .ZN(n15890) );
  OR2_X1 U18019 ( .A1(n15890), .A2(n16186), .ZN(n21985) );
  NAND2_X1 U18020 ( .A1(n22235), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n15891) );
  OAI211_X1 U18021 ( .C1(n21985), .C2(n22267), .A(n22092), .B(n15891), .ZN(
        n15894) );
  OAI22_X1 U18022 ( .A1(n15892), .A2(n22256), .B1(n22251), .B2(n16423), .ZN(
        n15893) );
  AOI211_X1 U18023 ( .C1(n15895), .C2(n22141), .A(n15894), .B(n15893), .ZN(
        n15896) );
  OAI21_X1 U18024 ( .B1(n16427), .B2(n22246), .A(n15896), .ZN(P1_U2830) );
  NAND2_X1 U18025 ( .A1(n11141), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n15900) );
  NAND2_X1 U18026 ( .A1(n15831), .A2(n15897), .ZN(n15898) );
  NAND2_X1 U18027 ( .A1(n15908), .A2(n15898), .ZN(n19019) );
  OR2_X1 U18028 ( .A1(n19019), .A2(n11141), .ZN(n15899) );
  OAI211_X1 U18029 ( .C1(n15901), .C2(n16740), .A(n15900), .B(n15899), .ZN(
        P2_U2869) );
  INV_X1 U18030 ( .A(n16212), .ZN(n15903) );
  OAI222_X1 U18031 ( .A1(n15917), .A2(n16238), .B1(n16268), .B2(n15903), .C1(
        n15902), .C2(n16265), .ZN(P1_U2895) );
  INV_X1 U18032 ( .A(n16208), .ZN(n15905) );
  OAI222_X1 U18033 ( .A1(n16427), .A2(n16238), .B1(n16268), .B2(n15905), .C1(
        n15904), .C2(n16265), .ZN(P1_U2894) );
  INV_X1 U18034 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n15906) );
  OAI222_X1 U18035 ( .A1(n21985), .A2(n20510), .B1(n15906), .B2(n20524), .C1(
        n16427), .C2(n16189), .ZN(P1_U2862) );
  AND2_X1 U18036 ( .A1(n15908), .A2(n15907), .ZN(n15909) );
  OR2_X1 U18037 ( .A1(n15909), .A2(n16737), .ZN(n17147) );
  AOI21_X1 U18038 ( .B1(n15911), .B2(n15875), .A(n15910), .ZN(n16812) );
  NAND2_X1 U18039 ( .A1(n16812), .A2(n16732), .ZN(n15913) );
  NAND2_X1 U18040 ( .A1(n11141), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n15912) );
  OAI211_X1 U18041 ( .C1(n17147), .C2(n11141), .A(n15913), .B(n15912), .ZN(
        P2_U2868) );
  OAI21_X1 U18042 ( .B1(n15915), .B2(n15914), .A(n16411), .ZN(n21978) );
  OAI22_X1 U18043 ( .A1(n16405), .A2(n15869), .B1(n22049), .B2(n15916), .ZN(
        n15919) );
  NOR2_X1 U18044 ( .A1(n15917), .A2(n16428), .ZN(n15918) );
  AOI211_X1 U18045 ( .C1(n20584), .C2(n15920), .A(n15919), .B(n15918), .ZN(
        n15921) );
  OAI21_X1 U18046 ( .B1(n21978), .B2(n22268), .A(n15921), .ZN(P1_U2990) );
  NAND2_X1 U18047 ( .A1(n15884), .A2(n15922), .ZN(n15923) );
  NAND2_X1 U18048 ( .A1(n15926), .A2(n15923), .ZN(n15928) );
  XOR2_X1 U18049 ( .A(n15927), .B(n15928), .Z(n22144) );
  INV_X1 U18050 ( .A(n22144), .ZN(n16190) );
  INV_X1 U18051 ( .A(n16204), .ZN(n15925) );
  OAI222_X1 U18052 ( .A1(n16238), .A2(n16190), .B1(n16268), .B2(n15925), .C1(
        n15924), .C2(n16265), .ZN(P1_U2893) );
  OAI21_X1 U18053 ( .B1(n15928), .B2(n15927), .A(n15926), .ZN(n15930) );
  AND2_X1 U18054 ( .A1(n15930), .A2(n15929), .ZN(n16135) );
  NOR2_X1 U18055 ( .A1(n15930), .A2(n15929), .ZN(n15931) );
  INV_X1 U18056 ( .A(n16201), .ZN(n15933) );
  OAI222_X1 U18057 ( .A1(n22159), .A2(n16238), .B1(n16268), .B2(n15933), .C1(
        n15932), .C2(n16265), .ZN(P1_U2892) );
  INV_X1 U18058 ( .A(n16260), .ZN(n15935) );
  AOI21_X1 U18059 ( .B1(n15936), .B2(n15934), .A(n15935), .ZN(n16395) );
  INV_X1 U18060 ( .A(n16395), .ZN(n16181) );
  INV_X1 U18061 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n15938) );
  INV_X1 U18062 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n22153) );
  INV_X1 U18063 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n22151) );
  NAND2_X1 U18064 ( .A1(n15976), .A2(n22236), .ZN(n22152) );
  NOR3_X1 U18065 ( .A1(n22153), .A2(n22151), .A3(n22152), .ZN(n16145) );
  NAND2_X1 U18066 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n16145), .ZN(n15937) );
  AOI211_X1 U18067 ( .C1(n15938), .C2(n15937), .A(n22167), .B(n22177), .ZN(
        n15944) );
  AND2_X1 U18068 ( .A1(n16139), .A2(n15939), .ZN(n15940) );
  OR2_X1 U18069 ( .A1(n15940), .A2(n20507), .ZN(n21906) );
  INV_X1 U18070 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n16182) );
  OAI22_X1 U18071 ( .A1(n21906), .A2(n22267), .B1(n22254), .B2(n16182), .ZN(
        n15943) );
  INV_X1 U18072 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n15941) );
  OAI22_X1 U18073 ( .A1(n16393), .A2(n22251), .B1(n22256), .B2(n15941), .ZN(
        n15942) );
  NOR4_X1 U18074 ( .A1(n15944), .A2(n22197), .A3(n15943), .A4(n15942), .ZN(
        n15945) );
  OAI21_X1 U18075 ( .B1(n16181), .B2(n22246), .A(n15945), .ZN(P1_U2826) );
  AOI22_X1 U18076 ( .A1(n15946), .A2(n16194), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n16252), .ZN(n15947) );
  OAI21_X1 U18077 ( .B1(n16181), .B2(n16238), .A(n15947), .ZN(P1_U2890) );
  OR2_X1 U18078 ( .A1(n16188), .A2(n15948), .ZN(n15949) );
  NAND2_X1 U18079 ( .A1(n16137), .A2(n15949), .ZN(n22149) );
  INV_X1 U18080 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n22148) );
  OAI222_X1 U18081 ( .A1(n22149), .A2(n20510), .B1(n22148), .B2(n20524), .C1(
        n16189), .C2(n22159), .ZN(P1_U2860) );
  INV_X1 U18082 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n21112) );
  INV_X1 U18083 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n15958) );
  NAND3_X1 U18084 ( .A1(n19470), .A2(n15950), .A3(n21197), .ZN(n15952) );
  NAND2_X1 U18085 ( .A1(n15951), .A2(n21813), .ZN(n15968) );
  NAND2_X1 U18086 ( .A1(n15952), .A2(n15968), .ZN(n21165) );
  INV_X1 U18087 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n20816) );
  NAND2_X1 U18088 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(P3_EBX_REG_4__SCAN_IN), 
        .ZN(n15956) );
  NAND4_X1 U18089 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(P3_EBX_REG_2__SCAN_IN), 
        .A3(P3_EBX_REG_0__SCAN_IN), .A4(P3_EBX_REG_1__SCAN_IN), .ZN(n17990) );
  INV_X1 U18090 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n15954) );
  NAND4_X1 U18091 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(P3_EBX_REG_12__SCAN_IN), 
        .A3(P3_EBX_REG_11__SCAN_IN), .A4(P3_EBX_REG_10__SCAN_IN), .ZN(n18031)
         );
  NAND4_X1 U18092 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(P3_EBX_REG_15__SCAN_IN), 
        .A3(P3_EBX_REG_14__SCAN_IN), .A4(P3_EBX_REG_9__SCAN_IN), .ZN(n15953)
         );
  NOR4_X1 U18093 ( .A1(n20816), .A2(n15956), .A3(n17990), .A4(n15955), .ZN(
        n18358) );
  NAND2_X1 U18094 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n18358), .ZN(n18357) );
  NOR2_X1 U18095 ( .A1(n18365), .A2(n18357), .ZN(n18320) );
  NAND2_X1 U18096 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n18320), .ZN(n18324) );
  NAND2_X1 U18097 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n18340), .ZN(n18241) );
  AND4_X1 U18098 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .A4(P3_EBX_REG_21__SCAN_IN), .ZN(n18243)
         );
  NAND4_X1 U18099 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(P3_EBX_REG_25__SCAN_IN), .A4(n18243), .ZN(n15957) );
  NOR4_X1 U18100 ( .A1(n21112), .A2(n15958), .A3(n18241), .A4(n15957), .ZN(
        n18227) );
  NAND2_X1 U18101 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n18227), .ZN(n15959) );
  NOR2_X1 U18102 ( .A1(n21267), .A2(n15959), .ZN(n15961) );
  NAND2_X1 U18103 ( .A1(n18362), .A2(n15959), .ZN(n18228) );
  INV_X1 U18104 ( .A(n18228), .ZN(n15960) );
  MUX2_X1 U18105 ( .A(n15961), .B(n15960), .S(P3_EBX_REG_31__SCAN_IN), .Z(
        P3_U2672) );
  NAND2_X1 U18106 ( .A1(n21855), .A2(n21354), .ZN(n17369) );
  INV_X1 U18107 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n21820) );
  NAND2_X1 U18108 ( .A1(n17747), .A2(n21820), .ZN(n15962) );
  NAND2_X1 U18109 ( .A1(n15964), .A2(n15962), .ZN(n21818) );
  NOR2_X1 U18110 ( .A1(n17369), .A2(n21818), .ZN(n15970) );
  INV_X1 U18111 ( .A(n15963), .ZN(n17756) );
  NOR2_X1 U18112 ( .A1(n22341), .A2(n21817), .ZN(n15967) );
  INV_X1 U18113 ( .A(n15967), .ZN(n15965) );
  AOI211_X1 U18114 ( .C1(n17755), .C2(n15967), .A(n21167), .B(n15966), .ZN(
        n15969) );
  NAND2_X1 U18115 ( .A1(n15969), .A2(n15968), .ZN(n21826) );
  NOR2_X1 U18116 ( .A1(n21862), .A2(n18371), .ZN(n17753) );
  AOI22_X1 U18117 ( .A1(n21845), .A2(n21826), .B1(P3_FLUSH_REG_SCAN_IN), .B2(
        n17753), .ZN(n21396) );
  NAND2_X1 U18118 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n21862), .ZN(n21852) );
  NAND2_X1 U18119 ( .A1(n21396), .A2(n21852), .ZN(n21393) );
  MUX2_X1 U18120 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n15970), .S(
        n21393), .Z(P3_U3284) );
  MUX2_X1 U18121 ( .A(n15971), .B(n14002), .S(n16052), .Z(n15975) );
  OAI22_X1 U18122 ( .A1(n15973), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        P1_EBX_REG_31__SCAN_IN), .B2(n15972), .ZN(n15974) );
  AOI22_X1 U18123 ( .A1(n22244), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B1(
        P1_EBX_REG_31__SCAN_IN), .B2(n22235), .ZN(n15984) );
  INV_X1 U18124 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n22225) );
  INV_X1 U18125 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n16113) );
  INV_X1 U18126 ( .A(n15976), .ZN(n15979) );
  INV_X1 U18127 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n22008) );
  INV_X1 U18128 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n22176) );
  NAND4_X1 U18129 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_14__SCAN_IN), 
        .A3(P1_REIP_REG_13__SCAN_IN), .A4(P1_REIP_REG_12__SCAN_IN), .ZN(n15977) );
  NOR4_X1 U18130 ( .A1(n22008), .A2(n22176), .A3(n22153), .A4(n15977), .ZN(
        n15978) );
  NAND3_X1 U18131 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .A3(n15978), .ZN(n16114) );
  NOR3_X1 U18132 ( .A1(n16113), .A2(n15979), .A3(n16114), .ZN(n22210) );
  NAND2_X1 U18133 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n22210), .ZN(n22221) );
  NOR2_X1 U18134 ( .A1(n22225), .A2(n22221), .ZN(n22237) );
  NAND2_X1 U18135 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n22237), .ZN(n22238) );
  INV_X1 U18136 ( .A(n22238), .ZN(n15980) );
  NAND2_X1 U18137 ( .A1(n22258), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n16101) );
  INV_X1 U18138 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n16310) );
  INV_X1 U18139 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20464) );
  INV_X1 U18140 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20467) );
  NOR2_X1 U18141 ( .A1(n16092), .A2(n20467), .ZN(n16076) );
  NAND2_X1 U18142 ( .A1(n16076), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n16064) );
  INV_X1 U18143 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n16281) );
  NOR2_X1 U18144 ( .A1(n16064), .A2(n16281), .ZN(n16054) );
  NAND2_X1 U18145 ( .A1(n16054), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n15982) );
  NAND2_X1 U18146 ( .A1(n22166), .A2(n15982), .ZN(n15981) );
  MUX2_X1 U18147 ( .A(n15982), .B(n15981), .S(P1_REIP_REG_31__SCAN_IN), .Z(
        n15983) );
  OAI211_X1 U18148 ( .C1(n16429), .C2(n22267), .A(n15984), .B(n15983), .ZN(
        n15985) );
  AOI21_X1 U18149 ( .B1(n15990), .B2(n22262), .A(n15985), .ZN(n15986) );
  INV_X1 U18150 ( .A(n15986), .ZN(P1_U2809) );
  NOR2_X1 U18151 ( .A1(n15992), .A2(n15987), .ZN(n15988) );
  NAND2_X1 U18152 ( .A1(n16265), .A2(n15988), .ZN(n16191) );
  AND2_X1 U18153 ( .A1(n16265), .A2(n16033), .ZN(n15989) );
  NAND2_X1 U18154 ( .A1(n15990), .A2(n15989), .ZN(n15995) );
  NOR3_X1 U18155 ( .A1(n16252), .A2(n15992), .A3(n15991), .ZN(n15993) );
  AOI22_X1 U18156 ( .A1(n16256), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P1_EAX_REG_31__SCAN_IN), .B2(n16252), .ZN(n15994) );
  OAI211_X1 U18157 ( .C1(n16191), .C2(n15086), .A(n15995), .B(n15994), .ZN(
        P1_U2873) );
  OAI22_X1 U18158 ( .A1(n16001), .A2(n17319), .B1(n15997), .B2(n15996), .ZN(
        n16007) );
  OAI21_X1 U18159 ( .B1(n16000), .B2(n15999), .A(n15998), .ZN(n17832) );
  OAI22_X1 U18160 ( .A1(n17832), .A2(n19178), .B1(n16001), .B2(n19176), .ZN(
        n16006) );
  AOI21_X1 U18161 ( .B1(n16004), .B2(n16003), .A(n16002), .ZN(n16005) );
  AOI211_X1 U18162 ( .C1(n17174), .C2(n16007), .A(n16006), .B(n16005), .ZN(
        n16013) );
  NOR2_X1 U18163 ( .A1(n18976), .A2(n17956), .ZN(n17834) );
  OAI21_X1 U18164 ( .B1(n16010), .B2(n16009), .A(n16008), .ZN(n17831) );
  NOR2_X1 U18165 ( .A1(n19187), .A2(n17831), .ZN(n16011) );
  AOI211_X1 U18166 ( .C1(n19208), .C2(n17889), .A(n17834), .B(n16011), .ZN(
        n16012) );
  OAI211_X1 U18167 ( .C1(n16014), .C2(n17283), .A(n16013), .B(n16012), .ZN(
        P2_U3044) );
  AOI22_X1 U18168 ( .A1(n20062), .A2(n19742), .B1(P2_EAX_REG_30__SCAN_IN), 
        .B2(n20060), .ZN(n16016) );
  NAND2_X1 U18169 ( .A1(n20063), .A2(BUF2_REG_30__SCAN_IN), .ZN(n16015) );
  OAI211_X1 U18170 ( .C1(n16017), .C2(n16818), .A(n16016), .B(n16015), .ZN(
        n16018) );
  AOI21_X1 U18171 ( .B1(BUF1_REG_30__SCAN_IN), .B2(n20064), .A(n16018), .ZN(
        n16019) );
  OAI21_X1 U18172 ( .B1(n16020), .B2(n20012), .A(n16019), .ZN(P2_U2889) );
  NAND4_X1 U18173 ( .A1(n12961), .A2(n16023), .A3(n16022), .A4(n16021), .ZN(
        n16025) );
  OAI21_X1 U18174 ( .B1(n16026), .B2(n16025), .A(n16024), .ZN(n16027) );
  NAND2_X1 U18175 ( .A1(n16027), .A2(n16036), .ZN(n16035) );
  INV_X1 U18176 ( .A(n16028), .ZN(n16031) );
  AOI22_X1 U18177 ( .A1(n16032), .A2(n16031), .B1(n16030), .B2(n16029), .ZN(
        n16034) );
  AOI21_X1 U18178 ( .B1(n16035), .B2(n16034), .A(n16033), .ZN(n17807) );
  AOI22_X1 U18179 ( .A1(n16039), .A2(n16038), .B1(n16037), .B2(n16036), .ZN(
        n20595) );
  OAI21_X1 U18180 ( .B1(n16041), .B2(n16040), .A(n21876), .ZN(n21879) );
  NAND2_X1 U18181 ( .A1(n20595), .A2(n21879), .ZN(n17800) );
  AND2_X1 U18182 ( .A1(n17800), .A2(n16042), .ZN(n22270) );
  MUX2_X1 U18183 ( .A(P1_MORE_REG_SCAN_IN), .B(n17807), .S(n22270), .Z(
        P1_U3484) );
  OAI22_X1 U18184 ( .A1(n22256), .A2(n16275), .B1(n16043), .B2(n22254), .ZN(
        n16047) );
  INV_X1 U18185 ( .A(n16273), .ZN(n16045) );
  XNOR2_X1 U18186 ( .A(n16054), .B(P1_REIP_REG_30__SCAN_IN), .ZN(n16044) );
  OAI22_X1 U18187 ( .A1(n22251), .A2(n16045), .B1(n22177), .B2(n16044), .ZN(
        n16046) );
  AOI211_X1 U18188 ( .C1(n16465), .C2(n22199), .A(n16047), .B(n16046), .ZN(
        n16048) );
  OAI21_X1 U18189 ( .B1(n16197), .B2(n22246), .A(n16048), .ZN(P1_U2810) );
  INV_X1 U18190 ( .A(n16285), .ZN(n16200) );
  OAI21_X1 U18191 ( .B1(n11210), .B2(n16053), .A(n16052), .ZN(n16148) );
  INV_X1 U18192 ( .A(n16148), .ZN(n16471) );
  NAND2_X1 U18193 ( .A1(n22166), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n16055) );
  AOI21_X1 U18194 ( .B1(n16055), .B2(n16064), .A(n16054), .ZN(n16058) );
  AOI22_X1 U18195 ( .A1(n22244), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B1(
        n22235), .B2(P1_EBX_REG_29__SCAN_IN), .ZN(n16056) );
  OAI21_X1 U18196 ( .B1(n22251), .B2(n16283), .A(n16056), .ZN(n16057) );
  AOI211_X1 U18197 ( .C1(n16471), .C2(n22199), .A(n16058), .B(n16057), .ZN(
        n16059) );
  OAI21_X1 U18198 ( .B1(n16200), .B2(n22246), .A(n16059), .ZN(P1_U2811) );
  AOI21_X1 U18199 ( .B1(n16062), .B2(n16075), .A(n11210), .ZN(n16480) );
  INV_X1 U18200 ( .A(n16063), .ZN(n16296) );
  INV_X1 U18201 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n16294) );
  NOR2_X1 U18202 ( .A1(n22177), .A2(n16294), .ZN(n16065) );
  OAI21_X1 U18203 ( .B1(n16065), .B2(n16076), .A(n16064), .ZN(n16067) );
  AOI22_X1 U18204 ( .A1(n22244), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B1(
        n22235), .B2(P1_EBX_REG_28__SCAN_IN), .ZN(n16066) );
  OAI211_X1 U18205 ( .C1(n22251), .C2(n16296), .A(n16067), .B(n16066), .ZN(
        n16068) );
  AOI21_X1 U18206 ( .B1(n16480), .B2(n22199), .A(n16068), .ZN(n16069) );
  OAI21_X1 U18207 ( .B1(n16293), .B2(n22246), .A(n16069), .ZN(P1_U2812) );
  AOI21_X1 U18208 ( .B1(n16071), .B2(n16070), .A(n16060), .ZN(n16305) );
  INV_X1 U18209 ( .A(n16305), .ZN(n16207) );
  NAND2_X1 U18210 ( .A1(n16072), .A2(n16073), .ZN(n16074) );
  NAND2_X1 U18211 ( .A1(n16075), .A2(n16074), .ZN(n16151) );
  INV_X1 U18212 ( .A(n16151), .ZN(n16489) );
  NAND2_X1 U18213 ( .A1(n22166), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n16077) );
  AOI21_X1 U18214 ( .B1(n16077), .B2(n16092), .A(n16076), .ZN(n16080) );
  AOI22_X1 U18215 ( .A1(n22244), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B1(
        n22235), .B2(P1_EBX_REG_27__SCAN_IN), .ZN(n16078) );
  OAI21_X1 U18216 ( .B1(n22251), .B2(n16303), .A(n16078), .ZN(n16079) );
  AOI211_X1 U18217 ( .C1(n16489), .C2(n22199), .A(n16080), .B(n16079), .ZN(
        n16081) );
  OAI21_X1 U18218 ( .B1(n16207), .B2(n22246), .A(n16081), .ZN(P1_U2813) );
  OR2_X1 U18219 ( .A1(n16104), .A2(n16082), .ZN(n16083) );
  NAND2_X1 U18220 ( .A1(n16072), .A2(n16083), .ZN(n16492) );
  NAND2_X1 U18221 ( .A1(n16084), .A2(n16158), .ZN(n16160) );
  INV_X1 U18222 ( .A(n16070), .ZN(n16085) );
  AOI21_X2 U18223 ( .B1(n16086), .B2(n16095), .A(n16085), .ZN(n16314) );
  NAND2_X1 U18224 ( .A1(n16314), .A2(n22262), .ZN(n16094) );
  NAND3_X1 U18225 ( .A1(n22258), .A2(P1_REIP_REG_24__SCAN_IN), .A3(
        P1_REIP_REG_25__SCAN_IN), .ZN(n16087) );
  OAI21_X1 U18226 ( .B1(n22177), .B2(n16310), .A(n16087), .ZN(n16091) );
  INV_X1 U18227 ( .A(n16088), .ZN(n16312) );
  AOI22_X1 U18228 ( .A1(n22244), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B1(
        n22235), .B2(P1_EBX_REG_26__SCAN_IN), .ZN(n16089) );
  OAI21_X1 U18229 ( .B1(n22251), .B2(n16312), .A(n16089), .ZN(n16090) );
  AOI21_X1 U18230 ( .B1(n16092), .B2(n16091), .A(n16090), .ZN(n16093) );
  OAI211_X1 U18231 ( .C1(n22267), .C2(n16492), .A(n16094), .B(n16093), .ZN(
        P1_U2814) );
  INV_X1 U18232 ( .A(n16095), .ZN(n16096) );
  AOI21_X1 U18233 ( .B1(n16097), .B2(n16160), .A(n16096), .ZN(n16321) );
  INV_X1 U18234 ( .A(n16321), .ZN(n16215) );
  AOI21_X1 U18235 ( .B1(n22238), .B2(n22236), .A(n16098), .ZN(n22242) );
  INV_X1 U18236 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n16327) );
  NAND2_X1 U18237 ( .A1(n22258), .A2(n16327), .ZN(n16099) );
  NAND2_X1 U18238 ( .A1(n22242), .A2(n16099), .ZN(n22259) );
  INV_X1 U18239 ( .A(n16100), .ZN(n16319) );
  INV_X1 U18240 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n16154) );
  OAI22_X1 U18241 ( .A1(n16101), .A2(P1_REIP_REG_25__SCAN_IN), .B1(n16154), 
        .B2(n22254), .ZN(n16102) );
  AOI21_X1 U18242 ( .B1(n22244), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16102), .ZN(n16103) );
  OAI21_X1 U18243 ( .B1(n22251), .B2(n16319), .A(n16103), .ZN(n16108) );
  INV_X1 U18244 ( .A(n16104), .ZN(n16105) );
  OAI21_X1 U18245 ( .B1(n16106), .B2(n16156), .A(n16105), .ZN(n16508) );
  NOR2_X1 U18246 ( .A1(n16508), .A2(n22267), .ZN(n16107) );
  AOI211_X1 U18247 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(n22259), .A(n16108), 
        .B(n16107), .ZN(n16109) );
  OAI21_X1 U18248 ( .B1(n16215), .B2(n22246), .A(n16109), .ZN(P1_U2815) );
  AOI21_X1 U18249 ( .B1(n16110), .B2(n16112), .A(n16111), .ZN(n16367) );
  INV_X1 U18250 ( .A(n16367), .ZN(n16239) );
  OAI21_X1 U18251 ( .B1(n22210), .B2(n22220), .A(n22104), .ZN(n22222) );
  OAI21_X1 U18252 ( .B1(n16114), .B2(n22152), .A(n16113), .ZN(n16121) );
  INV_X1 U18253 ( .A(n16115), .ZN(n16116) );
  OAI21_X1 U18254 ( .B1(n20522), .B2(n16117), .A(n16116), .ZN(n16565) );
  AOI22_X1 U18255 ( .A1(n22260), .A2(n16363), .B1(n22235), .B2(
        P1_EBX_REG_20__SCAN_IN), .ZN(n16119) );
  NAND2_X1 U18256 ( .A1(n22244), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16118) );
  OAI211_X1 U18257 ( .C1(n16565), .C2(n22267), .A(n16119), .B(n16118), .ZN(
        n16120) );
  AOI21_X1 U18258 ( .B1(n22222), .B2(n16121), .A(n16120), .ZN(n16122) );
  OAI21_X1 U18259 ( .B1(n16239), .B2(n22246), .A(n16122), .ZN(P1_U2820) );
  OAI21_X1 U18260 ( .B1(n16123), .B2(n16125), .A(n16124), .ZN(n20503) );
  INV_X1 U18261 ( .A(n16169), .ZN(n16126) );
  AOI21_X1 U18262 ( .B1(n16127), .B2(n16178), .A(n16126), .ZN(n22026) );
  INV_X1 U18263 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n20505) );
  AOI22_X1 U18264 ( .A1(n22244), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n22260), .B2(n20583), .ZN(n16128) );
  OAI211_X1 U18265 ( .C1(n22254), .C2(n20505), .A(n16128), .B(n22092), .ZN(
        n16129) );
  AOI21_X1 U18266 ( .B1(n22026), .B2(n22199), .A(n16129), .ZN(n16133) );
  INV_X1 U18267 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n16130) );
  NAND3_X1 U18268 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(n22167), .ZN(n22179) );
  NOR2_X1 U18269 ( .A1(n16130), .A2(n22179), .ZN(n22204) );
  NOR2_X1 U18270 ( .A1(n22177), .A2(n22204), .ZN(n22202) );
  NAND2_X1 U18271 ( .A1(n16130), .A2(n22179), .ZN(n16131) );
  NAND2_X1 U18272 ( .A1(n22202), .A2(n16131), .ZN(n16132) );
  OAI211_X1 U18273 ( .C1(n20503), .C2(n22246), .A(n16133), .B(n16132), .ZN(
        P1_U2823) );
  OAI21_X1 U18274 ( .B1(n16135), .B2(n16134), .A(n15934), .ZN(n16410) );
  INV_X1 U18275 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n17656) );
  NAND2_X1 U18276 ( .A1(n16137), .A2(n16136), .ZN(n16138) );
  AND2_X1 U18277 ( .A1(n16139), .A2(n16138), .ZN(n21895) );
  INV_X1 U18278 ( .A(n21895), .ZN(n16141) );
  NOR2_X1 U18279 ( .A1(n22177), .A2(n16145), .ZN(n22155) );
  AOI22_X1 U18280 ( .A1(n22235), .A2(P1_EBX_REG_13__SCAN_IN), .B1(
        P1_REIP_REG_13__SCAN_IN), .B2(n22155), .ZN(n16140) );
  OAI211_X1 U18281 ( .C1(n16141), .C2(n22267), .A(n16140), .B(n22092), .ZN(
        n16144) );
  INV_X1 U18282 ( .A(n16407), .ZN(n16142) );
  OAI22_X1 U18283 ( .A1(n16404), .A2(n22256), .B1(n22251), .B2(n16142), .ZN(
        n16143) );
  AOI211_X1 U18284 ( .C1(n16145), .C2(n17656), .A(n16144), .B(n16143), .ZN(
        n16146) );
  OAI21_X1 U18285 ( .B1(n16410), .B2(n22246), .A(n16146), .ZN(P1_U2827) );
  INV_X1 U18286 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n16147) );
  OAI22_X1 U18287 ( .A1(n16429), .A2(n20510), .B1(n16147), .B2(n20524), .ZN(
        P1_U2841) );
  INV_X1 U18288 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n16149) );
  OAI222_X1 U18289 ( .A1(n16149), .A2(n20524), .B1(n20510), .B2(n16148), .C1(
        n16200), .C2(n16189), .ZN(P1_U2843) );
  AOI22_X1 U18290 ( .A1(n16480), .A2(n20528), .B1(n16183), .B2(
        P1_EBX_REG_28__SCAN_IN), .ZN(n16150) );
  OAI21_X1 U18291 ( .B1(n16293), .B2(n16189), .A(n16150), .ZN(P1_U2844) );
  INV_X1 U18292 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n16152) );
  OAI222_X1 U18293 ( .A1(n16152), .A2(n20524), .B1(n20510), .B2(n16151), .C1(
        n16207), .C2(n16189), .ZN(P1_U2845) );
  INV_X1 U18294 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n16153) );
  INV_X1 U18295 ( .A(n16314), .ZN(n16211) );
  OAI222_X1 U18296 ( .A1(n16153), .A2(n20524), .B1(n20510), .B2(n16492), .C1(
        n16211), .C2(n16189), .ZN(P1_U2846) );
  OAI222_X1 U18297 ( .A1(n16154), .A2(n20524), .B1(n20510), .B2(n16508), .C1(
        n16215), .C2(n16189), .ZN(P1_U2847) );
  INV_X1 U18298 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n22253) );
  AND2_X1 U18299 ( .A1(n16527), .A2(n16155), .ZN(n16157) );
  OR2_X1 U18300 ( .A1(n16157), .A2(n16156), .ZN(n22266) );
  OR2_X1 U18301 ( .A1(n16084), .A2(n16158), .ZN(n16159) );
  OAI222_X1 U18302 ( .A1(n22253), .A2(n20524), .B1(n20510), .B2(n22266), .C1(
        n16219), .C2(n16189), .ZN(P1_U2848) );
  INV_X1 U18303 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n22224) );
  OR2_X1 U18304 ( .A1(n16560), .A2(n16161), .ZN(n16162) );
  NAND2_X1 U18305 ( .A1(n16525), .A2(n16162), .ZN(n22234) );
  AND2_X1 U18306 ( .A1(n16163), .A2(n16164), .ZN(n16165) );
  OR2_X1 U18307 ( .A1(n16165), .A2(n11214), .ZN(n22230) );
  OAI222_X1 U18308 ( .A1(n22224), .A2(n20524), .B1(n20510), .B2(n22234), .C1(
        n22230), .C2(n16189), .ZN(P1_U2850) );
  INV_X1 U18309 ( .A(n16565), .ZN(n16166) );
  AOI22_X1 U18310 ( .A1(n16166), .A2(n20528), .B1(n16183), .B2(
        P1_EBX_REG_20__SCAN_IN), .ZN(n16167) );
  OAI21_X1 U18311 ( .B1(n16239), .B2(n16189), .A(n16167), .ZN(P1_U2852) );
  NAND2_X1 U18312 ( .A1(n16169), .A2(n16168), .ZN(n16170) );
  NAND2_X1 U18313 ( .A1(n20520), .A2(n16170), .ZN(n22193) );
  INV_X1 U18314 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n16173) );
  AOI21_X1 U18315 ( .B1(n16172), .B2(n16124), .A(n16171), .ZN(n16373) );
  INV_X1 U18316 ( .A(n16373), .ZN(n22190) );
  OAI222_X1 U18317 ( .A1(n22193), .A2(n20510), .B1(n16173), .B2(n20524), .C1(
        n22190), .C2(n16189), .ZN(P1_U2854) );
  NOR2_X1 U18318 ( .A1(n11196), .A2(n16174), .ZN(n16175) );
  OR2_X1 U18319 ( .A1(n16123), .A2(n16175), .ZN(n16385) );
  INV_X1 U18320 ( .A(n16385), .ZN(n22180) );
  OR2_X1 U18321 ( .A1(n20509), .A2(n16176), .ZN(n16177) );
  NAND2_X1 U18322 ( .A1(n16178), .A2(n16177), .ZN(n22183) );
  OAI22_X1 U18323 ( .A1(n22183), .A2(n20510), .B1(n22171), .B2(n20524), .ZN(
        n16179) );
  AOI21_X1 U18324 ( .B1(n22180), .B2(n13916), .A(n16179), .ZN(n16180) );
  INV_X1 U18325 ( .A(n16180), .ZN(P1_U2856) );
  OAI222_X1 U18326 ( .A1(n21906), .A2(n20510), .B1(n16182), .B2(n20524), .C1(
        n16189), .C2(n16181), .ZN(P1_U2858) );
  AOI22_X1 U18327 ( .A1(n21895), .A2(n20528), .B1(n16183), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n16184) );
  OAI21_X1 U18328 ( .B1(n16410), .B2(n16189), .A(n16184), .ZN(P1_U2859) );
  INV_X1 U18329 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n22138) );
  NOR2_X1 U18330 ( .A1(n16186), .A2(n16185), .ZN(n16187) );
  OR2_X1 U18331 ( .A1(n16188), .A2(n16187), .ZN(n22142) );
  OAI222_X1 U18332 ( .A1(n22138), .A2(n20524), .B1(n20510), .B2(n22142), .C1(
        n16190), .C2(n16189), .ZN(P1_U2861) );
  AOI22_X1 U18333 ( .A1(n16253), .A2(DATAI_30_), .B1(P1_EAX_REG_30__SCAN_IN), 
        .B2(n16252), .ZN(n16196) );
  INV_X1 U18334 ( .A(n16192), .ZN(n16193) );
  NOR2_X2 U18335 ( .A1(n16252), .A2(n16193), .ZN(n16255) );
  AOI22_X1 U18336 ( .A1(n16256), .A2(BUF1_REG_30__SCAN_IN), .B1(n16255), .B2(
        n16194), .ZN(n16195) );
  OAI211_X1 U18337 ( .C1(n16197), .C2(n16238), .A(n16196), .B(n16195), .ZN(
        P1_U2874) );
  AOI22_X1 U18338 ( .A1(n16253), .A2(DATAI_29_), .B1(P1_EAX_REG_29__SCAN_IN), 
        .B2(n16252), .ZN(n16199) );
  AOI22_X1 U18339 ( .A1(n16256), .A2(BUF1_REG_29__SCAN_IN), .B1(n16255), .B2(
        n16264), .ZN(n16198) );
  OAI211_X1 U18340 ( .C1(n16200), .C2(n16238), .A(n16199), .B(n16198), .ZN(
        P1_U2875) );
  AOI22_X1 U18341 ( .A1(n16253), .A2(DATAI_28_), .B1(P1_EAX_REG_28__SCAN_IN), 
        .B2(n16252), .ZN(n16203) );
  AOI22_X1 U18342 ( .A1(n16256), .A2(BUF1_REG_28__SCAN_IN), .B1(n16255), .B2(
        n16201), .ZN(n16202) );
  OAI211_X1 U18343 ( .C1(n16293), .C2(n16238), .A(n16203), .B(n16202), .ZN(
        P1_U2876) );
  AOI22_X1 U18344 ( .A1(n16253), .A2(DATAI_27_), .B1(P1_EAX_REG_27__SCAN_IN), 
        .B2(n16252), .ZN(n16206) );
  AOI22_X1 U18345 ( .A1(n16256), .A2(BUF1_REG_27__SCAN_IN), .B1(n16255), .B2(
        n16204), .ZN(n16205) );
  OAI211_X1 U18346 ( .C1(n16207), .C2(n16238), .A(n16206), .B(n16205), .ZN(
        P1_U2877) );
  AOI22_X1 U18347 ( .A1(n16253), .A2(DATAI_26_), .B1(P1_EAX_REG_26__SCAN_IN), 
        .B2(n16252), .ZN(n16210) );
  AOI22_X1 U18348 ( .A1(n16256), .A2(BUF1_REG_26__SCAN_IN), .B1(n16255), .B2(
        n16208), .ZN(n16209) );
  OAI211_X1 U18349 ( .C1(n16211), .C2(n16238), .A(n16210), .B(n16209), .ZN(
        P1_U2878) );
  AOI22_X1 U18350 ( .A1(n16253), .A2(DATAI_25_), .B1(P1_EAX_REG_25__SCAN_IN), 
        .B2(n16252), .ZN(n16214) );
  AOI22_X1 U18351 ( .A1(n16256), .A2(BUF1_REG_25__SCAN_IN), .B1(n16255), .B2(
        n16212), .ZN(n16213) );
  OAI211_X1 U18352 ( .C1(n16215), .C2(n16238), .A(n16214), .B(n16213), .ZN(
        P1_U2879) );
  AOI22_X1 U18353 ( .A1(n16253), .A2(DATAI_24_), .B1(P1_EAX_REG_24__SCAN_IN), 
        .B2(n16252), .ZN(n16218) );
  AOI22_X1 U18354 ( .A1(n16256), .A2(BUF1_REG_24__SCAN_IN), .B1(n16255), .B2(
        n16216), .ZN(n16217) );
  OAI211_X1 U18355 ( .C1(n16219), .C2(n16238), .A(n16218), .B(n16217), .ZN(
        P1_U2880) );
  NOR2_X1 U18356 ( .A1(n11214), .A2(n16220), .ZN(n16221) );
  OR2_X1 U18357 ( .A1(n16084), .A2(n16221), .ZN(n22247) );
  AOI22_X1 U18358 ( .A1(n16253), .A2(DATAI_23_), .B1(P1_EAX_REG_23__SCAN_IN), 
        .B2(n16252), .ZN(n16224) );
  AOI22_X1 U18359 ( .A1(n16256), .A2(BUF1_REG_23__SCAN_IN), .B1(n16255), .B2(
        n16222), .ZN(n16223) );
  OAI211_X1 U18360 ( .C1(n22247), .C2(n16238), .A(n16224), .B(n16223), .ZN(
        P1_U2881) );
  AOI22_X1 U18361 ( .A1(n16253), .A2(DATAI_22_), .B1(P1_EAX_REG_22__SCAN_IN), 
        .B2(n16252), .ZN(n16227) );
  AOI22_X1 U18362 ( .A1(n16256), .A2(BUF1_REG_22__SCAN_IN), .B1(n16255), .B2(
        n16225), .ZN(n16226) );
  OAI211_X1 U18363 ( .C1(n22230), .C2(n16238), .A(n16227), .B(n16226), .ZN(
        P1_U2882) );
  NAND2_X1 U18364 ( .A1(n16229), .A2(n16228), .ZN(n16230) );
  AND2_X1 U18365 ( .A1(n16163), .A2(n16230), .ZN(n22216) );
  INV_X1 U18366 ( .A(n22216), .ZN(n16234) );
  AOI22_X1 U18367 ( .A1(n16253), .A2(DATAI_21_), .B1(P1_EAX_REG_21__SCAN_IN), 
        .B2(n16252), .ZN(n16233) );
  AOI22_X1 U18368 ( .A1(n16256), .A2(BUF1_REG_21__SCAN_IN), .B1(n16255), .B2(
        n16231), .ZN(n16232) );
  OAI211_X1 U18369 ( .C1(n16234), .C2(n16238), .A(n16233), .B(n16232), .ZN(
        P1_U2883) );
  AOI22_X1 U18370 ( .A1(n16253), .A2(DATAI_20_), .B1(P1_EAX_REG_20__SCAN_IN), 
        .B2(n16252), .ZN(n16237) );
  AOI22_X1 U18371 ( .A1(n16256), .A2(BUF1_REG_20__SCAN_IN), .B1(n16255), .B2(
        n16235), .ZN(n16236) );
  OAI211_X1 U18372 ( .C1(n16239), .C2(n16238), .A(n16237), .B(n16236), .ZN(
        P1_U2884) );
  OR2_X1 U18373 ( .A1(n16171), .A2(n16240), .ZN(n16241) );
  AND2_X1 U18374 ( .A1(n16110), .A2(n16241), .ZN(n22200) );
  INV_X1 U18375 ( .A(n22200), .ZN(n16245) );
  AOI22_X1 U18376 ( .A1(n16253), .A2(DATAI_19_), .B1(P1_EAX_REG_19__SCAN_IN), 
        .B2(n16252), .ZN(n16244) );
  AOI22_X1 U18377 ( .A1(n16256), .A2(BUF1_REG_19__SCAN_IN), .B1(n16255), .B2(
        n16242), .ZN(n16243) );
  OAI211_X1 U18378 ( .C1(n16245), .C2(n16238), .A(n16244), .B(n16243), .ZN(
        P1_U2885) );
  AOI22_X1 U18379 ( .A1(n16253), .A2(DATAI_18_), .B1(P1_EAX_REG_18__SCAN_IN), 
        .B2(n16252), .ZN(n16248) );
  AOI22_X1 U18380 ( .A1(n16256), .A2(BUF1_REG_18__SCAN_IN), .B1(n16255), .B2(
        n16246), .ZN(n16247) );
  OAI211_X1 U18381 ( .C1(n22190), .C2(n16238), .A(n16248), .B(n16247), .ZN(
        P1_U2886) );
  AOI22_X1 U18382 ( .A1(n16253), .A2(DATAI_17_), .B1(P1_EAX_REG_17__SCAN_IN), 
        .B2(n16252), .ZN(n16251) );
  AOI22_X1 U18383 ( .A1(n16256), .A2(BUF1_REG_17__SCAN_IN), .B1(n16255), .B2(
        n16249), .ZN(n16250) );
  OAI211_X1 U18384 ( .C1(n20503), .C2(n16238), .A(n16251), .B(n16250), .ZN(
        P1_U2887) );
  AOI22_X1 U18385 ( .A1(n16253), .A2(DATAI_16_), .B1(P1_EAX_REG_16__SCAN_IN), 
        .B2(n16252), .ZN(n16258) );
  AOI22_X1 U18386 ( .A1(n16256), .A2(BUF1_REG_16__SCAN_IN), .B1(n16255), .B2(
        n16254), .ZN(n16257) );
  OAI211_X1 U18387 ( .C1(n16385), .C2(n16238), .A(n16258), .B(n16257), .ZN(
        P1_U2888) );
  AND2_X1 U18388 ( .A1(n16260), .A2(n16259), .ZN(n16261) );
  OR2_X1 U18389 ( .A1(n16261), .A2(n11196), .ZN(n20569) );
  OAI222_X1 U18390 ( .A1(n20569), .A2(n16238), .B1(n16265), .B2(n16263), .C1(
        n16268), .C2(n16262), .ZN(P1_U2889) );
  INV_X1 U18391 ( .A(n16264), .ZN(n16267) );
  OAI222_X1 U18392 ( .A1(n16238), .A2(n16410), .B1(n16268), .B2(n16267), .C1(
        n16266), .C2(n16265), .ZN(P1_U2891) );
  INV_X1 U18393 ( .A(n16269), .ZN(n16270) );
  XNOR2_X1 U18394 ( .A(n11452), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16279) );
  OAI211_X1 U18395 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16271), .A(
        n16270), .B(n16279), .ZN(n16272) );
  XNOR2_X1 U18396 ( .A(n16272), .B(n16448), .ZN(n16467) );
  NAND2_X1 U18397 ( .A1(n20584), .A2(n16273), .ZN(n16274) );
  NAND2_X1 U18398 ( .A1(n22052), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n16460) );
  OAI211_X1 U18399 ( .C1(n16405), .C2(n16275), .A(n16274), .B(n16460), .ZN(
        n16276) );
  AOI21_X1 U18400 ( .B1(n16277), .B2(n20555), .A(n16276), .ZN(n16278) );
  OAI21_X1 U18401 ( .B1(n16467), .B2(n22268), .A(n16278), .ZN(P1_U2969) );
  XNOR2_X1 U18402 ( .A(n16280), .B(n16279), .ZN(n16474) );
  NOR2_X1 U18403 ( .A1(n22049), .A2(n16281), .ZN(n16469) );
  AOI21_X1 U18404 ( .B1(n20588), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n16469), .ZN(n16282) );
  OAI21_X1 U18405 ( .B1(n20594), .B2(n16283), .A(n16282), .ZN(n16284) );
  AOI21_X1 U18406 ( .B1(n16285), .B2(n20555), .A(n16284), .ZN(n16286) );
  OAI21_X1 U18407 ( .B1(n22268), .B2(n16474), .A(n16286), .ZN(P1_U2970) );
  NAND2_X1 U18408 ( .A1(n16412), .A2(n16493), .ZN(n16307) );
  NAND2_X1 U18409 ( .A1(n16334), .A2(n16307), .ZN(n16290) );
  NAND3_X1 U18410 ( .A1(n16513), .A2(n13990), .A3(n16494), .ZN(n16288) );
  MUX2_X1 U18411 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n16494), .S(
        n11452), .Z(n16287) );
  AOI21_X1 U18412 ( .B1(n16290), .B2(n16288), .A(n16287), .ZN(n16289) );
  OAI21_X1 U18413 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n16290), .A(
        n16289), .ZN(n16292) );
  XNOR2_X1 U18414 ( .A(n16292), .B(n16291), .ZN(n16483) );
  INV_X1 U18415 ( .A(n16293), .ZN(n16298) );
  NOR2_X1 U18416 ( .A1(n22049), .A2(n16294), .ZN(n16479) );
  AOI21_X1 U18417 ( .B1(n20588), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16479), .ZN(n16295) );
  OAI21_X1 U18418 ( .B1(n20594), .B2(n16296), .A(n16295), .ZN(n16297) );
  AOI21_X1 U18419 ( .B1(n16298), .B2(n20555), .A(n16297), .ZN(n16299) );
  OAI21_X1 U18420 ( .B1(n22268), .B2(n16483), .A(n16299), .ZN(P1_U2971) );
  XNOR2_X1 U18421 ( .A(n11452), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16301) );
  XNOR2_X1 U18422 ( .A(n16300), .B(n16301), .ZN(n16491) );
  NOR2_X1 U18423 ( .A1(n22049), .A2(n20467), .ZN(n16484) );
  AOI21_X1 U18424 ( .B1(n20588), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16484), .ZN(n16302) );
  OAI21_X1 U18425 ( .B1(n20594), .B2(n16303), .A(n16302), .ZN(n16304) );
  AOI21_X1 U18426 ( .B1(n16305), .B2(n20555), .A(n16304), .ZN(n16306) );
  OAI21_X1 U18427 ( .B1(n16491), .B2(n22268), .A(n16306), .ZN(P1_U2972) );
  NAND3_X1 U18428 ( .A1(n16308), .A2(n11465), .A3(n16307), .ZN(n16309) );
  XNOR2_X1 U18429 ( .A(n16309), .B(n16494), .ZN(n16503) );
  NOR2_X1 U18430 ( .A1(n22049), .A2(n16310), .ZN(n16497) );
  AOI21_X1 U18431 ( .B1(n20588), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16497), .ZN(n16311) );
  OAI21_X1 U18432 ( .B1(n20594), .B2(n16312), .A(n16311), .ZN(n16313) );
  AOI21_X1 U18433 ( .B1(n16314), .B2(n20555), .A(n16313), .ZN(n16315) );
  OAI21_X1 U18434 ( .B1(n22268), .B2(n16503), .A(n16315), .ZN(P1_U2973) );
  AND2_X1 U18435 ( .A1(n16412), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16336) );
  OAI21_X1 U18436 ( .B1(n16513), .B2(n16336), .A(n11465), .ZN(n16316) );
  AOI21_X1 U18437 ( .B1(n16334), .B2(n16325), .A(n16316), .ZN(n16317) );
  XNOR2_X1 U18438 ( .A(n16317), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16512) );
  NOR2_X1 U18439 ( .A1(n22049), .A2(n20464), .ZN(n16506) );
  AOI21_X1 U18440 ( .B1(n20588), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16506), .ZN(n16318) );
  OAI21_X1 U18441 ( .B1(n20594), .B2(n16319), .A(n16318), .ZN(n16320) );
  AOI21_X1 U18442 ( .B1(n16321), .B2(n20555), .A(n16320), .ZN(n16322) );
  OAI21_X1 U18443 ( .B1(n22268), .B2(n16512), .A(n16322), .ZN(P1_U2974) );
  INV_X1 U18444 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16323) );
  NAND2_X1 U18445 ( .A1(n16352), .A2(n16323), .ZN(n16332) );
  NOR2_X1 U18446 ( .A1(n16334), .A2(n16332), .ZN(n16337) );
  AOI21_X1 U18447 ( .B1(n16324), .B2(n16336), .A(n16337), .ZN(n16326) );
  XNOR2_X1 U18448 ( .A(n16326), .B(n16325), .ZN(n16523) );
  INV_X1 U18449 ( .A(n22261), .ZN(n16329) );
  NOR2_X1 U18450 ( .A1(n22049), .A2(n16327), .ZN(n16517) );
  AOI21_X1 U18451 ( .B1(n20588), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16517), .ZN(n16328) );
  OAI21_X1 U18452 ( .B1(n20594), .B2(n16329), .A(n16328), .ZN(n16330) );
  AOI21_X1 U18453 ( .B1(n22263), .B2(n20555), .A(n16330), .ZN(n16331) );
  OAI21_X1 U18454 ( .B1(n16523), .B2(n22268), .A(n16331), .ZN(P1_U2975) );
  INV_X1 U18455 ( .A(n16332), .ZN(n16333) );
  NOR2_X1 U18456 ( .A1(n16333), .A2(n16336), .ZN(n16335) );
  MUX2_X1 U18457 ( .A(n16336), .B(n16335), .S(n16334), .Z(n16338) );
  NOR2_X1 U18458 ( .A1(n16338), .A2(n16337), .ZN(n16535) );
  INV_X1 U18459 ( .A(n22247), .ZN(n16341) );
  INV_X1 U18460 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n22241) );
  NOR2_X1 U18461 ( .A1(n22049), .A2(n22241), .ZN(n16528) );
  AOI21_X1 U18462 ( .B1(n20588), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16528), .ZN(n16339) );
  OAI21_X1 U18463 ( .B1(n20594), .B2(n22252), .A(n16339), .ZN(n16340) );
  AOI21_X1 U18464 ( .B1(n16341), .B2(n20555), .A(n16340), .ZN(n16342) );
  OAI21_X1 U18465 ( .B1(n16535), .B2(n22268), .A(n16342), .ZN(P1_U2976) );
  INV_X1 U18466 ( .A(n16343), .ZN(n16344) );
  OAI21_X1 U18467 ( .B1(n16345), .B2(n16412), .A(n16344), .ZN(n16346) );
  XNOR2_X1 U18468 ( .A(n16346), .B(n16432), .ZN(n16554) );
  INV_X1 U18469 ( .A(n22230), .ZN(n16350) );
  INV_X1 U18470 ( .A(n16347), .ZN(n22229) );
  NOR2_X1 U18471 ( .A1(n22049), .A2(n22225), .ZN(n16549) );
  AOI21_X1 U18472 ( .B1(n20588), .B2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16549), .ZN(n16348) );
  OAI21_X1 U18473 ( .B1(n20594), .B2(n22229), .A(n16348), .ZN(n16349) );
  AOI21_X1 U18474 ( .B1(n16350), .B2(n20555), .A(n16349), .ZN(n16351) );
  OAI21_X1 U18475 ( .B1(n22268), .B2(n16554), .A(n16351), .ZN(P1_U2977) );
  INV_X1 U18476 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n22045) );
  XNOR2_X1 U18477 ( .A(n11452), .B(n22022), .ZN(n16369) );
  OR2_X1 U18478 ( .A1(n13238), .A2(n16369), .ZN(n16354) );
  NAND2_X1 U18479 ( .A1(n16352), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16353) );
  NAND2_X1 U18480 ( .A1(n16354), .A2(n16353), .ZN(n20590) );
  MUX2_X1 U18481 ( .A(n22045), .B(n20590), .S(n16352), .Z(n16360) );
  INV_X1 U18482 ( .A(n20590), .ZN(n16361) );
  MUX2_X1 U18483 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n16361), .S(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .Z(n16355) );
  NOR2_X1 U18484 ( .A1(n16360), .A2(n16355), .ZN(n16356) );
  XNOR2_X1 U18485 ( .A(n16356), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16564) );
  INV_X1 U18486 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n22223) );
  NOR2_X1 U18487 ( .A1(n22049), .A2(n22223), .ZN(n16556) );
  AOI21_X1 U18488 ( .B1(n20588), .B2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n16556), .ZN(n16357) );
  OAI21_X1 U18489 ( .B1(n20594), .B2(n22219), .A(n16357), .ZN(n16358) );
  AOI21_X1 U18490 ( .B1(n22216), .B2(n20555), .A(n16358), .ZN(n16359) );
  OAI21_X1 U18491 ( .B1(n16564), .B2(n22268), .A(n16359), .ZN(P1_U2978) );
  AOI21_X1 U18492 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n16361), .A(
        n16360), .ZN(n16362) );
  XNOR2_X1 U18493 ( .A(n16362), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16576) );
  NAND2_X1 U18494 ( .A1(n20584), .A2(n16363), .ZN(n16364) );
  NAND2_X1 U18495 ( .A1(n22052), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n16566) );
  OAI211_X1 U18496 ( .C1(n16405), .C2(n16365), .A(n16364), .B(n16566), .ZN(
        n16366) );
  AOI21_X1 U18497 ( .B1(n16367), .B2(n20555), .A(n16366), .ZN(n16368) );
  OAI21_X1 U18498 ( .B1(n22268), .B2(n16576), .A(n16368), .ZN(P1_U2979) );
  XNOR2_X1 U18499 ( .A(n13238), .B(n16369), .ZN(n22020) );
  INV_X1 U18500 ( .A(n16370), .ZN(n22184) );
  AOI22_X1 U18501 ( .A1(n20588), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n22052), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n16371) );
  OAI21_X1 U18502 ( .B1(n22184), .B2(n20594), .A(n16371), .ZN(n16372) );
  AOI21_X1 U18503 ( .B1(n16373), .B2(n20555), .A(n16372), .ZN(n16374) );
  OAI21_X1 U18504 ( .B1(n22020), .B2(n22268), .A(n16374), .ZN(P1_U2981) );
  INV_X1 U18505 ( .A(n16376), .ZN(n16378) );
  AOI21_X1 U18506 ( .B1(n16375), .B2(n16378), .A(n16377), .ZN(n20568) );
  NAND2_X1 U18507 ( .A1(n16412), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16380) );
  NAND3_X1 U18508 ( .A1(n20568), .A2(n16352), .A3(n22015), .ZN(n16379) );
  OAI21_X1 U18509 ( .B1(n20568), .B2(n16380), .A(n16379), .ZN(n16381) );
  XNOR2_X1 U18510 ( .A(n16381), .B(n22034), .ZN(n22037) );
  NAND2_X1 U18511 ( .A1(n22037), .A2(n20591), .ZN(n16384) );
  OAI22_X1 U18512 ( .A1(n16405), .A2(n22172), .B1(n22049), .B2(n22176), .ZN(
        n16382) );
  AOI21_X1 U18513 ( .B1(n22174), .B2(n20584), .A(n16382), .ZN(n16383) );
  OAI211_X1 U18514 ( .C1(n16428), .C2(n16385), .A(n16384), .B(n16383), .ZN(
        P1_U2983) );
  OAI21_X1 U18515 ( .B1(n16375), .B2(n16387), .A(n16386), .ZN(n16389) );
  NAND2_X1 U18516 ( .A1(n16389), .A2(n16388), .ZN(n16391) );
  MUX2_X1 U18517 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n13959), .S(
        n16412), .Z(n16390) );
  XNOR2_X1 U18518 ( .A(n16391), .B(n16390), .ZN(n21903) );
  INV_X1 U18519 ( .A(n21903), .ZN(n16397) );
  AOI22_X1 U18520 ( .A1(n20588), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n22052), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n16392) );
  OAI21_X1 U18521 ( .B1(n20594), .B2(n16393), .A(n16392), .ZN(n16394) );
  AOI21_X1 U18522 ( .B1(n16395), .B2(n20555), .A(n16394), .ZN(n16396) );
  OAI21_X1 U18523 ( .B1(n16397), .B2(n22268), .A(n16396), .ZN(P1_U2985) );
  INV_X1 U18524 ( .A(n16398), .ZN(n16399) );
  AOI21_X1 U18525 ( .B1(n16375), .B2(n16400), .A(n16399), .ZN(n20558) );
  OAI211_X1 U18526 ( .C1(n11452), .C2(n16401), .A(n20558), .B(n20560), .ZN(
        n20561) );
  NAND2_X1 U18527 ( .A1(n20561), .A2(n20560), .ZN(n16402) );
  XOR2_X1 U18528 ( .A(n16403), .B(n16402), .Z(n21894) );
  NAND2_X1 U18529 ( .A1(n21894), .A2(n20591), .ZN(n16409) );
  OAI22_X1 U18530 ( .A1(n16405), .A2(n16404), .B1(n22049), .B2(n17656), .ZN(
        n16406) );
  AOI21_X1 U18531 ( .B1(n20584), .B2(n16407), .A(n16406), .ZN(n16408) );
  OAI211_X1 U18532 ( .C1(n16428), .C2(n16410), .A(n16409), .B(n16408), .ZN(
        P1_U2986) );
  NOR2_X1 U18533 ( .A1(n16375), .A2(n16412), .ZN(n16413) );
  MUX2_X1 U18534 ( .A(n16411), .B(n16375), .S(n20578), .Z(n16421) );
  NOR2_X1 U18535 ( .A1(n16421), .A2(n21993), .ZN(n16420) );
  MUX2_X1 U18536 ( .A(n16413), .B(n16412), .S(n16420), .Z(n16415) );
  XNOR2_X1 U18537 ( .A(n16415), .B(n16414), .ZN(n16585) );
  INV_X1 U18538 ( .A(n16585), .ZN(n16419) );
  OR2_X1 U18539 ( .A1(n22049), .A2(n22153), .ZN(n16582) );
  NAND2_X1 U18540 ( .A1(n20588), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16416) );
  OAI211_X1 U18541 ( .C1(n20594), .C2(n22147), .A(n16582), .B(n16416), .ZN(
        n16417) );
  AOI21_X1 U18542 ( .B1(n22144), .B2(n20555), .A(n16417), .ZN(n16418) );
  OAI21_X1 U18543 ( .B1(n16419), .B2(n22268), .A(n16418), .ZN(P1_U2988) );
  AOI21_X1 U18544 ( .B1(n21993), .B2(n16421), .A(n16420), .ZN(n21988) );
  NAND2_X1 U18545 ( .A1(n21988), .A2(n20591), .ZN(n16426) );
  NOR2_X1 U18546 ( .A1(n22049), .A2(n16422), .ZN(n21987) );
  NOR2_X1 U18547 ( .A1(n20594), .A2(n16423), .ZN(n16424) );
  AOI211_X1 U18548 ( .C1(n20588), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n21987), .B(n16424), .ZN(n16425) );
  OAI211_X1 U18549 ( .C1(n16428), .C2(n16427), .A(n16426), .B(n16425), .ZN(
        P1_U2989) );
  NOR2_X1 U18550 ( .A1(n16429), .A2(n22033), .ZN(n16454) );
  NAND2_X1 U18551 ( .A1(n21908), .A2(n21892), .ZN(n22050) );
  NAND2_X1 U18552 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n22011) );
  INV_X1 U18553 ( .A(n22011), .ZN(n16430) );
  AND2_X1 U18554 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16430), .ZN(
        n16431) );
  AND2_X1 U18555 ( .A1(n22023), .A2(n16431), .ZN(n16538) );
  NAND2_X1 U18556 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21980) );
  NOR2_X1 U18557 ( .A1(n21930), .A2(n21937), .ZN(n21942) );
  NAND2_X1 U18558 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n21942), .ZN(
        n21945) );
  NAND2_X1 U18559 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21923) );
  NOR4_X1 U18560 ( .A1(n21949), .A2(n21980), .A3(n21945), .A4(n21923), .ZN(
        n21974) );
  NAND3_X1 U18561 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n21974), .ZN(n16580) );
  NOR3_X1 U18562 ( .A1(n16414), .A2(n16401), .A3(n16580), .ZN(n21887) );
  NAND2_X1 U18563 ( .A1(n16538), .A2(n21887), .ZN(n16438) );
  NOR2_X1 U18564 ( .A1(n22012), .A2(n16438), .ZN(n16540) );
  NOR2_X1 U18565 ( .A1(n16547), .A2(n16432), .ZN(n16441) );
  NAND2_X1 U18566 ( .A1(n16540), .A2(n16441), .ZN(n16437) );
  NAND2_X1 U18567 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n21989) );
  INV_X1 U18568 ( .A(n21945), .ZN(n16434) );
  OAI21_X1 U18569 ( .B1(n21908), .B2(n22064), .A(n16433), .ZN(n21924) );
  NAND2_X1 U18570 ( .A1(n16434), .A2(n21924), .ZN(n21940) );
  OR2_X1 U18571 ( .A1(n21949), .A2(n21940), .ZN(n21958) );
  OR2_X1 U18572 ( .A1(n21980), .A2(n21958), .ZN(n21976) );
  NOR2_X1 U18573 ( .A1(n21989), .A2(n21976), .ZN(n16579) );
  NAND2_X1 U18574 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16579), .ZN(
        n16577) );
  NOR2_X1 U18575 ( .A1(n16401), .A2(n16577), .ZN(n21886) );
  NAND2_X1 U18576 ( .A1(n16538), .A2(n21886), .ZN(n16542) );
  INV_X1 U18577 ( .A(n16542), .ZN(n16435) );
  AND2_X1 U18578 ( .A1(n16441), .A2(n16435), .ZN(n16443) );
  NAND2_X1 U18579 ( .A1(n22007), .A2(n16443), .ZN(n16436) );
  NOR3_X1 U18580 ( .A1(n16531), .A2(n16494), .A3(n16493), .ZN(n16477) );
  NAND3_X1 U18581 ( .A1(n16477), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n16458), .ZN(n16463) );
  NOR3_X1 U18582 ( .A1(n16463), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n16448), .ZN(n16453) );
  NAND2_X1 U18583 ( .A1(n21909), .A2(n16438), .ZN(n16440) );
  NAND2_X1 U18584 ( .A1(n16536), .A2(n21908), .ZN(n16439) );
  NAND2_X1 U18585 ( .A1(n16440), .A2(n22002), .ZN(n16544) );
  NOR2_X1 U18586 ( .A1(n22004), .A2(n16441), .ZN(n16442) );
  OR2_X1 U18587 ( .A1(n16544), .A2(n16442), .ZN(n16446) );
  INV_X1 U18588 ( .A(n16443), .ZN(n16444) );
  AND2_X1 U18589 ( .A1(n22007), .A2(n16444), .ZN(n16445) );
  NOR2_X1 U18590 ( .A1(n16446), .A2(n16445), .ZN(n16516) );
  INV_X1 U18591 ( .A(n22019), .ZN(n22051) );
  NAND2_X1 U18592 ( .A1(n22051), .A2(n16493), .ZN(n16447) );
  AND2_X1 U18593 ( .A1(n16516), .A2(n16447), .ZN(n16496) );
  AOI21_X1 U18594 ( .B1(n16496), .B2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n16545), .ZN(n16485) );
  NOR2_X1 U18595 ( .A1(n16485), .A2(n16448), .ZN(n16462) );
  NOR2_X1 U18596 ( .A1(n22019), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16459) );
  INV_X1 U18597 ( .A(n16458), .ZN(n16475) );
  NOR2_X1 U18598 ( .A1(n16459), .A2(n16475), .ZN(n16450) );
  AOI211_X1 U18599 ( .C1(n16462), .C2(n16450), .A(n16545), .B(n16449), .ZN(
        n16451) );
  OAI21_X1 U18600 ( .B1(n16456), .B2(n22031), .A(n16455), .ZN(P1_U3000) );
  INV_X1 U18601 ( .A(n16485), .ZN(n16457) );
  OAI21_X1 U18602 ( .B1(n16458), .B2(n16545), .A(n16457), .ZN(n16470) );
  OAI21_X1 U18603 ( .B1(n16470), .B2(n16459), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16461) );
  OAI211_X1 U18604 ( .C1(n16463), .C2(n16462), .A(n16461), .B(n16460), .ZN(
        n16464) );
  AOI21_X1 U18605 ( .B1(n16465), .B2(n22056), .A(n16464), .ZN(n16466) );
  OAI21_X1 U18606 ( .B1(n16467), .B2(n22031), .A(n16466), .ZN(P1_U3001) );
  INV_X1 U18607 ( .A(n16477), .ZN(n16487) );
  NOR3_X1 U18608 ( .A1(n16487), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n16475), .ZN(n16468) );
  AOI211_X1 U18609 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16470), .A(
        n16469), .B(n16468), .ZN(n16473) );
  NAND2_X1 U18610 ( .A1(n16471), .A2(n22056), .ZN(n16472) );
  OAI211_X1 U18611 ( .C1(n16474), .C2(n22031), .A(n16473), .B(n16472), .ZN(
        P1_U3002) );
  AND3_X1 U18612 ( .A1(n16477), .A2(n16476), .A3(n16475), .ZN(n16478) );
  AOI211_X1 U18613 ( .C1(n16485), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16479), .B(n16478), .ZN(n16482) );
  NAND2_X1 U18614 ( .A1(n16480), .A2(n22056), .ZN(n16481) );
  OAI211_X1 U18615 ( .C1(n16483), .C2(n22031), .A(n16482), .B(n16481), .ZN(
        P1_U3003) );
  AOI21_X1 U18616 ( .B1(n16485), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n16484), .ZN(n16486) );
  OAI21_X1 U18617 ( .B1(n16487), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n16486), .ZN(n16488) );
  AOI21_X1 U18618 ( .B1(n16489), .B2(n22056), .A(n16488), .ZN(n16490) );
  OAI21_X1 U18619 ( .B1(n16491), .B2(n22031), .A(n16490), .ZN(P1_U3004) );
  INV_X1 U18620 ( .A(n16492), .ZN(n16501) );
  INV_X1 U18621 ( .A(n16493), .ZN(n16495) );
  NAND2_X1 U18622 ( .A1(n16495), .A2(n16494), .ZN(n16499) );
  INV_X1 U18623 ( .A(n16496), .ZN(n16507) );
  AOI21_X1 U18624 ( .B1(n16507), .B2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n16497), .ZN(n16498) );
  OAI21_X1 U18625 ( .B1(n16531), .B2(n16499), .A(n16498), .ZN(n16500) );
  AOI21_X1 U18626 ( .B1(n16501), .B2(n22056), .A(n16500), .ZN(n16502) );
  OAI21_X1 U18627 ( .B1(n16503), .B2(n22031), .A(n16502), .ZN(P1_U3005) );
  INV_X1 U18628 ( .A(n16504), .ZN(n16514) );
  NOR3_X1 U18629 ( .A1(n16531), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n16514), .ZN(n16505) );
  AOI211_X1 U18630 ( .C1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n16507), .A(
        n16506), .B(n16505), .ZN(n16511) );
  INV_X1 U18631 ( .A(n16508), .ZN(n16509) );
  NAND2_X1 U18632 ( .A1(n16509), .A2(n22056), .ZN(n16510) );
  OAI211_X1 U18633 ( .C1(n16512), .C2(n22031), .A(n16511), .B(n16510), .ZN(
        P1_U3006) );
  INV_X1 U18634 ( .A(n22266), .ZN(n16521) );
  INV_X1 U18635 ( .A(n16513), .ZN(n16515) );
  NAND2_X1 U18636 ( .A1(n16515), .A2(n16514), .ZN(n16519) );
  INV_X1 U18637 ( .A(n16516), .ZN(n16529) );
  AOI21_X1 U18638 ( .B1(n16529), .B2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n16517), .ZN(n16518) );
  OAI21_X1 U18639 ( .B1(n16531), .B2(n16519), .A(n16518), .ZN(n16520) );
  AOI21_X1 U18640 ( .B1(n16521), .B2(n22056), .A(n16520), .ZN(n16522) );
  OAI21_X1 U18641 ( .B1(n16523), .B2(n22031), .A(n16522), .ZN(P1_U3007) );
  NAND2_X1 U18642 ( .A1(n16525), .A2(n16524), .ZN(n16526) );
  NAND2_X1 U18643 ( .A1(n16527), .A2(n16526), .ZN(n22245) );
  INV_X1 U18644 ( .A(n22245), .ZN(n16533) );
  AOI21_X1 U18645 ( .B1(n16529), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16528), .ZN(n16530) );
  OAI21_X1 U18646 ( .B1(n16531), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16530), .ZN(n16532) );
  AOI21_X1 U18647 ( .B1(n16533), .B2(n22056), .A(n16532), .ZN(n16534) );
  OAI21_X1 U18648 ( .B1(n16535), .B2(n22031), .A(n16534), .ZN(P1_U3008) );
  INV_X1 U18649 ( .A(n21887), .ZN(n22014) );
  NOR2_X1 U18650 ( .A1(n21908), .A2(n22014), .ZN(n21889) );
  NAND2_X1 U18651 ( .A1(n16536), .A2(n21889), .ZN(n16537) );
  NAND2_X1 U18652 ( .A1(n22007), .A2(n21886), .ZN(n22013) );
  INV_X1 U18653 ( .A(n16538), .ZN(n16539) );
  NOR2_X1 U18654 ( .A1(n21899), .A2(n16539), .ZN(n16568) );
  NOR2_X1 U18655 ( .A1(n16540), .A2(n16568), .ZN(n22043) );
  INV_X1 U18656 ( .A(n16546), .ZN(n16541) );
  NOR3_X1 U18657 ( .A1(n22043), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n16541), .ZN(n16555) );
  AND2_X1 U18658 ( .A1(n22007), .A2(n16542), .ZN(n16543) );
  NOR2_X1 U18659 ( .A1(n16544), .A2(n16543), .ZN(n22044) );
  AOI21_X1 U18660 ( .B1(n22044), .B2(n16546), .A(n16545), .ZN(n16557) );
  OR2_X1 U18661 ( .A1(n16555), .A2(n16557), .ZN(n16550) );
  NOR3_X1 U18662 ( .A1(n22043), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n16547), .ZN(n16548) );
  AOI211_X1 U18663 ( .C1(n16550), .C2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n16549), .B(n16548), .ZN(n16553) );
  INV_X1 U18664 ( .A(n22234), .ZN(n16551) );
  NAND2_X1 U18665 ( .A1(n16551), .A2(n22056), .ZN(n16552) );
  OAI211_X1 U18666 ( .C1(n16554), .C2(n22031), .A(n16553), .B(n16552), .ZN(
        P1_U3009) );
  AOI211_X1 U18667 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n16557), .A(
        n16556), .B(n16555), .ZN(n16563) );
  NOR2_X1 U18668 ( .A1(n16115), .A2(n16558), .ZN(n16559) );
  OR2_X1 U18669 ( .A1(n16560), .A2(n16559), .ZN(n22214) );
  INV_X1 U18670 ( .A(n22214), .ZN(n16561) );
  NAND2_X1 U18671 ( .A1(n16561), .A2(n22056), .ZN(n16562) );
  OAI211_X1 U18672 ( .C1(n16564), .C2(n22031), .A(n16563), .B(n16562), .ZN(
        P1_U3010) );
  NOR2_X1 U18673 ( .A1(n16565), .A2(n22033), .ZN(n16574) );
  NOR3_X1 U18674 ( .A1(n22043), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n22045), .ZN(n16573) );
  INV_X1 U18675 ( .A(n16566), .ZN(n16572) );
  INV_X1 U18676 ( .A(n21892), .ZN(n16567) );
  OAI21_X1 U18677 ( .B1(n16568), .B2(n16567), .A(n22045), .ZN(n16570) );
  AOI21_X1 U18678 ( .B1(n16570), .B2(n22044), .A(n16569), .ZN(n16571) );
  NOR4_X1 U18679 ( .A1(n16574), .A2(n16573), .A3(n16572), .A4(n16571), .ZN(
        n16575) );
  OAI21_X1 U18680 ( .B1(n16576), .B2(n22031), .A(n16575), .ZN(P1_U3011) );
  AOI22_X1 U18681 ( .A1(n22007), .A2(n16577), .B1(n21909), .B2(n16580), .ZN(
        n16578) );
  NAND2_X1 U18682 ( .A1(n22002), .A2(n16578), .ZN(n21997) );
  INV_X1 U18683 ( .A(n16579), .ZN(n16581) );
  OAI22_X1 U18684 ( .A1(n21907), .A2(n16581), .B1(n16580), .B2(n22012), .ZN(
        n21999) );
  AOI22_X1 U18685 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n21997), .B1(
        n21999), .B2(n16414), .ZN(n16583) );
  OAI211_X1 U18686 ( .C1(n22033), .C2(n22142), .A(n16583), .B(n16582), .ZN(
        n16584) );
  AOI21_X1 U18687 ( .B1(n16585), .B2(n22053), .A(n16584), .ZN(n16586) );
  INV_X1 U18688 ( .A(n16586), .ZN(P1_U3020) );
  INV_X1 U18689 ( .A(n16587), .ZN(n16588) );
  NOR2_X1 U18690 ( .A1(n16588), .A2(n22273), .ZN(n22281) );
  AOI21_X1 U18691 ( .B1(n13341), .B2(n16589), .A(n22281), .ZN(n16590) );
  OAI21_X1 U18692 ( .B1(n13338), .B2(n22424), .A(n16590), .ZN(n16591) );
  MUX2_X1 U18693 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n16591), .S(
        n17826), .Z(P1_U3478) );
  NOR3_X1 U18694 ( .A1(n16592), .A2(n14961), .A3(n14872), .ZN(n16594) );
  NOR2_X1 U18695 ( .A1(n14969), .A2(n16607), .ZN(n16593) );
  AOI211_X1 U18696 ( .C1(n16613), .C2(n16595), .A(n16594), .B(n16593), .ZN(
        n17789) );
  INV_X1 U18697 ( .A(n16596), .ZN(n16625) );
  NOR3_X1 U18698 ( .A1(n14961), .A2(n14872), .A3(n16623), .ZN(n16597) );
  AOI21_X1 U18699 ( .B1(n16599), .B2(n16598), .A(n16597), .ZN(n16600) );
  OAI21_X1 U18700 ( .B1(n17789), .B2(n16625), .A(n16600), .ZN(n16602) );
  MUX2_X1 U18701 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n16602), .S(
        n16601), .Z(P1_U3473) );
  INV_X1 U18702 ( .A(n14872), .ZN(n16609) );
  NAND2_X1 U18703 ( .A1(n16609), .A2(n16603), .ZN(n16618) );
  NOR2_X1 U18704 ( .A1(n14872), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n16604) );
  NOR2_X1 U18705 ( .A1(n16604), .A2(n12841), .ZN(n16606) );
  AND2_X1 U18706 ( .A1(n16606), .A2(n11167), .ZN(n16622) );
  NAND3_X1 U18707 ( .A1(n16607), .A2(n12975), .A3(n16622), .ZN(n16617) );
  NAND2_X1 U18708 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16608) );
  NAND2_X1 U18709 ( .A1(n16613), .A2(n16608), .ZN(n16615) );
  INV_X1 U18710 ( .A(n16608), .ZN(n16612) );
  NAND2_X1 U18711 ( .A1(n16609), .A2(n12838), .ZN(n16610) );
  AOI22_X1 U18712 ( .A1(n16613), .A2(n16612), .B1(n16611), .B2(n16610), .ZN(
        n16614) );
  MUX2_X1 U18713 ( .A(n16615), .B(n16614), .S(n12839), .Z(n16616) );
  NAND3_X1 U18714 ( .A1(n16618), .A2(n16617), .A3(n16616), .ZN(n16619) );
  AOI21_X1 U18715 ( .B1(n16621), .B2(n16620), .A(n16619), .ZN(n17786) );
  INV_X1 U18716 ( .A(n16622), .ZN(n16624) );
  OAI22_X1 U18717 ( .A1(n17786), .A2(n16625), .B1(n16624), .B2(n16623), .ZN(
        n16627) );
  MUX2_X1 U18718 ( .A(n16627), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n16626), .Z(P1_U3469) );
  NAND2_X1 U18719 ( .A1(n22557), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n16632) );
  AOI22_X1 U18720 ( .A1(n16628), .A2(n22551), .B1(n22433), .B2(n22553), .ZN(
        n16631) );
  NAND2_X1 U18721 ( .A1(n22556), .A2(n22442), .ZN(n16630) );
  NAND2_X1 U18722 ( .A1(n16653), .A2(n22434), .ZN(n16629) );
  NAND4_X1 U18723 ( .A1(n16632), .A2(n16631), .A3(n16630), .A4(n16629), .ZN(
        P1_U3145) );
  NAND2_X1 U18724 ( .A1(n22557), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n16637) );
  AOI22_X1 U18725 ( .A1(n16633), .A2(n22551), .B1(n22464), .B2(n22553), .ZN(
        n16636) );
  NAND2_X1 U18726 ( .A1(n22556), .A2(n22466), .ZN(n16635) );
  NAND2_X1 U18727 ( .A1(n16653), .A2(n22465), .ZN(n16634) );
  NAND4_X1 U18728 ( .A1(n16637), .A2(n16636), .A3(n16635), .A4(n16634), .ZN(
        P1_U3146) );
  NAND2_X1 U18729 ( .A1(n22557), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n16642) );
  AOI22_X1 U18730 ( .A1(n16638), .A2(n22551), .B1(n22487), .B2(n22553), .ZN(
        n16641) );
  NAND2_X1 U18731 ( .A1(n22556), .A2(n22489), .ZN(n16640) );
  NAND2_X1 U18732 ( .A1(n16653), .A2(n22488), .ZN(n16639) );
  NAND4_X1 U18733 ( .A1(n16642), .A2(n16641), .A3(n16640), .A4(n16639), .ZN(
        P1_U3147) );
  NAND2_X1 U18734 ( .A1(n22557), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n16647) );
  AOI22_X1 U18735 ( .A1(n16643), .A2(n22551), .B1(n22511), .B2(n22553), .ZN(
        n16646) );
  NAND2_X1 U18736 ( .A1(n22556), .A2(n22513), .ZN(n16645) );
  NAND2_X1 U18737 ( .A1(n16653), .A2(n22512), .ZN(n16644) );
  NAND4_X1 U18738 ( .A1(n16647), .A2(n16646), .A3(n16645), .A4(n16644), .ZN(
        P1_U3148) );
  NAND2_X1 U18739 ( .A1(n22557), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n16652) );
  AOI22_X1 U18740 ( .A1(n16648), .A2(n22551), .B1(n22608), .B2(n22553), .ZN(
        n16651) );
  NAND2_X1 U18741 ( .A1(n22556), .A2(n22610), .ZN(n16650) );
  NAND2_X1 U18742 ( .A1(n16653), .A2(n22609), .ZN(n16649) );
  NAND4_X1 U18743 ( .A1(n16652), .A2(n16651), .A3(n16650), .A4(n16649), .ZN(
        P1_U3151) );
  NAND2_X1 U18744 ( .A1(n22557), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n16657) );
  AOI22_X1 U18745 ( .A1(n22674), .A2(n22551), .B1(n22671), .B2(n22553), .ZN(
        n16656) );
  NAND2_X1 U18746 ( .A1(n22556), .A2(n22662), .ZN(n16655) );
  NAND2_X1 U18747 ( .A1(n16653), .A2(n22675), .ZN(n16654) );
  NAND4_X1 U18748 ( .A1(n16657), .A2(n16656), .A3(n16655), .A4(n16654), .ZN(
        P1_U3152) );
  INV_X1 U18749 ( .A(n16658), .ZN(n16674) );
  OAI211_X1 U18750 ( .C1(n16661), .C2(n16660), .A(n19127), .B(n16659), .ZN(
        n16673) );
  INV_X1 U18751 ( .A(n17052), .ZN(n16671) );
  INV_X1 U18752 ( .A(n16662), .ZN(n16666) );
  INV_X1 U18753 ( .A(n16663), .ZN(n16759) );
  NAND2_X1 U18754 ( .A1(n16759), .A2(n16664), .ZN(n16665) );
  NOR2_X1 U18755 ( .A1(n17050), .A2(n19133), .ZN(n16670) );
  INV_X1 U18756 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16668) );
  AOI22_X1 U18757 ( .A1(P2_EBX_REG_28__SCAN_IN), .A2(n19135), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n19134), .ZN(n16667) );
  OAI21_X1 U18758 ( .B1(n19121), .B2(n16668), .A(n16667), .ZN(n16669) );
  AOI211_X1 U18759 ( .C1(n16671), .C2(n19160), .A(n16670), .B(n16669), .ZN(
        n16672) );
  OAI211_X1 U18760 ( .C1(n19149), .C2(n16674), .A(n16673), .B(n16672), .ZN(
        P2_U2827) );
  MUX2_X1 U18761 ( .A(P2_EBX_REG_31__SCAN_IN), .B(n19161), .S(n16727), .Z(
        P2_U2856) );
  XNOR2_X1 U18762 ( .A(n16676), .B(n16675), .ZN(n16677) );
  XNOR2_X1 U18763 ( .A(n16678), .B(n16677), .ZN(n16750) );
  NAND2_X1 U18764 ( .A1(n11141), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n16682) );
  AOI21_X1 U18765 ( .B1(n16680), .B2(n12699), .A(n16679), .ZN(n19140) );
  NAND2_X1 U18766 ( .A1(n19140), .A2(n16727), .ZN(n16681) );
  OAI211_X1 U18767 ( .C1(n16750), .C2(n16740), .A(n16682), .B(n16681), .ZN(
        P2_U2858) );
  INV_X1 U18768 ( .A(n16683), .ZN(n16690) );
  NAND2_X1 U18769 ( .A1(n16690), .A2(n16684), .ZN(n16686) );
  XNOR2_X1 U18770 ( .A(n16686), .B(n16685), .ZN(n16755) );
  NOR2_X1 U18771 ( .A1(n17052), .A2(n11141), .ZN(n16687) );
  AOI21_X1 U18772 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n11141), .A(n16687), .ZN(
        n16688) );
  OAI21_X1 U18773 ( .B1(n16755), .B2(n16740), .A(n16688), .ZN(P2_U2859) );
  NAND2_X1 U18774 ( .A1(n16690), .A2(n16689), .ZN(n16691) );
  XOR2_X1 U18775 ( .A(n16692), .B(n16691), .Z(n16765) );
  INV_X1 U18776 ( .A(n12352), .ZN(n16693) );
  OAI21_X1 U18777 ( .B1(n12770), .B2(n16694), .A(n16693), .ZN(n19118) );
  NOR2_X1 U18778 ( .A1(n19118), .A2(n11141), .ZN(n16695) );
  AOI21_X1 U18779 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n11141), .A(n16695), .ZN(
        n16696) );
  OAI21_X1 U18780 ( .B1(n16765), .B2(n16740), .A(n16696), .ZN(P2_U2860) );
  INV_X1 U18781 ( .A(n19110), .ZN(n16702) );
  AOI21_X1 U18782 ( .B1(n16699), .B2(n16698), .A(n16697), .ZN(n16766) );
  NAND2_X1 U18783 ( .A1(n16766), .A2(n16732), .ZN(n16701) );
  NAND2_X1 U18784 ( .A1(n11141), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n16700) );
  OAI211_X1 U18785 ( .C1(n16702), .C2(n11141), .A(n16701), .B(n16700), .ZN(
        P2_U2861) );
  OAI21_X1 U18786 ( .B1(n16703), .B2(n16705), .A(n16704), .ZN(n16785) );
  NAND2_X1 U18787 ( .A1(n11238), .A2(n16706), .ZN(n16707) );
  NAND2_X1 U18788 ( .A1(n11515), .A2(n16707), .ZN(n19099) );
  NOR2_X1 U18789 ( .A1(n19099), .A2(n11141), .ZN(n16708) );
  AOI21_X1 U18790 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n11141), .A(n16708), .ZN(
        n16709) );
  OAI21_X1 U18791 ( .B1(n16785), .B2(n16740), .A(n16709), .ZN(P2_U2862) );
  OAI21_X1 U18792 ( .B1(n16712), .B2(n16711), .A(n16710), .ZN(n16793) );
  OR2_X1 U18793 ( .A1(n16719), .A2(n16713), .ZN(n16714) );
  NAND2_X1 U18794 ( .A1(n11238), .A2(n16714), .ZN(n19087) );
  NOR2_X1 U18795 ( .A1(n19087), .A2(n11141), .ZN(n16715) );
  AOI21_X1 U18796 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n11141), .A(n16715), .ZN(
        n16716) );
  OAI21_X1 U18797 ( .B1(n16793), .B2(n16740), .A(n16716), .ZN(P2_U2863) );
  XNOR2_X1 U18798 ( .A(n16717), .B(n16718), .ZN(n16804) );
  NAND2_X1 U18799 ( .A1(n11141), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n16722) );
  AOI21_X1 U18800 ( .B1(n16720), .B2(n16726), .A(n16719), .ZN(n19073) );
  NAND2_X1 U18801 ( .A1(n19073), .A2(n16727), .ZN(n16721) );
  OAI211_X1 U18802 ( .C1(n16804), .C2(n16740), .A(n16722), .B(n16721), .ZN(
        P2_U2864) );
  OAI21_X1 U18803 ( .B1(n11191), .B2(n16723), .A(n16717), .ZN(n19962) );
  NAND2_X1 U18804 ( .A1(n11141), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n16729) );
  NAND2_X1 U18805 ( .A1(n12331), .A2(n16724), .ZN(n16725) );
  NAND2_X1 U18806 ( .A1(n19065), .A2(n16727), .ZN(n16728) );
  OAI211_X1 U18807 ( .C1(n19962), .C2(n16740), .A(n16729), .B(n16728), .ZN(
        P2_U2865) );
  AOI21_X1 U18808 ( .B1(n16731), .B2(n16730), .A(n11191), .ZN(n16805) );
  NAND2_X1 U18809 ( .A1(n16805), .A2(n16732), .ZN(n16734) );
  NAND2_X1 U18810 ( .A1(n11141), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n16733) );
  OAI211_X1 U18811 ( .C1(n19054), .C2(n11141), .A(n16734), .B(n16733), .ZN(
        P2_U2866) );
  OAI21_X1 U18812 ( .B1(n15910), .B2(n16735), .A(n16730), .ZN(n20065) );
  OAI21_X1 U18813 ( .B1(n16737), .B2(n16736), .A(n12813), .ZN(n19042) );
  NOR2_X1 U18814 ( .A1(n19042), .A2(n11141), .ZN(n16738) );
  AOI21_X1 U18815 ( .B1(P2_EBX_REG_20__SCAN_IN), .B2(n11141), .A(n16738), .ZN(
        n16739) );
  OAI21_X1 U18816 ( .B1(n20065), .B2(n16740), .A(n16739), .ZN(P2_U2867) );
  NOR2_X1 U18817 ( .A1(n16819), .A2(n16741), .ZN(n16747) );
  INV_X1 U18818 ( .A(n16742), .ZN(n16743) );
  OAI21_X1 U18819 ( .B1(n16662), .B2(n16744), .A(n16743), .ZN(n19138) );
  OAI22_X1 U18820 ( .A1(n19138), .A2(n16818), .B1(n16817), .B2(n16745), .ZN(
        n16746) );
  AOI211_X1 U18821 ( .C1(BUF1_REG_29__SCAN_IN), .C2(n20064), .A(n16747), .B(
        n16746), .ZN(n16749) );
  NAND2_X1 U18822 ( .A1(n20063), .A2(BUF2_REG_29__SCAN_IN), .ZN(n16748) );
  OAI211_X1 U18823 ( .C1(n16750), .C2(n20012), .A(n16749), .B(n16748), .ZN(
        P2_U2890) );
  AOI22_X1 U18824 ( .A1(n20062), .A2(n19745), .B1(P2_EAX_REG_28__SCAN_IN), 
        .B2(n20060), .ZN(n16752) );
  NAND2_X1 U18825 ( .A1(n20063), .A2(BUF2_REG_28__SCAN_IN), .ZN(n16751) );
  OAI211_X1 U18826 ( .C1(n17050), .C2(n16818), .A(n16752), .B(n16751), .ZN(
        n16753) );
  AOI21_X1 U18827 ( .B1(n20064), .B2(BUF1_REG_28__SCAN_IN), .A(n16753), .ZN(
        n16754) );
  OAI21_X1 U18828 ( .B1(n16755), .B2(n20012), .A(n16754), .ZN(P2_U2891) );
  AND2_X1 U18829 ( .A1(n20062), .A2(n16756), .ZN(n16762) );
  NAND2_X1 U18830 ( .A1(n11198), .A2(n16757), .ZN(n16758) );
  NAND2_X1 U18831 ( .A1(n16759), .A2(n16758), .ZN(n19132) );
  OAI22_X1 U18832 ( .A1(n19132), .A2(n16818), .B1(n16817), .B2(n16760), .ZN(
        n16761) );
  AOI211_X1 U18833 ( .C1(BUF1_REG_27__SCAN_IN), .C2(n20064), .A(n16762), .B(
        n16761), .ZN(n16764) );
  NAND2_X1 U18834 ( .A1(n20063), .A2(BUF2_REG_27__SCAN_IN), .ZN(n16763) );
  OAI211_X1 U18835 ( .C1(n16765), .C2(n20012), .A(n16764), .B(n16763), .ZN(
        P2_U2892) );
  INV_X1 U18836 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n16774) );
  NAND2_X1 U18837 ( .A1(n16766), .A2(n20068), .ZN(n16773) );
  OR2_X1 U18838 ( .A1(n16776), .A2(n16767), .ZN(n16768) );
  NAND2_X1 U18839 ( .A1(n11198), .A2(n16768), .ZN(n17071) );
  INV_X1 U18840 ( .A(n17071), .ZN(n19109) );
  AOI22_X1 U18841 ( .A1(n19109), .A2(n20067), .B1(P2_EAX_REG_26__SCAN_IN), 
        .B2(n20060), .ZN(n16769) );
  OAI21_X1 U18842 ( .B1(n16770), .B2(n16819), .A(n16769), .ZN(n16771) );
  AOI21_X1 U18843 ( .B1(n20064), .B2(BUF1_REG_26__SCAN_IN), .A(n16771), .ZN(
        n16772) );
  OAI211_X1 U18844 ( .C1(n16824), .C2(n16774), .A(n16773), .B(n16772), .ZN(
        P2_U2893) );
  NOR2_X1 U18845 ( .A1(n16819), .A2(n16775), .ZN(n16782) );
  INV_X1 U18846 ( .A(n16776), .ZN(n16779) );
  NAND2_X1 U18847 ( .A1(n11245), .A2(n16777), .ZN(n16778) );
  NAND2_X1 U18848 ( .A1(n16779), .A2(n16778), .ZN(n19097) );
  OAI22_X1 U18849 ( .A1(n19097), .A2(n16818), .B1(n16817), .B2(n16780), .ZN(
        n16781) );
  AOI211_X1 U18850 ( .C1(BUF1_REG_25__SCAN_IN), .C2(n20064), .A(n16782), .B(
        n16781), .ZN(n16784) );
  NAND2_X1 U18851 ( .A1(n20063), .A2(BUF2_REG_25__SCAN_IN), .ZN(n16783) );
  OAI211_X1 U18852 ( .C1(n16785), .C2(n20012), .A(n16784), .B(n16783), .ZN(
        P2_U2894) );
  XNOR2_X1 U18853 ( .A(n16796), .B(n11559), .ZN(n17091) );
  INV_X1 U18854 ( .A(n17091), .ZN(n19086) );
  OAI22_X1 U18855 ( .A1(n19086), .A2(n16818), .B1(n16817), .B2(n16787), .ZN(
        n16790) );
  NOR2_X1 U18856 ( .A1(n16819), .A2(n16788), .ZN(n16789) );
  AOI211_X1 U18857 ( .C1(BUF1_REG_24__SCAN_IN), .C2(n20064), .A(n16790), .B(
        n16789), .ZN(n16792) );
  NAND2_X1 U18858 ( .A1(n20063), .A2(BUF2_REG_24__SCAN_IN), .ZN(n16791) );
  OAI211_X1 U18859 ( .C1(n16793), .C2(n20012), .A(n16792), .B(n16791), .ZN(
        P2_U2895) );
  INV_X1 U18860 ( .A(n16794), .ZN(n16798) );
  INV_X1 U18861 ( .A(n16795), .ZN(n16797) );
  OAI21_X1 U18862 ( .B1(n16798), .B2(n16797), .A(n16796), .ZN(n19084) );
  OAI22_X1 U18863 ( .A1(n16818), .A2(n19084), .B1(n16817), .B2(n16799), .ZN(
        n16801) );
  NOR2_X1 U18864 ( .A1(n16819), .A2(n19757), .ZN(n16800) );
  AOI211_X1 U18865 ( .C1(BUF1_REG_23__SCAN_IN), .C2(n20064), .A(n16801), .B(
        n16800), .ZN(n16803) );
  NAND2_X1 U18866 ( .A1(n20063), .A2(BUF2_REG_23__SCAN_IN), .ZN(n16802) );
  OAI211_X1 U18867 ( .C1(n16804), .C2(n20012), .A(n16803), .B(n16802), .ZN(
        P2_U2896) );
  INV_X1 U18868 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n16811) );
  NAND2_X1 U18869 ( .A1(n16805), .A2(n20068), .ZN(n16810) );
  OAI22_X1 U18870 ( .A1(n16818), .A2(n19053), .B1(n16817), .B2(n16806), .ZN(
        n16808) );
  NOR2_X1 U18871 ( .A1(n16819), .A2(n20019), .ZN(n16807) );
  AOI211_X1 U18872 ( .C1(BUF1_REG_21__SCAN_IN), .C2(n20064), .A(n16808), .B(
        n16807), .ZN(n16809) );
  OAI211_X1 U18873 ( .C1(n16824), .C2(n16811), .A(n16810), .B(n16809), .ZN(
        P2_U2898) );
  NAND2_X1 U18874 ( .A1(n16812), .A2(n20068), .ZN(n16823) );
  NAND2_X1 U18875 ( .A1(n16814), .A2(n16813), .ZN(n16815) );
  NAND2_X1 U18876 ( .A1(n17133), .A2(n16815), .ZN(n19036) );
  OAI22_X1 U18877 ( .A1(n16818), .A2(n19036), .B1(n16817), .B2(n16816), .ZN(
        n16821) );
  NOR2_X1 U18878 ( .A1(n16819), .A2(n20113), .ZN(n16820) );
  AOI211_X1 U18879 ( .C1(BUF1_REG_19__SCAN_IN), .C2(n20064), .A(n16821), .B(
        n16820), .ZN(n16822) );
  OAI211_X1 U18880 ( .C1(n16824), .C2(n19510), .A(n16823), .B(n16822), .ZN(
        P2_U2900) );
  NOR2_X1 U18881 ( .A1(n17883), .A2(n16825), .ZN(n16826) );
  AOI211_X1 U18882 ( .C1(n17866), .C2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n16827), .B(n16826), .ZN(n16828) );
  OAI21_X1 U18883 ( .B1(n16829), .B2(n17865), .A(n16828), .ZN(n16830) );
  AOI21_X1 U18884 ( .B1(n16831), .B2(n17879), .A(n16830), .ZN(n16832) );
  OAI21_X1 U18885 ( .B1(n16833), .B2(n17860), .A(n16832), .ZN(P2_U2984) );
  INV_X1 U18886 ( .A(n16834), .ZN(n16835) );
  NAND2_X1 U18887 ( .A1(n16835), .A2(n11155), .ZN(n17046) );
  NAND2_X1 U18888 ( .A1(n17850), .A2(n16836), .ZN(n16837) );
  NAND2_X1 U18889 ( .A1(n19213), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n17040) );
  OAI211_X1 U18890 ( .C1(n17029), .C2(n16838), .A(n16837), .B(n17040), .ZN(
        n16839) );
  AOI21_X1 U18891 ( .B1(n19140), .B2(n17878), .A(n16839), .ZN(n16845) );
  NAND2_X1 U18892 ( .A1(n16842), .A2(n16841), .ZN(n16843) );
  XNOR2_X1 U18893 ( .A(n16840), .B(n16843), .ZN(n17043) );
  NAND2_X1 U18894 ( .A1(n17043), .A2(n17879), .ZN(n16844) );
  OAI211_X1 U18895 ( .C1(n17046), .C2(n17860), .A(n16845), .B(n16844), .ZN(
        P2_U2985) );
  AOI21_X1 U18896 ( .B1(n16846), .B2(n16847), .A(n17058), .ZN(n16848) );
  OAI22_X1 U18897 ( .A1(n11220), .A2(n16848), .B1(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n16847), .ZN(n17065) );
  NOR2_X2 U18898 ( .A1(n16850), .A2(n16849), .ZN(n17055) );
  NOR2_X1 U18899 ( .A1(n18976), .A2(n17979), .ZN(n17056) );
  INV_X1 U18900 ( .A(n17056), .ZN(n16851) );
  OAI21_X1 U18901 ( .B1(n17029), .B2(n19120), .A(n16851), .ZN(n16853) );
  NOR2_X1 U18902 ( .A1(n19118), .A2(n17865), .ZN(n16852) );
  AOI211_X1 U18903 ( .C1(n17850), .C2(n16854), .A(n16853), .B(n16852), .ZN(
        n16855) );
  OAI211_X1 U18904 ( .C1(n17065), .C2(n17859), .A(n16856), .B(n16855), .ZN(
        P2_U2987) );
  NOR2_X1 U18905 ( .A1(n12765), .A2(n16858), .ZN(n16859) );
  XNOR2_X1 U18906 ( .A(n11631), .B(n16859), .ZN(n17088) );
  AOI21_X1 U18907 ( .B1(n17079), .B2(n16860), .A(n11154), .ZN(n17078) );
  NAND2_X1 U18908 ( .A1(n17078), .A2(n12415), .ZN(n16866) );
  NAND2_X1 U18909 ( .A1(n19213), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n17082) );
  OAI21_X1 U18910 ( .B1(n17029), .B2(n16861), .A(n17082), .ZN(n16863) );
  NOR2_X1 U18911 ( .A1(n19099), .A2(n17865), .ZN(n16862) );
  AOI211_X1 U18912 ( .C1(n17850), .C2(n16864), .A(n16863), .B(n16862), .ZN(
        n16865) );
  OAI211_X1 U18913 ( .C1(n17859), .C2(n17088), .A(n16866), .B(n16865), .ZN(
        P2_U2989) );
  OAI21_X1 U18914 ( .B1(n16867), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n16860), .ZN(n17098) );
  XNOR2_X1 U18915 ( .A(n16869), .B(n11610), .ZN(n16870) );
  XNOR2_X1 U18916 ( .A(n16868), .B(n16870), .ZN(n17096) );
  NOR2_X1 U18917 ( .A1(n18976), .A2(n17974), .ZN(n17089) );
  NOR2_X1 U18918 ( .A1(n17883), .A2(n19091), .ZN(n16871) );
  AOI211_X1 U18919 ( .C1(n17866), .C2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n17089), .B(n16871), .ZN(n16872) );
  OAI21_X1 U18920 ( .B1(n19087), .B2(n17865), .A(n16872), .ZN(n16873) );
  AOI21_X1 U18921 ( .B1(n17096), .B2(n17879), .A(n16873), .ZN(n16874) );
  OAI21_X1 U18922 ( .B1(n17098), .B2(n17860), .A(n16874), .ZN(P2_U2990) );
  INV_X1 U18923 ( .A(n16876), .ZN(n16878) );
  NAND2_X1 U18924 ( .A1(n16878), .A2(n16877), .ZN(n16879) );
  XNOR2_X1 U18925 ( .A(n16875), .B(n16879), .ZN(n17108) );
  AOI21_X1 U18926 ( .B1(n17100), .B2(n16880), .A(n16867), .ZN(n17099) );
  NAND2_X1 U18927 ( .A1(n17099), .A2(n12415), .ZN(n16885) );
  NAND2_X1 U18928 ( .A1(n17850), .A2(n16881), .ZN(n16882) );
  NAND2_X1 U18929 ( .A1(n19213), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n17102) );
  OAI211_X1 U18930 ( .C1(n17029), .C2(n19076), .A(n16882), .B(n17102), .ZN(
        n16883) );
  AOI21_X1 U18931 ( .B1(n19073), .B2(n17878), .A(n16883), .ZN(n16884) );
  OAI211_X1 U18932 ( .C1(n17859), .C2(n17108), .A(n16885), .B(n16884), .ZN(
        P2_U2991) );
  XNOR2_X1 U18933 ( .A(n16886), .B(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16887) );
  XNOR2_X1 U18934 ( .A(n16888), .B(n16887), .ZN(n17121) );
  NAND2_X1 U18935 ( .A1(n12812), .A2(n17110), .ZN(n17109) );
  NAND3_X1 U18936 ( .A1(n16880), .A2(n12415), .A3(n17109), .ZN(n16892) );
  NOR2_X1 U18937 ( .A1(n18976), .A2(n17972), .ZN(n17114) );
  AOI21_X1 U18938 ( .B1(n17866), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n17114), .ZN(n16889) );
  OAI21_X1 U18939 ( .B1(n17883), .B2(n19068), .A(n16889), .ZN(n16890) );
  AOI21_X1 U18940 ( .B1(n19065), .B2(n17878), .A(n16890), .ZN(n16891) );
  OAI211_X1 U18941 ( .C1(n17121), .C2(n17859), .A(n16892), .B(n16891), .ZN(
        P2_U2992) );
  XNOR2_X1 U18942 ( .A(n16893), .B(n17138), .ZN(n17146) );
  AOI21_X1 U18943 ( .B1(n17138), .B2(n17154), .A(n11232), .ZN(n17144) );
  NOR2_X1 U18944 ( .A1(n19042), .A2(n17865), .ZN(n16897) );
  NAND2_X1 U18945 ( .A1(n17016), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n17136) );
  NAND2_X1 U18946 ( .A1(n17866), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16895) );
  OAI211_X1 U18947 ( .C1(n17883), .C2(n19051), .A(n17136), .B(n16895), .ZN(
        n16896) );
  AOI211_X1 U18948 ( .C1(n17144), .C2(n12415), .A(n16897), .B(n16896), .ZN(
        n16898) );
  OAI21_X1 U18949 ( .B1(n17146), .B2(n17859), .A(n16898), .ZN(P2_U2994) );
  NAND2_X1 U18950 ( .A1(n16900), .A2(n16899), .ZN(n16903) );
  XNOR2_X1 U18951 ( .A(n16901), .B(n17159), .ZN(n16912) );
  OAI22_X1 U18952 ( .A1(n16912), .A2(n16911), .B1(n17159), .B2(n16901), .ZN(
        n16902) );
  XOR2_X1 U18953 ( .A(n16903), .B(n16902), .Z(n17158) );
  NAND2_X1 U18954 ( .A1(n17016), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n17150) );
  OAI21_X1 U18955 ( .B1(n17029), .B2(n16904), .A(n17150), .ZN(n16906) );
  NOR2_X1 U18956 ( .A1(n17147), .A2(n17865), .ZN(n16905) );
  AOI211_X1 U18957 ( .C1(n17850), .C2(n19030), .A(n16906), .B(n16905), .ZN(
        n16910) );
  AND2_X1 U18958 ( .A1(n16907), .A2(n17139), .ZN(n16913) );
  INV_X1 U18959 ( .A(n16913), .ZN(n16908) );
  NAND2_X1 U18960 ( .A1(n16908), .A2(n17148), .ZN(n17155) );
  NAND3_X1 U18961 ( .A1(n17155), .A2(n12415), .A3(n17154), .ZN(n16909) );
  OAI211_X1 U18962 ( .C1(n17158), .C2(n17859), .A(n16910), .B(n16909), .ZN(
        P2_U2995) );
  XNOR2_X1 U18963 ( .A(n16912), .B(n16911), .ZN(n17169) );
  INV_X1 U18964 ( .A(n17173), .ZN(n17188) );
  NAND2_X1 U18965 ( .A1(n16907), .A2(n17188), .ZN(n16938) );
  AOI21_X1 U18966 ( .B1(n17179), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16914) );
  NOR2_X1 U18967 ( .A1(n16914), .A2(n16913), .ZN(n17167) );
  NOR2_X1 U18968 ( .A1(n18976), .A2(n19011), .ZN(n17162) );
  NOR2_X1 U18969 ( .A1(n17883), .A2(n19017), .ZN(n16915) );
  AOI211_X1 U18970 ( .C1(n17866), .C2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n17162), .B(n16915), .ZN(n16916) );
  OAI21_X1 U18971 ( .B1(n19019), .B2(n17865), .A(n16916), .ZN(n16917) );
  AOI21_X1 U18972 ( .B1(n17167), .B2(n12415), .A(n16917), .ZN(n16918) );
  OAI21_X1 U18973 ( .B1(n17169), .B2(n17859), .A(n16918), .ZN(P2_U2996) );
  XNOR2_X1 U18974 ( .A(n17179), .B(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16927) );
  NAND2_X1 U18975 ( .A1(n16920), .A2(n16919), .ZN(n16921) );
  XNOR2_X1 U18976 ( .A(n16922), .B(n16921), .ZN(n17180) );
  AND2_X1 U18977 ( .A1(n19213), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n17181) );
  AOI21_X1 U18978 ( .B1(n17866), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n17181), .ZN(n16924) );
  NAND2_X1 U18979 ( .A1(n17850), .A2(n19001), .ZN(n16923) );
  OAI211_X1 U18980 ( .C1(n19005), .C2(n17865), .A(n16924), .B(n16923), .ZN(
        n16925) );
  AOI21_X1 U18981 ( .B1(n17180), .B2(n17879), .A(n16925), .ZN(n16926) );
  OAI21_X1 U18982 ( .B1(n17860), .B2(n16927), .A(n16926), .ZN(P2_U2997) );
  INV_X1 U18983 ( .A(n16938), .ZN(n17195) );
  OAI21_X1 U18984 ( .B1(n17195), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n12415), .ZN(n16936) );
  INV_X1 U18985 ( .A(n16928), .ZN(n18994) );
  NAND2_X1 U18986 ( .A1(n19213), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n17189) );
  NAND2_X1 U18987 ( .A1(n17866), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16929) );
  OAI211_X1 U18988 ( .C1(n17883), .C2(n18992), .A(n17189), .B(n16929), .ZN(
        n16934) );
  NOR2_X1 U18989 ( .A1(n16931), .A2(n16930), .ZN(n17191) );
  INV_X1 U18990 ( .A(n16932), .ZN(n17190) );
  NOR3_X1 U18991 ( .A1(n17191), .A2(n17190), .A3(n17859), .ZN(n16933) );
  AOI211_X1 U18992 ( .C1(n18994), .C2(n17878), .A(n16934), .B(n16933), .ZN(
        n16935) );
  OAI21_X1 U18993 ( .B1(n17179), .B2(n16936), .A(n16935), .ZN(P2_U2998) );
  INV_X1 U18994 ( .A(n16937), .ZN(n17242) );
  NAND2_X1 U18995 ( .A1(n16980), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16963) );
  INV_X1 U18996 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17215) );
  NOR2_X1 U18997 ( .A1(n16963), .A2(n17215), .ZN(n16956) );
  OAI21_X1 U18998 ( .B1(n16956), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n16938), .ZN(n17209) );
  INV_X1 U18999 ( .A(n16969), .ZN(n16940) );
  OAI21_X1 U19000 ( .B1(n16940), .B2(n16939), .A(n16968), .ZN(n16955) );
  INV_X1 U19001 ( .A(n16943), .ZN(n16942) );
  NAND2_X1 U19002 ( .A1(n16942), .A2(n16941), .ZN(n16954) );
  NOR2_X1 U19003 ( .A1(n16955), .A2(n16954), .ZN(n16953) );
  NOR2_X1 U19004 ( .A1(n16953), .A2(n16943), .ZN(n16947) );
  NAND2_X1 U19005 ( .A1(n16945), .A2(n16944), .ZN(n16946) );
  XNOR2_X1 U19006 ( .A(n16947), .B(n16946), .ZN(n17207) );
  NAND2_X1 U19007 ( .A1(n18982), .A2(n17878), .ZN(n16949) );
  INV_X1 U19008 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n17967) );
  NOR2_X1 U19009 ( .A1(n18976), .A2(n17967), .ZN(n17202) );
  AOI21_X1 U19010 ( .B1(n17866), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n17202), .ZN(n16948) );
  OAI211_X1 U19011 ( .C1(n17883), .C2(n16950), .A(n16949), .B(n16948), .ZN(
        n16951) );
  AOI21_X1 U19012 ( .B1(n17207), .B2(n17879), .A(n16951), .ZN(n16952) );
  OAI21_X1 U19013 ( .B1(n17209), .B2(n17860), .A(n16952), .ZN(P2_U2999) );
  AOI21_X1 U19014 ( .B1(n16955), .B2(n16954), .A(n16953), .ZN(n17225) );
  AOI21_X1 U19015 ( .B1(n17215), .B2(n16963), .A(n16956), .ZN(n17210) );
  NAND2_X1 U19016 ( .A1(n17210), .A2(n12415), .ZN(n16962) );
  NOR2_X1 U19017 ( .A1(n18976), .A2(n17966), .ZN(n17214) );
  AOI21_X1 U19018 ( .B1(n17866), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n17214), .ZN(n16957) );
  OAI21_X1 U19019 ( .B1(n17883), .B2(n16958), .A(n16957), .ZN(n16959) );
  AOI21_X1 U19020 ( .B1(n16960), .B2(n17878), .A(n16959), .ZN(n16961) );
  OAI211_X1 U19021 ( .C1(n17225), .C2(n17859), .A(n16962), .B(n16961), .ZN(
        P2_U3000) );
  OAI21_X1 U19022 ( .B1(n16980), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n16963), .ZN(n17238) );
  NAND2_X1 U19023 ( .A1(n17850), .A2(n18963), .ZN(n16964) );
  NAND2_X1 U19024 ( .A1(n17016), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n17227) );
  OAI211_X1 U19025 ( .C1(n17029), .C2(n16965), .A(n16964), .B(n17227), .ZN(
        n16966) );
  AOI21_X1 U19026 ( .B1(n18968), .B2(n17878), .A(n16966), .ZN(n16973) );
  NAND2_X1 U19027 ( .A1(n16968), .A2(n16967), .ZN(n16971) );
  NAND2_X1 U19028 ( .A1(n16969), .A2(n16975), .ZN(n16970) );
  XOR2_X1 U19029 ( .A(n16971), .B(n16970), .Z(n17236) );
  NAND2_X1 U19030 ( .A1(n17236), .A2(n17879), .ZN(n16972) );
  OAI211_X1 U19031 ( .C1(n17238), .C2(n17860), .A(n16973), .B(n16972), .ZN(
        P2_U3001) );
  NAND2_X1 U19032 ( .A1(n16975), .A2(n16974), .ZN(n16979) );
  NAND2_X1 U19033 ( .A1(n16977), .A2(n16976), .ZN(n16978) );
  XOR2_X1 U19034 ( .A(n16979), .B(n16978), .Z(n17252) );
  INV_X1 U19035 ( .A(n16980), .ZN(n17240) );
  NAND2_X1 U19036 ( .A1(n16987), .A2(n17228), .ZN(n17239) );
  NAND3_X1 U19037 ( .A1(n17240), .A2(n12415), .A3(n17239), .ZN(n16986) );
  NAND2_X1 U19038 ( .A1(n17016), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n17244) );
  NAND2_X1 U19039 ( .A1(n17866), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16981) );
  OAI211_X1 U19040 ( .C1(n17883), .C2(n16982), .A(n17244), .B(n16981), .ZN(
        n16983) );
  AOI21_X1 U19041 ( .B1(n16984), .B2(n17878), .A(n16983), .ZN(n16985) );
  OAI211_X1 U19042 ( .C1(n17252), .C2(n17859), .A(n16986), .B(n16985), .ZN(
        P2_U3002) );
  AND2_X1 U19043 ( .A1(n17014), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16988) );
  OAI21_X1 U19044 ( .B1(n16988), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n16987), .ZN(n17263) );
  NAND2_X1 U19045 ( .A1(n16990), .A2(n16989), .ZN(n16994) );
  NOR2_X1 U19046 ( .A1(n16992), .A2(n16991), .ZN(n16993) );
  XOR2_X1 U19047 ( .A(n16994), .B(n16993), .Z(n17260) );
  NOR2_X1 U19048 ( .A1(n18976), .A2(n17964), .ZN(n17255) );
  NOR2_X1 U19049 ( .A1(n17883), .A2(n18961), .ZN(n16995) );
  AOI211_X1 U19050 ( .C1(n17866), .C2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n17255), .B(n16995), .ZN(n16996) );
  OAI21_X1 U19051 ( .B1(n17865), .B2(n18947), .A(n16996), .ZN(n16997) );
  AOI21_X1 U19052 ( .B1(n17260), .B2(n17879), .A(n16997), .ZN(n16998) );
  OAI21_X1 U19053 ( .B1(n17263), .B2(n17860), .A(n16998), .ZN(P2_U3003) );
  NAND2_X1 U19054 ( .A1(n17000), .A2(n16999), .ZN(n17003) );
  NAND2_X1 U19055 ( .A1(n17001), .A2(n17011), .ZN(n17002) );
  XOR2_X1 U19056 ( .A(n17003), .B(n17002), .Z(n17276) );
  XNOR2_X1 U19057 ( .A(n17014), .B(n17270), .ZN(n17264) );
  NAND2_X1 U19058 ( .A1(n17264), .A2(n12415), .ZN(n17009) );
  INV_X1 U19059 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17004) );
  NAND2_X1 U19060 ( .A1(n17016), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n17265) );
  OAI21_X1 U19061 ( .B1(n17029), .B2(n17004), .A(n17265), .ZN(n17007) );
  NOR2_X1 U19062 ( .A1(n17883), .A2(n17005), .ZN(n17006) );
  AOI211_X1 U19063 ( .C1(n17267), .C2(n17878), .A(n17007), .B(n17006), .ZN(
        n17008) );
  OAI211_X1 U19064 ( .C1(n17276), .C2(n17859), .A(n17009), .B(n17008), .ZN(
        P2_U3004) );
  NAND2_X1 U19065 ( .A1(n17011), .A2(n17010), .ZN(n17013) );
  XOR2_X1 U19066 ( .A(n17013), .B(n17012), .Z(n17289) );
  INV_X1 U19067 ( .A(n17014), .ZN(n17278) );
  INV_X1 U19068 ( .A(n16907), .ZN(n17015) );
  NAND2_X1 U19069 ( .A1(n17015), .A2(n17279), .ZN(n17277) );
  NAND3_X1 U19070 ( .A1(n17278), .A2(n12415), .A3(n17277), .ZN(n17020) );
  NAND2_X1 U19071 ( .A1(n17016), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n17281) );
  OAI21_X1 U19072 ( .B1(n17029), .B2(n18933), .A(n17281), .ZN(n17018) );
  NOR2_X1 U19073 ( .A1(n17865), .A2(n18941), .ZN(n17017) );
  AOI211_X1 U19074 ( .C1(n17850), .C2(n18937), .A(n17018), .B(n17017), .ZN(
        n17019) );
  OAI211_X1 U19075 ( .C1(n17859), .C2(n17289), .A(n17020), .B(n17019), .ZN(
        P2_U3005) );
  NAND2_X1 U19076 ( .A1(n17023), .A2(n17022), .ZN(n17303) );
  XNOR2_X1 U19077 ( .A(n17021), .B(n11297), .ZN(n17302) );
  AND2_X1 U19078 ( .A1(n17303), .A2(n17302), .ZN(n17305) );
  AOI21_X1 U19079 ( .B1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17021), .A(
        n17305), .ZN(n17026) );
  NAND2_X1 U19080 ( .A1(n17873), .A2(n17024), .ZN(n17025) );
  XNOR2_X1 U19081 ( .A(n17026), .B(n17025), .ZN(n17301) );
  OR2_X1 U19082 ( .A1(n17027), .A2(n17028), .ZN(n17290) );
  NAND2_X1 U19083 ( .A1(n17027), .A2(n17028), .ZN(n17868) );
  NAND3_X1 U19084 ( .A1(n17290), .A2(n12415), .A3(n17868), .ZN(n17034) );
  NOR2_X1 U19085 ( .A1(n17865), .A2(n18927), .ZN(n17032) );
  OAI22_X1 U19086 ( .A1(n17030), .A2(n17029), .B1(n17958), .B2(n18976), .ZN(
        n17031) );
  AOI211_X1 U19087 ( .C1(n17850), .C2(n18923), .A(n17032), .B(n17031), .ZN(
        n17033) );
  OAI211_X1 U19088 ( .C1(n17301), .C2(n17859), .A(n17034), .B(n17033), .ZN(
        P2_U3007) );
  INV_X1 U19089 ( .A(n17035), .ZN(n17057) );
  NAND3_X1 U19090 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n17057), .ZN(n17038) );
  AOI21_X1 U19091 ( .B1(n17036), .B2(n17057), .A(n17062), .ZN(n17037) );
  AOI21_X1 U19092 ( .B1(n17039), .B2(n17038), .A(n17037), .ZN(n17042) );
  OAI21_X1 U19093 ( .B1(n19138), .B2(n19180), .A(n17040), .ZN(n17041) );
  AOI211_X1 U19094 ( .C1(n19140), .C2(n19202), .A(n17042), .B(n17041), .ZN(
        n17045) );
  NAND2_X1 U19095 ( .A1(n17043), .A2(n19211), .ZN(n17044) );
  OAI211_X1 U19096 ( .C1(n17046), .C2(n19187), .A(n17045), .B(n17044), .ZN(
        P2_U3017) );
  XNOR2_X1 U19097 ( .A(n17058), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n17047) );
  NAND2_X1 U19098 ( .A1(n17047), .A2(n17057), .ZN(n17048) );
  OAI211_X1 U19099 ( .C1(n17050), .C2(n19180), .A(n17049), .B(n17048), .ZN(
        n17051) );
  NAND2_X1 U19100 ( .A1(n17055), .A2(n12758), .ZN(n17064) );
  AOI21_X1 U19101 ( .B1(n17058), .B2(n17057), .A(n17056), .ZN(n17059) );
  OAI21_X1 U19102 ( .B1(n19132), .B2(n19180), .A(n17059), .ZN(n17061) );
  NOR2_X1 U19103 ( .A1(n19118), .A2(n17283), .ZN(n17060) );
  AOI211_X1 U19104 ( .C1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n17062), .A(
        n17061), .B(n17060), .ZN(n17063) );
  OAI211_X1 U19105 ( .C1(n19178), .C2(n17065), .A(n17064), .B(n17063), .ZN(
        P2_U3019) );
  NAND2_X1 U19106 ( .A1(n17079), .A2(n17067), .ZN(n17081) );
  AOI21_X1 U19107 ( .B1(n17080), .B2(n17081), .A(n17066), .ZN(n17073) );
  NAND3_X1 U19108 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17067), .A3(
        n17066), .ZN(n17070) );
  INV_X1 U19109 ( .A(n17068), .ZN(n17069) );
  OAI211_X1 U19110 ( .C1(n17071), .C2(n19180), .A(n17070), .B(n17069), .ZN(
        n17072) );
  AOI211_X1 U19111 ( .C1(n19110), .C2(n19202), .A(n17073), .B(n17072), .ZN(
        n17076) );
  OR2_X1 U19112 ( .A1(n17074), .A2(n19178), .ZN(n17075) );
  OAI211_X1 U19113 ( .C1(n17077), .C2(n19187), .A(n17076), .B(n17075), .ZN(
        P2_U3020) );
  NAND2_X1 U19114 ( .A1(n17078), .A2(n12758), .ZN(n17087) );
  INV_X1 U19115 ( .A(n19099), .ZN(n17085) );
  NOR2_X1 U19116 ( .A1(n17080), .A2(n17079), .ZN(n17084) );
  OAI211_X1 U19117 ( .C1(n19097), .C2(n19180), .A(n17082), .B(n17081), .ZN(
        n17083) );
  AOI211_X1 U19118 ( .C1(n17085), .C2(n19202), .A(n17084), .B(n17083), .ZN(
        n17086) );
  OAI211_X1 U19119 ( .C1(n17088), .C2(n19178), .A(n17087), .B(n17086), .ZN(
        P2_U3021) );
  AOI211_X1 U19120 ( .C1(n19208), .C2(n17091), .A(n17090), .B(n17089), .ZN(
        n17094) );
  NAND2_X1 U19121 ( .A1(n17092), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17093) );
  OAI211_X1 U19122 ( .C1(n19087), .C2(n17283), .A(n17094), .B(n17093), .ZN(
        n17095) );
  AOI21_X1 U19123 ( .B1(n17096), .B2(n19211), .A(n17095), .ZN(n17097) );
  OAI21_X1 U19124 ( .B1(n17098), .B2(n19187), .A(n17097), .ZN(P2_U3022) );
  NAND2_X1 U19125 ( .A1(n17099), .A2(n12758), .ZN(n17107) );
  NAND2_X1 U19126 ( .A1(n17110), .A2(n17101), .ZN(n17115) );
  AOI21_X1 U19127 ( .B1(n17111), .B2(n17115), .A(n17100), .ZN(n17105) );
  NAND3_X1 U19128 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17101), .A3(
        n17100), .ZN(n17103) );
  OAI211_X1 U19129 ( .C1(n19180), .C2(n19084), .A(n17103), .B(n17102), .ZN(
        n17104) );
  AOI211_X1 U19130 ( .C1(n19073), .C2(n19202), .A(n17105), .B(n17104), .ZN(
        n17106) );
  OAI211_X1 U19131 ( .C1(n17108), .C2(n19178), .A(n17107), .B(n17106), .ZN(
        P2_U3023) );
  NAND3_X1 U19132 ( .A1(n16880), .A2(n12758), .A3(n17109), .ZN(n17120) );
  NOR2_X1 U19133 ( .A1(n17111), .A2(n17110), .ZN(n17118) );
  OR2_X1 U19134 ( .A1(n12826), .A2(n17112), .ZN(n17113) );
  NAND2_X1 U19135 ( .A1(n16794), .A2(n17113), .ZN(n19963) );
  INV_X1 U19136 ( .A(n17114), .ZN(n17116) );
  OAI211_X1 U19137 ( .C1(n19180), .C2(n19963), .A(n17116), .B(n17115), .ZN(
        n17117) );
  AOI211_X1 U19138 ( .C1(n19065), .C2(n19202), .A(n17118), .B(n17117), .ZN(
        n17119) );
  OAI211_X1 U19139 ( .C1(n17121), .C2(n19178), .A(n17120), .B(n17119), .ZN(
        P2_U3024) );
  NAND2_X1 U19140 ( .A1(n17188), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n17122) );
  NOR2_X1 U19141 ( .A1(n17211), .A2(n17122), .ZN(n17170) );
  AND2_X1 U19142 ( .A1(n17159), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17123) );
  NAND2_X1 U19143 ( .A1(n17170), .A2(n17123), .ZN(n17164) );
  NAND3_X1 U19144 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17127) );
  OR2_X1 U19145 ( .A1(n17125), .A2(n17124), .ZN(n17126) );
  OAI211_X1 U19146 ( .C1(n17174), .C2(n17127), .A(n19183), .B(n17126), .ZN(
        n17128) );
  NAND2_X1 U19147 ( .A1(n17171), .A2(n17200), .ZN(n17172) );
  AND2_X1 U19148 ( .A1(n17128), .A2(n17172), .ZN(n17129) );
  AND2_X1 U19149 ( .A1(n17130), .A2(n17129), .ZN(n17160) );
  AND2_X1 U19150 ( .A1(n17164), .A2(n17160), .ZN(n17149) );
  NAND2_X1 U19151 ( .A1(n17131), .A2(n17148), .ZN(n17151) );
  AOI21_X1 U19152 ( .B1(n17149), .B2(n17151), .A(n17138), .ZN(n17143) );
  AND2_X1 U19153 ( .A1(n17133), .A2(n17132), .ZN(n17134) );
  NOR2_X1 U19154 ( .A1(n17135), .A2(n17134), .ZN(n20066) );
  INV_X1 U19155 ( .A(n17136), .ZN(n17137) );
  AOI21_X1 U19156 ( .B1(n19208), .B2(n20066), .A(n17137), .ZN(n17141) );
  INV_X1 U19157 ( .A(n17211), .ZN(n17280) );
  NAND4_X1 U19158 ( .A1(n17280), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n17139), .A4(n17138), .ZN(n17140) );
  OAI211_X1 U19159 ( .C1(n19042), .C2(n17283), .A(n17141), .B(n17140), .ZN(
        n17142) );
  AOI211_X1 U19160 ( .C1(n17144), .C2(n12758), .A(n17143), .B(n17142), .ZN(
        n17145) );
  OAI21_X1 U19161 ( .B1(n17146), .B2(n19178), .A(n17145), .ZN(P2_U3026) );
  INV_X1 U19162 ( .A(n17147), .ZN(n19032) );
  NOR2_X1 U19163 ( .A1(n17149), .A2(n17148), .ZN(n17153) );
  OAI211_X1 U19164 ( .C1(n19180), .C2(n19036), .A(n17151), .B(n17150), .ZN(
        n17152) );
  AOI211_X1 U19165 ( .C1(n19032), .C2(n19202), .A(n17153), .B(n17152), .ZN(
        n17157) );
  NAND3_X1 U19166 ( .A1(n17155), .A2(n12758), .A3(n17154), .ZN(n17156) );
  OAI211_X1 U19167 ( .C1(n17158), .C2(n19178), .A(n17157), .B(n17156), .ZN(
        P2_U3027) );
  NOR2_X1 U19168 ( .A1(n17160), .A2(n17159), .ZN(n17161) );
  AOI211_X1 U19169 ( .C1(n19208), .C2(n17163), .A(n17162), .B(n17161), .ZN(
        n17165) );
  OAI211_X1 U19170 ( .C1(n19019), .C2(n17283), .A(n17165), .B(n17164), .ZN(
        n17166) );
  AOI21_X1 U19171 ( .B1(n17167), .B2(n12758), .A(n17166), .ZN(n17168) );
  OAI21_X1 U19172 ( .B1(n17169), .B2(n19178), .A(n17168), .ZN(P2_U3028) );
  AOI21_X1 U19173 ( .B1(n17179), .B2(n12758), .A(n17170), .ZN(n17187) );
  NOR2_X1 U19174 ( .A1(n12758), .A2(n17171), .ZN(n17194) );
  INV_X1 U19175 ( .A(n17172), .ZN(n17176) );
  AND2_X1 U19176 ( .A1(n17174), .A2(n17173), .ZN(n17175) );
  OR3_X1 U19177 ( .A1(n17286), .A2(n17176), .A3(n17175), .ZN(n17203) );
  AOI21_X1 U19178 ( .B1(n17177), .B2(n19183), .A(n17203), .ZN(n17178) );
  OAI21_X1 U19179 ( .B1(n17179), .B2(n17194), .A(n17178), .ZN(n17185) );
  NAND2_X1 U19180 ( .A1(n17180), .A2(n19211), .ZN(n17183) );
  AOI21_X1 U19181 ( .B1(n19208), .B2(n19006), .A(n17181), .ZN(n17182) );
  OAI211_X1 U19182 ( .C1(n19005), .C2(n17283), .A(n17183), .B(n17182), .ZN(
        n17184) );
  AOI21_X1 U19183 ( .B1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17185), .A(
        n17184), .ZN(n17186) );
  OAI21_X1 U19184 ( .B1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17187), .A(
        n17186), .ZN(P2_U3029) );
  AOI22_X1 U19185 ( .A1(n17195), .A2(n12758), .B1(n17188), .B2(n17280), .ZN(
        n17199) );
  OAI21_X1 U19186 ( .B1(n19180), .B2(n18998), .A(n17189), .ZN(n17193) );
  NOR3_X1 U19187 ( .A1(n17191), .A2(n17190), .A3(n19178), .ZN(n17192) );
  AOI211_X1 U19188 ( .C1(n19202), .C2(n18994), .A(n17193), .B(n17192), .ZN(
        n17198) );
  NOR2_X1 U19189 ( .A1(n17195), .A2(n17194), .ZN(n17196) );
  OAI21_X1 U19190 ( .B1(n17196), .B2(n17203), .A(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17197) );
  OAI211_X1 U19191 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n17199), .A(
        n17198), .B(n17197), .ZN(P2_U3030) );
  NOR3_X1 U19192 ( .A1(n17211), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        n17200), .ZN(n17201) );
  AOI211_X1 U19193 ( .C1(n18982), .C2(n19202), .A(n17202), .B(n17201), .ZN(
        n17205) );
  NAND2_X1 U19194 ( .A1(n17203), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17204) );
  OAI211_X1 U19195 ( .C1(n18986), .C2(n19180), .A(n17205), .B(n17204), .ZN(
        n17206) );
  AOI21_X1 U19196 ( .B1(n17207), .B2(n19211), .A(n17206), .ZN(n17208) );
  OAI21_X1 U19197 ( .B1(n17209), .B2(n19187), .A(n17208), .ZN(P2_U3031) );
  NAND2_X1 U19198 ( .A1(n17210), .A2(n12758), .ZN(n17224) );
  INV_X1 U19199 ( .A(n19744), .ZN(n17222) );
  NOR2_X1 U19200 ( .A1(n17211), .A2(n17279), .ZN(n17253) );
  NAND2_X1 U19201 ( .A1(n17253), .A2(n17242), .ZN(n17213) );
  NOR2_X1 U19202 ( .A1(n17213), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17248) );
  AOI21_X1 U19203 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17242), .A(
        n17318), .ZN(n17212) );
  NOR3_X1 U19204 ( .A1(n17248), .A2(n17212), .A3(n17286), .ZN(n17234) );
  OR2_X1 U19205 ( .A1(n17213), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17229) );
  AOI21_X1 U19206 ( .B1(n17234), .B2(n17229), .A(n17215), .ZN(n17221) );
  INV_X1 U19207 ( .A(n17214), .ZN(n17218) );
  NAND3_X1 U19208 ( .A1(n17280), .A2(n17216), .A3(n17215), .ZN(n17217) );
  OAI211_X1 U19209 ( .C1(n17219), .C2(n17283), .A(n17218), .B(n17217), .ZN(
        n17220) );
  AOI211_X1 U19210 ( .C1(n17222), .C2(n19208), .A(n17221), .B(n17220), .ZN(
        n17223) );
  OAI211_X1 U19211 ( .C1(n17225), .C2(n19178), .A(n17224), .B(n17223), .ZN(
        P2_U3032) );
  NAND2_X1 U19212 ( .A1(n17226), .A2(n19208), .ZN(n17232) );
  OAI21_X1 U19213 ( .B1(n17229), .B2(n17228), .A(n17227), .ZN(n17230) );
  AOI21_X1 U19214 ( .B1(n18968), .B2(n19202), .A(n17230), .ZN(n17231) );
  OAI211_X1 U19215 ( .C1(n17234), .C2(n17233), .A(n17232), .B(n17231), .ZN(
        n17235) );
  AOI21_X1 U19216 ( .B1(n17236), .B2(n19211), .A(n17235), .ZN(n17237) );
  OAI21_X1 U19217 ( .B1(n17238), .B2(n19187), .A(n17237), .ZN(P2_U3033) );
  NAND3_X1 U19218 ( .A1(n17240), .A2(n12758), .A3(n17239), .ZN(n17251) );
  AND2_X1 U19219 ( .A1(n19183), .A2(n17279), .ZN(n17241) );
  NOR2_X1 U19220 ( .A1(n17286), .A2(n17241), .ZN(n17271) );
  OAI21_X1 U19221 ( .B1(n17242), .B2(n17318), .A(n17271), .ZN(n17243) );
  NAND2_X1 U19222 ( .A1(n17243), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17245) );
  OAI211_X1 U19223 ( .C1(n17246), .C2(n17283), .A(n17245), .B(n17244), .ZN(
        n17247) );
  AOI211_X1 U19224 ( .C1(n17249), .C2(n19208), .A(n17248), .B(n17247), .ZN(
        n17250) );
  OAI211_X1 U19225 ( .C1(n17252), .C2(n19178), .A(n17251), .B(n17250), .ZN(
        P2_U3034) );
  NAND2_X1 U19226 ( .A1(n17253), .A2(n17270), .ZN(n17268) );
  AOI21_X1 U19227 ( .B1(n17268), .B2(n17271), .A(n17254), .ZN(n17259) );
  NAND4_X1 U19228 ( .A1(n17280), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A4(n17254), .ZN(n17257) );
  INV_X1 U19229 ( .A(n17255), .ZN(n17256) );
  OAI211_X1 U19230 ( .C1(n18947), .C2(n17283), .A(n17257), .B(n17256), .ZN(
        n17258) );
  AOI211_X1 U19231 ( .C1(n18955), .C2(n19208), .A(n17259), .B(n17258), .ZN(
        n17262) );
  NAND2_X1 U19232 ( .A1(n17260), .A2(n19211), .ZN(n17261) );
  OAI211_X1 U19233 ( .C1(n17263), .C2(n19187), .A(n17262), .B(n17261), .ZN(
        P2_U3035) );
  NAND2_X1 U19234 ( .A1(n17264), .A2(n12758), .ZN(n17275) );
  INV_X1 U19235 ( .A(n17265), .ZN(n17266) );
  AOI21_X1 U19236 ( .B1(n17267), .B2(n19202), .A(n17266), .ZN(n17269) );
  OAI211_X1 U19237 ( .C1(n17271), .C2(n17270), .A(n17269), .B(n17268), .ZN(
        n17272) );
  AOI21_X1 U19238 ( .B1(n17273), .B2(n19208), .A(n17272), .ZN(n17274) );
  OAI211_X1 U19239 ( .C1(n17276), .C2(n19178), .A(n17275), .B(n17274), .ZN(
        P2_U3036) );
  NAND3_X1 U19240 ( .A1(n17278), .A2(n12758), .A3(n17277), .ZN(n17288) );
  NAND2_X1 U19241 ( .A1(n17280), .A2(n17279), .ZN(n17282) );
  OAI211_X1 U19242 ( .C1(n18941), .C2(n17283), .A(n17282), .B(n17281), .ZN(
        n17285) );
  NOR2_X1 U19243 ( .A1(n18946), .A2(n19180), .ZN(n17284) );
  AOI211_X1 U19244 ( .C1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n17286), .A(
        n17285), .B(n17284), .ZN(n17287) );
  OAI211_X1 U19245 ( .C1(n17289), .C2(n19178), .A(n17288), .B(n17287), .ZN(
        P2_U3037) );
  NAND3_X1 U19246 ( .A1(n17290), .A2(n12758), .A3(n17868), .ZN(n17300) );
  INV_X1 U19247 ( .A(n17291), .ZN(n17292) );
  NOR2_X1 U19248 ( .A1(n17309), .A2(n17292), .ZN(n19195) );
  AND2_X1 U19249 ( .A1(n19183), .A2(n17292), .ZN(n17293) );
  NOR2_X1 U19250 ( .A1(n17294), .A2(n17293), .ZN(n19189) );
  INV_X1 U19251 ( .A(n18927), .ZN(n17296) );
  OAI22_X1 U19252 ( .A1(n19180), .A2(n18928), .B1(n17958), .B2(n18976), .ZN(
        n17295) );
  AOI21_X1 U19253 ( .B1(n19202), .B2(n17296), .A(n17295), .ZN(n17297) );
  OAI21_X1 U19254 ( .B1(n19189), .B2(n19196), .A(n17297), .ZN(n17298) );
  AOI21_X1 U19255 ( .B1(n19195), .B2(n19196), .A(n17298), .ZN(n17299) );
  OAI211_X1 U19256 ( .C1(n17301), .C2(n19178), .A(n17300), .B(n17299), .ZN(
        P2_U3039) );
  NOR2_X1 U19257 ( .A1(n17303), .A2(n17302), .ZN(n17304) );
  OAI21_X1 U19258 ( .B1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17307), .A(
        n17306), .ZN(n17861) );
  OR2_X1 U19259 ( .A1(n17861), .A2(n19187), .ZN(n17317) );
  NOR2_X1 U19260 ( .A1(n17309), .A2(n17308), .ZN(n17315) );
  INV_X1 U19261 ( .A(n18916), .ZN(n17310) );
  AOI22_X1 U19262 ( .A1(n19202), .A2(n17310), .B1(n19213), .B2(
        P2_REIP_REG_6__SCAN_IN), .ZN(n17313) );
  NAND2_X1 U19263 ( .A1(n19208), .A2(n17311), .ZN(n17312) );
  OAI211_X1 U19264 ( .C1(n19189), .C2(n11297), .A(n17313), .B(n17312), .ZN(
        n17314) );
  AOI21_X1 U19265 ( .B1(n17315), .B2(n11297), .A(n17314), .ZN(n17316) );
  OAI211_X1 U19266 ( .C1(n17858), .C2(n19178), .A(n17317), .B(n17316), .ZN(
        P2_U3040) );
  NOR2_X1 U19267 ( .A1(n19176), .A2(n14746), .ZN(n17321) );
  AOI211_X1 U19268 ( .C1(n14746), .C2(n19184), .A(n17319), .B(n17318), .ZN(
        n17320) );
  AOI211_X1 U19269 ( .C1(n12758), .C2(n17322), .A(n17321), .B(n17320), .ZN(
        n17328) );
  AOI22_X1 U19270 ( .A1(n19208), .A2(n17323), .B1(n19202), .B2(n18879), .ZN(
        n17327) );
  NAND2_X1 U19271 ( .A1(n19211), .A2(n17324), .ZN(n17325) );
  NAND4_X1 U19272 ( .A1(n17328), .A2(n17327), .A3(n17326), .A4(n17325), .ZN(
        P2_U3045) );
  INV_X1 U19273 ( .A(n17329), .ZN(n17333) );
  INV_X1 U19274 ( .A(n11892), .ZN(n17331) );
  INV_X1 U19275 ( .A(n11893), .ZN(n17330) );
  NAND2_X1 U19276 ( .A1(n17331), .A2(n17330), .ZN(n17332) );
  AOI22_X1 U19277 ( .A1(n17333), .A2(n17332), .B1(n12709), .B2(n11298), .ZN(
        n17334) );
  OAI21_X1 U19278 ( .B1(n17336), .B2(n17335), .A(n17334), .ZN(n19218) );
  NOR2_X1 U19279 ( .A1(n17337), .A2(n19256), .ZN(n17342) );
  AOI211_X1 U19280 ( .C1(n18857), .C2(n17339), .A(n19015), .B(n17338), .ZN(
        n18881) );
  AOI21_X1 U19281 ( .B1(n19015), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n18881), .ZN(n17350) );
  AOI22_X1 U19282 ( .A1(n19218), .A2(n19170), .B1(n17342), .B2(n17350), .ZN(
        n17340) );
  OAI21_X1 U19283 ( .B1(n19820), .B2(n17365), .A(n17340), .ZN(n17341) );
  MUX2_X1 U19284 ( .A(n17341), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n19166), .Z(P2_U3600) );
  INV_X1 U19285 ( .A(n17342), .ZN(n17351) );
  AND2_X1 U19286 ( .A1(n19241), .A2(n17343), .ZN(n17359) );
  NOR2_X1 U19287 ( .A1(n11890), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n17358) );
  NOR2_X1 U19288 ( .A1(n17358), .A2(n11883), .ZN(n17348) );
  AND2_X1 U19289 ( .A1(n11816), .A2(n17344), .ZN(n17355) );
  INV_X1 U19290 ( .A(n17355), .ZN(n17346) );
  AOI22_X1 U19291 ( .A1(n17346), .A2(n17348), .B1(n12709), .B2(n17345), .ZN(
        n17347) );
  OAI21_X1 U19292 ( .B1(n17359), .B2(n17348), .A(n17347), .ZN(n17349) );
  AOI21_X1 U19293 ( .B1(n17838), .B2(n17364), .A(n17349), .ZN(n19224) );
  OAI222_X1 U19294 ( .A1(n17365), .A2(n19879), .B1(n17351), .B2(n17350), .C1(
        n19263), .C2(n19224), .ZN(n17352) );
  MUX2_X1 U19295 ( .A(n17352), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n19166), .Z(P2_U3599) );
  INV_X1 U19296 ( .A(n12255), .ZN(n17356) );
  NAND2_X1 U19297 ( .A1(n12709), .A2(n17356), .ZN(n17354) );
  INV_X1 U19298 ( .A(n17358), .ZN(n17353) );
  OAI211_X1 U19299 ( .C1(n11883), .C2(n17355), .A(n17354), .B(n17353), .ZN(
        n17361) );
  OAI22_X1 U19300 ( .A1(n17359), .A2(n17358), .B1(n17357), .B2(n17356), .ZN(
        n17360) );
  MUX2_X1 U19301 ( .A(n17361), .B(n17360), .S(n11716), .Z(n17362) );
  AOI211_X1 U19302 ( .C1(n15441), .C2(n17364), .A(n17363), .B(n17362), .ZN(
        n19228) );
  OAI22_X1 U19303 ( .A1(n19880), .A2(n17365), .B1(n19228), .B2(n19263), .ZN(
        n17366) );
  MUX2_X1 U19304 ( .A(n17366), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n19166), .Z(P2_U3596) );
  INV_X1 U19305 ( .A(n21367), .ZN(n21864) );
  NOR2_X1 U19306 ( .A1(n17367), .A2(n21576), .ZN(n21351) );
  AOI22_X1 U19307 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21795), .B1(
        n21351), .B2(n17368), .ZN(n21828) );
  INV_X1 U19308 ( .A(n17369), .ZN(n21390) );
  AOI22_X1 U19309 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n21508), .B1(n21828), 
        .B2(n21390), .ZN(n17370) );
  OAI21_X1 U19310 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21864), .A(
        n17370), .ZN(n17371) );
  MUX2_X1 U19311 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n17371), .S(
        n21393), .Z(n17746) );
  XOR2_X1 U19312 ( .A(DATAI_29_), .B(keyinput_3), .Z(n17375) );
  XOR2_X1 U19313 ( .A(DATAI_30_), .B(keyinput_2), .Z(n17374) );
  XNOR2_X1 U19314 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(keyinput_0), .ZN(n17373) );
  XNOR2_X1 U19315 ( .A(DATAI_31_), .B(keyinput_1), .ZN(n17372) );
  NOR4_X1 U19316 ( .A1(n17375), .A2(n17374), .A3(n17373), .A4(n17372), .ZN(
        n17378) );
  XOR2_X1 U19317 ( .A(DATAI_28_), .B(keyinput_4), .Z(n17377) );
  XOR2_X1 U19318 ( .A(DATAI_27_), .B(keyinput_5), .Z(n17376) );
  NOR3_X1 U19319 ( .A1(n17378), .A2(n17377), .A3(n17376), .ZN(n17384) );
  XNOR2_X1 U19320 ( .A(DATAI_26_), .B(keyinput_6), .ZN(n17383) );
  XOR2_X1 U19321 ( .A(DATAI_24_), .B(keyinput_8), .Z(n17381) );
  XOR2_X1 U19322 ( .A(DATAI_23_), .B(keyinput_9), .Z(n17380) );
  XNOR2_X1 U19323 ( .A(DATAI_25_), .B(keyinput_7), .ZN(n17379) );
  NOR3_X1 U19324 ( .A1(n17381), .A2(n17380), .A3(n17379), .ZN(n17382) );
  OAI21_X1 U19325 ( .B1(n17384), .B2(n17383), .A(n17382), .ZN(n17387) );
  XOR2_X1 U19326 ( .A(DATAI_22_), .B(keyinput_10), .Z(n17386) );
  XOR2_X1 U19327 ( .A(DATAI_21_), .B(keyinput_11), .Z(n17385) );
  AOI21_X1 U19328 ( .B1(n17387), .B2(n17386), .A(n17385), .ZN(n17391) );
  XOR2_X1 U19329 ( .A(DATAI_19_), .B(keyinput_13), .Z(n17390) );
  XOR2_X1 U19330 ( .A(DATAI_18_), .B(keyinput_14), .Z(n17389) );
  XNOR2_X1 U19331 ( .A(DATAI_20_), .B(keyinput_12), .ZN(n17388) );
  NOR4_X1 U19332 ( .A1(n17391), .A2(n17390), .A3(n17389), .A4(n17388), .ZN(
        n17395) );
  XOR2_X1 U19333 ( .A(DATAI_17_), .B(keyinput_15), .Z(n17394) );
  XOR2_X1 U19334 ( .A(DATAI_16_), .B(keyinput_16), .Z(n17393) );
  XNOR2_X1 U19335 ( .A(DATAI_15_), .B(keyinput_17), .ZN(n17392) );
  NOR4_X1 U19336 ( .A1(n17395), .A2(n17394), .A3(n17393), .A4(n17392), .ZN(
        n17398) );
  XOR2_X1 U19337 ( .A(DATAI_14_), .B(keyinput_18), .Z(n17397) );
  XOR2_X1 U19338 ( .A(DATAI_13_), .B(keyinput_19), .Z(n17396) );
  OAI21_X1 U19339 ( .B1(n17398), .B2(n17397), .A(n17396), .ZN(n17404) );
  XOR2_X1 U19340 ( .A(DATAI_12_), .B(keyinput_20), .Z(n17403) );
  XOR2_X1 U19341 ( .A(DATAI_10_), .B(keyinput_22), .Z(n17401) );
  XOR2_X1 U19342 ( .A(DATAI_11_), .B(keyinput_21), .Z(n17400) );
  XOR2_X1 U19343 ( .A(DATAI_9_), .B(keyinput_23), .Z(n17399) );
  NAND3_X1 U19344 ( .A1(n17401), .A2(n17400), .A3(n17399), .ZN(n17402) );
  AOI21_X1 U19345 ( .B1(n17404), .B2(n17403), .A(n17402), .ZN(n17408) );
  XOR2_X1 U19346 ( .A(DATAI_8_), .B(keyinput_24), .Z(n17407) );
  XOR2_X1 U19347 ( .A(DATAI_7_), .B(keyinput_25), .Z(n17406) );
  XNOR2_X1 U19348 ( .A(DATAI_6_), .B(keyinput_26), .ZN(n17405) );
  NOR4_X1 U19349 ( .A1(n17408), .A2(n17407), .A3(n17406), .A4(n17405), .ZN(
        n17411) );
  XOR2_X1 U19350 ( .A(DATAI_5_), .B(keyinput_27), .Z(n17410) );
  XOR2_X1 U19351 ( .A(DATAI_4_), .B(keyinput_28), .Z(n17409) );
  NOR3_X1 U19352 ( .A1(n17411), .A2(n17410), .A3(n17409), .ZN(n17414) );
  XOR2_X1 U19353 ( .A(DATAI_3_), .B(keyinput_29), .Z(n17413) );
  XNOR2_X1 U19354 ( .A(DATAI_2_), .B(keyinput_30), .ZN(n17412) );
  OAI21_X1 U19355 ( .B1(n17414), .B2(n17413), .A(n17412), .ZN(n17417) );
  XOR2_X1 U19356 ( .A(DATAI_0_), .B(keyinput_32), .Z(n17416) );
  XNOR2_X1 U19357 ( .A(DATAI_1_), .B(keyinput_31), .ZN(n17415) );
  NAND3_X1 U19358 ( .A1(n17417), .A2(n17416), .A3(n17415), .ZN(n17421) );
  XNOR2_X1 U19359 ( .A(HOLD), .B(keyinput_33), .ZN(n17420) );
  XNOR2_X1 U19360 ( .A(NA), .B(keyinput_34), .ZN(n17419) );
  XNOR2_X1 U19361 ( .A(BS16), .B(keyinput_35), .ZN(n17418) );
  NAND4_X1 U19362 ( .A1(n17421), .A2(n17420), .A3(n17419), .A4(n17418), .ZN(
        n17430) );
  XOR2_X1 U19363 ( .A(READY1), .B(keyinput_36), .Z(n17429) );
  INV_X1 U19364 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n17829) );
  INV_X1 U19365 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n17423) );
  OAI22_X1 U19366 ( .A1(n17829), .A2(keyinput_39), .B1(n17423), .B2(
        keyinput_38), .ZN(n17422) );
  AOI221_X1 U19367 ( .B1(n17829), .B2(keyinput_39), .C1(keyinput_38), .C2(
        n17423), .A(n17422), .ZN(n17427) );
  XOR2_X1 U19368 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(keyinput_41), .Z(n17426) );
  INV_X1 U19369 ( .A(READY2), .ZN(n17607) );
  OAI22_X1 U19370 ( .A1(n17607), .A2(keyinput_37), .B1(
        P1_CODEFETCH_REG_SCAN_IN), .B2(keyinput_40), .ZN(n17424) );
  AOI221_X1 U19371 ( .B1(n17607), .B2(keyinput_37), .C1(keyinput_40), .C2(
        P1_CODEFETCH_REG_SCAN_IN), .A(n17424), .ZN(n17425) );
  NAND3_X1 U19372 ( .A1(n17427), .A2(n17426), .A3(n17425), .ZN(n17428) );
  AOI21_X1 U19373 ( .B1(n17430), .B2(n17429), .A(n17428), .ZN(n17434) );
  XNOR2_X1 U19374 ( .A(n22286), .B(keyinput_44), .ZN(n17433) );
  INV_X1 U19375 ( .A(P1_D_C_N_REG_SCAN_IN), .ZN(n20600) );
  XNOR2_X1 U19376 ( .A(n20600), .B(keyinput_42), .ZN(n17432) );
  XNOR2_X1 U19377 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .B(keyinput_43), .ZN(
        n17431) );
  NOR4_X1 U19378 ( .A1(n17434), .A2(n17433), .A3(n17432), .A4(n17431), .ZN(
        n17441) );
  XNOR2_X1 U19379 ( .A(P1_MORE_REG_SCAN_IN), .B(keyinput_45), .ZN(n17440) );
  INV_X1 U19380 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20494) );
  XNOR2_X1 U19381 ( .A(n20494), .B(keyinput_49), .ZN(n17438) );
  XNOR2_X1 U19382 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .B(keyinput_48), .ZN(
        n17437) );
  XNOR2_X1 U19383 ( .A(P1_FLUSH_REG_SCAN_IN), .B(keyinput_46), .ZN(n17436) );
  XNOR2_X1 U19384 ( .A(P1_W_R_N_REG_SCAN_IN), .B(keyinput_47), .ZN(n17435) );
  NOR4_X1 U19385 ( .A1(n17438), .A2(n17437), .A3(n17436), .A4(n17435), .ZN(
        n17439) );
  OAI21_X1 U19386 ( .B1(n17441), .B2(n17440), .A(n17439), .ZN(n17445) );
  INV_X1 U19387 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20490) );
  XNOR2_X1 U19388 ( .A(n20490), .B(keyinput_50), .ZN(n17444) );
  XNOR2_X1 U19389 ( .A(P1_REIP_REG_31__SCAN_IN), .B(keyinput_52), .ZN(n17443)
         );
  XNOR2_X1 U19390 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .B(keyinput_51), .ZN(
        n17442) );
  AOI211_X1 U19391 ( .C1(n17445), .C2(n17444), .A(n17443), .B(n17442), .ZN(
        n17449) );
  XOR2_X1 U19392 ( .A(P1_REIP_REG_30__SCAN_IN), .B(keyinput_53), .Z(n17448) );
  XOR2_X1 U19393 ( .A(P1_REIP_REG_29__SCAN_IN), .B(keyinput_54), .Z(n17447) );
  XNOR2_X1 U19394 ( .A(P1_REIP_REG_28__SCAN_IN), .B(keyinput_55), .ZN(n17446)
         );
  OAI211_X1 U19395 ( .C1(n17449), .C2(n17448), .A(n17447), .B(n17446), .ZN(
        n17453) );
  XOR2_X1 U19396 ( .A(P1_REIP_REG_25__SCAN_IN), .B(keyinput_58), .Z(n17452) );
  XNOR2_X1 U19397 ( .A(P1_REIP_REG_27__SCAN_IN), .B(keyinput_56), .ZN(n17451)
         );
  XNOR2_X1 U19398 ( .A(P1_REIP_REG_26__SCAN_IN), .B(keyinput_57), .ZN(n17450)
         );
  NAND4_X1 U19399 ( .A1(n17453), .A2(n17452), .A3(n17451), .A4(n17450), .ZN(
        n17459) );
  XNOR2_X1 U19400 ( .A(P1_REIP_REG_24__SCAN_IN), .B(keyinput_59), .ZN(n17458)
         );
  XOR2_X1 U19401 ( .A(P1_REIP_REG_22__SCAN_IN), .B(keyinput_61), .Z(n17456) );
  XNOR2_X1 U19402 ( .A(P1_REIP_REG_21__SCAN_IN), .B(keyinput_62), .ZN(n17455)
         );
  XNOR2_X1 U19403 ( .A(P1_REIP_REG_23__SCAN_IN), .B(keyinput_60), .ZN(n17454)
         );
  NAND3_X1 U19404 ( .A1(n17456), .A2(n17455), .A3(n17454), .ZN(n17457) );
  AOI21_X1 U19405 ( .B1(n17459), .B2(n17458), .A(n17457), .ZN(n17462) );
  XOR2_X1 U19406 ( .A(P1_REIP_REG_20__SCAN_IN), .B(keyinput_63), .Z(n17461) );
  XNOR2_X1 U19407 ( .A(P1_REIP_REG_19__SCAN_IN), .B(keyinput_64), .ZN(n17460)
         );
  NOR3_X1 U19408 ( .A1(n17462), .A2(n17461), .A3(n17460), .ZN(n17465) );
  XOR2_X1 U19409 ( .A(P1_REIP_REG_18__SCAN_IN), .B(keyinput_65), .Z(n17464) );
  XOR2_X1 U19410 ( .A(P1_REIP_REG_17__SCAN_IN), .B(keyinput_66), .Z(n17463) );
  NOR3_X1 U19411 ( .A1(n17465), .A2(n17464), .A3(n17463), .ZN(n17468) );
  XOR2_X1 U19412 ( .A(P1_REIP_REG_16__SCAN_IN), .B(keyinput_67), .Z(n17467) );
  XNOR2_X1 U19413 ( .A(P1_REIP_REG_15__SCAN_IN), .B(keyinput_68), .ZN(n17466)
         );
  NOR3_X1 U19414 ( .A1(n17468), .A2(n17467), .A3(n17466), .ZN(n17480) );
  XNOR2_X1 U19415 ( .A(P1_REIP_REG_14__SCAN_IN), .B(keyinput_69), .ZN(n17470)
         );
  XNOR2_X1 U19416 ( .A(P1_REIP_REG_13__SCAN_IN), .B(keyinput_70), .ZN(n17469)
         );
  NOR2_X1 U19417 ( .A1(n17470), .A2(n17469), .ZN(n17476) );
  XNOR2_X1 U19418 ( .A(P1_REIP_REG_11__SCAN_IN), .B(keyinput_72), .ZN(n17472)
         );
  XNOR2_X1 U19419 ( .A(P1_REIP_REG_10__SCAN_IN), .B(keyinput_73), .ZN(n17471)
         );
  NOR2_X1 U19420 ( .A1(n17472), .A2(n17471), .ZN(n17475) );
  XNOR2_X1 U19421 ( .A(P1_REIP_REG_9__SCAN_IN), .B(keyinput_74), .ZN(n17474)
         );
  XNOR2_X1 U19422 ( .A(P1_REIP_REG_12__SCAN_IN), .B(keyinput_71), .ZN(n17473)
         );
  NAND4_X1 U19423 ( .A1(n17476), .A2(n17475), .A3(n17474), .A4(n17473), .ZN(
        n17479) );
  XOR2_X1 U19424 ( .A(P1_REIP_REG_8__SCAN_IN), .B(keyinput_75), .Z(n17478) );
  XNOR2_X1 U19425 ( .A(P1_REIP_REG_7__SCAN_IN), .B(keyinput_76), .ZN(n17477)
         );
  OAI211_X1 U19426 ( .C1(n17480), .C2(n17479), .A(n17478), .B(n17477), .ZN(
        n17484) );
  XNOR2_X1 U19427 ( .A(n17481), .B(keyinput_77), .ZN(n17483) );
  XOR2_X1 U19428 ( .A(P1_REIP_REG_5__SCAN_IN), .B(keyinput_78), .Z(n17482) );
  AOI21_X1 U19429 ( .B1(n17484), .B2(n17483), .A(n17482), .ZN(n17487) );
  XOR2_X1 U19430 ( .A(P1_REIP_REG_3__SCAN_IN), .B(keyinput_80), .Z(n17486) );
  XNOR2_X1 U19431 ( .A(P1_REIP_REG_4__SCAN_IN), .B(keyinput_79), .ZN(n17485)
         );
  NOR3_X1 U19432 ( .A1(n17487), .A2(n17486), .A3(n17485), .ZN(n17498) );
  XOR2_X1 U19433 ( .A(P1_EBX_REG_30__SCAN_IN), .B(keyinput_85), .Z(n17490) );
  XNOR2_X1 U19434 ( .A(P1_REIP_REG_2__SCAN_IN), .B(keyinput_81), .ZN(n17489)
         );
  XNOR2_X1 U19435 ( .A(P1_REIP_REG_1__SCAN_IN), .B(keyinput_82), .ZN(n17488)
         );
  NOR3_X1 U19436 ( .A1(n17490), .A2(n17489), .A3(n17488), .ZN(n17493) );
  XOR2_X1 U19437 ( .A(P1_EBX_REG_31__SCAN_IN), .B(keyinput_84), .Z(n17492) );
  XOR2_X1 U19438 ( .A(P1_REIP_REG_0__SCAN_IN), .B(keyinput_83), .Z(n17491) );
  NAND3_X1 U19439 ( .A1(n17493), .A2(n17492), .A3(n17491), .ZN(n17497) );
  XNOR2_X1 U19440 ( .A(n17494), .B(keyinput_87), .ZN(n17496) );
  XNOR2_X1 U19441 ( .A(P1_EBX_REG_29__SCAN_IN), .B(keyinput_86), .ZN(n17495)
         );
  OAI211_X1 U19442 ( .C1(n17498), .C2(n17497), .A(n17496), .B(n17495), .ZN(
        n17502) );
  XNOR2_X1 U19443 ( .A(P1_EBX_REG_27__SCAN_IN), .B(keyinput_88), .ZN(n17501)
         );
  XOR2_X1 U19444 ( .A(P1_EBX_REG_25__SCAN_IN), .B(keyinput_90), .Z(n17500) );
  XNOR2_X1 U19445 ( .A(P1_EBX_REG_26__SCAN_IN), .B(keyinput_89), .ZN(n17499)
         );
  AOI211_X1 U19446 ( .C1(n17502), .C2(n17501), .A(n17500), .B(n17499), .ZN(
        n17505) );
  XOR2_X1 U19447 ( .A(P1_EBX_REG_24__SCAN_IN), .B(keyinput_91), .Z(n17504) );
  XOR2_X1 U19448 ( .A(P1_EBX_REG_23__SCAN_IN), .B(keyinput_92), .Z(n17503) );
  OAI21_X1 U19449 ( .B1(n17505), .B2(n17504), .A(n17503), .ZN(n17512) );
  XOR2_X1 U19450 ( .A(P1_EBX_REG_22__SCAN_IN), .B(keyinput_93), .Z(n17511) );
  XOR2_X1 U19451 ( .A(P1_EBX_REG_18__SCAN_IN), .B(keyinput_97), .Z(n17509) );
  XOR2_X1 U19452 ( .A(P1_EBX_REG_20__SCAN_IN), .B(keyinput_95), .Z(n17508) );
  XOR2_X1 U19453 ( .A(P1_EBX_REG_19__SCAN_IN), .B(keyinput_96), .Z(n17507) );
  XNOR2_X1 U19454 ( .A(P1_EBX_REG_21__SCAN_IN), .B(keyinput_94), .ZN(n17506)
         );
  NAND4_X1 U19455 ( .A1(n17509), .A2(n17508), .A3(n17507), .A4(n17506), .ZN(
        n17510) );
  AOI21_X1 U19456 ( .B1(n17512), .B2(n17511), .A(n17510), .ZN(n17515) );
  XOR2_X1 U19457 ( .A(P1_EBX_REG_17__SCAN_IN), .B(keyinput_98), .Z(n17514) );
  XNOR2_X1 U19458 ( .A(P1_EBX_REG_16__SCAN_IN), .B(keyinput_99), .ZN(n17513)
         );
  NOR3_X1 U19459 ( .A1(n17515), .A2(n17514), .A3(n17513), .ZN(n17521) );
  XOR2_X1 U19460 ( .A(P1_EBX_REG_15__SCAN_IN), .B(keyinput_100), .Z(n17520) );
  XOR2_X1 U19461 ( .A(P1_EBX_REG_13__SCAN_IN), .B(keyinput_102), .Z(n17518) );
  XOR2_X1 U19462 ( .A(P1_EBX_REG_14__SCAN_IN), .B(keyinput_101), .Z(n17517) );
  XNOR2_X1 U19463 ( .A(P1_EBX_REG_12__SCAN_IN), .B(keyinput_103), .ZN(n17516)
         );
  NOR3_X1 U19464 ( .A1(n17518), .A2(n17517), .A3(n17516), .ZN(n17519) );
  OAI21_X1 U19465 ( .B1(n17521), .B2(n17520), .A(n17519), .ZN(n17524) );
  XNOR2_X1 U19466 ( .A(P1_EBX_REG_11__SCAN_IN), .B(keyinput_104), .ZN(n17523)
         );
  XOR2_X1 U19467 ( .A(P1_EBX_REG_10__SCAN_IN), .B(keyinput_105), .Z(n17522) );
  AOI21_X1 U19468 ( .B1(n17524), .B2(n17523), .A(n17522), .ZN(n17527) );
  XNOR2_X1 U19469 ( .A(P1_EBX_REG_9__SCAN_IN), .B(keyinput_106), .ZN(n17526)
         );
  XNOR2_X1 U19470 ( .A(P1_EBX_REG_8__SCAN_IN), .B(keyinput_107), .ZN(n17525)
         );
  OAI21_X1 U19471 ( .B1(n17527), .B2(n17526), .A(n17525), .ZN(n17530) );
  XOR2_X1 U19472 ( .A(P1_EBX_REG_7__SCAN_IN), .B(keyinput_108), .Z(n17529) );
  XNOR2_X1 U19473 ( .A(P1_EBX_REG_6__SCAN_IN), .B(keyinput_109), .ZN(n17528)
         );
  AOI21_X1 U19474 ( .B1(n17530), .B2(n17529), .A(n17528), .ZN(n17533) );
  XOR2_X1 U19475 ( .A(P1_EBX_REG_5__SCAN_IN), .B(keyinput_110), .Z(n17532) );
  XNOR2_X1 U19476 ( .A(P1_EBX_REG_4__SCAN_IN), .B(keyinput_111), .ZN(n17531)
         );
  NOR3_X1 U19477 ( .A1(n17533), .A2(n17532), .A3(n17531), .ZN(n17539) );
  XNOR2_X1 U19478 ( .A(P1_EBX_REG_3__SCAN_IN), .B(keyinput_112), .ZN(n17538)
         );
  XOR2_X1 U19479 ( .A(P1_EBX_REG_2__SCAN_IN), .B(keyinput_113), .Z(n17536) );
  XNOR2_X1 U19480 ( .A(P1_EBX_REG_0__SCAN_IN), .B(keyinput_115), .ZN(n17535)
         );
  XNOR2_X1 U19481 ( .A(P1_EBX_REG_1__SCAN_IN), .B(keyinput_114), .ZN(n17534)
         );
  NOR3_X1 U19482 ( .A1(n17536), .A2(n17535), .A3(n17534), .ZN(n17537) );
  OAI21_X1 U19483 ( .B1(n17539), .B2(n17538), .A(n17537), .ZN(n17542) );
  XNOR2_X1 U19484 ( .A(P1_EAX_REG_30__SCAN_IN), .B(keyinput_117), .ZN(n17541)
         );
  XNOR2_X1 U19485 ( .A(P1_EAX_REG_31__SCAN_IN), .B(keyinput_116), .ZN(n17540)
         );
  NAND3_X1 U19486 ( .A1(n17542), .A2(n17541), .A3(n17540), .ZN(n17545) );
  XNOR2_X1 U19487 ( .A(P1_EAX_REG_29__SCAN_IN), .B(keyinput_118), .ZN(n17544)
         );
  XOR2_X1 U19488 ( .A(P1_EAX_REG_28__SCAN_IN), .B(keyinput_119), .Z(n17543) );
  AOI21_X1 U19489 ( .B1(n17545), .B2(n17544), .A(n17543), .ZN(n17555) );
  XOR2_X1 U19490 ( .A(P1_EAX_REG_27__SCAN_IN), .B(keyinput_120), .Z(n17549) );
  XOR2_X1 U19491 ( .A(P1_EAX_REG_24__SCAN_IN), .B(keyinput_123), .Z(n17548) );
  XNOR2_X1 U19492 ( .A(P1_EAX_REG_25__SCAN_IN), .B(keyinput_122), .ZN(n17547)
         );
  XNOR2_X1 U19493 ( .A(P1_EAX_REG_26__SCAN_IN), .B(keyinput_121), .ZN(n17546)
         );
  NAND4_X1 U19494 ( .A1(n17549), .A2(n17548), .A3(n17547), .A4(n17546), .ZN(
        n17554) );
  XOR2_X1 U19495 ( .A(P1_EAX_REG_21__SCAN_IN), .B(keyinput_126), .Z(n17552) );
  XOR2_X1 U19496 ( .A(P1_EAX_REG_22__SCAN_IN), .B(keyinput_125), .Z(n17551) );
  XNOR2_X1 U19497 ( .A(P1_EAX_REG_23__SCAN_IN), .B(keyinput_124), .ZN(n17550)
         );
  NOR3_X1 U19498 ( .A1(n17552), .A2(n17551), .A3(n17550), .ZN(n17553) );
  OAI21_X1 U19499 ( .B1(n17555), .B2(n17554), .A(n17553), .ZN(n17744) );
  XOR2_X1 U19500 ( .A(keyinput_255), .B(keyinput_127), .Z(n17743) );
  XOR2_X1 U19501 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(keyinput_128), .Z(n17559) );
  XNOR2_X1 U19502 ( .A(n15086), .B(keyinput_129), .ZN(n17558) );
  XNOR2_X1 U19503 ( .A(DATAI_29_), .B(keyinput_131), .ZN(n17557) );
  XNOR2_X1 U19504 ( .A(DATAI_30_), .B(keyinput_130), .ZN(n17556) );
  NAND4_X1 U19505 ( .A1(n17559), .A2(n17558), .A3(n17557), .A4(n17556), .ZN(
        n17562) );
  XOR2_X1 U19506 ( .A(DATAI_28_), .B(keyinput_132), .Z(n17561) );
  XOR2_X1 U19507 ( .A(DATAI_27_), .B(keyinput_133), .Z(n17560) );
  NAND3_X1 U19508 ( .A1(n17562), .A2(n17561), .A3(n17560), .ZN(n17568) );
  XOR2_X1 U19509 ( .A(DATAI_26_), .B(keyinput_134), .Z(n17567) );
  XOR2_X1 U19510 ( .A(DATAI_24_), .B(keyinput_136), .Z(n17565) );
  XNOR2_X1 U19511 ( .A(DATAI_25_), .B(keyinput_135), .ZN(n17564) );
  XNOR2_X1 U19512 ( .A(DATAI_23_), .B(keyinput_137), .ZN(n17563) );
  NAND3_X1 U19513 ( .A1(n17565), .A2(n17564), .A3(n17563), .ZN(n17566) );
  AOI21_X1 U19514 ( .B1(n17568), .B2(n17567), .A(n17566), .ZN(n17571) );
  XNOR2_X1 U19515 ( .A(DATAI_22_), .B(keyinput_138), .ZN(n17570) );
  XNOR2_X1 U19516 ( .A(DATAI_21_), .B(keyinput_139), .ZN(n17569) );
  OAI21_X1 U19517 ( .B1(n17571), .B2(n17570), .A(n17569), .ZN(n17575) );
  XOR2_X1 U19518 ( .A(DATAI_20_), .B(keyinput_140), .Z(n17574) );
  XOR2_X1 U19519 ( .A(DATAI_19_), .B(keyinput_141), .Z(n17573) );
  XNOR2_X1 U19520 ( .A(DATAI_18_), .B(keyinput_142), .ZN(n17572) );
  NAND4_X1 U19521 ( .A1(n17575), .A2(n17574), .A3(n17573), .A4(n17572), .ZN(
        n17579) );
  XOR2_X1 U19522 ( .A(DATAI_16_), .B(keyinput_144), .Z(n17578) );
  XOR2_X1 U19523 ( .A(DATAI_17_), .B(keyinput_143), .Z(n17577) );
  XNOR2_X1 U19524 ( .A(DATAI_15_), .B(keyinput_145), .ZN(n17576) );
  NAND4_X1 U19525 ( .A1(n17579), .A2(n17578), .A3(n17577), .A4(n17576), .ZN(
        n17582) );
  XNOR2_X1 U19526 ( .A(DATAI_14_), .B(keyinput_146), .ZN(n17581) );
  XNOR2_X1 U19527 ( .A(DATAI_13_), .B(keyinput_147), .ZN(n17580) );
  AOI21_X1 U19528 ( .B1(n17582), .B2(n17581), .A(n17580), .ZN(n17588) );
  XNOR2_X1 U19529 ( .A(DATAI_12_), .B(keyinput_148), .ZN(n17587) );
  XOR2_X1 U19530 ( .A(DATAI_11_), .B(keyinput_149), .Z(n17585) );
  XNOR2_X1 U19531 ( .A(DATAI_9_), .B(keyinput_151), .ZN(n17584) );
  XNOR2_X1 U19532 ( .A(DATAI_10_), .B(keyinput_150), .ZN(n17583) );
  NOR3_X1 U19533 ( .A1(n17585), .A2(n17584), .A3(n17583), .ZN(n17586) );
  OAI21_X1 U19534 ( .B1(n17588), .B2(n17587), .A(n17586), .ZN(n17592) );
  XOR2_X1 U19535 ( .A(DATAI_7_), .B(keyinput_153), .Z(n17591) );
  XOR2_X1 U19536 ( .A(DATAI_8_), .B(keyinput_152), .Z(n17590) );
  XNOR2_X1 U19537 ( .A(DATAI_6_), .B(keyinput_154), .ZN(n17589) );
  NAND4_X1 U19538 ( .A1(n17592), .A2(n17591), .A3(n17590), .A4(n17589), .ZN(
        n17595) );
  XOR2_X1 U19539 ( .A(DATAI_4_), .B(keyinput_156), .Z(n17594) );
  XNOR2_X1 U19540 ( .A(DATAI_5_), .B(keyinput_155), .ZN(n17593) );
  NAND3_X1 U19541 ( .A1(n17595), .A2(n17594), .A3(n17593), .ZN(n17598) );
  XOR2_X1 U19542 ( .A(DATAI_3_), .B(keyinput_157), .Z(n17597) );
  XNOR2_X1 U19543 ( .A(DATAI_2_), .B(keyinput_158), .ZN(n17596) );
  AOI21_X1 U19544 ( .B1(n17598), .B2(n17597), .A(n17596), .ZN(n17601) );
  XNOR2_X1 U19545 ( .A(DATAI_0_), .B(keyinput_160), .ZN(n17600) );
  XNOR2_X1 U19546 ( .A(DATAI_1_), .B(keyinput_159), .ZN(n17599) );
  NOR3_X1 U19547 ( .A1(n17601), .A2(n17600), .A3(n17599), .ZN(n17605) );
  XOR2_X1 U19548 ( .A(HOLD), .B(keyinput_161), .Z(n17604) );
  INV_X1 U19549 ( .A(BS16), .ZN(n17763) );
  XNOR2_X1 U19550 ( .A(n17763), .B(keyinput_163), .ZN(n17603) );
  XNOR2_X1 U19551 ( .A(NA), .B(keyinput_162), .ZN(n17602) );
  NOR4_X1 U19552 ( .A1(n17605), .A2(n17604), .A3(n17603), .A4(n17602), .ZN(
        n17615) );
  XOR2_X1 U19553 ( .A(READY1), .B(keyinput_164), .Z(n17614) );
  AOI22_X1 U19554 ( .A1(n17829), .A2(keyinput_167), .B1(keyinput_165), .B2(
        n17607), .ZN(n17606) );
  OAI221_X1 U19555 ( .B1(n17829), .B2(keyinput_167), .C1(n17607), .C2(
        keyinput_165), .A(n17606), .ZN(n17612) );
  INV_X1 U19556 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n17609) );
  AOI22_X1 U19557 ( .A1(P1_READREQUEST_REG_SCAN_IN), .A2(keyinput_166), .B1(
        n17609), .B2(keyinput_168), .ZN(n17608) );
  OAI221_X1 U19558 ( .B1(P1_READREQUEST_REG_SCAN_IN), .B2(keyinput_166), .C1(
        n17609), .C2(keyinput_168), .A(n17608), .ZN(n17611) );
  XNOR2_X1 U19559 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(keyinput_169), .ZN(n17610)
         );
  NOR3_X1 U19560 ( .A1(n17612), .A2(n17611), .A3(n17610), .ZN(n17613) );
  OAI21_X1 U19561 ( .B1(n17615), .B2(n17614), .A(n17613), .ZN(n17619) );
  XNOR2_X1 U19562 ( .A(n22286), .B(keyinput_172), .ZN(n17618) );
  XNOR2_X1 U19563 ( .A(n20600), .B(keyinput_170), .ZN(n17617) );
  XNOR2_X1 U19564 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .B(keyinput_171), .ZN(
        n17616) );
  NAND4_X1 U19565 ( .A1(n17619), .A2(n17618), .A3(n17617), .A4(n17616), .ZN(
        n17627) );
  XNOR2_X1 U19566 ( .A(P1_MORE_REG_SCAN_IN), .B(keyinput_173), .ZN(n17626) );
  INV_X1 U19567 ( .A(keyinput_174), .ZN(n17620) );
  XNOR2_X1 U19568 ( .A(n17620), .B(P1_FLUSH_REG_SCAN_IN), .ZN(n17624) );
  XNOR2_X1 U19569 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .B(keyinput_176), .ZN(
        n17623) );
  XNOR2_X1 U19570 ( .A(P1_W_R_N_REG_SCAN_IN), .B(keyinput_175), .ZN(n17622) );
  XNOR2_X1 U19571 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .B(keyinput_177), .ZN(
        n17621) );
  NAND4_X1 U19572 ( .A1(n17624), .A2(n17623), .A3(n17622), .A4(n17621), .ZN(
        n17625) );
  AOI21_X1 U19573 ( .B1(n17627), .B2(n17626), .A(n17625), .ZN(n17632) );
  XNOR2_X1 U19574 ( .A(n20490), .B(keyinput_178), .ZN(n17631) );
  XNOR2_X1 U19575 ( .A(n17628), .B(keyinput_180), .ZN(n17630) );
  XNOR2_X1 U19576 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .B(keyinput_179), .ZN(
        n17629) );
  OAI211_X1 U19577 ( .C1(n17632), .C2(n17631), .A(n17630), .B(n17629), .ZN(
        n17636) );
  XOR2_X1 U19578 ( .A(P1_REIP_REG_30__SCAN_IN), .B(keyinput_181), .Z(n17635)
         );
  XOR2_X1 U19579 ( .A(P1_REIP_REG_29__SCAN_IN), .B(keyinput_182), .Z(n17634)
         );
  XNOR2_X1 U19580 ( .A(P1_REIP_REG_28__SCAN_IN), .B(keyinput_183), .ZN(n17633)
         );
  AOI211_X1 U19581 ( .C1(n17636), .C2(n17635), .A(n17634), .B(n17633), .ZN(
        n17640) );
  XOR2_X1 U19582 ( .A(P1_REIP_REG_25__SCAN_IN), .B(keyinput_186), .Z(n17639)
         );
  XNOR2_X1 U19583 ( .A(P1_REIP_REG_26__SCAN_IN), .B(keyinput_185), .ZN(n17638)
         );
  XNOR2_X1 U19584 ( .A(P1_REIP_REG_27__SCAN_IN), .B(keyinput_184), .ZN(n17637)
         );
  NOR4_X1 U19585 ( .A1(n17640), .A2(n17639), .A3(n17638), .A4(n17637), .ZN(
        n17642) );
  XOR2_X1 U19586 ( .A(P1_REIP_REG_24__SCAN_IN), .B(keyinput_187), .Z(n17641)
         );
  NOR2_X1 U19587 ( .A1(n17642), .A2(n17641), .ZN(n17646) );
  XOR2_X1 U19588 ( .A(P1_REIP_REG_22__SCAN_IN), .B(keyinput_189), .Z(n17645)
         );
  XNOR2_X1 U19589 ( .A(P1_REIP_REG_23__SCAN_IN), .B(keyinput_188), .ZN(n17644)
         );
  XNOR2_X1 U19590 ( .A(P1_REIP_REG_21__SCAN_IN), .B(keyinput_190), .ZN(n17643)
         );
  NOR4_X1 U19591 ( .A1(n17646), .A2(n17645), .A3(n17644), .A4(n17643), .ZN(
        n17649) );
  XOR2_X1 U19592 ( .A(P1_REIP_REG_20__SCAN_IN), .B(keyinput_191), .Z(n17648)
         );
  XOR2_X1 U19593 ( .A(P1_REIP_REG_19__SCAN_IN), .B(keyinput_192), .Z(n17647)
         );
  NOR3_X1 U19594 ( .A1(n17649), .A2(n17648), .A3(n17647), .ZN(n17652) );
  XOR2_X1 U19595 ( .A(P1_REIP_REG_18__SCAN_IN), .B(keyinput_193), .Z(n17651)
         );
  XNOR2_X1 U19596 ( .A(P1_REIP_REG_17__SCAN_IN), .B(keyinput_194), .ZN(n17650)
         );
  NOR3_X1 U19597 ( .A1(n17652), .A2(n17651), .A3(n17650), .ZN(n17655) );
  XOR2_X1 U19598 ( .A(P1_REIP_REG_16__SCAN_IN), .B(keyinput_195), .Z(n17654)
         );
  XOR2_X1 U19599 ( .A(P1_REIP_REG_15__SCAN_IN), .B(keyinput_196), .Z(n17653)
         );
  NOR3_X1 U19600 ( .A1(n17655), .A2(n17654), .A3(n17653), .ZN(n17664) );
  XNOR2_X1 U19601 ( .A(n17656), .B(keyinput_198), .ZN(n17663) );
  XNOR2_X1 U19602 ( .A(P1_REIP_REG_12__SCAN_IN), .B(keyinput_199), .ZN(n17662)
         );
  XNOR2_X1 U19603 ( .A(P1_REIP_REG_9__SCAN_IN), .B(keyinput_202), .ZN(n17660)
         );
  XNOR2_X1 U19604 ( .A(P1_REIP_REG_11__SCAN_IN), .B(keyinput_200), .ZN(n17659)
         );
  XNOR2_X1 U19605 ( .A(P1_REIP_REG_10__SCAN_IN), .B(keyinput_201), .ZN(n17658)
         );
  XNOR2_X1 U19606 ( .A(P1_REIP_REG_14__SCAN_IN), .B(keyinput_197), .ZN(n17657)
         );
  NAND4_X1 U19607 ( .A1(n17660), .A2(n17659), .A3(n17658), .A4(n17657), .ZN(
        n17661) );
  NOR4_X1 U19608 ( .A1(n17664), .A2(n17663), .A3(n17662), .A4(n17661), .ZN(
        n17669) );
  XOR2_X1 U19609 ( .A(P1_REIP_REG_8__SCAN_IN), .B(keyinput_203), .Z(n17666) );
  XNOR2_X1 U19610 ( .A(P1_REIP_REG_7__SCAN_IN), .B(keyinput_204), .ZN(n17665)
         );
  NAND2_X1 U19611 ( .A1(n17666), .A2(n17665), .ZN(n17668) );
  XNOR2_X1 U19612 ( .A(P1_REIP_REG_6__SCAN_IN), .B(keyinput_205), .ZN(n17667)
         );
  OAI21_X1 U19613 ( .B1(n17669), .B2(n17668), .A(n17667), .ZN(n17673) );
  XNOR2_X1 U19614 ( .A(P1_REIP_REG_5__SCAN_IN), .B(keyinput_206), .ZN(n17672)
         );
  XOR2_X1 U19615 ( .A(P1_REIP_REG_3__SCAN_IN), .B(keyinput_208), .Z(n17671) );
  XOR2_X1 U19616 ( .A(P1_REIP_REG_4__SCAN_IN), .B(keyinput_207), .Z(n17670) );
  AOI211_X1 U19617 ( .C1(n17673), .C2(n17672), .A(n17671), .B(n17670), .ZN(
        n17680) );
  XNOR2_X1 U19618 ( .A(P1_REIP_REG_2__SCAN_IN), .B(keyinput_209), .ZN(n17679)
         );
  XNOR2_X1 U19619 ( .A(P1_REIP_REG_1__SCAN_IN), .B(keyinput_210), .ZN(n17678)
         );
  XOR2_X1 U19620 ( .A(P1_EBX_REG_31__SCAN_IN), .B(keyinput_212), .Z(n17676) );
  XNOR2_X1 U19621 ( .A(P1_REIP_REG_0__SCAN_IN), .B(keyinput_211), .ZN(n17675)
         );
  XNOR2_X1 U19622 ( .A(P1_EBX_REG_30__SCAN_IN), .B(keyinput_213), .ZN(n17674)
         );
  NAND3_X1 U19623 ( .A1(n17676), .A2(n17675), .A3(n17674), .ZN(n17677) );
  NOR4_X1 U19624 ( .A1(n17680), .A2(n17679), .A3(n17678), .A4(n17677), .ZN(
        n17683) );
  XOR2_X1 U19625 ( .A(P1_EBX_REG_29__SCAN_IN), .B(keyinput_214), .Z(n17682) );
  XNOR2_X1 U19626 ( .A(P1_EBX_REG_28__SCAN_IN), .B(keyinput_215), .ZN(n17681)
         );
  NOR3_X1 U19627 ( .A1(n17683), .A2(n17682), .A3(n17681), .ZN(n17687) );
  XOR2_X1 U19628 ( .A(P1_EBX_REG_27__SCAN_IN), .B(keyinput_216), .Z(n17686) );
  XOR2_X1 U19629 ( .A(P1_EBX_REG_25__SCAN_IN), .B(keyinput_218), .Z(n17685) );
  XNOR2_X1 U19630 ( .A(P1_EBX_REG_26__SCAN_IN), .B(keyinput_217), .ZN(n17684)
         );
  OAI211_X1 U19631 ( .C1(n17687), .C2(n17686), .A(n17685), .B(n17684), .ZN(
        n17690) );
  XOR2_X1 U19632 ( .A(P1_EBX_REG_24__SCAN_IN), .B(keyinput_219), .Z(n17689) );
  XNOR2_X1 U19633 ( .A(P1_EBX_REG_23__SCAN_IN), .B(keyinput_220), .ZN(n17688)
         );
  AOI21_X1 U19634 ( .B1(n17690), .B2(n17689), .A(n17688), .ZN(n17697) );
  XOR2_X1 U19635 ( .A(P1_EBX_REG_22__SCAN_IN), .B(keyinput_221), .Z(n17696) );
  XOR2_X1 U19636 ( .A(P1_EBX_REG_19__SCAN_IN), .B(keyinput_224), .Z(n17694) );
  XOR2_X1 U19637 ( .A(P1_EBX_REG_18__SCAN_IN), .B(keyinput_225), .Z(n17693) );
  XNOR2_X1 U19638 ( .A(n20518), .B(keyinput_222), .ZN(n17692) );
  XNOR2_X1 U19639 ( .A(P1_EBX_REG_20__SCAN_IN), .B(keyinput_223), .ZN(n17691)
         );
  NOR4_X1 U19640 ( .A1(n17694), .A2(n17693), .A3(n17692), .A4(n17691), .ZN(
        n17695) );
  OAI21_X1 U19641 ( .B1(n17697), .B2(n17696), .A(n17695), .ZN(n17700) );
  XOR2_X1 U19642 ( .A(P1_EBX_REG_16__SCAN_IN), .B(keyinput_227), .Z(n17699) );
  XOR2_X1 U19643 ( .A(P1_EBX_REG_17__SCAN_IN), .B(keyinput_226), .Z(n17698) );
  NAND3_X1 U19644 ( .A1(n17700), .A2(n17699), .A3(n17698), .ZN(n17706) );
  XNOR2_X1 U19645 ( .A(P1_EBX_REG_15__SCAN_IN), .B(keyinput_228), .ZN(n17705)
         );
  XNOR2_X1 U19646 ( .A(P1_EBX_REG_14__SCAN_IN), .B(keyinput_229), .ZN(n17703)
         );
  XNOR2_X1 U19647 ( .A(P1_EBX_REG_12__SCAN_IN), .B(keyinput_231), .ZN(n17702)
         );
  XNOR2_X1 U19648 ( .A(P1_EBX_REG_13__SCAN_IN), .B(keyinput_230), .ZN(n17701)
         );
  NAND3_X1 U19649 ( .A1(n17703), .A2(n17702), .A3(n17701), .ZN(n17704) );
  AOI21_X1 U19650 ( .B1(n17706), .B2(n17705), .A(n17704), .ZN(n17709) );
  XOR2_X1 U19651 ( .A(P1_EBX_REG_11__SCAN_IN), .B(keyinput_232), .Z(n17708) );
  XOR2_X1 U19652 ( .A(P1_EBX_REG_10__SCAN_IN), .B(keyinput_233), .Z(n17707) );
  OAI21_X1 U19653 ( .B1(n17709), .B2(n17708), .A(n17707), .ZN(n17712) );
  XNOR2_X1 U19654 ( .A(P1_EBX_REG_9__SCAN_IN), .B(keyinput_234), .ZN(n17711)
         );
  XOR2_X1 U19655 ( .A(P1_EBX_REG_8__SCAN_IN), .B(keyinput_235), .Z(n17710) );
  AOI21_X1 U19656 ( .B1(n17712), .B2(n17711), .A(n17710), .ZN(n17715) );
  XOR2_X1 U19657 ( .A(P1_EBX_REG_7__SCAN_IN), .B(keyinput_236), .Z(n17714) );
  XNOR2_X1 U19658 ( .A(P1_EBX_REG_6__SCAN_IN), .B(keyinput_237), .ZN(n17713)
         );
  OAI21_X1 U19659 ( .B1(n17715), .B2(n17714), .A(n17713), .ZN(n17718) );
  XOR2_X1 U19660 ( .A(P1_EBX_REG_4__SCAN_IN), .B(keyinput_239), .Z(n17717) );
  XNOR2_X1 U19661 ( .A(P1_EBX_REG_5__SCAN_IN), .B(keyinput_238), .ZN(n17716)
         );
  NAND3_X1 U19662 ( .A1(n17718), .A2(n17717), .A3(n17716), .ZN(n17724) );
  XNOR2_X1 U19663 ( .A(P1_EBX_REG_3__SCAN_IN), .B(keyinput_240), .ZN(n17723)
         );
  XOR2_X1 U19664 ( .A(P1_EBX_REG_1__SCAN_IN), .B(keyinput_242), .Z(n17721) );
  XOR2_X1 U19665 ( .A(P1_EBX_REG_0__SCAN_IN), .B(keyinput_243), .Z(n17720) );
  XOR2_X1 U19666 ( .A(P1_EBX_REG_2__SCAN_IN), .B(keyinput_241), .Z(n17719) );
  NAND3_X1 U19667 ( .A1(n17721), .A2(n17720), .A3(n17719), .ZN(n17722) );
  AOI21_X1 U19668 ( .B1(n17724), .B2(n17723), .A(n17722), .ZN(n17727) );
  XOR2_X1 U19669 ( .A(P1_EAX_REG_30__SCAN_IN), .B(keyinput_245), .Z(n17726) );
  XOR2_X1 U19670 ( .A(P1_EAX_REG_31__SCAN_IN), .B(keyinput_244), .Z(n17725) );
  NOR3_X1 U19671 ( .A1(n17727), .A2(n17726), .A3(n17725), .ZN(n17730) );
  XNOR2_X1 U19672 ( .A(P1_EAX_REG_29__SCAN_IN), .B(keyinput_246), .ZN(n17729)
         );
  XNOR2_X1 U19673 ( .A(P1_EAX_REG_28__SCAN_IN), .B(keyinput_247), .ZN(n17728)
         );
  OAI21_X1 U19674 ( .B1(n17730), .B2(n17729), .A(n17728), .ZN(n17740) );
  XOR2_X1 U19675 ( .A(P1_EAX_REG_24__SCAN_IN), .B(keyinput_251), .Z(n17734) );
  XNOR2_X1 U19676 ( .A(P1_EAX_REG_26__SCAN_IN), .B(keyinput_249), .ZN(n17733)
         );
  XNOR2_X1 U19677 ( .A(P1_EAX_REG_27__SCAN_IN), .B(keyinput_248), .ZN(n17732)
         );
  XNOR2_X1 U19678 ( .A(P1_EAX_REG_25__SCAN_IN), .B(keyinput_250), .ZN(n17731)
         );
  NOR4_X1 U19679 ( .A1(n17734), .A2(n17733), .A3(n17732), .A4(n17731), .ZN(
        n17739) );
  XOR2_X1 U19680 ( .A(P1_EAX_REG_22__SCAN_IN), .B(keyinput_253), .Z(n17737) );
  XOR2_X1 U19681 ( .A(P1_EAX_REG_23__SCAN_IN), .B(keyinput_252), .Z(n17736) );
  XOR2_X1 U19682 ( .A(P1_EAX_REG_21__SCAN_IN), .B(keyinput_254), .Z(n17735) );
  NAND3_X1 U19683 ( .A1(n17737), .A2(n17736), .A3(n17735), .ZN(n17738) );
  AOI21_X1 U19684 ( .B1(n17740), .B2(n17739), .A(n17738), .ZN(n17742) );
  XNOR2_X1 U19685 ( .A(P1_EAX_REG_20__SCAN_IN), .B(keyinput_255), .ZN(n17741)
         );
  AOI211_X1 U19686 ( .C1(n17744), .C2(n17743), .A(n17742), .B(n17741), .ZN(
        n17745) );
  XOR2_X1 U19687 ( .A(n17746), .B(n17745), .Z(P3_U3290) );
  NAND2_X1 U19688 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19337) );
  NOR2_X1 U19689 ( .A1(n21354), .A2(n22296), .ZN(n18626) );
  NOR2_X1 U19690 ( .A1(n18626), .A2(n20674), .ZN(n17749) );
  NOR2_X1 U19691 ( .A1(n21855), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18373) );
  INV_X1 U19692 ( .A(n18373), .ZN(n19318) );
  NAND3_X1 U19693 ( .A1(n11190), .A2(n17747), .A3(n21820), .ZN(n18372) );
  NOR2_X1 U19694 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18372), .ZN(n17748) );
  INV_X1 U19695 ( .A(n17753), .ZN(n21853) );
  OAI21_X1 U19696 ( .B1(n17748), .B2(n21853), .A(n19552), .ZN(n18375) );
  NAND2_X1 U19697 ( .A1(n19318), .A2(n18375), .ZN(n18762) );
  AOI221_X1 U19698 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n19337), .C1(n17749), 
        .C2(n19337), .A(n18762), .ZN(n18761) );
  NOR2_X1 U19699 ( .A1(n21855), .A2(n21825), .ZN(n19322) );
  OAI21_X1 U19700 ( .B1(n17749), .B2(n19322), .A(n18375), .ZN(n18764) );
  INV_X1 U19701 ( .A(n18764), .ZN(n17750) );
  AOI22_X1 U19702 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n17750), .B1(
        n19355), .B2(n18375), .ZN(n18760) );
  AOI22_X1 U19703 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18761), .B1(
        n18760), .B2(n21834), .ZN(P3_U2865) );
  INV_X1 U19704 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n22346) );
  OAI21_X1 U19705 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(n22346), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n18827) );
  INV_X1 U19706 ( .A(n17752), .ZN(n22299) );
  NOR2_X1 U19707 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(P3_STATE_REG_0__SCAN_IN), 
        .ZN(n22340) );
  OAI21_X1 U19708 ( .B1(BS16), .B2(n22340), .A(n22299), .ZN(n22297) );
  OAI21_X1 U19709 ( .B1(P3_DATAWIDTH_REG_0__SCAN_IN), .B2(n22299), .A(n22297), 
        .ZN(n17751) );
  INV_X1 U19710 ( .A(n17751), .ZN(P3_U3280) );
  AND2_X1 U19711 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n17752), .ZN(P3_U3028) );
  AND2_X1 U19712 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n17752), .ZN(P3_U3027) );
  AND2_X1 U19713 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n17752), .ZN(P3_U3026) );
  AND2_X1 U19714 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n17752), .ZN(P3_U3025) );
  AND2_X1 U19715 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n17752), .ZN(P3_U3024) );
  AND2_X1 U19716 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n17752), .ZN(P3_U3023) );
  AND2_X1 U19717 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n17752), .ZN(P3_U3022) );
  AND2_X1 U19718 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n17752), .ZN(P3_U3021) );
  AND2_X1 U19719 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n17752), .ZN(
        P3_U3020) );
  AND2_X1 U19720 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n17752), .ZN(
        P3_U3019) );
  AND2_X1 U19721 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n17752), .ZN(
        P3_U3018) );
  AND2_X1 U19722 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n17752), .ZN(
        P3_U3017) );
  AND2_X1 U19723 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n17752), .ZN(
        P3_U3016) );
  AND2_X1 U19724 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n17752), .ZN(
        P3_U3015) );
  AND2_X1 U19725 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n17752), .ZN(
        P3_U3014) );
  AND2_X1 U19726 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n17752), .ZN(
        P3_U3013) );
  AND2_X1 U19727 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n17752), .ZN(
        P3_U3012) );
  AND2_X1 U19728 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n17752), .ZN(
        P3_U3011) );
  AND2_X1 U19729 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n17752), .ZN(
        P3_U3010) );
  AND2_X1 U19730 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n17752), .ZN(
        P3_U3009) );
  AND2_X1 U19731 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n17752), .ZN(
        P3_U3008) );
  AND2_X1 U19732 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n17752), .ZN(
        P3_U3007) );
  AND2_X1 U19733 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n17752), .ZN(
        P3_U3006) );
  AND2_X1 U19734 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n17752), .ZN(
        P3_U3005) );
  AND2_X1 U19735 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n17752), .ZN(
        P3_U3004) );
  AND2_X1 U19736 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n17752), .ZN(
        P3_U3003) );
  AND2_X1 U19737 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n17752), .ZN(
        P3_U3002) );
  AND2_X1 U19738 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n17752), .ZN(
        P3_U3001) );
  AND2_X1 U19739 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n17752), .ZN(
        P3_U3000) );
  AND2_X1 U19740 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n17752), .ZN(
        P3_U2999) );
  INV_X1 U19741 ( .A(n18626), .ZN(n18715) );
  AOI21_X1 U19742 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n17754)
         );
  NOR4_X1 U19743 ( .A1(n21354), .A2(n21862), .A3(n22352), .A4(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n21806) );
  AOI211_X1 U19744 ( .C1(n18715), .C2(n17754), .A(n17753), .B(n21806), .ZN(
        P3_U2998) );
  NOR2_X1 U19745 ( .A1(n21838), .A2(n18375), .ZN(P3_U2867) );
  NOR2_X4 U19746 ( .A1(n21805), .A2(n18808), .ZN(n18817) );
  AND2_X1 U19747 ( .A1(n18817), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NAND2_X1 U19748 ( .A1(n17757), .A2(n17756), .ZN(n21807) );
  NAND2_X1 U19749 ( .A1(n17758), .A2(n20745), .ZN(n17760) );
  OAI22_X1 U19750 ( .A1(n17760), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n20745), 
        .B2(n20671), .ZN(n17759) );
  INV_X1 U19751 ( .A(n17759), .ZN(P3_U3298) );
  NOR2_X1 U19752 ( .A1(n18807), .A2(n20745), .ZN(n20781) );
  INV_X1 U19753 ( .A(n20781), .ZN(n21164) );
  OAI21_X1 U19754 ( .B1(n17760), .B2(P3_MEMORYFETCH_REG_SCAN_IN), .A(n21164), 
        .ZN(n17761) );
  INV_X1 U19755 ( .A(n17761), .ZN(P3_U3299) );
  INV_X1 U19756 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n17762) );
  NOR2_X1 U19757 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n17762), .ZN(n22329) );
  AOI21_X1 U19758 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n22329), .A(n22322), 
        .ZN(n17764) );
  INV_X1 U19759 ( .A(n17764), .ZN(n22295) );
  INV_X1 U19760 ( .A(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17780) );
  NAND2_X1 U19761 ( .A1(n22328), .A2(n17762), .ZN(n22324) );
  AOI21_X1 U19762 ( .B1(n17763), .B2(n22324), .A(n17765), .ZN(n22291) );
  AOI21_X1 U19763 ( .B1(n17765), .B2(n17780), .A(n22291), .ZN(P2_U3591) );
  AND2_X1 U19764 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n17765), .ZN(P2_U3208) );
  AND2_X1 U19765 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n17765), .ZN(P2_U3207) );
  AND2_X1 U19766 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n17765), .ZN(P2_U3206) );
  AND2_X1 U19767 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n17765), .ZN(P2_U3205) );
  AND2_X1 U19768 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n17765), .ZN(P2_U3204) );
  AND2_X1 U19769 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n17765), .ZN(P2_U3203) );
  AND2_X1 U19770 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n17765), .ZN(P2_U3202) );
  AND2_X1 U19771 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n17765), .ZN(P2_U3201) );
  AND2_X1 U19772 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n17765), .ZN(
        P2_U3200) );
  AND2_X1 U19773 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n17765), .ZN(
        P2_U3199) );
  AND2_X1 U19774 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n17765), .ZN(
        P2_U3198) );
  AND2_X1 U19775 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n17765), .ZN(
        P2_U3197) );
  AND2_X1 U19776 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n17765), .ZN(
        P2_U3196) );
  AND2_X1 U19777 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n17765), .ZN(
        P2_U3195) );
  AND2_X1 U19778 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n17765), .ZN(
        P2_U3194) );
  AND2_X1 U19779 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n17764), .ZN(
        P2_U3193) );
  AND2_X1 U19780 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n17764), .ZN(
        P2_U3192) );
  AND2_X1 U19781 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n17764), .ZN(
        P2_U3191) );
  AND2_X1 U19782 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n17764), .ZN(
        P2_U3190) );
  AND2_X1 U19783 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n17764), .ZN(
        P2_U3189) );
  AND2_X1 U19784 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n17764), .ZN(
        P2_U3188) );
  AND2_X1 U19785 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n17764), .ZN(
        P2_U3187) );
  AND2_X1 U19786 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n17764), .ZN(
        P2_U3186) );
  AND2_X1 U19787 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n17764), .ZN(
        P2_U3185) );
  AND2_X1 U19788 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n17764), .ZN(
        P2_U3184) );
  AND2_X1 U19789 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n17764), .ZN(
        P2_U3183) );
  AND2_X1 U19790 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n17764), .ZN(
        P2_U3182) );
  AND2_X1 U19791 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n17765), .ZN(
        P2_U3181) );
  AND2_X1 U19792 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n17765), .ZN(
        P2_U3180) );
  AND2_X1 U19793 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n17765), .ZN(
        P2_U3179) );
  NAND2_X1 U19794 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19281), .ZN(n19262) );
  AOI21_X1 U19795 ( .B1(n17766), .B2(n19270), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n17767) );
  AOI221_X1 U19796 ( .B1(n19262), .B2(n17767), .C1(n19256), .C2(n17767), .A(
        n19269), .ZN(P2_U3178) );
  INV_X1 U19797 ( .A(n19269), .ZN(n19274) );
  AOI21_X1 U19798 ( .B1(n19256), .B2(n19833), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n19282) );
  OAI221_X1 U19799 ( .B1(n12257), .B2(n19274), .C1(n19272), .C2(n19274), .A(
        n20244), .ZN(n17904) );
  NOR2_X1 U19800 ( .A1(n17769), .A2(n17904), .ZN(P2_U3047) );
  AND2_X1 U19801 ( .A1(n17928), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  NOR4_X1 U19802 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n17773) );
  NOR4_X1 U19803 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n17772) );
  NOR4_X1 U19804 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n17771) );
  NOR4_X1 U19805 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n17770) );
  NAND4_X1 U19806 ( .A1(n17773), .A2(n17772), .A3(n17771), .A4(n17770), .ZN(
        n17779) );
  NOR4_X1 U19807 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n17777) );
  AOI211_X1 U19808 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_31__SCAN_IN), .B(
        P2_DATAWIDTH_REG_30__SCAN_IN), .ZN(n17776) );
  NOR4_X1 U19809 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n17775) );
  NOR4_X1 U19810 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n17774) );
  NAND4_X1 U19811 ( .A1(n17777), .A2(n17776), .A3(n17775), .A4(n17774), .ZN(
        n17778) );
  NOR2_X1 U19812 ( .A1(n17779), .A2(n17778), .ZN(n17914) );
  INV_X1 U19813 ( .A(n17914), .ZN(n17912) );
  NOR2_X1 U19814 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n17912), .ZN(n17907) );
  INV_X1 U19815 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n22294) );
  NAND3_X1 U19816 ( .A1(n18861), .A2(n22294), .A3(n17780), .ZN(n17911) );
  INV_X1 U19817 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n17781) );
  AOI22_X1 U19818 ( .A1(n17907), .A2(n17911), .B1(n17912), .B2(n17781), .ZN(
        P2_U2821) );
  INV_X1 U19819 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n17782) );
  AOI22_X1 U19820 ( .A1(n17907), .A2(n18861), .B1(n17912), .B2(n17782), .ZN(
        P2_U2820) );
  INV_X1 U19821 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17783) );
  NOR2_X1 U19822 ( .A1(n22311), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n22682) );
  AOI21_X1 U19823 ( .B1(n22304), .B2(P1_STATE_REG_0__SCAN_IN), .A(n22682), 
        .ZN(n22287) );
  OAI221_X1 U19824 ( .B1(n22311), .B2(BS16), .C1(n22312), .C2(BS16), .A(n22287), .ZN(n22285) );
  INV_X1 U19825 ( .A(n22285), .ZN(n22288) );
  AOI21_X1 U19826 ( .B1(n17783), .B2(n22289), .A(n22288), .ZN(P1_U3464) );
  AND2_X1 U19827 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n22289), .ZN(P1_U3193) );
  AND2_X1 U19828 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n22289), .ZN(P1_U3192) );
  AND2_X1 U19829 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n22289), .ZN(P1_U3191) );
  AND2_X1 U19830 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n22289), .ZN(P1_U3190) );
  AND2_X1 U19831 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n22289), .ZN(P1_U3189) );
  AND2_X1 U19832 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n22289), .ZN(P1_U3188) );
  AND2_X1 U19833 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n22289), .ZN(P1_U3187) );
  AND2_X1 U19834 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n22289), .ZN(P1_U3186) );
  AND2_X1 U19835 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n22289), .ZN(
        P1_U3185) );
  AND2_X1 U19836 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n22289), .ZN(
        P1_U3184) );
  AND2_X1 U19837 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n22289), .ZN(
        P1_U3183) );
  AND2_X1 U19838 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n22289), .ZN(
        P1_U3182) );
  AND2_X1 U19839 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n22289), .ZN(
        P1_U3181) );
  AND2_X1 U19840 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n22289), .ZN(
        P1_U3180) );
  AND2_X1 U19841 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n22289), .ZN(
        P1_U3179) );
  AND2_X1 U19842 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n22289), .ZN(
        P1_U3178) );
  AND2_X1 U19843 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n22289), .ZN(
        P1_U3177) );
  AND2_X1 U19844 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n22289), .ZN(
        P1_U3176) );
  AND2_X1 U19845 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n22289), .ZN(
        P1_U3175) );
  AND2_X1 U19846 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n22289), .ZN(
        P1_U3174) );
  AND2_X1 U19847 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n22289), .ZN(
        P1_U3173) );
  AND2_X1 U19848 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n22289), .ZN(
        P1_U3172) );
  AND2_X1 U19849 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n22289), .ZN(
        P1_U3171) );
  AND2_X1 U19850 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n22289), .ZN(
        P1_U3170) );
  AND2_X1 U19851 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n22289), .ZN(
        P1_U3169) );
  AND2_X1 U19852 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n22289), .ZN(
        P1_U3168) );
  AND2_X1 U19853 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n22289), .ZN(
        P1_U3167) );
  AND2_X1 U19854 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n22289), .ZN(
        P1_U3166) );
  AND2_X1 U19855 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n22289), .ZN(
        P1_U3165) );
  AND2_X1 U19856 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n22289), .ZN(
        P1_U3164) );
  MUX2_X1 U19857 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n17784), .S(
        n17803), .Z(n17813) );
  NOR2_X1 U19858 ( .A1(n17803), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n17785) );
  AOI21_X1 U19859 ( .B1(n17786), .B2(n17803), .A(n17785), .ZN(n17812) );
  INV_X1 U19860 ( .A(n17812), .ZN(n17798) );
  NOR3_X1 U19861 ( .A1(n17788), .A2(n17787), .A3(n22415), .ZN(n17793) );
  INV_X1 U19862 ( .A(n17793), .ZN(n17791) );
  INV_X1 U19863 ( .A(n17789), .ZN(n17790) );
  OAI211_X1 U19864 ( .C1(n22374), .C2(n17791), .A(n17790), .B(n17803), .ZN(
        n17792) );
  OAI21_X1 U19865 ( .B1(n17793), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n17792), .ZN(n17794) );
  AOI222_X1 U19866 ( .A1(n17813), .A2(n17795), .B1(n17813), .B2(n17794), .C1(
        n17795), .C2(n17794), .ZN(n17796) );
  OR2_X1 U19867 ( .A1(n17796), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n17797) );
  AOI221_X1 U19868 ( .B1(n17798), .B2(n17797), .C1(n17796), .C2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17811) );
  NAND2_X1 U19869 ( .A1(n17799), .A2(n22075), .ZN(n17809) );
  INV_X1 U19870 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n17801) );
  AOI21_X1 U19871 ( .B1(n17801), .B2(n22269), .A(n17800), .ZN(n17806) );
  NOR2_X1 U19872 ( .A1(n17803), .A2(n17802), .ZN(n17805) );
  NOR4_X1 U19873 ( .A1(n17807), .A2(n17806), .A3(n17805), .A4(n17804), .ZN(
        n17808) );
  NAND2_X1 U19874 ( .A1(n17809), .A2(n17808), .ZN(n17810) );
  AOI211_X1 U19875 ( .C1(n17813), .C2(n17812), .A(n17811), .B(n17810), .ZN(
        n22284) );
  INV_X1 U19876 ( .A(n22284), .ZN(n17818) );
  INV_X1 U19877 ( .A(n17814), .ZN(n17815) );
  NAND3_X1 U19878 ( .A1(n14828), .A2(n21878), .A3(n17815), .ZN(n17817) );
  OAI21_X1 U19879 ( .B1(n17825), .B2(n22274), .A(P1_STATE2_REG_2__SCAN_IN), 
        .ZN(n22272) );
  INV_X1 U19880 ( .A(n22272), .ZN(n17816) );
  NAND2_X1 U19881 ( .A1(n21876), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n17820) );
  NAND3_X1 U19882 ( .A1(n17817), .A2(n17816), .A3(n17820), .ZN(n17824) );
  AOI221_X1 U19883 ( .B1(n22274), .B2(n17825), .C1(n17818), .C2(n17825), .A(
        n17824), .ZN(n22276) );
  NOR2_X1 U19884 ( .A1(n22276), .A2(n22274), .ZN(n22275) );
  OAI211_X1 U19885 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n21876), .A(n22275), 
        .B(n17819), .ZN(n22280) );
  NOR3_X1 U19886 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n22274), .A3(n17820), 
        .ZN(n17822) );
  NOR2_X1 U19887 ( .A1(n17822), .A2(n17821), .ZN(n22271) );
  NAND2_X1 U19888 ( .A1(n22271), .A2(n22273), .ZN(n17823) );
  AOI22_X1 U19889 ( .A1(n17825), .A2(n22280), .B1(n17824), .B2(n17823), .ZN(
        P1_U3162) );
  NOR2_X1 U19890 ( .A1(n17827), .A2(n17826), .ZN(P1_U3032) );
  AND2_X1 U19891 ( .A1(n20429), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  INV_X1 U19892 ( .A(n22304), .ZN(n17828) );
  NOR2_X1 U19893 ( .A1(n17828), .A2(n14846), .ZN(n17830) );
  AOI21_X1 U19894 ( .B1(n17830), .B2(n17829), .A(n22682), .ZN(P1_U2802) );
  OAI22_X1 U19895 ( .A1(n17832), .A2(n17859), .B1(n17860), .B2(n17831), .ZN(
        n17833) );
  INV_X1 U19896 ( .A(n17833), .ZN(n17840) );
  AOI21_X1 U19897 ( .B1(n17866), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n17834), .ZN(n17835) );
  OAI21_X1 U19898 ( .B1(n17883), .B2(n17836), .A(n17835), .ZN(n17837) );
  AOI21_X1 U19899 ( .B1(n17838), .B2(n17878), .A(n17837), .ZN(n17839) );
  NAND2_X1 U19900 ( .A1(n17840), .A2(n17839), .ZN(P2_U3012) );
  OAI22_X1 U19901 ( .A1(n12525), .A2(n18976), .B1(n17883), .B2(n18888), .ZN(
        n17841) );
  AOI21_X1 U19902 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17866), .A(
        n17841), .ZN(n17849) );
  AOI21_X1 U19903 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n17843), .A(
        n17842), .ZN(n17846) );
  XNOR2_X1 U19904 ( .A(n17844), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17845) );
  XNOR2_X1 U19905 ( .A(n17846), .B(n17845), .ZN(n19212) );
  XNOR2_X1 U19906 ( .A(n17847), .B(n19204), .ZN(n19210) );
  AOI22_X1 U19907 ( .A1(n19212), .A2(n17879), .B1(n12415), .B2(n19210), .ZN(
        n17848) );
  OAI211_X1 U19908 ( .C1(n17865), .C2(n19201), .A(n17849), .B(n17848), .ZN(
        P2_U3010) );
  AOI22_X1 U19909 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n17866), .B1(
        n17850), .B2(n18898), .ZN(n17856) );
  AOI22_X1 U19910 ( .A1(n17851), .A2(n12415), .B1(n17878), .B2(n18903), .ZN(
        n17855) );
  OR2_X1 U19911 ( .A1(n17852), .A2(n17859), .ZN(n17854) );
  NAND4_X1 U19912 ( .A1(n17856), .A2(n17855), .A3(n17854), .A4(n17853), .ZN(
        P2_U3009) );
  OAI22_X1 U19913 ( .A1(n17957), .A2(n18976), .B1(n17883), .B2(n18911), .ZN(
        n17857) );
  AOI21_X1 U19914 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17866), .A(
        n17857), .ZN(n17864) );
  OAI22_X1 U19915 ( .A1(n17861), .A2(n17860), .B1(n17859), .B2(n17858), .ZN(
        n17862) );
  INV_X1 U19916 ( .A(n17862), .ZN(n17863) );
  OAI211_X1 U19917 ( .C1(n17865), .C2(n18916), .A(n17864), .B(n17863), .ZN(
        P2_U3008) );
  AOI22_X1 U19918 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17866), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19213), .ZN(n17881) );
  NAND2_X1 U19919 ( .A1(n17868), .A2(n17867), .ZN(n17871) );
  OAI21_X1 U19920 ( .B1(n17871), .B2(n17870), .A(n17869), .ZN(n17872) );
  INV_X1 U19921 ( .A(n17872), .ZN(n19194) );
  NAND2_X1 U19922 ( .A1(n17874), .A2(n17873), .ZN(n17877) );
  XNOR2_X1 U19923 ( .A(n17875), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17876) );
  XNOR2_X1 U19924 ( .A(n17877), .B(n17876), .ZN(n19193) );
  AOI222_X1 U19925 ( .A1(n19194), .A2(n12415), .B1(n17879), .B2(n19193), .C1(
        n17878), .C2(n19192), .ZN(n17880) );
  OAI211_X1 U19926 ( .C1(n17883), .C2(n17882), .A(n17881), .B(n17880), .ZN(
        P2_U3006) );
  INV_X1 U19927 ( .A(n17904), .ZN(n17906) );
  INV_X1 U19928 ( .A(n17884), .ZN(n18853) );
  OAI22_X1 U19929 ( .A1(n19925), .A2(n18853), .B1(n19833), .B2(n17885), .ZN(
        n17886) );
  AOI21_X1 U19930 ( .B1(n19927), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n17886), 
        .ZN(n17887) );
  OAI22_X1 U19931 ( .A1(n19927), .A2(n17904), .B1(n17906), .B2(n17887), .ZN(
        P2_U3605) );
  OR2_X1 U19932 ( .A1(n19820), .A2(n22292), .ZN(n19844) );
  INV_X1 U19933 ( .A(n19844), .ZN(n17888) );
  NAND2_X1 U19934 ( .A1(n19879), .A2(n17888), .ZN(n19898) );
  NAND2_X1 U19935 ( .A1(n19844), .A2(n19932), .ZN(n17894) );
  NAND2_X1 U19936 ( .A1(n17894), .A2(n19263), .ZN(n17903) );
  NAND2_X1 U19937 ( .A1(n17899), .A2(n17903), .ZN(n17891) );
  NAND2_X1 U19938 ( .A1(n17889), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17890) );
  OAI211_X1 U19939 ( .C1(n19898), .C2(n19942), .A(n17891), .B(n17890), .ZN(
        n17892) );
  INV_X1 U19940 ( .A(n17892), .ZN(n17893) );
  AOI22_X1 U19941 ( .A1(n17906), .A2(n19832), .B1(n17893), .B2(n17904), .ZN(
        P2_U3603) );
  AOI21_X1 U19942 ( .B1(n22292), .B2(n19820), .A(n17894), .ZN(n17896) );
  OAI22_X1 U19943 ( .A1(n19820), .A2(n19263), .B1(n18873), .B2(n19916), .ZN(
        n17895) );
  NOR2_X1 U19944 ( .A1(n17896), .A2(n17895), .ZN(n17897) );
  AOI22_X1 U19945 ( .A1(n17906), .A2(n19926), .B1(n17897), .B2(n17904), .ZN(
        P2_U3604) );
  INV_X1 U19946 ( .A(n19880), .ZN(n19899) );
  NOR2_X1 U19947 ( .A1(n17898), .A2(n19916), .ZN(n17902) );
  AOI21_X1 U19948 ( .B1(n19913), .B2(n19866), .A(n19819), .ZN(n17900) );
  NOR3_X1 U19949 ( .A1(n17900), .A2(n19942), .A3(n22292), .ZN(n17901) );
  AOI211_X1 U19950 ( .C1(n19899), .C2(n17903), .A(n17902), .B(n17901), .ZN(
        n17905) );
  AOI22_X1 U19951 ( .A1(n17906), .A2(n19809), .B1(n17905), .B2(n17904), .ZN(
        P2_U3602) );
  NAND2_X1 U19952 ( .A1(n17907), .A2(n22294), .ZN(n17910) );
  OAI21_X1 U19953 ( .B1(n18870), .B2(n18861), .A(n17914), .ZN(n17908) );
  OAI21_X1 U19954 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n17914), .A(n17908), 
        .ZN(n17909) );
  OAI221_X1 U19955 ( .B1(n17910), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n17910), .C2(P2_REIP_REG_0__SCAN_IN), .A(n17909), .ZN(P2_U2822) );
  INV_X1 U19956 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n17913) );
  OAI221_X1 U19957 ( .B1(n17914), .B2(n17913), .C1(n17912), .C2(n17911), .A(
        n17910), .ZN(P2_U2823) );
  OAI22_X1 U19958 ( .A1(n17988), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n17987), .ZN(n17915) );
  INV_X1 U19959 ( .A(n17915), .ZN(P2_U3611) );
  INV_X1 U19960 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n17916) );
  AOI22_X1 U19961 ( .A1(n17987), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n17916), 
        .B2(n17988), .ZN(P2_U3608) );
  AOI21_X1 U19962 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n22295), .ZN(n17917) );
  INV_X1 U19963 ( .A(n17917), .ZN(P2_U2815) );
  AOI22_X1 U19964 ( .A1(n17949), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n17948), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n17919) );
  OAI21_X1 U19965 ( .B1(n14822), .B2(n17951), .A(n17919), .ZN(P2_U2951) );
  AOI22_X1 U19966 ( .A1(n17949), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n17948), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n17920) );
  OAI21_X1 U19967 ( .B1(n12500), .B2(n17951), .A(n17920), .ZN(P2_U2950) );
  INV_X1 U19968 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n17922) );
  AOI22_X1 U19969 ( .A1(n17949), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n17928), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n17921) );
  OAI21_X1 U19970 ( .B1(n17922), .B2(n17951), .A(n17921), .ZN(P2_U2949) );
  INV_X1 U19971 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n17924) );
  AOI22_X1 U19972 ( .A1(n17937), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n17948), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n17923) );
  OAI21_X1 U19973 ( .B1(n17924), .B2(n17951), .A(n17923), .ZN(P2_U2948) );
  INV_X1 U19974 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n17926) );
  AOI22_X1 U19975 ( .A1(n17949), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n17948), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n17925) );
  OAI21_X1 U19976 ( .B1(n17926), .B2(n17951), .A(n17925), .ZN(P2_U2947) );
  AOI22_X1 U19977 ( .A1(n17937), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n17928), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n17927) );
  OAI21_X1 U19978 ( .B1(n12536), .B2(n17951), .A(n17927), .ZN(P2_U2946) );
  AOI22_X1 U19979 ( .A1(n17937), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n17928), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n17929) );
  OAI21_X1 U19980 ( .B1(n17930), .B2(n17951), .A(n17929), .ZN(P2_U2945) );
  AOI22_X1 U19981 ( .A1(n17937), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n17948), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n17931) );
  OAI21_X1 U19982 ( .B1(n17932), .B2(n17951), .A(n17931), .ZN(P2_U2944) );
  AOI22_X1 U19983 ( .A1(n17937), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n17948), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n17933) );
  OAI21_X1 U19984 ( .B1(n17934), .B2(n17951), .A(n17933), .ZN(P2_U2943) );
  AOI22_X1 U19985 ( .A1(n17949), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n17948), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n17935) );
  OAI21_X1 U19986 ( .B1(n17936), .B2(n17951), .A(n17935), .ZN(P2_U2942) );
  AOI22_X1 U19987 ( .A1(n17937), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n17948), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n17938) );
  OAI21_X1 U19988 ( .B1(n17939), .B2(n17951), .A(n17938), .ZN(P2_U2941) );
  AOI22_X1 U19989 ( .A1(n17949), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n17948), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n17940) );
  OAI21_X1 U19990 ( .B1(n17941), .B2(n17951), .A(n17940), .ZN(P2_U2940) );
  AOI22_X1 U19991 ( .A1(n17949), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n17948), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n17942) );
  OAI21_X1 U19992 ( .B1(n17943), .B2(n17951), .A(n17942), .ZN(P2_U2939) );
  AOI22_X1 U19993 ( .A1(n17949), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n17948), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n17944) );
  OAI21_X1 U19994 ( .B1(n17945), .B2(n17951), .A(n17944), .ZN(P2_U2938) );
  AOI22_X1 U19995 ( .A1(n17949), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n17948), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n17946) );
  OAI21_X1 U19996 ( .B1(n17947), .B2(n17951), .A(n17946), .ZN(P2_U2937) );
  AOI22_X1 U19997 ( .A1(n17949), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n17948), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n17950) );
  OAI21_X1 U19998 ( .B1(n17952), .B2(n17951), .A(n17950), .ZN(P2_U2936) );
  AOI21_X1 U19999 ( .B1(n17954), .B2(n17953), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n17955) );
  AOI21_X1 U20000 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n17987), .A(n17955), 
        .ZN(P2_U2817) );
  NOR2_X1 U20001 ( .A1(n22328), .A2(n17988), .ZN(n22327) );
  INV_X2 U20002 ( .A(n22327), .ZN(n17981) );
  OAI222_X1 U20003 ( .A1(n17984), .A2(n17956), .B1(n20360), .B2(n17987), .C1(
        n18870), .C2(n17981), .ZN(P2_U3212) );
  INV_X1 U20004 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20362) );
  OAI222_X1 U20005 ( .A1(n17984), .A2(n12520), .B1(n20362), .B2(n17987), .C1(
        n17956), .C2(n17981), .ZN(P2_U3213) );
  INV_X1 U20006 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20364) );
  OAI222_X1 U20007 ( .A1(n17984), .A2(n12525), .B1(n20364), .B2(n17987), .C1(
        n12520), .C2(n17981), .ZN(P2_U3214) );
  INV_X1 U20008 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20366) );
  OAI222_X1 U20009 ( .A1(n17984), .A2(n12530), .B1(n20366), .B2(n17987), .C1(
        n12525), .C2(n17981), .ZN(P2_U3215) );
  INV_X1 U20010 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20368) );
  OAI222_X1 U20011 ( .A1(n17984), .A2(n17957), .B1(n20368), .B2(n17987), .C1(
        n12530), .C2(n17981), .ZN(P2_U3216) );
  INV_X1 U20012 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20370) );
  OAI222_X1 U20013 ( .A1(n17984), .A2(n17958), .B1(n20370), .B2(n17987), .C1(
        n17957), .C2(n17981), .ZN(P2_U3217) );
  INV_X1 U20014 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n17959) );
  OAI222_X1 U20015 ( .A1(n17984), .A2(n12542), .B1(n17959), .B2(n17987), .C1(
        n17958), .C2(n17981), .ZN(P2_U3218) );
  INV_X1 U20016 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n17960) );
  OAI222_X1 U20017 ( .A1(n17984), .A2(n17962), .B1(n17960), .B2(n17987), .C1(
        n12542), .C2(n17981), .ZN(P2_U3219) );
  INV_X1 U20018 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n17961) );
  OAI222_X1 U20019 ( .A1(n17981), .A2(n17962), .B1(n17961), .B2(n17987), .C1(
        n12571), .C2(n17984), .ZN(P2_U3220) );
  INV_X1 U20020 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n17963) );
  OAI222_X1 U20021 ( .A1(n17981), .A2(n12571), .B1(n17963), .B2(n17987), .C1(
        n17964), .C2(n17984), .ZN(P2_U3221) );
  INV_X1 U20022 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20376) );
  OAI222_X1 U20023 ( .A1(n17981), .A2(n17964), .B1(n20376), .B2(n17987), .C1(
        n17965), .C2(n17984), .ZN(P2_U3222) );
  INV_X1 U20024 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20378) );
  OAI222_X1 U20025 ( .A1(n17981), .A2(n17965), .B1(n20378), .B2(n17987), .C1(
        n12612), .C2(n17984), .ZN(P2_U3223) );
  INV_X1 U20026 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20380) );
  OAI222_X1 U20027 ( .A1(n17981), .A2(n12612), .B1(n20380), .B2(n17987), .C1(
        n17966), .C2(n17984), .ZN(P2_U3224) );
  INV_X1 U20028 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20382) );
  OAI222_X1 U20029 ( .A1(n17981), .A2(n17966), .B1(n20382), .B2(n17987), .C1(
        n17967), .C2(n17984), .ZN(P2_U3225) );
  INV_X1 U20030 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20384) );
  OAI222_X1 U20031 ( .A1(n17981), .A2(n17967), .B1(n20384), .B2(n17987), .C1(
        n18989), .C2(n17984), .ZN(P2_U3226) );
  INV_X1 U20032 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20386) );
  OAI222_X1 U20033 ( .A1(n17981), .A2(n18989), .B1(n20386), .B2(n17987), .C1(
        n17969), .C2(n17984), .ZN(P2_U3227) );
  INV_X1 U20034 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n17968) );
  OAI222_X1 U20035 ( .A1(n17981), .A2(n17969), .B1(n17968), .B2(n17987), .C1(
        n19011), .C2(n17984), .ZN(P2_U3228) );
  INV_X1 U20036 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n17970) );
  OAI222_X1 U20037 ( .A1(n17984), .A2(n19026), .B1(n17970), .B2(n17987), .C1(
        n19011), .C2(n17981), .ZN(P2_U3229) );
  INV_X1 U20038 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20390) );
  OAI222_X1 U20039 ( .A1(n17981), .A2(n19026), .B1(n20390), .B2(n17987), .C1(
        n19040), .C2(n17984), .ZN(P2_U3230) );
  INV_X1 U20040 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20392) );
  OAI222_X1 U20041 ( .A1(n17984), .A2(n17971), .B1(n20392), .B2(n17987), .C1(
        n19040), .C2(n17981), .ZN(P2_U3231) );
  INV_X1 U20042 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20394) );
  OAI222_X1 U20043 ( .A1(n17984), .A2(n17972), .B1(n20394), .B2(n17987), .C1(
        n17971), .C2(n17981), .ZN(P2_U3232) );
  INV_X1 U20044 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20396) );
  OAI222_X1 U20045 ( .A1(n17984), .A2(n17973), .B1(n20396), .B2(n17987), .C1(
        n17972), .C2(n17981), .ZN(P2_U3233) );
  INV_X1 U20046 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20398) );
  OAI222_X1 U20047 ( .A1(n17984), .A2(n17974), .B1(n20398), .B2(n17987), .C1(
        n17973), .C2(n17981), .ZN(P2_U3234) );
  INV_X1 U20048 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20400) );
  OAI222_X1 U20049 ( .A1(n17984), .A2(n17976), .B1(n20400), .B2(n17987), .C1(
        n17974), .C2(n17981), .ZN(P2_U3235) );
  INV_X1 U20050 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n17975) );
  OAI222_X1 U20051 ( .A1(n17981), .A2(n17976), .B1(n17975), .B2(n17987), .C1(
        n17977), .C2(n17984), .ZN(P2_U3236) );
  INV_X1 U20052 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n17978) );
  OAI222_X1 U20053 ( .A1(n17984), .A2(n17979), .B1(n17978), .B2(n17987), .C1(
        n17977), .C2(n17981), .ZN(P2_U3237) );
  INV_X1 U20054 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20404) );
  INV_X1 U20055 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n17980) );
  OAI222_X1 U20056 ( .A1(n17981), .A2(n17979), .B1(n20404), .B2(n17987), .C1(
        n17980), .C2(n17984), .ZN(P2_U3238) );
  INV_X1 U20057 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20406) );
  OAI222_X1 U20058 ( .A1(n17981), .A2(n17980), .B1(n20406), .B2(n17987), .C1(
        n17982), .C2(n17984), .ZN(P2_U3239) );
  INV_X1 U20059 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20408) );
  OAI222_X1 U20060 ( .A1(n17981), .A2(n17982), .B1(n20408), .B2(n17987), .C1(
        n17983), .C2(n17984), .ZN(P2_U3240) );
  INV_X1 U20061 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20411) );
  OAI222_X1 U20062 ( .A1(n17984), .A2(n19152), .B1(n20411), .B2(n17987), .C1(
        n17983), .C2(n17981), .ZN(P2_U3241) );
  OAI22_X1 U20063 ( .A1(n17988), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n17987), .ZN(n17985) );
  INV_X1 U20064 ( .A(n17985), .ZN(P2_U3588) );
  OAI22_X1 U20065 ( .A1(n17988), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n17987), .ZN(n17986) );
  INV_X1 U20066 ( .A(n17986), .ZN(P2_U3587) );
  MUX2_X1 U20067 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n17988), .Z(P2_U3586) );
  OAI22_X1 U20068 ( .A1(n17988), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n17987), .ZN(n17989) );
  INV_X1 U20069 ( .A(n17989), .ZN(P2_U3585) );
  NAND2_X1 U20070 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17998), .ZN(n18018) );
  OAI21_X1 U20071 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17998), .A(n18018), .ZN(
        n17991) );
  AOI22_X1 U20072 ( .A1(n18366), .A2(n18296), .B1(n17991), .B2(n18362), .ZN(
        P3_U2699) );
  NOR2_X1 U20073 ( .A1(n21267), .A2(n18365), .ZN(n18364) );
  NAND4_X1 U20074 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .A4(n18364), .ZN(n17995) );
  INV_X1 U20075 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17993) );
  NAND3_X1 U20076 ( .A1(n17995), .A2(P3_EBX_REG_3__SCAN_IN), .A3(n18362), .ZN(
        n17992) );
  OAI221_X1 U20077 ( .B1(n17995), .B2(P3_EBX_REG_3__SCAN_IN), .C1(n18362), 
        .C2(n17993), .A(n17992), .ZN(P3_U2700) );
  NAND2_X1 U20078 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17994) );
  INV_X1 U20079 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n20753) );
  OAI21_X1 U20080 ( .B1(n18365), .B2(n17994), .A(n20753), .ZN(n17996) );
  NAND3_X1 U20081 ( .A1(n18362), .A2(n17996), .A3(n17995), .ZN(n17997) );
  OAI21_X1 U20082 ( .B1(n18362), .B2(n18195), .A(n17997), .ZN(P3_U2701) );
  NAND3_X1 U20083 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(P3_EBX_REG_4__SCAN_IN), 
        .A3(n17998), .ZN(n18015) );
  NOR2_X1 U20084 ( .A1(n20816), .A2(n18015), .ZN(n18011) );
  INV_X1 U20085 ( .A(n18011), .ZN(n18012) );
  NOR2_X1 U20086 ( .A1(n20825), .A2(n18012), .ZN(n17999) );
  OAI21_X1 U20087 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17999), .A(n18362), .ZN(
        n18010) );
  AOI22_X1 U20088 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18165), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18003) );
  AOI22_X1 U20089 ( .A1(n18288), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18130), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n18002) );
  AOI22_X1 U20090 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18326), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18001) );
  AOI22_X1 U20091 ( .A1(n11147), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11175), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18000) );
  NAND4_X1 U20092 ( .A1(n18003), .A2(n18002), .A3(n18001), .A4(n18000), .ZN(
        n18009) );
  AOI22_X1 U20093 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18007) );
  AOI22_X1 U20094 ( .A1(n18342), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n18006) );
  AOI22_X1 U20095 ( .A1(n18332), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11144), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18005) );
  AOI22_X1 U20096 ( .A1(n11145), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18347), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n18004) );
  NAND4_X1 U20097 ( .A1(n18007), .A2(n18006), .A3(n18005), .A4(n18004), .ZN(
        n18008) );
  NOR2_X1 U20098 ( .A1(n18009), .A2(n18008), .ZN(n21336) );
  OAI22_X1 U20099 ( .A1(n18128), .A2(n18010), .B1(n21336), .B2(n18362), .ZN(
        P3_U2695) );
  OAI33_X1 U20100 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n21267), .A3(n18012), .B1(
        n20825), .B2(n18366), .B3(n18011), .ZN(n18013) );
  INV_X1 U20101 ( .A(n18013), .ZN(n18014) );
  OAI21_X1 U20102 ( .B1(n18184), .B2(n18362), .A(n18014), .ZN(P3_U2696) );
  NAND2_X1 U20103 ( .A1(n18362), .A2(n18015), .ZN(n18019) );
  NOR3_X1 U20104 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n21267), .A3(n18015), .ZN(
        n18016) );
  AOI21_X1 U20105 ( .B1(n18366), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n18016), .ZN(n18017) );
  OAI21_X1 U20106 ( .B1(n20816), .B2(n18019), .A(n18017), .ZN(P3_U2697) );
  AND2_X1 U20107 ( .A1(n20798), .A2(n18018), .ZN(n18020) );
  OAI22_X1 U20108 ( .A1(n18020), .A2(n18019), .B1(n18048), .B2(n18362), .ZN(
        P3_U2698) );
  AOI22_X1 U20109 ( .A1(n18288), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18332), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n18024) );
  AOI22_X1 U20110 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11144), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n18023) );
  AOI22_X1 U20111 ( .A1(n11147), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n18022) );
  AOI22_X1 U20112 ( .A1(n18326), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n18055), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18021) );
  NAND4_X1 U20113 ( .A1(n18024), .A2(n18023), .A3(n18022), .A4(n18021), .ZN(
        n18030) );
  AOI22_X1 U20114 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n18130), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n18028) );
  AOI22_X1 U20115 ( .A1(n11145), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18165), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n18027) );
  AOI22_X1 U20116 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n18347), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n18026) );
  AOI22_X1 U20117 ( .A1(n18342), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n18025) );
  NAND4_X1 U20118 ( .A1(n18028), .A2(n18027), .A3(n18026), .A4(n18025), .ZN(
        n18029) );
  NOR2_X1 U20119 ( .A1(n18030), .A2(n18029), .ZN(n21317) );
  INV_X1 U20120 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n20930) );
  NOR2_X1 U20121 ( .A1(n18031), .A2(n18127), .ZN(n18061) );
  NAND2_X1 U20122 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n18061), .ZN(n18033) );
  NOR2_X1 U20123 ( .A1(n20930), .A2(n18033), .ZN(n18046) );
  XNOR2_X1 U20124 ( .A(P3_EBX_REG_16__SCAN_IN), .B(n18046), .ZN(n18032) );
  AOI22_X1 U20125 ( .A1(n18366), .A2(n21317), .B1(n18032), .B2(n18362), .ZN(
        P3_U2687) );
  AOI21_X1 U20126 ( .B1(n20930), .B2(n18033), .A(n18366), .ZN(n18034) );
  INV_X1 U20127 ( .A(n18034), .ZN(n18045) );
  AOI22_X1 U20128 ( .A1(n11144), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n18038) );
  AOI22_X1 U20129 ( .A1(n18342), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n18165), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n18037) );
  AOI22_X1 U20130 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11147), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n18036) );
  AOI22_X1 U20131 ( .A1(n18326), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n18055), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n18035) );
  NAND4_X1 U20132 ( .A1(n18038), .A2(n18037), .A3(n18036), .A4(n18035), .ZN(
        n18044) );
  AOI22_X1 U20133 ( .A1(n18288), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n18332), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n18042) );
  AOI22_X1 U20134 ( .A1(n11145), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18313), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n18041) );
  AOI22_X1 U20135 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18130), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n18040) );
  AOI22_X1 U20136 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18347), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n18039) );
  NAND4_X1 U20137 ( .A1(n18042), .A2(n18041), .A3(n18040), .A4(n18039), .ZN(
        n18043) );
  NOR2_X1 U20138 ( .A1(n18044), .A2(n18043), .ZN(n21329) );
  OAI22_X1 U20139 ( .A1(n18046), .A2(n18045), .B1(n21329), .B2(n18362), .ZN(
        P3_U2688) );
  AOI22_X1 U20140 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n18332), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n18058) );
  AOI22_X1 U20141 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n11144), .B1(
        n18234), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n18057) );
  AOI22_X1 U20142 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n11147), .B1(
        P3_INSTQUEUE_REG_6__5__SCAN_IN), .B2(n18165), .ZN(n18047) );
  OAI21_X1 U20143 ( .B1(n18103), .B2(n18048), .A(n18047), .ZN(n18054) );
  AOI22_X1 U20144 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n11145), .B1(
        P3_INSTQUEUE_REG_2__5__SCAN_IN), .B2(n18349), .ZN(n18052) );
  AOI22_X1 U20145 ( .A1(n18342), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18347), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n18051) );
  AOI22_X1 U20146 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18288), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n18050) );
  AOI22_X1 U20147 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18350), .B1(
        n18130), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n18049) );
  NAND4_X1 U20148 ( .A1(n18052), .A2(n18051), .A3(n18050), .A4(n18049), .ZN(
        n18053) );
  AOI211_X1 U20149 ( .C1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .C2(n18055), .A(
        n18054), .B(n18053), .ZN(n18056) );
  NAND3_X1 U20150 ( .A1(n18058), .A2(n18057), .A3(n18056), .ZN(n21172) );
  INV_X1 U20151 ( .A(n21172), .ZN(n18060) );
  INV_X1 U20152 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n20892) );
  INV_X1 U20153 ( .A(n18127), .ZN(n18113) );
  NAND3_X1 U20154 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_10__SCAN_IN), 
        .A3(n18113), .ZN(n18098) );
  NOR2_X1 U20155 ( .A1(n20892), .A2(n18098), .ZN(n18087) );
  NOR2_X1 U20156 ( .A1(n18366), .A2(n18061), .ZN(n18072) );
  OAI21_X1 U20157 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n18087), .A(n18072), .ZN(
        n18059) );
  OAI21_X1 U20158 ( .B1(n18060), .B2(n18362), .A(n18059), .ZN(P3_U2690) );
  NAND2_X1 U20159 ( .A1(n21197), .A2(n18061), .ZN(n18074) );
  AOI22_X1 U20160 ( .A1(n18288), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n18071) );
  AOI22_X1 U20161 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18070) );
  AOI22_X1 U20162 ( .A1(n11147), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18055), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n18062) );
  OAI21_X1 U20163 ( .B1(n18103), .B2(n18281), .A(n18062), .ZN(n18068) );
  AOI22_X1 U20164 ( .A1(n18130), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18347), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n18066) );
  AOI22_X1 U20165 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n18065) );
  AOI22_X1 U20166 ( .A1(n18332), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11144), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n18064) );
  AOI22_X1 U20167 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18063) );
  NAND4_X1 U20168 ( .A1(n18066), .A2(n18065), .A3(n18064), .A4(n18063), .ZN(
        n18067) );
  AOI211_X1 U20169 ( .C1(n18165), .C2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A(
        n18068), .B(n18067), .ZN(n18069) );
  NAND3_X1 U20170 ( .A1(n18071), .A2(n18070), .A3(n18069), .ZN(n21319) );
  AOI22_X1 U20171 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n18072), .B1(n18366), 
        .B2(n21319), .ZN(n18073) );
  OAI21_X1 U20172 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n18074), .A(n18073), .ZN(
        P3_U2689) );
  INV_X1 U20173 ( .A(n18098), .ZN(n18075) );
  OAI21_X1 U20174 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n18075), .A(n18362), .ZN(
        n18086) );
  AOI22_X1 U20175 ( .A1(n18342), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n18079) );
  AOI22_X1 U20176 ( .A1(n18288), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n18234), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n18078) );
  AOI22_X1 U20177 ( .A1(n18347), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11147), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n18077) );
  AOI22_X1 U20178 ( .A1(n18326), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11175), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n18076) );
  NAND4_X1 U20179 ( .A1(n18079), .A2(n18078), .A3(n18077), .A4(n18076), .ZN(
        n18085) );
  AOI22_X1 U20180 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18165), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18083) );
  AOI22_X1 U20181 ( .A1(n18332), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18130), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n18082) );
  AOI22_X1 U20182 ( .A1(n11144), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n18081) );
  AOI22_X1 U20183 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n18080) );
  NAND4_X1 U20184 ( .A1(n18083), .A2(n18082), .A3(n18081), .A4(n18080), .ZN(
        n18084) );
  NOR2_X1 U20185 ( .A1(n18085), .A2(n18084), .ZN(n21176) );
  OAI22_X1 U20186 ( .A1(n18087), .A2(n18086), .B1(n21176), .B2(n18362), .ZN(
        P3_U2691) );
  AOI22_X1 U20187 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n18091) );
  AOI22_X1 U20188 ( .A1(n18130), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18347), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n18090) );
  AOI22_X1 U20189 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n18326), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18089) );
  AOI22_X1 U20190 ( .A1(n11147), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18055), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18088) );
  NAND4_X1 U20191 ( .A1(n18091), .A2(n18090), .A3(n18089), .A4(n18088), .ZN(
        n18097) );
  AOI22_X1 U20192 ( .A1(n11145), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n18095) );
  AOI22_X1 U20193 ( .A1(n18288), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18165), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n18094) );
  AOI22_X1 U20194 ( .A1(n11144), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18093) );
  AOI22_X1 U20195 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18332), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n18092) );
  NAND4_X1 U20196 ( .A1(n18095), .A2(n18094), .A3(n18093), .A4(n18092), .ZN(
        n18096) );
  NOR2_X1 U20197 ( .A1(n18097), .A2(n18096), .ZN(n21181) );
  INV_X1 U20198 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n18114) );
  NOR2_X1 U20199 ( .A1(n18114), .A2(n18127), .ZN(n18099) );
  OAI21_X1 U20200 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n18099), .A(n18098), .ZN(
        n18100) );
  AOI22_X1 U20201 ( .A1(n18366), .A2(n21181), .B1(n18100), .B2(n18362), .ZN(
        P3_U2692) );
  AOI22_X1 U20202 ( .A1(n18288), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n18101), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n18112) );
  AOI22_X1 U20203 ( .A1(n11144), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18347), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18111) );
  AOI22_X1 U20204 ( .A1(n11147), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n18055), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18102) );
  OAI21_X1 U20205 ( .B1(n18103), .B2(n18195), .A(n18102), .ZN(n18109) );
  AOI22_X1 U20206 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n18107) );
  AOI22_X1 U20207 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14341), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n18106) );
  AOI22_X1 U20208 ( .A1(n18130), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18105) );
  AOI22_X1 U20209 ( .A1(n18165), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18104) );
  NAND4_X1 U20210 ( .A1(n18107), .A2(n18106), .A3(n18105), .A4(n18104), .ZN(
        n18108) );
  AOI211_X1 U20211 ( .C1(n11164), .C2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n18109), .B(n18108), .ZN(n18110) );
  NAND3_X1 U20212 ( .A1(n18112), .A2(n18111), .A3(n18110), .ZN(n21185) );
  OAI33_X1 U20213 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n21267), .A3(n18127), 
        .B1(n18114), .B2(n18366), .B3(n18113), .ZN(n18115) );
  AOI21_X1 U20214 ( .B1(n18366), .B2(n21185), .A(n18115), .ZN(n18116) );
  INV_X1 U20215 ( .A(n18116), .ZN(P3_U2693) );
  AOI22_X1 U20216 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n18165), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n18120) );
  AOI22_X1 U20217 ( .A1(n18288), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n18313), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n18119) );
  AOI22_X1 U20218 ( .A1(n18342), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11147), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n18118) );
  AOI22_X1 U20219 ( .A1(n18326), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n18055), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n18117) );
  NAND4_X1 U20220 ( .A1(n18120), .A2(n18119), .A3(n18118), .A4(n18117), .ZN(
        n18126) );
  AOI22_X1 U20221 ( .A1(n11145), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n18347), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n18124) );
  AOI22_X1 U20222 ( .A1(n11144), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n18123) );
  AOI22_X1 U20223 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n18130), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n18122) );
  AOI22_X1 U20224 ( .A1(n18332), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n18234), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n18121) );
  NAND4_X1 U20225 ( .A1(n18124), .A2(n18123), .A3(n18122), .A4(n18121), .ZN(
        n18125) );
  NOR2_X1 U20226 ( .A1(n18126), .A2(n18125), .ZN(n21192) );
  OAI211_X1 U20227 ( .C1(P3_EBX_REG_9__SCAN_IN), .C2(n18128), .A(n18127), .B(
        n18362), .ZN(n18129) );
  OAI21_X1 U20228 ( .B1(n21192), .B2(n18362), .A(n18129), .ZN(P3_U2694) );
  AOI22_X1 U20229 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11144), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n18134) );
  AOI22_X1 U20230 ( .A1(n18332), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18347), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n18133) );
  AOI22_X1 U20231 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n18130), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18132) );
  AOI22_X1 U20232 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18165), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n18131) );
  NAND4_X1 U20233 ( .A1(n18134), .A2(n18133), .A3(n18132), .A4(n18131), .ZN(
        n18140) );
  AOI22_X1 U20234 ( .A1(n18342), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n18138) );
  AOI22_X1 U20235 ( .A1(n18288), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18313), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n18137) );
  AOI22_X1 U20236 ( .A1(n11145), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11175), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n18136) );
  AOI22_X1 U20237 ( .A1(n11147), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n18326), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n18135) );
  NAND4_X1 U20238 ( .A1(n18138), .A2(n18137), .A3(n18136), .A4(n18135), .ZN(
        n18139) );
  NOR2_X1 U20239 ( .A1(n18140), .A2(n18139), .ZN(n18226) );
  AOI22_X1 U20240 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18234), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n18144) );
  AOI22_X1 U20241 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18342), .B1(
        P3_INSTQUEUE_REG_1__5__SCAN_IN), .B2(n11164), .ZN(n18143) );
  AOI22_X1 U20242 ( .A1(n18288), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__5__SCAN_IN), .B2(n11147), .ZN(n18142) );
  AOI22_X1 U20243 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n11175), .B1(
        P3_INSTQUEUE_REG_2__5__SCAN_IN), .B2(n18326), .ZN(n18141) );
  NAND4_X1 U20244 ( .A1(n18144), .A2(n18143), .A3(n18142), .A4(n18141), .ZN(
        n18150) );
  AOI22_X1 U20245 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18347), .B1(
        P3_INSTQUEUE_REG_12__5__SCAN_IN), .B2(n11144), .ZN(n18148) );
  AOI22_X1 U20246 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18165), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n18147) );
  AOI22_X1 U20247 ( .A1(n18130), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__5__SCAN_IN), .B2(n18349), .ZN(n18146) );
  AOI22_X1 U20248 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n18332), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n18145) );
  NAND4_X1 U20249 ( .A1(n18148), .A2(n18147), .A3(n18146), .A4(n18145), .ZN(
        n18149) );
  NOR2_X1 U20250 ( .A1(n18150), .A2(n18149), .ZN(n18254) );
  AOI22_X1 U20251 ( .A1(n18342), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18165), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n18154) );
  AOI22_X1 U20252 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18234), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n18153) );
  AOI22_X1 U20253 ( .A1(n18130), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11147), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n18152) );
  AOI22_X1 U20254 ( .A1(n18326), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11175), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n18151) );
  NAND4_X1 U20255 ( .A1(n18154), .A2(n18153), .A3(n18152), .A4(n18151), .ZN(
        n18160) );
  AOI22_X1 U20256 ( .A1(n11144), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18158) );
  AOI22_X1 U20257 ( .A1(n11145), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18313), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n18157) );
  AOI22_X1 U20258 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n18332), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18156) );
  AOI22_X1 U20259 ( .A1(n18288), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18347), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n18155) );
  NAND4_X1 U20260 ( .A1(n18158), .A2(n18157), .A3(n18156), .A4(n18155), .ZN(
        n18159) );
  NOR2_X1 U20261 ( .A1(n18160), .A2(n18159), .ZN(n18259) );
  AOI22_X1 U20262 ( .A1(n18342), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n18313), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n18164) );
  AOI22_X1 U20263 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n18163) );
  AOI22_X1 U20264 ( .A1(n11144), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n18326), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n18162) );
  AOI22_X1 U20265 ( .A1(n11147), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n18055), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n18161) );
  NAND4_X1 U20266 ( .A1(n18164), .A2(n18163), .A3(n18162), .A4(n18161), .ZN(
        n18171) );
  AOI22_X1 U20267 ( .A1(n18332), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n18130), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18169) );
  AOI22_X1 U20268 ( .A1(n18350), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n18165), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n18168) );
  AOI22_X1 U20269 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n18234), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n18167) );
  AOI22_X1 U20270 ( .A1(n18288), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n18347), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n18166) );
  NAND4_X1 U20271 ( .A1(n18169), .A2(n18168), .A3(n18167), .A4(n18166), .ZN(
        n18170) );
  NOR2_X1 U20272 ( .A1(n18171), .A2(n18170), .ZN(n18269) );
  AOI22_X1 U20273 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n18130), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18182) );
  AOI22_X1 U20274 ( .A1(n11145), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18347), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18181) );
  INV_X1 U20275 ( .A(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n18173) );
  AOI22_X1 U20276 ( .A1(n11144), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n18172) );
  OAI21_X1 U20277 ( .B1(n11209), .B2(n18173), .A(n18172), .ZN(n18179) );
  AOI22_X1 U20278 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n18332), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n18177) );
  AOI22_X1 U20279 ( .A1(n18288), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18176) );
  AOI22_X1 U20280 ( .A1(n18165), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11147), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n18175) );
  AOI22_X1 U20281 ( .A1(n18326), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n18055), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n18174) );
  NAND4_X1 U20282 ( .A1(n18177), .A2(n18176), .A3(n18175), .A4(n18174), .ZN(
        n18178) );
  AOI211_X1 U20283 ( .C1(n18341), .C2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A(
        n18179), .B(n18178), .ZN(n18180) );
  NAND3_X1 U20284 ( .A1(n18182), .A2(n18181), .A3(n18180), .ZN(n18275) );
  AOI22_X1 U20285 ( .A1(n18165), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n18313), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n18193) );
  AOI22_X1 U20286 ( .A1(n18288), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18347), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n18192) );
  AOI22_X1 U20287 ( .A1(n18332), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n18183) );
  OAI21_X1 U20288 ( .B1(n11190), .B2(n18184), .A(n18183), .ZN(n18190) );
  AOI22_X1 U20289 ( .A1(n18130), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n18188) );
  AOI22_X1 U20290 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n18187) );
  AOI22_X1 U20291 ( .A1(n11144), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11175), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n18186) );
  AOI22_X1 U20292 ( .A1(n11147), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n18326), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n18185) );
  NAND4_X1 U20293 ( .A1(n18188), .A2(n18187), .A3(n18186), .A4(n18185), .ZN(
        n18189) );
  AOI211_X1 U20294 ( .C1(n11143), .C2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n18190), .B(n18189), .ZN(n18191) );
  NAND3_X1 U20295 ( .A1(n18193), .A2(n18192), .A3(n18191), .ZN(n18276) );
  NAND2_X1 U20296 ( .A1(n18275), .A2(n18276), .ZN(n18274) );
  NOR2_X1 U20297 ( .A1(n18269), .A2(n18274), .ZN(n18268) );
  AOI22_X1 U20298 ( .A1(n18342), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18204) );
  AOI22_X1 U20299 ( .A1(n11144), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18331), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n18203) );
  AOI22_X1 U20300 ( .A1(n18347), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18313), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18194) );
  OAI21_X1 U20301 ( .B1(n18216), .B2(n18195), .A(n18194), .ZN(n18201) );
  AOI22_X1 U20302 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n18199) );
  AOI22_X1 U20303 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11164), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18198) );
  AOI22_X1 U20304 ( .A1(n18332), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11147), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n18197) );
  AOI22_X1 U20305 ( .A1(n18326), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11175), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n18196) );
  NAND4_X1 U20306 ( .A1(n18199), .A2(n18198), .A3(n18197), .A4(n18196), .ZN(
        n18200) );
  AOI211_X1 U20307 ( .C1(n18288), .C2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A(
        n18201), .B(n18200), .ZN(n18202) );
  NAND3_X1 U20308 ( .A1(n18204), .A2(n18203), .A3(n18202), .ZN(n18265) );
  NAND2_X1 U20309 ( .A1(n18268), .A2(n18265), .ZN(n18264) );
  NOR2_X1 U20310 ( .A1(n18259), .A2(n18264), .ZN(n18258) );
  AOI22_X1 U20311 ( .A1(n18342), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18347), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18214) );
  AOI22_X1 U20312 ( .A1(n18348), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n18331), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n18213) );
  AOI22_X1 U20313 ( .A1(n11144), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n18205) );
  OAI21_X1 U20314 ( .B1(n18216), .B2(n18296), .A(n18205), .ZN(n18211) );
  AOI22_X1 U20315 ( .A1(n18332), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n18209) );
  AOI22_X1 U20316 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18313), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n18208) );
  AOI22_X1 U20317 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11147), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n18207) );
  AOI22_X1 U20318 ( .A1(n18326), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n18055), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n18206) );
  NAND4_X1 U20319 ( .A1(n18209), .A2(n18208), .A3(n18207), .A4(n18206), .ZN(
        n18210) );
  AOI211_X1 U20320 ( .C1(n11143), .C2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n18211), .B(n18210), .ZN(n18212) );
  NAND3_X1 U20321 ( .A1(n18214), .A2(n18213), .A3(n18212), .ZN(n18244) );
  NAND2_X1 U20322 ( .A1(n18258), .A2(n18244), .ZN(n18253) );
  NOR2_X1 U20323 ( .A1(n18254), .A2(n18253), .ZN(n18252) );
  AOI22_X1 U20324 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18225) );
  AOI22_X1 U20325 ( .A1(n18348), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18331), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n18224) );
  AOI22_X1 U20326 ( .A1(n18332), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18347), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18215) );
  OAI21_X1 U20327 ( .B1(n18216), .B2(n18281), .A(n18215), .ZN(n18222) );
  AOI22_X1 U20328 ( .A1(n11144), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18220) );
  AOI22_X1 U20329 ( .A1(n18342), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18313), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n18219) );
  AOI22_X1 U20330 ( .A1(n18341), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18055), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n18218) );
  AOI22_X1 U20331 ( .A1(n11147), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n18326), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18217) );
  NAND4_X1 U20332 ( .A1(n18220), .A2(n18219), .A3(n18218), .A4(n18217), .ZN(
        n18221) );
  AOI211_X1 U20333 ( .C1(n11143), .C2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A(
        n18222), .B(n18221), .ZN(n18223) );
  NAND3_X1 U20334 ( .A1(n18225), .A2(n18224), .A3(n18223), .ZN(n18247) );
  NAND2_X1 U20335 ( .A1(n18252), .A2(n18247), .ZN(n18246) );
  XNOR2_X1 U20336 ( .A(n18226), .B(n18246), .ZN(n21284) );
  NOR2_X1 U20337 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n18227), .ZN(n18229) );
  OAI22_X1 U20338 ( .A1(n21284), .A2(n18362), .B1(n18229), .B2(n18228), .ZN(
        P3_U2673) );
  AOI22_X1 U20339 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__5__SCAN_IN), .B2(n11145), .ZN(n18233) );
  AOI22_X1 U20340 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18349), .B1(
        n18331), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n18232) );
  AOI22_X1 U20341 ( .A1(n18348), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__5__SCAN_IN), .B2(n11147), .ZN(n18231) );
  AOI22_X1 U20342 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18326), .B1(
        P3_INSTQUEUE_REG_10__5__SCAN_IN), .B2(n11175), .ZN(n18230) );
  NAND4_X1 U20343 ( .A1(n18233), .A2(n18232), .A3(n18231), .A4(n18230), .ZN(
        n18240) );
  AOI22_X1 U20344 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18332), .B1(
        n18130), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n18238) );
  AOI22_X1 U20345 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18234), .B1(
        n11164), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18237) );
  AOI22_X1 U20346 ( .A1(n11144), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__5__SCAN_IN), .B2(n18342), .ZN(n18236) );
  AOI22_X1 U20347 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18347), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n18235) );
  NAND4_X1 U20348 ( .A1(n18238), .A2(n18237), .A3(n18236), .A4(n18235), .ZN(
        n18239) );
  NOR2_X1 U20349 ( .A1(n18240), .A2(n18239), .ZN(n21233) );
  AND2_X1 U20350 ( .A1(n18362), .A2(n18241), .ZN(n18306) );
  INV_X1 U20351 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n21018) );
  AOI22_X1 U20352 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n18306), .B1(n18279), 
        .B2(n21018), .ZN(n18242) );
  OAI21_X1 U20353 ( .B1(n21233), .B2(n18362), .A(n18242), .ZN(P3_U2682) );
  INV_X1 U20354 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n21068) );
  NAND2_X1 U20355 ( .A1(n18279), .A2(n18243), .ZN(n18263) );
  NAND2_X1 U20356 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n18262), .ZN(n18257) );
  INV_X1 U20357 ( .A(n18257), .ZN(n18248) );
  AOI21_X1 U20358 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n18362), .A(n18262), .ZN(
        n18245) );
  OAI21_X1 U20359 ( .B1(n18258), .B2(n18244), .A(n18253), .ZN(n21299) );
  OAI22_X1 U20360 ( .A1(n18248), .A2(n18245), .B1(n21299), .B2(n18362), .ZN(
        P3_U2676) );
  OAI21_X1 U20361 ( .B1(n18252), .B2(n18247), .A(n18246), .ZN(n21288) );
  NOR2_X1 U20362 ( .A1(n18366), .A2(n18248), .ZN(n18255) );
  INV_X1 U20363 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n18249) );
  OAI221_X1 U20364 ( .B1(n18255), .B2(n18364), .C1(n18255), .C2(n18249), .A(
        P3_EBX_REG_29__SCAN_IN), .ZN(n18251) );
  NAND4_X1 U20365 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(n18262), .A4(n21112), .ZN(n18250) );
  OAI211_X1 U20366 ( .C1(n18362), .C2(n21288), .A(n18251), .B(n18250), .ZN(
        P3_U2674) );
  AOI21_X1 U20367 ( .B1(n18254), .B2(n18253), .A(n18252), .ZN(n21289) );
  AOI22_X1 U20368 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n18255), .B1(n21289), 
        .B2(n18366), .ZN(n18256) );
  OAI21_X1 U20369 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n18257), .A(n18256), .ZN(
        P3_U2675) );
  AOI21_X1 U20370 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n18362), .A(n18267), .ZN(
        n18261) );
  AOI21_X1 U20371 ( .B1(n18259), .B2(n18264), .A(n18258), .ZN(n21272) );
  INV_X1 U20372 ( .A(n21272), .ZN(n18260) );
  OAI22_X1 U20373 ( .A1(n18262), .A2(n18261), .B1(n18260), .B2(n18362), .ZN(
        P3_U2677) );
  INV_X1 U20374 ( .A(n18263), .ZN(n18272) );
  AOI21_X1 U20375 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n18362), .A(n18272), .ZN(
        n18266) );
  OAI21_X1 U20376 ( .B1(n18268), .B2(n18265), .A(n18264), .ZN(n21271) );
  OAI22_X1 U20377 ( .A1(n18267), .A2(n18266), .B1(n21271), .B2(n18362), .ZN(
        P3_U2678) );
  INV_X1 U20378 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n21045) );
  NAND3_X1 U20379 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .A3(n18279), .ZN(n18273) );
  NOR2_X1 U20380 ( .A1(n21045), .A2(n18273), .ZN(n18278) );
  AOI21_X1 U20381 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n18362), .A(n18278), .ZN(
        n18271) );
  AOI21_X1 U20382 ( .B1(n18269), .B2(n18274), .A(n18268), .ZN(n21300) );
  INV_X1 U20383 ( .A(n21300), .ZN(n18270) );
  OAI22_X1 U20384 ( .A1(n18272), .A2(n18271), .B1(n18270), .B2(n18362), .ZN(
        P3_U2679) );
  INV_X1 U20385 ( .A(n18273), .ZN(n18294) );
  AOI21_X1 U20386 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n18362), .A(n18294), .ZN(
        n18277) );
  OAI21_X1 U20387 ( .B1(n18276), .B2(n18275), .A(n18274), .ZN(n21311) );
  OAI22_X1 U20388 ( .A1(n18278), .A2(n18277), .B1(n21311), .B2(n18362), .ZN(
        P3_U2680) );
  AOI22_X1 U20389 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n18362), .B1(
        P3_EBX_REG_21__SCAN_IN), .B2(n18279), .ZN(n18293) );
  AOI22_X1 U20390 ( .A1(n11144), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18313), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18291) );
  AOI22_X1 U20391 ( .A1(n18350), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18347), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n18290) );
  AOI22_X1 U20392 ( .A1(n18341), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18331), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18280) );
  OAI21_X1 U20393 ( .B1(n11190), .B2(n18281), .A(n18280), .ZN(n18287) );
  AOI22_X1 U20394 ( .A1(n18342), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18285) );
  AOI22_X1 U20395 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18130), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18284) );
  AOI22_X1 U20396 ( .A1(n18332), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11147), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18283) );
  AOI22_X1 U20397 ( .A1(n18326), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18055), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n18282) );
  NAND4_X1 U20398 ( .A1(n18285), .A2(n18284), .A3(n18283), .A4(n18282), .ZN(
        n18286) );
  AOI211_X1 U20399 ( .C1(n18288), .C2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A(
        n18287), .B(n18286), .ZN(n18289) );
  NAND3_X1 U20400 ( .A1(n18291), .A2(n18290), .A3(n18289), .ZN(n21244) );
  INV_X1 U20401 ( .A(n21244), .ZN(n18292) );
  OAI22_X1 U20402 ( .A1(n18294), .A2(n18293), .B1(n18292), .B2(n18362), .ZN(
        P3_U2681) );
  AOI22_X1 U20403 ( .A1(n18341), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n18305) );
  AOI22_X1 U20404 ( .A1(n18348), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18130), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n18304) );
  AOI22_X1 U20405 ( .A1(n11144), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18313), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n18295) );
  OAI21_X1 U20406 ( .B1(n11190), .B2(n18296), .A(n18295), .ZN(n18302) );
  AOI22_X1 U20407 ( .A1(n11145), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18347), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n18300) );
  AOI22_X1 U20408 ( .A1(n18332), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n18299) );
  AOI22_X1 U20409 ( .A1(n18165), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11175), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18298) );
  AOI22_X1 U20410 ( .A1(n11147), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n18326), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n18297) );
  NAND4_X1 U20411 ( .A1(n18300), .A2(n18299), .A3(n18298), .A4(n18297), .ZN(
        n18301) );
  AOI211_X1 U20412 ( .C1(n11143), .C2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A(
        n18302), .B(n18301), .ZN(n18303) );
  NAND3_X1 U20413 ( .A1(n18305), .A2(n18304), .A3(n18303), .ZN(n21237) );
  INV_X1 U20414 ( .A(n21237), .ZN(n18308) );
  OAI21_X1 U20415 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n18340), .A(n18306), .ZN(
        n18307) );
  OAI21_X1 U20416 ( .B1(n18308), .B2(n18362), .A(n18307), .ZN(P3_U2683) );
  AOI22_X1 U20417 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n18312) );
  AOI22_X1 U20418 ( .A1(n18341), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n18311) );
  AOI22_X1 U20419 ( .A1(n18130), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18326), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18310) );
  AOI22_X1 U20420 ( .A1(n11147), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n18055), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n18309) );
  NAND4_X1 U20421 ( .A1(n18312), .A2(n18311), .A3(n18310), .A4(n18309), .ZN(
        n18319) );
  AOI22_X1 U20422 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18347), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18317) );
  AOI22_X1 U20423 ( .A1(n11144), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18331), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n18316) );
  AOI22_X1 U20424 ( .A1(n18348), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n18313), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n18315) );
  AOI22_X1 U20425 ( .A1(n18332), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n18314) );
  NAND4_X1 U20426 ( .A1(n18317), .A2(n18316), .A3(n18315), .A4(n18314), .ZN(
        n18318) );
  NOR2_X1 U20427 ( .A1(n18319), .A2(n18318), .ZN(n21259) );
  NOR2_X1 U20428 ( .A1(n18366), .A2(n18320), .ZN(n18322) );
  NOR2_X1 U20429 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n18357), .ZN(n18321) );
  AOI22_X1 U20430 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n18322), .B1(n18364), 
        .B2(n18321), .ZN(n18323) );
  OAI21_X1 U20431 ( .B1(n21259), .B2(n18362), .A(n18323), .ZN(P3_U2685) );
  AOI21_X1 U20432 ( .B1(n20992), .B2(n18324), .A(n18366), .ZN(n18325) );
  INV_X1 U20433 ( .A(n18325), .ZN(n18339) );
  AOI22_X1 U20434 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11164), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18330) );
  AOI22_X1 U20435 ( .A1(n18341), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n18329) );
  AOI22_X1 U20436 ( .A1(n11144), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11175), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n18328) );
  AOI22_X1 U20437 ( .A1(n11147), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n18326), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n18327) );
  NAND4_X1 U20438 ( .A1(n18330), .A2(n18329), .A3(n18328), .A4(n18327), .ZN(
        n18338) );
  AOI22_X1 U20439 ( .A1(n11145), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18336) );
  AOI22_X1 U20440 ( .A1(n18348), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18347), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n18335) );
  AOI22_X1 U20441 ( .A1(n18332), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n18331), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n18334) );
  AOI22_X1 U20442 ( .A1(n18130), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n18333) );
  NAND4_X1 U20443 ( .A1(n18336), .A2(n18335), .A3(n18334), .A4(n18333), .ZN(
        n18337) );
  NOR2_X1 U20444 ( .A1(n18338), .A2(n18337), .ZN(n21253) );
  OAI22_X1 U20445 ( .A1(n18340), .A2(n18339), .B1(n21253), .B2(n18362), .ZN(
        P3_U2684) );
  AOI22_X1 U20446 ( .A1(n18341), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n18346) );
  AOI22_X1 U20447 ( .A1(n11143), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n18345) );
  AOI22_X1 U20448 ( .A1(n18165), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11147), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n18344) );
  AOI22_X1 U20449 ( .A1(n18326), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11175), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n18343) );
  NAND4_X1 U20450 ( .A1(n18346), .A2(n18345), .A3(n18344), .A4(n18343), .ZN(
        n18356) );
  AOI22_X1 U20451 ( .A1(n18332), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11144), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n18354) );
  AOI22_X1 U20452 ( .A1(n18348), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n18347), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n18353) );
  AOI22_X1 U20453 ( .A1(n18130), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18352) );
  AOI22_X1 U20454 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n18350), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n18351) );
  NAND4_X1 U20455 ( .A1(n18354), .A2(n18353), .A3(n18352), .A4(n18351), .ZN(
        n18355) );
  NOR2_X1 U20456 ( .A1(n18356), .A2(n18355), .ZN(n21264) );
  NAND2_X1 U20457 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n18365), .ZN(n18360) );
  OAI211_X1 U20458 ( .C1(P3_EBX_REG_17__SCAN_IN), .C2(n18358), .A(n18364), .B(
        n18357), .ZN(n18359) );
  OAI211_X1 U20459 ( .C1(n21264), .C2(n18362), .A(n18360), .B(n18359), .ZN(
        P3_U2686) );
  INV_X1 U20460 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18363) );
  NOR2_X1 U20461 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n20754) );
  AOI21_X1 U20462 ( .B1(P3_EBX_REG_1__SCAN_IN), .B2(P3_EBX_REG_0__SCAN_IN), 
        .A(n20754), .ZN(n20743) );
  AOI22_X1 U20463 ( .A1(P3_EBX_REG_1__SCAN_IN), .A2(n18365), .B1(n18364), .B2(
        n20743), .ZN(n18361) );
  OAI21_X1 U20464 ( .B1(n18363), .B2(n18362), .A(n18361), .ZN(P3_U2702) );
  INV_X1 U20465 ( .A(n18364), .ZN(n18368) );
  AOI22_X1 U20466 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18366), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n18365), .ZN(n18367) );
  OAI21_X1 U20467 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n18368), .A(n18367), .ZN(
        P3_U2703) );
  INV_X1 U20468 ( .A(n20681), .ZN(n20680) );
  OAI21_X1 U20469 ( .B1(n21816), .B2(n20680), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n18369) );
  OAI21_X1 U20470 ( .B1(n18370), .B2(n21857), .A(n18369), .ZN(P3_U2634) );
  INV_X1 U20471 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n21872) );
  AOI21_X1 U20472 ( .B1(n21872), .B2(n18372), .A(n18371), .ZN(n21860) );
  OAI21_X1 U20473 ( .B1(n21860), .B2(n18373), .A(n18375), .ZN(n18374) );
  OAI221_X1 U20474 ( .B1(n21825), .B2(n20674), .C1(n21825), .C2(n18375), .A(
        n18374), .ZN(P3_U2863) );
  OAI21_X1 U20475 ( .B1(n18393), .B2(n21668), .A(n18394), .ZN(n18377) );
  XNOR2_X1 U20476 ( .A(n18377), .B(n18376), .ZN(n21743) );
  INV_X1 U20477 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n18381) );
  NAND2_X1 U20478 ( .A1(n18378), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18379) );
  INV_X1 U20479 ( .A(n18379), .ZN(n18599) );
  XNOR2_X1 U20480 ( .A(n18381), .B(n18599), .ZN(n20976) );
  NAND2_X1 U20481 ( .A1(n18378), .A2(n18549), .ZN(n18388) );
  OAI21_X1 U20482 ( .B1(n18378), .B2(n18715), .A(n18753), .ZN(n18603) );
  AOI21_X1 U20483 ( .B1(n11315), .B2(n18379), .A(n18603), .ZN(n18389) );
  NAND2_X1 U20484 ( .A1(n14606), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18380) );
  OAI221_X1 U20485 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18388), .C1(
        n18381), .C2(n18389), .A(n18380), .ZN(n18382) );
  AOI21_X1 U20486 ( .B1(n18593), .B2(n20976), .A(n18382), .ZN(n18384) );
  NAND2_X1 U20487 ( .A1(n18645), .A2(n21725), .ZN(n18416) );
  AOI22_X1 U20488 ( .A1(n18672), .A2(n21567), .B1(n18748), .B2(n11422), .ZN(
        n18422) );
  OAI21_X1 U20489 ( .B1(n21730), .B2(n18416), .A(n18422), .ZN(n18606) );
  NOR2_X1 U20490 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n21398), .ZN(
        n21726) );
  AOI22_X1 U20491 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18606), .B1(
        n18607), .B2(n21726), .ZN(n18383) );
  OAI211_X1 U20492 ( .C1(n18675), .C2(n21743), .A(n18384), .B(n18383), .ZN(
        P3_U2812) );
  NAND2_X1 U20493 ( .A1(n21403), .A2(n18607), .ZN(n18474) );
  INV_X1 U20494 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n20996) );
  NAND2_X1 U20495 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18599), .ZN(
        n18385) );
  AOI22_X1 U20496 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18478), .B1(
        n20996), .B2(n18385), .ZN(n20986) );
  INV_X1 U20497 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n20998) );
  NOR2_X1 U20498 ( .A1(n11142), .A2(n20998), .ZN(n18391) );
  OAI21_X1 U20499 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n18386), .ZN(n18387) );
  OAI22_X1 U20500 ( .A1(n18389), .A2(n20996), .B1(n18388), .B2(n18387), .ZN(
        n18390) );
  AOI211_X1 U20501 ( .C1(n20986), .C2(n18593), .A(n18391), .B(n18390), .ZN(
        n18397) );
  NAND2_X1 U20502 ( .A1(n21403), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n21404) );
  NOR2_X1 U20503 ( .A1(n21567), .A2(n21404), .ZN(n21706) );
  NOR2_X1 U20504 ( .A1(n11422), .A2(n21404), .ZN(n21705) );
  OAI22_X1 U20505 ( .A1(n21706), .A2(n18589), .B1(n21705), .B2(n18758), .ZN(
        n18476) );
  NOR3_X1 U20506 ( .A1(n21668), .A2(n18393), .A3(n18392), .ZN(n18463) );
  NOR2_X1 U20507 ( .A1(n18604), .A2(n18394), .ZN(n18469) );
  NOR2_X1 U20508 ( .A1(n18463), .A2(n18469), .ZN(n18395) );
  XOR2_X1 U20509 ( .A(n18395), .B(n21714), .Z(n21712) );
  AOI22_X1 U20510 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18476), .B1(
        n18661), .B2(n21712), .ZN(n18396) );
  OAI211_X1 U20511 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n18474), .A(
        n18397), .B(n18396), .ZN(P3_U2811) );
  NOR2_X1 U20512 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21565), .ZN(
        n18409) );
  NAND2_X1 U20513 ( .A1(n18398), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20932) );
  INV_X1 U20514 ( .A(n20932), .ZN(n18616) );
  OAI22_X1 U20515 ( .A1(n18411), .A2(n20932), .B1(n18616), .B2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n20934) );
  INV_X1 U20516 ( .A(n20934), .ZN(n20935) );
  NAND4_X1 U20517 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n20900), .A3(
        n18399), .A4(n18549), .ZN(n18410) );
  OAI21_X1 U20518 ( .B1(n18398), .B2(n18715), .A(n18753), .ZN(n18620) );
  AOI21_X1 U20519 ( .B1(n11315), .B2(n20932), .A(n18620), .ZN(n18413) );
  NAND2_X1 U20520 ( .A1(n14606), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n21570) );
  OAI221_X1 U20521 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18410), .C1(
        n18411), .C2(n18413), .A(n21570), .ZN(n18400) );
  AOI21_X1 U20522 ( .B1(n18593), .B2(n20935), .A(n18400), .ZN(n18408) );
  NOR2_X1 U20523 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21555), .ZN(
        n18406) );
  INV_X1 U20524 ( .A(n21522), .ZN(n18436) );
  NAND4_X1 U20525 ( .A1(n18548), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A4(n18401), .ZN(n18651) );
  NOR3_X1 U20526 ( .A1(n18436), .A2(n21543), .A3(n18651), .ZN(n18613) );
  NOR2_X1 U20527 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18402), .ZN(
        n18640) );
  INV_X1 U20528 ( .A(n18640), .ZN(n18652) );
  NOR2_X1 U20529 ( .A1(n18403), .A2(n18652), .ZN(n18614) );
  AOI22_X1 U20530 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18613), .B1(
        n18614), .B2(n21544), .ZN(n18404) );
  XOR2_X1 U20531 ( .A(n18405), .B(n18404), .Z(n21568) );
  AOI22_X1 U20532 ( .A1(n18748), .A2(n18406), .B1(n18661), .B2(n21568), .ZN(
        n18407) );
  OAI211_X1 U20533 ( .C1(n18422), .C2(n18409), .A(n18408), .B(n18407), .ZN(
        P3_U2815) );
  INV_X1 U20534 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n20943) );
  NOR2_X1 U20535 ( .A1(n11142), .A2(n20943), .ZN(n18420) );
  AOI211_X1 U20536 ( .C1(n18411), .C2(n20955), .A(n20966), .B(n18410), .ZN(
        n18419) );
  NOR2_X1 U20537 ( .A1(n18411), .A2(n20932), .ZN(n18412) );
  OR2_X1 U20538 ( .A1(n18601), .A2(n20757), .ZN(n18600) );
  OAI21_X1 U20539 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n18412), .A(
        n18600), .ZN(n20951) );
  OAI22_X1 U20540 ( .A1(n18413), .A2(n20955), .B1(n18571), .B2(n20951), .ZN(
        n18418) );
  AOI22_X1 U20541 ( .A1(n18548), .A2(n21752), .B1(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n21668), .ZN(n18414) );
  XNOR2_X1 U20542 ( .A(n18415), .B(n18414), .ZN(n21760) );
  OAI22_X1 U20543 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18416), .B1(
        n21760), .B2(n18675), .ZN(n18417) );
  NOR4_X1 U20544 ( .A1(n18420), .A2(n18419), .A3(n18418), .A4(n18417), .ZN(
        n18421) );
  OAI21_X1 U20545 ( .B1(n18422), .B2(n21752), .A(n18421), .ZN(P3_U2814) );
  NAND2_X1 U20546 ( .A1(n21732), .A2(n21522), .ZN(n21523) );
  NAND2_X1 U20547 ( .A1(n21522), .A2(n11416), .ZN(n21528) );
  AOI22_X1 U20548 ( .A1(n18672), .A2(n21523), .B1(n18748), .B2(n21528), .ZN(
        n18439) );
  NAND2_X1 U20549 ( .A1(n18399), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18628) );
  NOR2_X1 U20550 ( .A1(n20893), .A2(n18628), .ZN(n20902) );
  AOI21_X1 U20551 ( .B1(n20893), .B2(n18628), .A(n20902), .ZN(n20890) );
  NAND2_X1 U20552 ( .A1(n18399), .A2(n18549), .ZN(n18433) );
  OAI21_X1 U20553 ( .B1(n18399), .B2(n18715), .A(n18754), .ZN(n18423) );
  AOI21_X1 U20554 ( .B1(n18628), .B2(n18423), .A(n18730), .ZN(n18444) );
  NAND2_X1 U20555 ( .A1(n14606), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n21534) );
  OAI221_X1 U20556 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18433), .C1(
        n20893), .C2(n18444), .A(n21534), .ZN(n18424) );
  AOI21_X1 U20557 ( .B1(n18593), .B2(n20890), .A(n18424), .ZN(n18431) );
  NOR2_X1 U20558 ( .A1(n21513), .A2(n21763), .ZN(n21532) );
  NAND2_X1 U20559 ( .A1(n18548), .A2(n21532), .ZN(n18427) );
  OR2_X1 U20560 ( .A1(n18646), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18426) );
  OAI22_X1 U20561 ( .A1(n18425), .A2(n18427), .B1(n18426), .B2(n18652), .ZN(
        n18428) );
  XNOR2_X1 U20562 ( .A(n21762), .B(n18428), .ZN(n21533) );
  INV_X1 U20563 ( .A(n18645), .ZN(n18664) );
  NOR2_X1 U20564 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18664), .ZN(
        n18429) );
  AOI22_X1 U20565 ( .A1(n18661), .A2(n21533), .B1(n21532), .B2(n18429), .ZN(
        n18430) );
  OAI211_X1 U20566 ( .C1(n18439), .C2(n21762), .A(n18431), .B(n18430), .ZN(
        P3_U2818) );
  INV_X1 U20567 ( .A(n20902), .ZN(n18432) );
  AOI22_X1 U20568 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n20902), .B1(
        n18432), .B2(n18443), .ZN(n20908) );
  AOI211_X1 U20569 ( .C1(n20893), .C2(n18443), .A(n20900), .B(n18433), .ZN(
        n18435) );
  INV_X1 U20570 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n20914) );
  NOR2_X1 U20571 ( .A1(n11142), .A2(n20914), .ZN(n18434) );
  AOI211_X1 U20572 ( .C1(n18593), .C2(n20908), .A(n18435), .B(n18434), .ZN(
        n18442) );
  NOR2_X1 U20573 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18436), .ZN(
        n21761) );
  INV_X1 U20574 ( .A(n18651), .ZN(n18641) );
  AOI22_X1 U20575 ( .A1(n21522), .A2(n18641), .B1(n18437), .B2(n18640), .ZN(
        n18438) );
  XOR2_X1 U20576 ( .A(n18438), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .Z(
        n21771) );
  OAI22_X1 U20577 ( .A1(n21771), .A2(n18675), .B1(n18439), .B2(n21543), .ZN(
        n18440) );
  AOI21_X1 U20578 ( .B1(n21761), .B2(n18645), .A(n18440), .ZN(n18441) );
  OAI211_X1 U20579 ( .C1(n18444), .C2(n18443), .A(n18442), .B(n18441), .ZN(
        P3_U2817) );
  INV_X1 U20580 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n21679) );
  AOI21_X1 U20581 ( .B1(n18446), .B2(n11429), .A(n18445), .ZN(n18493) );
  XOR2_X1 U20582 ( .A(n21679), .B(n18493), .Z(n21582) );
  NOR2_X1 U20583 ( .A1(n18447), .A2(n18474), .ZN(n18524) );
  NOR2_X1 U20584 ( .A1(n21573), .A2(n11422), .ZN(n21408) );
  NOR2_X1 U20585 ( .A1(n21573), .A2(n21567), .ZN(n21407) );
  OAI22_X1 U20586 ( .A1(n21408), .A2(n18758), .B1(n21407), .B2(n18589), .ZN(
        n18466) );
  INV_X1 U20587 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n18480) );
  NAND2_X1 U20588 ( .A1(n18478), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18479) );
  AOI21_X1 U20589 ( .B1(n11315), .B2(n18479), .A(n18730), .ZN(n18448) );
  OAI21_X1 U20590 ( .B1(n18451), .B2(n18715), .A(n18448), .ZN(n18477) );
  AOI21_X1 U20591 ( .B1(n18562), .B2(n18480), .A(n18477), .ZN(n18458) );
  INV_X1 U20592 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18454) );
  NAND2_X1 U20593 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n18449), .ZN(
        n18450) );
  INV_X1 U20594 ( .A(n18485), .ZN(n18486) );
  AOI21_X1 U20595 ( .B1(n18454), .B2(n18450), .A(n18486), .ZN(n21027) );
  AOI22_X1 U20596 ( .A1(n21774), .A2(P3_REIP_REG_22__SCAN_IN), .B1(n18593), 
        .B2(n21027), .ZN(n18453) );
  INV_X1 U20597 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n21022) );
  AND2_X1 U20598 ( .A1(n18549), .A2(n18451), .ZN(n18461) );
  OAI221_X1 U20599 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C1(n18454), .C2(n21022), .A(
        n18461), .ZN(n18452) );
  OAI211_X1 U20600 ( .C1(n18458), .C2(n18454), .A(n18453), .B(n18452), .ZN(
        n18455) );
  AOI221_X1 U20601 ( .B1(n18524), .B2(n21679), .C1(n18466), .C2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n18455), .ZN(n18456) );
  OAI21_X1 U20602 ( .B1(n18675), .B2(n21582), .A(n18456), .ZN(P3_U2808) );
  INV_X1 U20603 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18465) );
  NAND2_X1 U20604 ( .A1(n21411), .A2(n18465), .ZN(n21415) );
  INV_X1 U20605 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n21023) );
  NOR2_X1 U20606 ( .A1(n11142), .A2(n21023), .ZN(n18460) );
  INV_X1 U20607 ( .A(n18449), .ZN(n18457) );
  OAI22_X1 U20608 ( .A1(n21022), .A2(n18457), .B1(n18449), .B2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n21011) );
  OAI22_X1 U20609 ( .A1(n18458), .A2(n21022), .B1(n18571), .B2(n21011), .ZN(
        n18459) );
  AOI211_X1 U20610 ( .C1(n18461), .C2(n21022), .A(n18460), .B(n18459), .ZN(
        n18468) );
  NOR2_X1 U20611 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18462) );
  AOI22_X1 U20612 ( .A1(n21411), .A2(n18463), .B1(n18462), .B2(n18469), .ZN(
        n18464) );
  XOR2_X1 U20613 ( .A(n18465), .B(n18464), .Z(n21402) );
  AOI22_X1 U20614 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18466), .B1(
        n18661), .B2(n21402), .ZN(n18467) );
  OAI211_X1 U20615 ( .C1(n18474), .C2(n21415), .A(n18468), .B(n18467), .ZN(
        P3_U2809) );
  AOI21_X1 U20616 ( .B1(n18548), .B2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n18469), .ZN(n18470) );
  AOI21_X1 U20617 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18471), .A(
        n18470), .ZN(n18472) );
  XOR2_X1 U20618 ( .A(n18473), .B(n18472), .Z(n21718) );
  NAND2_X1 U20619 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18473), .ZN(
        n21724) );
  OAI22_X1 U20620 ( .A1(n18675), .A2(n21718), .B1(n18474), .B2(n21724), .ZN(
        n18475) );
  AOI21_X1 U20621 ( .B1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n18476), .A(
        n18475), .ZN(n18483) );
  NAND2_X1 U20622 ( .A1(n21774), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n21721) );
  OAI221_X1 U20623 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18478), .C1(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n19639), .A(n18477), .ZN(
        n18482) );
  AOI21_X1 U20624 ( .B1(n18480), .B2(n18479), .A(n18449), .ZN(n21003) );
  OAI21_X1 U20625 ( .B1(n18593), .B2(n18562), .A(n21003), .ZN(n18481) );
  NAND4_X1 U20626 ( .A1(n18483), .A2(n21721), .A3(n18482), .A4(n18481), .ZN(
        P3_U2810) );
  NOR2_X1 U20627 ( .A1(n21682), .A2(n18589), .ZN(n18484) );
  NOR2_X1 U20628 ( .A1(n21683), .A2(n18758), .ZN(n18491) );
  AOI22_X1 U20629 ( .A1(n18484), .A2(n21407), .B1(n18491), .B2(n21408), .ZN(
        n18500) );
  AOI21_X1 U20630 ( .B1(n21041), .B2(n18485), .A(n18516), .ZN(n21040) );
  INV_X1 U20631 ( .A(n18740), .ZN(n18490) );
  OAI22_X1 U20632 ( .A1(n18504), .A2(n19551), .B1(n18486), .B2(n18754), .ZN(
        n18487) );
  NOR2_X1 U20633 ( .A1(n18730), .A2(n18487), .ZN(n18505) );
  AOI221_X1 U20634 ( .B1(n18488), .B2(n21041), .C1(n19551), .C2(n21041), .A(
        n18505), .ZN(n18489) );
  INV_X1 U20635 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n21036) );
  NOR2_X1 U20636 ( .A1(n11142), .A2(n21036), .ZN(n21688) );
  AOI211_X1 U20637 ( .C1(n21040), .C2(n18490), .A(n18489), .B(n21688), .ZN(
        n18499) );
  INV_X1 U20638 ( .A(n21682), .ZN(n18492) );
  AOI21_X1 U20639 ( .B1(n18492), .B2(n18672), .A(n18491), .ZN(n18527) );
  INV_X1 U20640 ( .A(n18527), .ZN(n18497) );
  OAI221_X1 U20641 ( .B1(n18494), .B2(n18548), .C1(n18494), .C2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n18493), .ZN(n18495) );
  XOR2_X1 U20642 ( .A(n18496), .B(n18495), .Z(n21689) );
  AOI22_X1 U20643 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n18497), .B1(
        n18661), .B2(n21689), .ZN(n18498) );
  OAI211_X1 U20644 ( .C1(n18500), .C2(n21679), .A(n18499), .B(n18498), .ZN(
        P3_U2807) );
  OAI21_X1 U20645 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n18502), .A(
        n18501), .ZN(n21591) );
  NAND2_X1 U20646 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n18516), .ZN(
        n18503) );
  AOI21_X1 U20647 ( .B1(n21064), .B2(n18503), .A(n18561), .ZN(n21062) );
  NAND2_X1 U20648 ( .A1(n18504), .A2(n18549), .ZN(n18519) );
  AOI221_X1 U20649 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C1(n21064), .C2(n21058), .A(
        n18519), .ZN(n18508) );
  OAI21_X1 U20650 ( .B1(n18529), .B2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n18505), .ZN(n18506) );
  INV_X1 U20651 ( .A(n18506), .ZN(n18518) );
  INV_X1 U20652 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n21074) );
  OAI22_X1 U20653 ( .A1(n18518), .A2(n21064), .B1(n11142), .B2(n21074), .ZN(
        n18507) );
  AOI211_X1 U20654 ( .C1(n21062), .C2(n18593), .A(n18508), .B(n18507), .ZN(
        n18515) );
  AOI21_X1 U20655 ( .B1(n21598), .B2(n18510), .A(n18509), .ZN(n21590) );
  AOI21_X1 U20656 ( .B1(n18548), .B2(n18512), .A(n18511), .ZN(n18513) );
  XOR2_X1 U20657 ( .A(n18513), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n21595) );
  AOI22_X1 U20658 ( .A1(n18672), .A2(n21590), .B1(n18661), .B2(n21595), .ZN(
        n18514) );
  OAI211_X1 U20659 ( .C1(n18758), .C2(n21591), .A(n18515), .B(n18514), .ZN(
        P3_U2805) );
  AOI22_X1 U20660 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n18516), .B1(
        n11345), .B2(n21058), .ZN(n21053) );
  NAND2_X1 U20661 ( .A1(n14606), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n18517) );
  OAI221_X1 U20662 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n18519), .C1(
        n21058), .C2(n18518), .A(n18517), .ZN(n18520) );
  AOI21_X1 U20663 ( .B1(n18593), .B2(n21053), .A(n18520), .ZN(n18526) );
  OAI21_X1 U20664 ( .B1(n18522), .B2(n21696), .A(n18521), .ZN(n21700) );
  NOR2_X1 U20665 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n21692), .ZN(
        n18523) );
  AOI22_X1 U20666 ( .A1(n18661), .A2(n21700), .B1(n18524), .B2(n18523), .ZN(
        n18525) );
  OAI211_X1 U20667 ( .C1(n18527), .C2(n21696), .A(n18526), .B(n18525), .ZN(
        P3_U2806) );
  OAI21_X1 U20668 ( .B1(n18550), .B2(n18715), .A(n18753), .ZN(n18528) );
  AOI21_X1 U20669 ( .B1(n11315), .B2(n14616), .A(n18528), .ZN(n18558) );
  OAI21_X1 U20670 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18529), .A(
        n18558), .ZN(n18545) );
  INV_X1 U20671 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n21676) );
  NOR2_X1 U20672 ( .A1(n11142), .A2(n21676), .ZN(n18533) );
  OAI211_X1 U20673 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(n18550), .B(n18549), .ZN(n18530) );
  NOR2_X1 U20674 ( .A1(n21093), .A2(n18560), .ZN(n18544) );
  OAI21_X1 U20675 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n18544), .A(
        n14619), .ZN(n21101) );
  OAI22_X1 U20676 ( .A1(n18531), .A2(n18530), .B1(n21101), .B2(n18571), .ZN(
        n18532) );
  AOI211_X1 U20677 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n18545), .A(
        n18533), .B(n18532), .ZN(n18543) );
  AOI22_X1 U20678 ( .A1(n18672), .A2(n21631), .B1(n18748), .B2(n21605), .ZN(
        n18566) );
  NAND2_X1 U20679 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18566), .ZN(
        n18552) );
  OAI211_X1 U20680 ( .C1(n18672), .C2(n18748), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18552), .ZN(n18542) );
  NAND2_X1 U20681 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21586) );
  NOR2_X1 U20682 ( .A1(n21586), .A2(n21598), .ZN(n21600) );
  NAND3_X1 U20683 ( .A1(n18534), .A2(n21600), .A3(n18607), .ZN(n18567) );
  NOR2_X1 U20684 ( .A1(n21599), .A2(n18567), .ZN(n18578) );
  INV_X1 U20685 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n18535) );
  NAND3_X1 U20686 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18578), .A3(
        n18535), .ZN(n18541) );
  AOI21_X1 U20687 ( .B1(n18548), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n18536), .ZN(n21673) );
  NOR2_X1 U20688 ( .A1(n18538), .A2(n18537), .ZN(n18547) );
  NAND2_X1 U20689 ( .A1(n18547), .A2(n18548), .ZN(n18546) );
  NAND2_X1 U20690 ( .A1(n21674), .A2(n18546), .ZN(n18539) );
  OAI211_X1 U20691 ( .C1(n21673), .C2(n18539), .A(n18661), .B(n21652), .ZN(
        n18540) );
  NAND4_X1 U20692 ( .A1(n18543), .A2(n18542), .A3(n18541), .A4(n18540), .ZN(
        P3_U2802) );
  AOI21_X1 U20693 ( .B1(n21093), .B2(n18560), .A(n18544), .ZN(n21092) );
  AOI22_X1 U20694 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n18545), .B1(
        n18593), .B2(n21092), .ZN(n18555) );
  OAI21_X1 U20695 ( .B1(n18548), .B2(n18547), .A(n18546), .ZN(n21622) );
  AND2_X1 U20696 ( .A1(n18550), .A2(n18549), .ZN(n18551) );
  AOI22_X1 U20697 ( .A1(n18661), .A2(n21622), .B1(n18551), .B2(n21093), .ZN(
        n18554) );
  OAI21_X1 U20698 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18578), .A(
        n18552), .ZN(n18553) );
  NAND2_X1 U20699 ( .A1(n21774), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n21623) );
  NAND4_X1 U20700 ( .A1(n18555), .A2(n18554), .A3(n18553), .A4(n21623), .ZN(
        P3_U2803) );
  OAI21_X1 U20701 ( .B1(n18557), .B2(n21599), .A(n18556), .ZN(n21608) );
  AOI221_X1 U20702 ( .B1(n18559), .B2(n11362), .C1(n19551), .C2(n11362), .A(
        n18558), .ZN(n18564) );
  OAI21_X1 U20703 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18561), .A(
        n18560), .ZN(n21080) );
  NAND2_X1 U20704 ( .A1(n21774), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n21610) );
  OAI221_X1 U20705 ( .B1(n21080), .B2(n18571), .C1(n21080), .C2(n18529), .A(
        n21610), .ZN(n18563) );
  AOI211_X1 U20706 ( .C1(n18661), .C2(n21608), .A(n18564), .B(n18563), .ZN(
        n18565) );
  OAI221_X1 U20707 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n18567), 
        .C1(n21599), .C2(n18566), .A(n18565), .ZN(P3_U2804) );
  AOI21_X1 U20708 ( .B1(n18569), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n18568), .ZN(n21651) );
  OAI22_X1 U20709 ( .A1(n21626), .A2(n18758), .B1(n21627), .B2(n18589), .ZN(
        n18577) );
  INV_X1 U20710 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n18572) );
  OAI21_X1 U20711 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n18591), .A(
        n18570), .ZN(n21130) );
  OAI22_X1 U20712 ( .A1(n18573), .A2(n18572), .B1(n18571), .B2(n21130), .ZN(
        n18576) );
  INV_X1 U20713 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n21152) );
  OAI22_X1 U20714 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n18574), .B1(
        n11142), .B2(n21152), .ZN(n18575) );
  AOI211_X1 U20715 ( .C1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n18577), .A(
        n18576), .B(n18575), .ZN(n18581) );
  INV_X1 U20716 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21643) );
  NAND3_X1 U20717 ( .A1(n18579), .A2(n18578), .A3(n21643), .ZN(n18580) );
  OAI211_X1 U20718 ( .C1(n21651), .C2(n18675), .A(n18581), .B(n18580), .ZN(
        P3_U2800) );
  INV_X2 U20719 ( .A(n11142), .ZN(n21774) );
  OAI21_X1 U20720 ( .B1(n18582), .B2(n19551), .A(n18592), .ZN(n18583) );
  AOI22_X1 U20721 ( .A1(n21774), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n18584), 
        .B2(n18583), .ZN(n18598) );
  INV_X1 U20722 ( .A(n21654), .ZN(n18585) );
  NOR2_X1 U20723 ( .A1(n18586), .A2(n18585), .ZN(n18587) );
  XOR2_X1 U20724 ( .A(n18587), .B(n21641), .Z(n21637) );
  OR2_X1 U20725 ( .A1(n21605), .A2(n21636), .ZN(n21655) );
  AOI211_X1 U20726 ( .C1(n21655), .C2(n21641), .A(n21626), .B(n18758), .ZN(
        n18588) );
  AOI21_X1 U20727 ( .B1(n18661), .B2(n21637), .A(n18588), .ZN(n18597) );
  NOR2_X1 U20728 ( .A1(n21636), .A2(n21631), .ZN(n21661) );
  NOR2_X1 U20729 ( .A1(n21627), .A2(n18589), .ZN(n18590) );
  OAI21_X1 U20730 ( .B1(n21661), .B2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n18590), .ZN(n18596) );
  AOI21_X1 U20731 ( .B1(n18592), .B2(n14619), .A(n18591), .ZN(n21118) );
  OAI21_X1 U20732 ( .B1(n18594), .B2(n18593), .A(n21118), .ZN(n18595) );
  NAND4_X1 U20733 ( .A1(n18598), .A2(n18597), .A3(n18596), .A4(n18595), .ZN(
        P3_U2801) );
  AOI21_X1 U20734 ( .B1(n20973), .B2(n18600), .A(n18599), .ZN(n20968) );
  OAI21_X1 U20735 ( .B1(n18601), .B2(n19551), .A(n20973), .ZN(n18602) );
  AOI22_X1 U20736 ( .A1(n20968), .A2(n18490), .B1(n18603), .B2(n18602), .ZN(
        n18610) );
  OAI21_X1 U20737 ( .B1(n18605), .B2(n21750), .A(n18604), .ZN(n21747) );
  AOI22_X1 U20738 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18606), .B1(
        n18661), .B2(n21747), .ZN(n18609) );
  NAND2_X1 U20739 ( .A1(n21774), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n21748) );
  NOR2_X1 U20740 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n21752), .ZN(
        n21746) );
  NAND2_X1 U20741 ( .A1(n18607), .A2(n21746), .ZN(n18608) );
  NAND4_X1 U20742 ( .A1(n18610), .A2(n18609), .A3(n21748), .A4(n18608), .ZN(
        P3_U2813) );
  OAI21_X1 U20743 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18611), .A(
        n21555), .ZN(n21549) );
  AOI21_X1 U20744 ( .B1(n21544), .B2(n18612), .A(n21565), .ZN(n21548) );
  NOR2_X1 U20745 ( .A1(n18614), .A2(n18613), .ZN(n18615) );
  XOR2_X1 U20746 ( .A(n18615), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(
        n21550) );
  INV_X1 U20747 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n20923) );
  NAND2_X1 U20748 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n20902), .ZN(
        n18617) );
  AOI21_X1 U20749 ( .B1(n20923), .B2(n18617), .A(n18616), .ZN(n20916) );
  INV_X1 U20750 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n20919) );
  NOR2_X1 U20751 ( .A1(n11142), .A2(n20919), .ZN(n21552) );
  AOI21_X1 U20752 ( .B1(n20916), .B2(n18490), .A(n21552), .ZN(n18622) );
  NAND3_X1 U20753 ( .A1(n18618), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A3(
        n19639), .ZN(n18680) );
  NOR2_X1 U20754 ( .A1(n18619), .A2(n18680), .ZN(n18630) );
  OAI221_X1 U20755 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n20900), .C1(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .C2(n18630), .A(n18620), .ZN(
        n18621) );
  OAI211_X1 U20756 ( .C1(n21550), .C2(n18675), .A(n18622), .B(n18621), .ZN(
        n18623) );
  AOI21_X1 U20757 ( .B1(n18672), .B2(n21548), .A(n18623), .ZN(n18624) );
  OAI21_X1 U20758 ( .B1(n18758), .B2(n21549), .A(n18624), .ZN(P3_U2816) );
  OAI22_X1 U20759 ( .A1(n21513), .A2(n18651), .B1(n18646), .B2(n18652), .ZN(
        n18625) );
  XOR2_X1 U20760 ( .A(n21763), .B(n18625), .Z(n21521) );
  AOI22_X1 U20761 ( .A1(n21509), .A2(n18672), .B1(n18748), .B2(n21397), .ZN(
        n18663) );
  INV_X1 U20762 ( .A(n18663), .ZN(n18644) );
  INV_X1 U20763 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n20878) );
  NOR2_X1 U20764 ( .A1(n11142), .A2(n20878), .ZN(n21518) );
  NOR2_X1 U20765 ( .A1(n18730), .A2(n18626), .ZN(n18695) );
  INV_X1 U20766 ( .A(n18695), .ZN(n18749) );
  INV_X1 U20767 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18636) );
  INV_X1 U20768 ( .A(n18680), .ZN(n18655) );
  NAND3_X1 U20769 ( .A1(n18656), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        n18655), .ZN(n18654) );
  NOR2_X1 U20770 ( .A1(n18636), .A2(n18654), .ZN(n18635) );
  AOI21_X1 U20771 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18749), .A(
        n18635), .ZN(n18629) );
  INV_X1 U20772 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n20841) );
  INV_X1 U20773 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20829) );
  NOR2_X1 U20774 ( .A1(n20829), .A2(n18627), .ZN(n20834) );
  NAND2_X1 U20775 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n20834), .ZN(
        n18679) );
  NOR2_X1 U20776 ( .A1(n20841), .A2(n18679), .ZN(n20848) );
  NAND2_X1 U20777 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n20848), .ZN(
        n20863) );
  NOR2_X1 U20778 ( .A1(n18636), .A2(n20863), .ZN(n20874) );
  OAI21_X1 U20779 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n20874), .A(
        n18628), .ZN(n20875) );
  OAI22_X1 U20780 ( .A1(n18630), .A2(n18629), .B1(n18740), .B2(n20875), .ZN(
        n18631) );
  AOI211_X1 U20781 ( .C1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n18644), .A(
        n21518), .B(n18631), .ZN(n18634) );
  INV_X1 U20782 ( .A(n21513), .ZN(n21517) );
  INV_X1 U20783 ( .A(n21532), .ZN(n18632) );
  OAI211_X1 U20784 ( .C1(n21517), .C2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n18632), .B(n18645), .ZN(n18633) );
  OAI211_X1 U20785 ( .C1(n21521), .C2(n18675), .A(n18634), .B(n18633), .ZN(
        P3_U2819) );
  AOI21_X1 U20786 ( .B1(n18636), .B2(n20863), .A(n20874), .ZN(n20867) );
  AOI211_X1 U20787 ( .C1(n18654), .C2(n18636), .A(n18695), .B(n18635), .ZN(
        n18637) );
  AOI21_X1 U20788 ( .B1(n20867), .B2(n18490), .A(n18637), .ZN(n18650) );
  AOI21_X1 U20789 ( .B1(n21668), .B2(n21798), .A(n18641), .ZN(n18638) );
  AOI21_X1 U20790 ( .B1(n21798), .B2(n18639), .A(n18638), .ZN(n18643) );
  AOI221_X1 U20791 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18641), .C1(
        n21798), .C2(n18640), .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n18642) );
  AOI21_X1 U20792 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n18643), .A(
        n18642), .ZN(n21773) );
  AOI22_X1 U20793 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18644), .B1(
        n18661), .B2(n21773), .ZN(n18649) );
  NAND2_X1 U20794 ( .A1(n21774), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n18648) );
  NAND3_X1 U20795 ( .A1(n21513), .A2(n18646), .A3(n18645), .ZN(n18647) );
  NAND4_X1 U20796 ( .A1(n18650), .A2(n18649), .A3(n18648), .A4(n18647), .ZN(
        P3_U2820) );
  NAND2_X1 U20797 ( .A1(n18652), .A2(n18651), .ZN(n18653) );
  XOR2_X1 U20798 ( .A(n18653), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(
        n21800) );
  INV_X1 U20799 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n21803) );
  NOR2_X1 U20800 ( .A1(n11142), .A2(n21803), .ZN(n18660) );
  INV_X1 U20801 ( .A(n18654), .ZN(n18658) );
  AOI22_X1 U20802 ( .A1(n18656), .A2(n18655), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18749), .ZN(n18657) );
  OAI21_X1 U20803 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n20848), .A(
        n20863), .ZN(n20850) );
  OAI22_X1 U20804 ( .A1(n18658), .A2(n18657), .B1(n18740), .B2(n20850), .ZN(
        n18659) );
  AOI211_X1 U20805 ( .C1(n18661), .C2(n21800), .A(n18660), .B(n18659), .ZN(
        n18662) );
  OAI221_X1 U20806 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18664), .C1(
        n21798), .C2(n18663), .A(n18662), .ZN(P3_U2821) );
  OAI21_X1 U20807 ( .B1(n18666), .B2(n18665), .A(n18425), .ZN(n21503) );
  AOI21_X1 U20808 ( .B1(n20841), .B2(n18679), .A(n20848), .ZN(n20836) );
  OAI21_X1 U20809 ( .B1(n18730), .B2(n18627), .A(n18749), .ZN(n18683) );
  NAND2_X1 U20810 ( .A1(n14606), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n21501) );
  OAI211_X1 U20811 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n20834), .A(
        n19639), .B(n18667), .ZN(n18668) );
  OAI211_X1 U20812 ( .C1(n20841), .C2(n18683), .A(n21501), .B(n18668), .ZN(
        n18669) );
  AOI21_X1 U20813 ( .B1(n20836), .B2(n18490), .A(n18669), .ZN(n18674) );
  AOI21_X1 U20814 ( .B1(n18671), .B2(n21495), .A(n18670), .ZN(n21494) );
  AOI22_X1 U20815 ( .A1(n18672), .A2(n21503), .B1(n18748), .B2(n21494), .ZN(
        n18673) );
  OAI211_X1 U20816 ( .C1(n18675), .C2(n21503), .A(n18674), .B(n18673), .ZN(
        P3_U2822) );
  NAND2_X1 U20817 ( .A1(n18677), .A2(n18676), .ZN(n18678) );
  XOR2_X1 U20818 ( .A(n18678), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n21487) );
  NOR2_X1 U20819 ( .A1(n18627), .A2(n20757), .ZN(n18687) );
  OAI21_X1 U20820 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18687), .A(
        n18679), .ZN(n20820) );
  OAI22_X1 U20821 ( .A1(n18740), .A2(n20820), .B1(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18680), .ZN(n18685) );
  OAI21_X1 U20822 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n18682), .A(
        n18681), .ZN(n21488) );
  OAI22_X1 U20823 ( .A1(n18757), .A2(n21488), .B1(n20829), .B2(n18683), .ZN(
        n18684) );
  AOI211_X1 U20824 ( .C1(n14606), .C2(P3_REIP_REG_7__SCAN_IN), .A(n18685), .B(
        n18684), .ZN(n18686) );
  OAI21_X1 U20825 ( .B1(n18758), .B2(n21487), .A(n18686), .ZN(P3_U2823) );
  AND2_X1 U20826 ( .A1(n18618), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20809) );
  INV_X1 U20827 ( .A(n18687), .ZN(n20818) );
  OAI21_X1 U20828 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n20809), .A(
        n20818), .ZN(n20812) );
  NAND2_X1 U20829 ( .A1(n18618), .A2(n19639), .ZN(n18691) );
  OAI21_X1 U20830 ( .B1(n18690), .B2(n18689), .A(n18688), .ZN(n21484) );
  OAI22_X1 U20831 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18691), .B1(
        n18757), .B2(n21484), .ZN(n18692) );
  AOI21_X1 U20832 ( .B1(n21774), .B2(P3_REIP_REG_6__SCAN_IN), .A(n18692), .ZN(
        n18697) );
  AOI21_X1 U20833 ( .B1(n21787), .B2(n18694), .A(n18693), .ZN(n21479) );
  AOI21_X1 U20834 ( .B1(n19639), .B2(n18618), .A(n18695), .ZN(n18704) );
  AOI22_X1 U20835 ( .A1(n18748), .A2(n21479), .B1(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18704), .ZN(n18696) );
  OAI211_X1 U20836 ( .C1(n18740), .C2(n20812), .A(n18697), .B(n18696), .ZN(
        P3_U2824) );
  OAI21_X1 U20837 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n18699), .A(
        n18698), .ZN(n21475) );
  AOI21_X1 U20838 ( .B1(n18702), .B2(n18701), .A(n18700), .ZN(n21473) );
  AOI22_X1 U20839 ( .A1(n14606), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n18748), 
        .B2(n21473), .ZN(n18706) );
  OAI21_X1 U20840 ( .B1(n18730), .B2(n20795), .A(n20793), .ZN(n18703) );
  OR2_X1 U20841 ( .A1(n20795), .A2(n20757), .ZN(n18718) );
  AOI21_X1 U20842 ( .B1(n20793), .B2(n18718), .A(n20809), .ZN(n20797) );
  AOI22_X1 U20843 ( .A1(n18704), .A2(n18703), .B1(n20797), .B2(n18490), .ZN(
        n18705) );
  OAI211_X1 U20844 ( .C1(n18757), .C2(n21475), .A(n18706), .B(n18705), .ZN(
        P3_U2825) );
  OAI21_X1 U20845 ( .B1(n18709), .B2(n18708), .A(n18707), .ZN(n21458) );
  AOI21_X1 U20846 ( .B1(n18712), .B2(n18711), .A(n18710), .ZN(n21459) );
  NAND2_X1 U20847 ( .A1(n21774), .A2(P3_REIP_REG_4__SCAN_IN), .ZN(n21461) );
  INV_X1 U20848 ( .A(n21461), .ZN(n18714) );
  NOR3_X1 U20849 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18717), .A3(
        n19551), .ZN(n18713) );
  AOI211_X1 U20850 ( .C1(n18748), .C2(n21459), .A(n18714), .B(n18713), .ZN(
        n18720) );
  OAI21_X1 U20851 ( .B1(n18716), .B2(n18715), .A(n18753), .ZN(n18731) );
  NOR2_X1 U20852 ( .A1(n18717), .A2(n20757), .ZN(n18721) );
  OAI21_X1 U20853 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18721), .A(
        n18718), .ZN(n20782) );
  INV_X1 U20854 ( .A(n20782), .ZN(n20779) );
  AOI22_X1 U20855 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18731), .B1(
        n20779), .B2(n18490), .ZN(n18719) );
  OAI211_X1 U20856 ( .C1(n18757), .C2(n21458), .A(n18720), .B(n18719), .ZN(
        P3_U2826) );
  NAND2_X1 U20857 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20767) );
  INV_X1 U20858 ( .A(n20767), .ZN(n18722) );
  INV_X1 U20859 ( .A(n18721), .ZN(n20777) );
  OAI21_X1 U20860 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18722), .A(
        n20777), .ZN(n20769) );
  AOI21_X1 U20861 ( .B1(n18725), .B2(n18724), .A(n18723), .ZN(n21442) );
  OAI21_X1 U20862 ( .B1(n18728), .B2(n18727), .A(n18726), .ZN(n21453) );
  OAI22_X1 U20863 ( .A1(n11142), .A2(n21440), .B1(n18757), .B2(n21453), .ZN(
        n18729) );
  AOI21_X1 U20864 ( .B1(n18748), .B2(n21442), .A(n18729), .ZN(n18733) );
  INV_X1 U20865 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n20764) );
  NOR2_X1 U20866 ( .A1(n18730), .A2(n20764), .ZN(n18744) );
  OAI21_X1 U20867 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18744), .A(
        n18731), .ZN(n18732) );
  OAI211_X1 U20868 ( .C1(n18740), .C2(n20769), .A(n18733), .B(n18732), .ZN(
        P3_U2827) );
  AOI21_X1 U20869 ( .B1(n18736), .B2(n18735), .A(n18734), .ZN(n21431) );
  NAND2_X1 U20870 ( .A1(n21774), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n21437) );
  INV_X1 U20871 ( .A(n21437), .ZN(n18742) );
  OAI21_X1 U20872 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n20767), .ZN(n20758) );
  OAI21_X1 U20873 ( .B1(n18739), .B2(n18738), .A(n18737), .ZN(n21439) );
  OAI22_X1 U20874 ( .A1(n18740), .A2(n20758), .B1(n18757), .B2(n21439), .ZN(
        n18741) );
  AOI211_X1 U20875 ( .C1(n18748), .C2(n21431), .A(n18742), .B(n18741), .ZN(
        n18743) );
  OAI221_X1 U20876 ( .B1(n18744), .B2(n20764), .C1(n18744), .C2(n19551), .A(
        n18743), .ZN(P3_U2828) );
  OAI21_X1 U20877 ( .B1(n18746), .B2(n18752), .A(n18745), .ZN(n21424) );
  NAND2_X1 U20878 ( .A1(n21508), .A2(n21350), .ZN(n18747) );
  XNOR2_X1 U20879 ( .A(n18747), .B(n18746), .ZN(n21422) );
  AOI22_X1 U20880 ( .A1(n14606), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n18748), 
        .B2(n21422), .ZN(n18751) );
  AOI22_X1 U20881 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18749), .B1(
        n18490), .B2(n20757), .ZN(n18750) );
  OAI211_X1 U20882 ( .C1(n18757), .C2(n21424), .A(n18751), .B(n18750), .ZN(
        P3_U2829) );
  AOI21_X1 U20883 ( .B1(n21350), .B2(n21508), .A(n18752), .ZN(n21421) );
  INV_X1 U20884 ( .A(n21421), .ZN(n21420) );
  NAND3_X1 U20885 ( .A1(n21354), .A2(n18754), .A3(n18753), .ZN(n18755) );
  AOI22_X1 U20886 ( .A1(n21774), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18755), .ZN(n18756) );
  OAI221_X1 U20887 ( .B1(n21421), .B2(n18758), .C1(n21420), .C2(n18757), .A(
        n18756), .ZN(P3_U2830) );
  INV_X1 U20888 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21837) );
  NAND2_X1 U20889 ( .A1(n21837), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19358) );
  INV_X1 U20890 ( .A(n19358), .ZN(n19359) );
  NAND2_X1 U20891 ( .A1(n21834), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19341) );
  NOR2_X1 U20892 ( .A1(n19359), .A2(n19342), .ZN(n18759) );
  OAI22_X1 U20893 ( .A1(n18761), .A2(n21837), .B1(n18760), .B2(n18759), .ZN(
        P3_U2866) );
  OAI21_X1 U20894 ( .B1(n18762), .B2(n19355), .A(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18763) );
  OAI21_X1 U20895 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18764), .A(
        n18763), .ZN(P3_U2864) );
  NOR4_X1 U20896 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18768) );
  NOR4_X1 U20897 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18767) );
  NOR4_X1 U20898 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18766) );
  NOR4_X1 U20899 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18765) );
  NAND4_X1 U20900 ( .A1(n18768), .A2(n18767), .A3(n18766), .A4(n18765), .ZN(
        n18774) );
  NOR4_X1 U20901 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n18772) );
  AOI211_X1 U20902 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_31__SCAN_IN), .B(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n18771) );
  NOR4_X1 U20903 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18770) );
  NOR4_X1 U20904 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18769) );
  NAND4_X1 U20905 ( .A1(n18772), .A2(n18771), .A3(n18770), .A4(n18769), .ZN(
        n18773) );
  NOR2_X1 U20906 ( .A1(n18774), .A2(n18773), .ZN(n18782) );
  INV_X1 U20907 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18776) );
  OAI21_X1 U20908 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18782), .ZN(n18775) );
  OAI21_X1 U20909 ( .B1(n18782), .B2(n18776), .A(n18775), .ZN(P3_U3293) );
  INV_X1 U20910 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n21416) );
  NOR2_X1 U20911 ( .A1(P3_DATAWIDTH_REG_1__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18780) );
  AOI21_X1 U20912 ( .B1(P3_DATAWIDTH_REG_0__SCAN_IN), .B2(n21416), .A(n18780), 
        .ZN(n18779) );
  INV_X1 U20913 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n21429) );
  NAND2_X1 U20914 ( .A1(n18782), .A2(n21429), .ZN(n18786) );
  OAI21_X1 U20915 ( .B1(n21416), .B2(n21429), .A(n18782), .ZN(n18777) );
  OAI21_X1 U20916 ( .B1(P3_BYTEENABLE_REG_2__SCAN_IN), .B2(n18782), .A(n18777), 
        .ZN(n18778) );
  OAI21_X1 U20917 ( .B1(n18779), .B2(n18786), .A(n18778), .ZN(P3_U3292) );
  OAI21_X1 U20918 ( .B1(n18782), .B2(P3_BYTEENABLE_REG_1__SCAN_IN), .A(n18786), 
        .ZN(n18781) );
  NAND3_X1 U20919 ( .A1(n18782), .A2(n18780), .A3(n21416), .ZN(n18784) );
  NAND2_X1 U20920 ( .A1(n18781), .A2(n18784), .ZN(P3_U2638) );
  INV_X1 U20921 ( .A(n18782), .ZN(n18783) );
  NAND2_X1 U20922 ( .A1(P3_BYTEENABLE_REG_3__SCAN_IN), .A2(n18783), .ZN(n18785) );
  OAI211_X1 U20923 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(n18786), .A(n18785), 
        .B(n18784), .ZN(P3_U2639) );
  INV_X1 U20924 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18787) );
  INV_X1 U20925 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n18844) );
  AOI22_X1 U20926 ( .A1(n22303), .A2(n18787), .B1(n18844), .B2(n18843), .ZN(
        P3_U3297) );
  INV_X1 U20927 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18788) );
  AOI22_X1 U20928 ( .A1(n22303), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18788), 
        .B2(n18843), .ZN(P3_U3294) );
  OAI21_X1 U20929 ( .B1(n22340), .B2(P3_D_C_N_REG_SCAN_IN), .A(n18843), .ZN(
        n18789) );
  OAI21_X1 U20930 ( .B1(P3_CODEFETCH_REG_SCAN_IN), .B2(n18843), .A(n18789), 
        .ZN(P3_U2635) );
  INV_X1 U20931 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n21198) );
  AOI22_X1 U20932 ( .A1(n21805), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18817), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18790) );
  OAI21_X1 U20933 ( .B1(n21198), .B2(n18806), .A(n18790), .ZN(P3_U2767) );
  INV_X1 U20934 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n20709) );
  AOI22_X1 U20935 ( .A1(n21805), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18817), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18791) );
  OAI21_X1 U20936 ( .B1(n20709), .B2(n18806), .A(n18791), .ZN(P3_U2766) );
  INV_X1 U20937 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n21222) );
  AOI22_X1 U20938 ( .A1(n21805), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18817), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18792) );
  OAI21_X1 U20939 ( .B1(n21222), .B2(n18806), .A(n18792), .ZN(P3_U2765) );
  INV_X1 U20940 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n20712) );
  AOI22_X1 U20941 ( .A1(n21805), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18817), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18793) );
  OAI21_X1 U20942 ( .B1(n20712), .B2(n18806), .A(n18793), .ZN(P3_U2764) );
  INV_X1 U20943 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n21199) );
  AOI22_X1 U20944 ( .A1(n21805), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18817), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18794) );
  OAI21_X1 U20945 ( .B1(n21199), .B2(n18806), .A(n18794), .ZN(P3_U2763) );
  INV_X1 U20946 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n20715) );
  AOI22_X1 U20947 ( .A1(n21805), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18817), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18795) );
  OAI21_X1 U20948 ( .B1(n20715), .B2(n18806), .A(n18795), .ZN(P3_U2762) );
  INV_X1 U20949 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n21200) );
  AOI22_X1 U20950 ( .A1(n21805), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18817), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18796) );
  OAI21_X1 U20951 ( .B1(n21200), .B2(n18806), .A(n18796), .ZN(P3_U2761) );
  INV_X1 U20952 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n20718) );
  AOI22_X1 U20953 ( .A1(n21805), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18817), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18797) );
  OAI21_X1 U20954 ( .B1(n20718), .B2(n18806), .A(n18797), .ZN(P3_U2760) );
  INV_X1 U20955 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n21330) );
  AOI22_X1 U20956 ( .A1(n18824), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18817), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18798) );
  OAI21_X1 U20957 ( .B1(n21330), .B2(n18806), .A(n18798), .ZN(P3_U2759) );
  INV_X1 U20958 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n21190) );
  AOI22_X1 U20959 ( .A1(n21805), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18817), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18799) );
  OAI21_X1 U20960 ( .B1(n21190), .B2(n18806), .A(n18799), .ZN(P3_U2758) );
  INV_X1 U20961 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n20722) );
  AOI22_X1 U20962 ( .A1(n21805), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18817), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18800) );
  OAI21_X1 U20963 ( .B1(n20722), .B2(n18806), .A(n18800), .ZN(P3_U2757) );
  INV_X1 U20964 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n21179) );
  AOI22_X1 U20965 ( .A1(n21805), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18817), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18801) );
  OAI21_X1 U20966 ( .B1(n21179), .B2(n18806), .A(n18801), .ZN(P3_U2756) );
  INV_X1 U20967 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n20725) );
  AOI22_X1 U20968 ( .A1(n21805), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18817), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18802) );
  OAI21_X1 U20969 ( .B1(n20725), .B2(n18806), .A(n18802), .ZN(P3_U2755) );
  INV_X1 U20970 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n20727) );
  AOI22_X1 U20971 ( .A1(n21805), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18817), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18803) );
  OAI21_X1 U20972 ( .B1(n20727), .B2(n18806), .A(n18803), .ZN(P3_U2754) );
  INV_X1 U20973 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n20730) );
  AOI22_X1 U20974 ( .A1(n21805), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18817), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18804) );
  OAI21_X1 U20975 ( .B1(n20730), .B2(n18806), .A(n18804), .ZN(P3_U2753) );
  INV_X1 U20976 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n21325) );
  AOI22_X1 U20977 ( .A1(n21805), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18817), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18805) );
  OAI21_X1 U20978 ( .B1(n21325), .B2(n18806), .A(n18805), .ZN(P3_U2752) );
  INV_X1 U20979 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n20685) );
  AOI22_X1 U20980 ( .A1(n21805), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18817), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18809) );
  OAI21_X1 U20981 ( .B1(n20685), .B2(n18826), .A(n18809), .ZN(P3_U2751) );
  INV_X1 U20982 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n20687) );
  AOI22_X1 U20983 ( .A1(n21805), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18817), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18810) );
  OAI21_X1 U20984 ( .B1(n20687), .B2(n18826), .A(n18810), .ZN(P3_U2750) );
  INV_X1 U20985 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n21255) );
  AOI22_X1 U20986 ( .A1(n21805), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18817), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18811) );
  OAI21_X1 U20987 ( .B1(n21255), .B2(n18826), .A(n18811), .ZN(P3_U2749) );
  INV_X1 U20988 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n21229) );
  AOI22_X1 U20989 ( .A1(n21805), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18817), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18812) );
  OAI21_X1 U20990 ( .B1(n21229), .B2(n18826), .A(n18812), .ZN(P3_U2748) );
  INV_X1 U20991 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n21242) );
  AOI22_X1 U20992 ( .A1(n18824), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18817), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18813) );
  OAI21_X1 U20993 ( .B1(n21242), .B2(n18826), .A(n18813), .ZN(P3_U2747) );
  INV_X1 U20994 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n21236) );
  AOI22_X1 U20995 ( .A1(n18824), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18817), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18814) );
  OAI21_X1 U20996 ( .B1(n21236), .B2(n18826), .A(n18814), .ZN(P3_U2746) );
  INV_X1 U20997 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n21265) );
  AOI22_X1 U20998 ( .A1(n18824), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18817), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18815) );
  OAI21_X1 U20999 ( .B1(n21265), .B2(n18826), .A(n18815), .ZN(P3_U2745) );
  INV_X1 U21000 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n20694) );
  AOI22_X1 U21001 ( .A1(n18824), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18817), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18816) );
  OAI21_X1 U21002 ( .B1(n20694), .B2(n18826), .A(n18816), .ZN(P3_U2744) );
  INV_X1 U21003 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n20696) );
  AOI22_X1 U21004 ( .A1(n21805), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18817), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18818) );
  OAI21_X1 U21005 ( .B1(n20696), .B2(n18826), .A(n18818), .ZN(P3_U2743) );
  INV_X1 U21006 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n20698) );
  AOI22_X1 U21007 ( .A1(n18824), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18817), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18819) );
  OAI21_X1 U21008 ( .B1(n20698), .B2(n18826), .A(n18819), .ZN(P3_U2742) );
  INV_X1 U21009 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n21274) );
  AOI22_X1 U21010 ( .A1(n18824), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18817), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18820) );
  OAI21_X1 U21011 ( .B1(n21274), .B2(n18826), .A(n18820), .ZN(P3_U2741) );
  INV_X1 U21012 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n20701) );
  AOI22_X1 U21013 ( .A1(n18824), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18817), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18821) );
  OAI21_X1 U21014 ( .B1(n20701), .B2(n18826), .A(n18821), .ZN(P3_U2740) );
  INV_X1 U21015 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n21290) );
  AOI22_X1 U21016 ( .A1(n18824), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18817), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18822) );
  OAI21_X1 U21017 ( .B1(n21290), .B2(n18826), .A(n18822), .ZN(P3_U2739) );
  INV_X1 U21018 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n20704) );
  AOI22_X1 U21019 ( .A1(n18824), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18817), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18823) );
  OAI21_X1 U21020 ( .B1(n20704), .B2(n18826), .A(n18823), .ZN(P3_U2738) );
  INV_X1 U21021 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n20706) );
  AOI22_X1 U21022 ( .A1(n18824), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18817), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18825) );
  OAI21_X1 U21023 ( .B1(n20706), .B2(n18826), .A(n18825), .ZN(P3_U2737) );
  NOR2_X1 U21024 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(n18827), .ZN(n18828) );
  NOR2_X1 U21025 ( .A1(n22303), .A2(n18828), .ZN(P3_U2633) );
  NOR2_X1 U21026 ( .A1(n18843), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18835) );
  INV_X1 U21027 ( .A(n18835), .ZN(n18841) );
  INV_X1 U21028 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n20755) );
  INV_X1 U21029 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n20361) );
  OAI222_X1 U21030 ( .A1(n18841), .A2(n20755), .B1(n20361), .B2(n22303), .C1(
        n21429), .C2(n18840), .ZN(P3_U3032) );
  INV_X1 U21031 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n20363) );
  OAI222_X1 U21032 ( .A1(n18841), .A2(n21440), .B1(n20363), .B2(n22303), .C1(
        n20755), .C2(n18840), .ZN(P3_U3033) );
  INV_X1 U21033 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n20790) );
  INV_X1 U21034 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n20365) );
  OAI222_X1 U21035 ( .A1(n18841), .A2(n20790), .B1(n20365), .B2(n22303), .C1(
        n21440), .C2(n18840), .ZN(P3_U3034) );
  INV_X1 U21036 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n20367) );
  OAI222_X1 U21037 ( .A1(n18841), .A2(n21464), .B1(n20367), .B2(n22303), .C1(
        n20790), .C2(n18840), .ZN(P3_U3035) );
  INV_X1 U21038 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n21476) );
  INV_X1 U21039 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n20369) );
  OAI222_X1 U21040 ( .A1(n18841), .A2(n21476), .B1(n20369), .B2(n22303), .C1(
        n21464), .C2(n18840), .ZN(P3_U3036) );
  INV_X1 U21041 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n20839) );
  INV_X1 U21042 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n20371) );
  OAI222_X1 U21043 ( .A1(n18841), .A2(n20839), .B1(n20371), .B2(n22303), .C1(
        n21476), .C2(n18840), .ZN(P3_U3037) );
  AOI22_X1 U21044 ( .A1(n18835), .A2(P3_REIP_REG_8__SCAN_IN), .B1(
        P3_ADDRESS_REG_6__SCAN_IN), .B2(n18843), .ZN(n18829) );
  OAI21_X1 U21045 ( .B1(n18840), .B2(n20839), .A(n18829), .ZN(P3_U3038) );
  AOI22_X1 U21046 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n18837), .B1(
        P3_ADDRESS_REG_7__SCAN_IN), .B2(n18843), .ZN(n18830) );
  OAI21_X1 U21047 ( .B1(n21803), .B2(n18841), .A(n18830), .ZN(P3_U3039) );
  AOI22_X1 U21048 ( .A1(n18835), .A2(P3_REIP_REG_10__SCAN_IN), .B1(
        P3_ADDRESS_REG_8__SCAN_IN), .B2(n18843), .ZN(n18831) );
  OAI21_X1 U21049 ( .B1(n18840), .B2(n21803), .A(n18831), .ZN(P3_U3040) );
  AOI22_X1 U21050 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n18837), .B1(
        P3_ADDRESS_REG_9__SCAN_IN), .B2(n18843), .ZN(n18832) );
  OAI21_X1 U21051 ( .B1(n20878), .B2(n18841), .A(n18832), .ZN(P3_U3041) );
  INV_X1 U21052 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n20377) );
  INV_X1 U21053 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n20898) );
  OAI222_X1 U21054 ( .A1(n20878), .A2(n18840), .B1(n20377), .B2(n22303), .C1(
        n20898), .C2(n18841), .ZN(P3_U3042) );
  INV_X1 U21055 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n20379) );
  OAI222_X1 U21056 ( .A1(n18841), .A2(n20914), .B1(n20379), .B2(n22303), .C1(
        n20898), .C2(n18840), .ZN(P3_U3043) );
  INV_X1 U21057 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n20381) );
  OAI222_X1 U21058 ( .A1(n18841), .A2(n20919), .B1(n20381), .B2(n22303), .C1(
        n20914), .C2(n18840), .ZN(P3_U3044) );
  INV_X1 U21059 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n20941) );
  INV_X1 U21060 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n20383) );
  OAI222_X1 U21061 ( .A1(n18841), .A2(n20941), .B1(n20383), .B2(n22303), .C1(
        n20919), .C2(n18840), .ZN(P3_U3045) );
  INV_X1 U21062 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n20385) );
  OAI222_X1 U21063 ( .A1(n18841), .A2(n20943), .B1(n20385), .B2(n22303), .C1(
        n20941), .C2(n18840), .ZN(P3_U3046) );
  INV_X1 U21064 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n20960) );
  INV_X1 U21065 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n20387) );
  OAI222_X1 U21066 ( .A1(n18841), .A2(n20960), .B1(n20387), .B2(n22303), .C1(
        n20943), .C2(n18840), .ZN(P3_U3047) );
  AOI22_X1 U21067 ( .A1(n18835), .A2(P3_REIP_REG_18__SCAN_IN), .B1(
        P3_ADDRESS_REG_16__SCAN_IN), .B2(n18843), .ZN(n18833) );
  OAI21_X1 U21068 ( .B1(n18840), .B2(n20960), .A(n18833), .ZN(P3_U3048) );
  AOI22_X1 U21069 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n18837), .B1(
        P3_ADDRESS_REG_17__SCAN_IN), .B2(n18843), .ZN(n18834) );
  OAI21_X1 U21070 ( .B1(n20998), .B2(n18841), .A(n18834), .ZN(P3_U3049) );
  INV_X1 U21071 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n21009) );
  INV_X1 U21072 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n20391) );
  OAI222_X1 U21073 ( .A1(n18841), .A2(n21009), .B1(n20391), .B2(n22303), .C1(
        n20998), .C2(n18840), .ZN(P3_U3050) );
  INV_X1 U21074 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n20393) );
  OAI222_X1 U21075 ( .A1(n21009), .A2(n18840), .B1(n20393), .B2(n22303), .C1(
        n21023), .C2(n18841), .ZN(P3_U3051) );
  INV_X1 U21076 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n21033) );
  INV_X1 U21077 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n20395) );
  OAI222_X1 U21078 ( .A1(n18841), .A2(n21033), .B1(n20395), .B2(n22303), .C1(
        n21023), .C2(n18840), .ZN(P3_U3052) );
  INV_X1 U21079 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n20397) );
  OAI222_X1 U21080 ( .A1(n18841), .A2(n21036), .B1(n20397), .B2(n22303), .C1(
        n21033), .C2(n18840), .ZN(P3_U3053) );
  INV_X1 U21081 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n21702) );
  INV_X1 U21082 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n20399) );
  OAI222_X1 U21083 ( .A1(n18841), .A2(n21702), .B1(n20399), .B2(n22303), .C1(
        n21036), .C2(n18840), .ZN(P3_U3054) );
  INV_X1 U21084 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n20401) );
  OAI222_X1 U21085 ( .A1(n18841), .A2(n21074), .B1(n20401), .B2(n22303), .C1(
        n21702), .C2(n18840), .ZN(P3_U3055) );
  AOI22_X1 U21086 ( .A1(n18835), .A2(P3_REIP_REG_26__SCAN_IN), .B1(
        P3_ADDRESS_REG_24__SCAN_IN), .B2(n18843), .ZN(n18836) );
  OAI21_X1 U21087 ( .B1(n18840), .B2(n21074), .A(n18836), .ZN(P3_U3056) );
  INV_X1 U21088 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18839) );
  AOI22_X1 U21089 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n18837), .B1(
        P3_ADDRESS_REG_25__SCAN_IN), .B2(n18843), .ZN(n18838) );
  OAI21_X1 U21090 ( .B1(n18839), .B2(n18841), .A(n18838), .ZN(P3_U3057) );
  INV_X1 U21091 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n20405) );
  OAI222_X1 U21092 ( .A1(n18841), .A2(n21676), .B1(n20405), .B2(n22303), .C1(
        n18839), .C2(n18840), .ZN(P3_U3058) );
  INV_X1 U21093 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n20407) );
  INV_X1 U21094 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n21124) );
  OAI222_X1 U21095 ( .A1(n21676), .A2(n18840), .B1(n20407), .B2(n22303), .C1(
        n21124), .C2(n18841), .ZN(P3_U3059) );
  INV_X1 U21096 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n20409) );
  OAI222_X1 U21097 ( .A1(n18841), .A2(n21152), .B1(n20409), .B2(n22303), .C1(
        n21124), .C2(n18840), .ZN(P3_U3060) );
  INV_X1 U21098 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n21153) );
  INV_X1 U21099 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n20412) );
  OAI222_X1 U21100 ( .A1(n18841), .A2(n21153), .B1(n20412), .B2(n22303), .C1(
        n21152), .C2(n18840), .ZN(P3_U3061) );
  OAI22_X1 U21101 ( .A1(n18843), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n22303), .ZN(n18842) );
  INV_X1 U21102 ( .A(n18842), .ZN(P3_U3277) );
  MUX2_X1 U21103 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .B(P3_BE_N_REG_1__SCAN_IN), .S(n18843), .Z(P3_U3276) );
  MUX2_X1 U21104 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .B(P3_BE_N_REG_2__SCAN_IN), .S(n18843), .Z(P3_U3275) );
  MUX2_X1 U21105 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .B(P3_BE_N_REG_3__SCAN_IN), .S(n18843), .Z(P3_U3274) );
  NOR4_X1 U21106 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_BE_N_REG_2__SCAN_IN), .A4(P3_BE_N_REG_0__SCAN_IN), .ZN(n18846)
         );
  NOR4_X1 U21107 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(P3_D_C_N_REG_SCAN_IN), .A3(
        P3_W_R_N_REG_SCAN_IN), .A4(n18844), .ZN(n18845) );
  INV_X2 U21108 ( .A(n19593), .ZN(U215) );
  NAND3_X1 U21109 ( .A1(n18846), .A2(n18845), .A3(U215), .ZN(U213) );
  NOR2_X1 U21110 ( .A1(n22321), .A2(n19833), .ZN(n18850) );
  NAND3_X1 U21111 ( .A1(n22332), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n11785), 
        .ZN(n18848) );
  OAI21_X1 U21112 ( .B1(n22332), .B2(n22292), .A(n11768), .ZN(n18847) );
  MUX2_X1 U21113 ( .A(n18848), .B(n18847), .S(n14673), .Z(n18849) );
  OAI21_X1 U21114 ( .B1(n18850), .B2(n19282), .A(n18849), .ZN(n18856) );
  NAND4_X1 U21115 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .A3(n19270), .A4(n19281), .ZN(n18851) );
  OAI211_X1 U21116 ( .C1(n18854), .C2(n18853), .A(n18852), .B(n18851), .ZN(
        n18855) );
  MUX2_X1 U21117 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .B(n18856), .S(n18855), 
        .Z(P2_U3610) );
  INV_X1 U21118 ( .A(n18857), .ZN(n18869) );
  INV_X1 U21119 ( .A(n18858), .ZN(n19174) );
  INV_X1 U21120 ( .A(n18859), .ZN(n18860) );
  OAI22_X1 U21121 ( .A1(n19133), .A2(n19179), .B1(n19149), .B2(n18860), .ZN(
        n18864) );
  OAI22_X1 U21122 ( .A1(n19153), .A2(n18862), .B1(n18861), .B2(n19151), .ZN(
        n18863) );
  AOI211_X1 U21123 ( .C1(n19174), .C2(n19160), .A(n18864), .B(n18863), .ZN(
        n18868) );
  NOR2_X1 U21124 ( .A1(n19121), .A2(n18865), .ZN(n18866) );
  AOI21_X1 U21125 ( .B1(n18880), .B2(n19915), .A(n18866), .ZN(n18867) );
  OAI211_X1 U21126 ( .C1(n19267), .C2(n18869), .A(n18868), .B(n18867), .ZN(
        P2_U2855) );
  NAND2_X1 U21127 ( .A1(n19127), .A2(n19015), .ZN(n19050) );
  OAI22_X1 U21128 ( .A1(n19153), .A2(n18871), .B1(n18870), .B2(n19151), .ZN(
        n18875) );
  OAI22_X1 U21129 ( .A1(n19133), .A2(n18873), .B1(n19149), .B2(n18872), .ZN(
        n18874) );
  NOR2_X1 U21130 ( .A1(n18875), .A2(n18874), .ZN(n18876) );
  OAI21_X1 U21131 ( .B1(n18877), .B2(n19121), .A(n18876), .ZN(n18878) );
  AOI21_X1 U21132 ( .B1(n19160), .B2(n18879), .A(n18878), .ZN(n18883) );
  AOI22_X1 U21133 ( .A1(n18881), .A2(n19127), .B1(n19913), .B2(n18880), .ZN(
        n18882) );
  OAI211_X1 U21134 ( .C1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n19050), .A(
        n18883), .B(n18882), .ZN(P2_U2854) );
  OAI22_X1 U21135 ( .A1(n12275), .A2(n19153), .B1(n12525), .B2(n19151), .ZN(
        n18884) );
  AOI211_X1 U21136 ( .C1(n19159), .C2(n19207), .A(n19213), .B(n18884), .ZN(
        n18896) );
  AOI22_X1 U21137 ( .A1(n19157), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n19136), .B2(n18885), .ZN(n18895) );
  OAI22_X1 U21138 ( .A1(n20013), .A2(n18886), .B1(n19098), .B2(n19201), .ZN(
        n18887) );
  INV_X1 U21139 ( .A(n18887), .ZN(n18894) );
  INV_X1 U21140 ( .A(n18888), .ZN(n18892) );
  NOR2_X1 U21141 ( .A1(n19015), .A2(n18889), .ZN(n18891) );
  AOI21_X1 U21142 ( .B1(n18892), .B2(n18891), .A(n19267), .ZN(n18890) );
  OAI21_X1 U21143 ( .B1(n18892), .B2(n18891), .A(n18890), .ZN(n18893) );
  NAND4_X1 U21144 ( .A1(n18896), .A2(n18895), .A3(n18894), .A4(n18893), .ZN(
        P2_U2851) );
  NAND2_X1 U21145 ( .A1(n19029), .A2(n18897), .ZN(n18899) );
  XOR2_X1 U21146 ( .A(n18899), .B(n18898), .Z(n18908) );
  INV_X1 U21147 ( .A(n18900), .ZN(n18901) );
  AOI22_X1 U21148 ( .A1(n19134), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n19136), 
        .B2(n18901), .ZN(n18902) );
  OAI211_X1 U21149 ( .C1(n12046), .C2(n19153), .A(n18902), .B(n18976), .ZN(
        n18906) );
  INV_X1 U21150 ( .A(n18903), .ZN(n18904) );
  OAI22_X1 U21151 ( .A1(n19098), .A2(n18904), .B1(n19133), .B2(n20017), .ZN(
        n18905) );
  AOI211_X1 U21152 ( .C1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n19157), .A(
        n18906), .B(n18905), .ZN(n18907) );
  OAI21_X1 U21153 ( .B1(n18908), .B2(n19267), .A(n18907), .ZN(P2_U2850) );
  NOR2_X1 U21154 ( .A1(n19015), .A2(n18909), .ZN(n18910) );
  XOR2_X1 U21155 ( .A(n18911), .B(n18910), .Z(n18921) );
  INV_X1 U21156 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n18915) );
  INV_X1 U21157 ( .A(n18912), .ZN(n18913) );
  AOI22_X1 U21158 ( .A1(n18913), .A2(n19136), .B1(n19134), .B2(
        P2_REIP_REG_6__SCAN_IN), .ZN(n18914) );
  OAI211_X1 U21159 ( .C1(n18915), .C2(n19153), .A(n18914), .B(n18976), .ZN(
        n18919) );
  OAI22_X1 U21160 ( .A1(n19133), .A2(n18917), .B1(n19098), .B2(n18916), .ZN(
        n18918) );
  AOI211_X1 U21161 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n19157), .A(
        n18919), .B(n18918), .ZN(n18920) );
  OAI21_X1 U21162 ( .B1(n19267), .B2(n18921), .A(n18920), .ZN(P2_U2849) );
  NAND2_X1 U21163 ( .A1(n19029), .A2(n18922), .ZN(n18924) );
  XOR2_X1 U21164 ( .A(n18924), .B(n18923), .Z(n18932) );
  AOI22_X1 U21165 ( .A1(n18925), .A2(n19136), .B1(n19134), .B2(
        P2_REIP_REG_7__SCAN_IN), .ZN(n18926) );
  OAI211_X1 U21166 ( .C1(n12285), .C2(n19153), .A(n18926), .B(n18976), .ZN(
        n18930) );
  OAI22_X1 U21167 ( .A1(n19133), .A2(n18928), .B1(n19098), .B2(n18927), .ZN(
        n18929) );
  AOI211_X1 U21168 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19157), .A(
        n18930), .B(n18929), .ZN(n18931) );
  OAI21_X1 U21169 ( .B1(n18932), .B2(n19267), .A(n18931), .ZN(P2_U2848) );
  OAI21_X1 U21170 ( .B1(n12132), .B2(n19153), .A(n18976), .ZN(n18936) );
  OAI22_X1 U21171 ( .A1(n18934), .A2(n19149), .B1(n18933), .B2(n19121), .ZN(
        n18935) );
  AOI211_X1 U21172 ( .C1(P2_REIP_REG_9__SCAN_IN), .C2(n19134), .A(n18936), .B(
        n18935), .ZN(n18945) );
  INV_X1 U21173 ( .A(n18937), .ZN(n18940) );
  NAND2_X1 U21174 ( .A1(n19029), .A2(n18938), .ZN(n18939) );
  XOR2_X1 U21175 ( .A(n18940), .B(n18939), .Z(n18943) );
  INV_X1 U21176 ( .A(n18941), .ZN(n18942) );
  AOI22_X1 U21177 ( .A1(n18943), .A2(n19127), .B1(n18942), .B2(n19160), .ZN(
        n18944) );
  OAI211_X1 U21178 ( .C1(n18946), .C2(n19133), .A(n18945), .B(n18944), .ZN(
        P2_U2846) );
  INV_X1 U21179 ( .A(n18947), .ZN(n18951) );
  INV_X1 U21180 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n18949) );
  AOI22_X1 U21181 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n19135), .B1(
        P2_REIP_REG_11__SCAN_IN), .B2(n19134), .ZN(n18948) );
  OAI211_X1 U21182 ( .C1(n19121), .C2(n18949), .A(n18948), .B(n18976), .ZN(
        n18950) );
  AOI21_X1 U21183 ( .B1(n18951), .B2(n19160), .A(n18950), .ZN(n18952) );
  OAI21_X1 U21184 ( .B1(n18953), .B2(n19149), .A(n18952), .ZN(n18954) );
  AOI21_X1 U21185 ( .B1(n18955), .B2(n19159), .A(n18954), .ZN(n18960) );
  INV_X1 U21186 ( .A(n18956), .ZN(n18958) );
  OAI211_X1 U21187 ( .C1(n18958), .C2(n18961), .A(n19127), .B(n18957), .ZN(
        n18959) );
  OAI211_X1 U21188 ( .C1(n19050), .C2(n18961), .A(n18960), .B(n18959), .ZN(
        P2_U2844) );
  NAND2_X1 U21189 ( .A1(n19029), .A2(n18962), .ZN(n18964) );
  XOR2_X1 U21190 ( .A(n18964), .B(n18963), .Z(n18974) );
  AOI22_X1 U21191 ( .A1(n18965), .A2(n19136), .B1(n19134), .B2(
        P2_REIP_REG_13__SCAN_IN), .ZN(n18966) );
  OAI211_X1 U21192 ( .C1(n18967), .C2(n19153), .A(n18966), .B(n18976), .ZN(
        n18972) );
  INV_X1 U21193 ( .A(n18968), .ZN(n18969) );
  OAI22_X1 U21194 ( .A1(n18970), .A2(n19133), .B1(n18969), .B2(n19098), .ZN(
        n18971) );
  AOI211_X1 U21195 ( .C1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n19157), .A(
        n18972), .B(n18971), .ZN(n18973) );
  OAI21_X1 U21196 ( .B1(n18974), .B2(n19267), .A(n18973), .ZN(P2_U2842) );
  AOI22_X1 U21197 ( .A1(n18975), .A2(n19136), .B1(n19157), .B2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18977) );
  OAI211_X1 U21198 ( .C1(n12144), .C2(n19153), .A(n18977), .B(n18976), .ZN(
        n18978) );
  AOI21_X1 U21199 ( .B1(P2_REIP_REG_15__SCAN_IN), .B2(n19134), .A(n18978), 
        .ZN(n18985) );
  NAND2_X1 U21200 ( .A1(n19029), .A2(n18979), .ZN(n18981) );
  XNOR2_X1 U21201 ( .A(n18981), .B(n18980), .ZN(n18983) );
  AOI22_X1 U21202 ( .A1(n18983), .A2(n19127), .B1(n18982), .B2(n19160), .ZN(
        n18984) );
  OAI211_X1 U21203 ( .C1(n18986), .C2(n19133), .A(n18985), .B(n18984), .ZN(
        P2_U2840) );
  AOI22_X1 U21204 ( .A1(n18987), .A2(n19136), .B1(n19157), .B2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18988) );
  OAI21_X1 U21205 ( .B1(n18989), .B2(n19151), .A(n18988), .ZN(n18990) );
  AOI211_X1 U21206 ( .C1(P2_EBX_REG_16__SCAN_IN), .C2(n19135), .A(n19213), .B(
        n18990), .ZN(n18997) );
  NOR2_X1 U21207 ( .A1(n19015), .A2(n18991), .ZN(n18993) );
  XNOR2_X1 U21208 ( .A(n18993), .B(n18992), .ZN(n18995) );
  AOI22_X1 U21209 ( .A1(n18995), .A2(n19127), .B1(n18994), .B2(n19160), .ZN(
        n18996) );
  OAI211_X1 U21210 ( .C1(n18998), .C2(n19133), .A(n18997), .B(n18996), .ZN(
        P2_U2839) );
  INV_X1 U21211 ( .A(n19001), .ZN(n19010) );
  AOI22_X1 U21212 ( .A1(P2_EBX_REG_17__SCAN_IN), .A2(n19135), .B1(
        P2_REIP_REG_17__SCAN_IN), .B2(n19134), .ZN(n18999) );
  OAI211_X1 U21213 ( .C1(n19121), .C2(n12358), .A(n18999), .B(n18976), .ZN(
        n19003) );
  NOR2_X1 U21214 ( .A1(n19267), .A2(n19015), .ZN(n19046) );
  INV_X1 U21215 ( .A(n19046), .ZN(n19165) );
  AOI211_X1 U21216 ( .C1(n19001), .C2(n19000), .A(n19014), .B(n19165), .ZN(
        n19002) );
  AOI211_X1 U21217 ( .C1(n19136), .C2(n19004), .A(n19003), .B(n19002), .ZN(
        n19009) );
  INV_X1 U21218 ( .A(n19005), .ZN(n19007) );
  AOI22_X1 U21219 ( .A1(n19007), .A2(n19160), .B1(n19159), .B2(n19006), .ZN(
        n19008) );
  OAI211_X1 U21220 ( .C1(n19010), .C2(n19050), .A(n19009), .B(n19008), .ZN(
        P2_U2838) );
  OAI22_X1 U21221 ( .A1(n19012), .A2(n19149), .B1(n19011), .B2(n19151), .ZN(
        n19013) );
  AOI211_X1 U21222 ( .C1(P2_EBX_REG_18__SCAN_IN), .C2(n19135), .A(n19213), .B(
        n19013), .ZN(n19023) );
  NOR2_X1 U21223 ( .A1(n19015), .A2(n19014), .ZN(n19016) );
  XNOR2_X1 U21224 ( .A(n19017), .B(n19016), .ZN(n19021) );
  OAI22_X1 U21225 ( .A1(n19019), .A2(n19098), .B1(n19018), .B2(n19133), .ZN(
        n19020) );
  AOI21_X1 U21226 ( .B1(n19021), .B2(n19127), .A(n19020), .ZN(n19022) );
  OAI211_X1 U21227 ( .C1(n11539), .C2(n19121), .A(n19023), .B(n19022), .ZN(
        P2_U2837) );
  AOI22_X1 U21228 ( .A1(n19024), .A2(n19136), .B1(n19157), .B2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n19025) );
  OAI21_X1 U21229 ( .B1(n19026), .B2(n19151), .A(n19025), .ZN(n19027) );
  AOI211_X1 U21230 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n19135), .A(n19213), .B(
        n19027), .ZN(n19035) );
  NAND2_X1 U21231 ( .A1(n19029), .A2(n19028), .ZN(n19031) );
  XNOR2_X1 U21232 ( .A(n19031), .B(n19030), .ZN(n19033) );
  AOI22_X1 U21233 ( .A1(n19033), .A2(n19127), .B1(n19032), .B2(n19160), .ZN(
        n19034) );
  OAI211_X1 U21234 ( .C1(n19036), .C2(n19133), .A(n19035), .B(n19034), .ZN(
        P2_U2836) );
  INV_X1 U21235 ( .A(n19037), .ZN(n19038) );
  OAI222_X1 U21236 ( .A1(n19151), .A2(n19040), .B1(n19153), .B2(n19039), .C1(
        n19149), .C2(n19038), .ZN(n19044) );
  INV_X1 U21237 ( .A(n20066), .ZN(n19041) );
  OAI22_X1 U21238 ( .A1(n19042), .A2(n19098), .B1(n19041), .B2(n19133), .ZN(
        n19043) );
  AOI211_X1 U21239 ( .C1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n19157), .A(
        n19044), .B(n19043), .ZN(n19049) );
  OAI211_X1 U21240 ( .C1(n19047), .C2(n19051), .A(n19046), .B(n19045), .ZN(
        n19048) );
  OAI211_X1 U21241 ( .C1(n19051), .C2(n19050), .A(n19049), .B(n19048), .ZN(
        P2_U2835) );
  AOI22_X1 U21242 ( .A1(P2_EBX_REG_21__SCAN_IN), .A2(n19135), .B1(
        P2_REIP_REG_21__SCAN_IN), .B2(n19134), .ZN(n19062) );
  AOI22_X1 U21243 ( .A1(n19052), .A2(n19136), .B1(n19157), .B2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n19061) );
  OAI22_X1 U21244 ( .A1(n19054), .A2(n19098), .B1(n19053), .B2(n19133), .ZN(
        n19055) );
  INV_X1 U21245 ( .A(n19055), .ZN(n19060) );
  OAI211_X1 U21246 ( .C1(n19058), .C2(n19057), .A(n19127), .B(n19056), .ZN(
        n19059) );
  NAND4_X1 U21247 ( .A1(n19062), .A2(n19061), .A3(n19060), .A4(n19059), .ZN(
        P2_U2834) );
  AOI22_X1 U21248 ( .A1(P2_EBX_REG_22__SCAN_IN), .A2(n19135), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19134), .ZN(n19072) );
  AOI22_X1 U21249 ( .A1(n19063), .A2(n19136), .B1(n19157), .B2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n19071) );
  NOR2_X1 U21250 ( .A1(n19963), .A2(n19133), .ZN(n19064) );
  AOI21_X1 U21251 ( .B1(n19065), .B2(n19160), .A(n19064), .ZN(n19070) );
  OAI211_X1 U21252 ( .C1(n19068), .C2(n19067), .A(n19127), .B(n19066), .ZN(
        n19069) );
  NAND4_X1 U21253 ( .A1(n19072), .A2(n19071), .A3(n19070), .A4(n19069), .ZN(
        P2_U2833) );
  NAND2_X1 U21254 ( .A1(n19073), .A2(n19160), .ZN(n19075) );
  AOI22_X1 U21255 ( .A1(n19134), .A2(P2_REIP_REG_23__SCAN_IN), .B1(n19135), 
        .B2(P2_EBX_REG_23__SCAN_IN), .ZN(n19074) );
  OAI211_X1 U21256 ( .C1(n19121), .C2(n19076), .A(n19075), .B(n19074), .ZN(
        n19077) );
  AOI21_X1 U21257 ( .B1(n19078), .B2(n19136), .A(n19077), .ZN(n19083) );
  OAI211_X1 U21258 ( .C1(n19081), .C2(n19080), .A(n19127), .B(n19079), .ZN(
        n19082) );
  OAI211_X1 U21259 ( .C1(n19133), .C2(n19084), .A(n19083), .B(n19082), .ZN(
        P2_U2832) );
  AOI22_X1 U21260 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(n19135), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19134), .ZN(n19095) );
  AOI22_X1 U21261 ( .A1(n19085), .A2(n19136), .B1(n19157), .B2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n19094) );
  OAI22_X1 U21262 ( .A1(n19087), .A2(n19098), .B1(n19086), .B2(n19133), .ZN(
        n19088) );
  INV_X1 U21263 ( .A(n19088), .ZN(n19093) );
  OAI211_X1 U21264 ( .C1(n19091), .C2(n19090), .A(n19127), .B(n19089), .ZN(
        n19092) );
  NAND4_X1 U21265 ( .A1(n19095), .A2(n19094), .A3(n19093), .A4(n19092), .ZN(
        P2_U2831) );
  AOI22_X1 U21266 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(n19135), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n19134), .ZN(n19107) );
  AOI22_X1 U21267 ( .A1(n19096), .A2(n19136), .B1(n19157), .B2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n19106) );
  OAI22_X1 U21268 ( .A1(n19099), .A2(n19098), .B1(n19097), .B2(n19133), .ZN(
        n19100) );
  INV_X1 U21269 ( .A(n19100), .ZN(n19105) );
  OAI211_X1 U21270 ( .C1(n19103), .C2(n19102), .A(n19127), .B(n19101), .ZN(
        n19104) );
  NAND4_X1 U21271 ( .A1(n19107), .A2(n19106), .A3(n19105), .A4(n19104), .ZN(
        P2_U2830) );
  AOI22_X1 U21272 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n19135), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n19134), .ZN(n19117) );
  AOI22_X1 U21273 ( .A1(n19108), .A2(n19136), .B1(n19157), .B2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n19116) );
  AOI22_X1 U21274 ( .A1(n19110), .A2(n19160), .B1(n19109), .B2(n19159), .ZN(
        n19115) );
  OAI211_X1 U21275 ( .C1(n19113), .C2(n19112), .A(n19127), .B(n19111), .ZN(
        n19114) );
  NAND4_X1 U21276 ( .A1(n19117), .A2(n19116), .A3(n19115), .A4(n19114), .ZN(
        P2_U2829) );
  INV_X1 U21277 ( .A(n19118), .ZN(n19125) );
  AOI22_X1 U21278 ( .A1(n19134), .A2(P2_REIP_REG_27__SCAN_IN), .B1(n19135), 
        .B2(P2_EBX_REG_27__SCAN_IN), .ZN(n19119) );
  OAI21_X1 U21279 ( .B1(n19121), .B2(n19120), .A(n19119), .ZN(n19124) );
  NOR2_X1 U21280 ( .A1(n19122), .A2(n19149), .ZN(n19123) );
  AOI211_X1 U21281 ( .C1(n19160), .C2(n19125), .A(n19124), .B(n19123), .ZN(
        n19131) );
  OAI211_X1 U21282 ( .C1(n19129), .C2(n19128), .A(n19127), .B(n19126), .ZN(
        n19130) );
  OAI211_X1 U21283 ( .C1(n19133), .C2(n19132), .A(n19131), .B(n19130), .ZN(
        P2_U2828) );
  AOI22_X1 U21284 ( .A1(P2_EBX_REG_29__SCAN_IN), .A2(n19135), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n19134), .ZN(n19147) );
  AOI22_X1 U21285 ( .A1(n19137), .A2(n19136), .B1(n19157), .B2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n19146) );
  INV_X1 U21286 ( .A(n19138), .ZN(n19139) );
  AOI22_X1 U21287 ( .A1(n19140), .A2(n19160), .B1(n19139), .B2(n19159), .ZN(
        n19145) );
  OAI211_X1 U21288 ( .C1(n19143), .C2(n19142), .A(n19127), .B(n19141), .ZN(
        n19144) );
  NAND4_X1 U21289 ( .A1(n19147), .A2(n19146), .A3(n19145), .A4(n19144), .ZN(
        P2_U2826) );
  INV_X1 U21290 ( .A(n19148), .ZN(n19150) );
  NOR2_X1 U21291 ( .A1(n19150), .A2(n19149), .ZN(n19156) );
  OAI22_X1 U21292 ( .A1(n19154), .A2(n19153), .B1(n19152), .B2(n19151), .ZN(
        n19155) );
  AOI211_X1 U21293 ( .C1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n19157), .A(
        n19156), .B(n19155), .ZN(n19163) );
  AOI22_X1 U21294 ( .A1(n19161), .A2(n19160), .B1(n19159), .B2(n19158), .ZN(
        n19162) );
  OAI211_X1 U21295 ( .C1(n19165), .C2(n19164), .A(n19163), .B(n19162), .ZN(
        P2_U2824) );
  INV_X1 U21296 ( .A(n19166), .ZN(n19173) );
  AND3_X1 U21297 ( .A1(n19169), .A2(n19168), .A3(n19167), .ZN(n19244) );
  NAND3_X1 U21298 ( .A1(n19173), .A2(n19170), .A3(n19244), .ZN(n19171) );
  OAI21_X1 U21299 ( .B1(n19173), .B2(n19172), .A(n19171), .ZN(P2_U3595) );
  NAND2_X1 U21300 ( .A1(n19202), .A2(n19174), .ZN(n19175) );
  OAI21_X1 U21301 ( .B1(n19184), .B2(n19176), .A(n19175), .ZN(n19182) );
  OAI22_X1 U21302 ( .A1(n19180), .A2(n19179), .B1(n19178), .B2(n19177), .ZN(
        n19181) );
  AOI211_X1 U21303 ( .C1(n19184), .C2(n19183), .A(n19182), .B(n19181), .ZN(
        n19186) );
  OAI211_X1 U21304 ( .C1(n19188), .C2(n19187), .A(n19186), .B(n19185), .ZN(
        P2_U3046) );
  INV_X1 U21305 ( .A(n19189), .ZN(n19191) );
  AOI22_X1 U21306 ( .A1(n19191), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n19208), .B2(n19190), .ZN(n19200) );
  AOI222_X1 U21307 ( .A1(n19194), .A2(n12758), .B1(n19211), .B2(n19193), .C1(
        n19202), .C2(n19192), .ZN(n19199) );
  NAND2_X1 U21308 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19213), .ZN(n19198) );
  OAI221_X1 U21309 ( .B1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n12125), .C2(n19196), .A(
        n19195), .ZN(n19197) );
  NAND4_X1 U21310 ( .A1(n19200), .A2(n19199), .A3(n19198), .A4(n19197), .ZN(
        P2_U3038) );
  INV_X1 U21311 ( .A(n19201), .ZN(n19203) );
  AOI22_X1 U21312 ( .A1(n19205), .A2(n19204), .B1(n19203), .B2(n19202), .ZN(
        n19217) );
  INV_X1 U21313 ( .A(n19206), .ZN(n19209) );
  AOI22_X1 U21314 ( .A1(n19209), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n19208), .B2(n19207), .ZN(n19216) );
  AOI22_X1 U21315 ( .A1(n19212), .A2(n19211), .B1(n12758), .B2(n19210), .ZN(
        n19215) );
  NAND2_X1 U21316 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19213), .ZN(n19214) );
  NAND4_X1 U21317 ( .A1(n19217), .A2(n19216), .A3(n19215), .A4(n19214), .ZN(
        P2_U3042) );
  INV_X1 U21318 ( .A(n19218), .ZN(n19223) );
  NOR2_X1 U21319 ( .A1(n19219), .A2(n19927), .ZN(n19220) );
  OR2_X1 U21320 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19220), .ZN(
        n19222) );
  AND2_X1 U21321 ( .A1(n19220), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19221) );
  AOI211_X1 U21322 ( .C1(n19223), .C2(n19222), .A(n19255), .B(n19221), .ZN(
        n19227) );
  INV_X1 U21323 ( .A(n19255), .ZN(n19230) );
  MUX2_X1 U21324 ( .A(n19225), .B(n19224), .S(n19230), .Z(n19252) );
  INV_X1 U21325 ( .A(n19252), .ZN(n19226) );
  AOI222_X1 U21326 ( .A1(n19227), .A2(n19832), .B1(n19227), .B2(n19226), .C1(
        n19832), .C2(n19226), .ZN(n19231) );
  NAND2_X1 U21327 ( .A1(n19228), .A2(n19230), .ZN(n19229) );
  OAI21_X1 U21328 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19230), .A(
        n19229), .ZN(n19251) );
  OR2_X1 U21329 ( .A1(n19231), .A2(n19251), .ZN(n19232) );
  AOI221_X1 U21330 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n19232), 
        .C1(n19231), .C2(n19251), .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n19254) );
  INV_X1 U21331 ( .A(n19233), .ZN(n19237) );
  AOI22_X1 U21332 ( .A1(n19235), .A2(n19234), .B1(n19248), .B2(n19245), .ZN(
        n19236) );
  OAI21_X1 U21333 ( .B1(n19272), .B2(n19237), .A(n19236), .ZN(n19238) );
  AOI21_X1 U21334 ( .B1(n19239), .B2(n19242), .A(n19238), .ZN(n19240) );
  OAI21_X1 U21335 ( .B1(n19242), .B2(n19241), .A(n19240), .ZN(n19289) );
  NOR3_X1 U21336 ( .A1(n19289), .A2(n19244), .A3(n19243), .ZN(n19250) );
  NOR4_X1 U21337 ( .A1(n19248), .A2(n11157), .A3(n19247), .A4(n19246), .ZN(
        n19288) );
  OAI21_X1 U21338 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n19288), .ZN(n19249) );
  OAI211_X1 U21339 ( .C1(n19252), .C2(n19251), .A(n19250), .B(n19249), .ZN(
        n19253) );
  AOI211_X1 U21340 ( .C1(n19255), .C2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n19254), .B(n19253), .ZN(n19286) );
  NAND3_X1 U21341 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19286), .A3(n19256), 
        .ZN(n19260) );
  INV_X1 U21342 ( .A(n19257), .ZN(n19258) );
  AOI21_X1 U21343 ( .B1(n19260), .B2(n19259), .A(n19258), .ZN(n19278) );
  NAND2_X1 U21344 ( .A1(n19278), .A2(n19261), .ZN(n19280) );
  OAI21_X1 U21345 ( .B1(n19263), .B2(n19262), .A(n19287), .ZN(n19266) );
  NAND2_X1 U21346 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n22321), .ZN(n19264) );
  AOI21_X1 U21347 ( .B1(n19273), .B2(n19280), .A(n19264), .ZN(n19265) );
  AOI21_X1 U21348 ( .B1(n19280), .B2(n19266), .A(n19265), .ZN(n19268) );
  NAND2_X1 U21349 ( .A1(n19268), .A2(n19267), .ZN(P2_U3177) );
  AOI221_X1 U21350 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19270), .C1(
        P2_STATE2_REG_3__SCAN_IN), .C2(n19278), .A(n19269), .ZN(n19271) );
  INV_X1 U21351 ( .A(n19271), .ZN(P2_U3593) );
  INV_X1 U21352 ( .A(n19272), .ZN(n19275) );
  OAI22_X1 U21353 ( .A1(n19275), .A2(n19274), .B1(n19273), .B2(n19281), .ZN(
        n19276) );
  AOI211_X1 U21354 ( .C1(P2_STATE2_REG_0__SCAN_IN), .C2(n19278), .A(n19277), 
        .B(n19276), .ZN(n19285) );
  NOR2_X1 U21355 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19279), .ZN(n19283) );
  OAI22_X1 U21356 ( .A1(n19283), .A2(n19282), .B1(n19281), .B2(n19280), .ZN(
        n19284) );
  OAI211_X1 U21357 ( .C1(n19286), .C2(n19287), .A(n19285), .B(n19284), .ZN(
        P2_U3176) );
  NOR2_X1 U21358 ( .A1(n19288), .A2(n19287), .ZN(n19291) );
  MUX2_X1 U21359 ( .A(P2_MORE_REG_SCAN_IN), .B(n19289), .S(n19291), .Z(
        P2_U3609) );
  OAI21_X1 U21360 ( .B1(n19291), .B2(n12257), .A(n19290), .ZN(P2_U2819) );
  INV_X1 U21361 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n20666) );
  INV_X1 U21362 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19753) );
  AOI22_X1 U21363 ( .A1(n19593), .A2(n20666), .B1(n19753), .B2(U215), .ZN(U282) );
  OAI22_X1 U21364 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19593), .ZN(n19292) );
  INV_X1 U21365 ( .A(n19292), .ZN(U281) );
  OAI22_X1 U21366 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19593), .ZN(n19293) );
  INV_X1 U21367 ( .A(n19293), .ZN(U280) );
  OAI22_X1 U21368 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19593), .ZN(n19294) );
  INV_X1 U21369 ( .A(n19294), .ZN(U279) );
  OAI22_X1 U21370 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19593), .ZN(n19295) );
  INV_X1 U21371 ( .A(n19295), .ZN(U278) );
  OAI22_X1 U21372 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19593), .ZN(n19296) );
  INV_X1 U21373 ( .A(n19296), .ZN(U277) );
  OAI22_X1 U21374 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19593), .ZN(n19297) );
  INV_X1 U21375 ( .A(n19297), .ZN(U276) );
  OAI22_X1 U21376 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19593), .ZN(n19298) );
  INV_X1 U21377 ( .A(n19298), .ZN(U275) );
  OAI22_X1 U21378 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19593), .ZN(n19299) );
  INV_X1 U21379 ( .A(n19299), .ZN(U274) );
  OAI22_X1 U21380 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19593), .ZN(n19300) );
  INV_X1 U21381 ( .A(n19300), .ZN(U273) );
  OAI22_X1 U21382 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19636), .ZN(n19301) );
  INV_X1 U21383 ( .A(n19301), .ZN(U272) );
  OAI22_X1 U21384 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19636), .ZN(n19302) );
  INV_X1 U21385 ( .A(n19302), .ZN(U271) );
  OAI22_X1 U21386 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19593), .ZN(n19303) );
  INV_X1 U21387 ( .A(n19303), .ZN(U270) );
  OAI22_X1 U21388 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19636), .ZN(n19304) );
  INV_X1 U21389 ( .A(n19304), .ZN(U269) );
  OAI22_X1 U21390 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19593), .ZN(n19305) );
  INV_X1 U21391 ( .A(n19305), .ZN(U268) );
  OAI22_X1 U21392 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19593), .ZN(n19306) );
  INV_X1 U21393 ( .A(n19306), .ZN(U267) );
  OAI22_X1 U21394 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19636), .ZN(n19307) );
  INV_X1 U21395 ( .A(n19307), .ZN(U266) );
  OAI22_X1 U21396 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n19636), .ZN(n19308) );
  INV_X1 U21397 ( .A(n19308), .ZN(U265) );
  OAI22_X1 U21398 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n19636), .ZN(n19309) );
  INV_X1 U21399 ( .A(n19309), .ZN(U264) );
  OAI22_X1 U21400 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n19636), .ZN(n19310) );
  INV_X1 U21401 ( .A(n19310), .ZN(U263) );
  OAI22_X1 U21402 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n19636), .ZN(n19311) );
  INV_X1 U21403 ( .A(n19311), .ZN(U262) );
  INV_X1 U21404 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n19313) );
  INV_X1 U21405 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n19312) );
  AOI22_X1 U21406 ( .A1(n19593), .A2(n19313), .B1(n19312), .B2(U215), .ZN(U261) );
  OAI22_X1 U21407 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n19636), .ZN(n19314) );
  INV_X1 U21408 ( .A(n19314), .ZN(U260) );
  OAI22_X1 U21409 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n19593), .ZN(n19315) );
  INV_X1 U21410 ( .A(n19315), .ZN(U259) );
  OAI22_X1 U21411 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n19593), .ZN(n19316) );
  INV_X1 U21412 ( .A(n19316), .ZN(U258) );
  NOR2_X1 U21413 ( .A1(n21837), .A2(n19337), .ZN(n19378) );
  NAND2_X1 U21414 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19378), .ZN(
        n19721) );
  NOR2_X1 U21415 ( .A1(n19317), .A2(n21852), .ZN(n19429) );
  NAND2_X1 U21416 ( .A1(n19429), .A2(n21267), .ZN(n19389) );
  NAND2_X1 U21417 ( .A1(n21827), .A2(n21825), .ZN(n21830) );
  NOR2_X1 U21418 ( .A1(n21834), .A2(n21837), .ZN(n19327) );
  INV_X1 U21419 ( .A(n19327), .ZN(n19325) );
  NOR2_X2 U21420 ( .A1(n21830), .A2(n19325), .ZN(n19658) );
  NOR2_X2 U21421 ( .A1(n19551), .A2(n19753), .ZN(n19386) );
  NOR2_X1 U21422 ( .A1(n21855), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n21848) );
  INV_X1 U21423 ( .A(n21848), .ZN(n21856) );
  AND2_X1 U21424 ( .A1(n21856), .A2(n19378), .ZN(n19641) );
  INV_X1 U21425 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n21202) );
  NOR2_X2 U21426 ( .A1(n19552), .A2(n21202), .ZN(n19381) );
  AOI22_X1 U21427 ( .A1(n19658), .A2(n19386), .B1(n19641), .B2(n19381), .ZN(
        n19321) );
  NAND2_X1 U21428 ( .A1(n19640), .A2(n19318), .ZN(n19326) );
  OAI21_X1 U21429 ( .B1(n21827), .B2(n19326), .A(n19551), .ZN(n19368) );
  NAND2_X1 U21430 ( .A1(n19327), .A2(n19368), .ZN(n19643) );
  NOR2_X1 U21431 ( .A1(n21825), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19345) );
  NAND2_X1 U21432 ( .A1(n19345), .A2(n19327), .ZN(n19739) );
  INV_X1 U21433 ( .A(n19739), .ZN(n19652) );
  INV_X1 U21434 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n19319) );
  NOR2_X2 U21435 ( .A1(n19551), .A2(n19319), .ZN(n19382) );
  AOI22_X1 U21436 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19643), .B1(
        n19652), .B2(n19382), .ZN(n19320) );
  OAI211_X1 U21437 ( .C1(n19721), .C2(n19389), .A(n19321), .B(n19320), .ZN(
        P3_U2995) );
  NAND2_X1 U21438 ( .A1(n19378), .A2(n21825), .ZN(n19728) );
  NAND2_X1 U21439 ( .A1(n19739), .A2(n19728), .ZN(n19385) );
  AND2_X1 U21440 ( .A1(n21856), .A2(n19385), .ZN(n19646) );
  AOI22_X1 U21441 ( .A1(n19382), .A2(n19658), .B1(n19381), .B2(n19646), .ZN(
        n19324) );
  NAND2_X1 U21442 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19342), .ZN(
        n19334) );
  NOR2_X2 U21443 ( .A1(n21825), .A2(n19334), .ZN(n19663) );
  NAND2_X1 U21444 ( .A1(n19556), .A2(n19650), .ZN(n19331) );
  NOR2_X1 U21445 ( .A1(n19552), .A2(n19322), .ZN(n19384) );
  OAI221_X1 U21446 ( .B1(n19385), .B2(n19355), .C1(n19385), .C2(n19331), .A(
        n19384), .ZN(n19647) );
  AOI22_X1 U21447 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19647), .B1(
        n19386), .B2(n19663), .ZN(n19323) );
  OAI211_X1 U21448 ( .C1(n19389), .C2(n19728), .A(n19324), .B(n19323), .ZN(
        P3_U2987) );
  INV_X1 U21449 ( .A(n19334), .ZN(n19328) );
  NAND2_X1 U21450 ( .A1(n21825), .A2(n19328), .ZN(n19656) );
  NAND2_X1 U21451 ( .A1(n21827), .A2(n21856), .ZN(n19375) );
  NOR2_X1 U21452 ( .A1(n19325), .A2(n19375), .ZN(n19651) );
  AOI22_X1 U21453 ( .A1(n19386), .A2(n19669), .B1(n19381), .B2(n19651), .ZN(
        n19330) );
  NOR2_X1 U21454 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19326), .ZN(
        n19377) );
  AOI22_X1 U21455 ( .A1(n19639), .A2(n19328), .B1(n19327), .B2(n19377), .ZN(
        n19653) );
  AOI22_X1 U21456 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19653), .B1(
        n19382), .B2(n19663), .ZN(n19329) );
  OAI211_X1 U21457 ( .C1(n19739), .C2(n19389), .A(n19330), .B(n19329), .ZN(
        P3_U2979) );
  NAND2_X1 U21458 ( .A1(n19342), .A2(n19345), .ZN(n19667) );
  INV_X1 U21459 ( .A(n19667), .ZN(n19675) );
  AND2_X1 U21460 ( .A1(n21856), .A2(n19331), .ZN(n19657) );
  AOI22_X1 U21461 ( .A1(n19386), .A2(n19675), .B1(n19381), .B2(n19657), .ZN(
        n19333) );
  NAND2_X1 U21462 ( .A1(n19656), .A2(n19667), .ZN(n19338) );
  AOI22_X1 U21463 ( .A1(n19639), .A2(n19338), .B1(n19384), .B2(n19331), .ZN(
        n19659) );
  AOI22_X1 U21464 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19659), .B1(
        n19382), .B2(n19669), .ZN(n19332) );
  OAI211_X1 U21465 ( .C1(n19389), .C2(n19556), .A(n19333), .B(n19332), .ZN(
        P3_U2971) );
  NOR2_X1 U21466 ( .A1(n21848), .A2(n19334), .ZN(n19662) );
  AOI22_X1 U21467 ( .A1(n19382), .A2(n19675), .B1(n19381), .B2(n19662), .ZN(
        n19336) );
  NAND2_X1 U21468 ( .A1(n19342), .A2(n19368), .ZN(n19664) );
  NOR2_X2 U21469 ( .A1(n21830), .A2(n19341), .ZN(n19681) );
  AOI22_X1 U21470 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19664), .B1(
        n19386), .B2(n19681), .ZN(n19335) );
  OAI211_X1 U21471 ( .C1(n19389), .C2(n19650), .A(n19336), .B(n19335), .ZN(
        P3_U2963) );
  NOR2_X1 U21472 ( .A1(n19337), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19349) );
  NAND2_X1 U21473 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19349), .ZN(
        n19609) );
  AND2_X1 U21474 ( .A1(n21856), .A2(n19338), .ZN(n19668) );
  AOI22_X1 U21475 ( .A1(n19386), .A2(n19686), .B1(n19381), .B2(n19668), .ZN(
        n19340) );
  NAND2_X1 U21476 ( .A1(n19673), .A2(n19609), .ZN(n19346) );
  OAI221_X1 U21477 ( .B1(n19338), .B2(n19355), .C1(n19338), .C2(n19346), .A(
        n19384), .ZN(n19670) );
  AOI22_X1 U21478 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19670), .B1(
        n19382), .B2(n19681), .ZN(n19339) );
  OAI211_X1 U21479 ( .C1(n19389), .C2(n19656), .A(n19340), .B(n19339), .ZN(
        P3_U2955) );
  NAND2_X1 U21480 ( .A1(n21825), .A2(n19349), .ZN(n19679) );
  NOR2_X1 U21481 ( .A1(n19341), .A2(n19375), .ZN(n19674) );
  AOI22_X1 U21482 ( .A1(n19386), .A2(n19692), .B1(n19381), .B2(n19674), .ZN(
        n19344) );
  AOI22_X1 U21483 ( .A1(n19639), .A2(n19349), .B1(n19342), .B2(n19377), .ZN(
        n19676) );
  AOI22_X1 U21484 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19676), .B1(
        n19382), .B2(n19686), .ZN(n19343) );
  OAI211_X1 U21485 ( .C1(n19389), .C2(n19667), .A(n19344), .B(n19343), .ZN(
        P3_U2947) );
  AND2_X1 U21486 ( .A1(n21856), .A2(n19346), .ZN(n19680) );
  AOI22_X1 U21487 ( .A1(n19382), .A2(n19692), .B1(n19381), .B2(n19680), .ZN(
        n19348) );
  INV_X1 U21488 ( .A(n19345), .ZN(n19363) );
  NOR2_X2 U21489 ( .A1(n19358), .A2(n19363), .ZN(n19698) );
  NAND2_X1 U21490 ( .A1(n19679), .A2(n19690), .ZN(n19354) );
  AOI22_X1 U21491 ( .A1(n19639), .A2(n19354), .B1(n19384), .B2(n19346), .ZN(
        n19682) );
  AOI22_X1 U21492 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19682), .B1(
        n19386), .B2(n19698), .ZN(n19347) );
  OAI211_X1 U21493 ( .C1(n19389), .C2(n19673), .A(n19348), .B(n19347), .ZN(
        P3_U2939) );
  INV_X1 U21494 ( .A(n19349), .ZN(n19350) );
  NOR2_X1 U21495 ( .A1(n21848), .A2(n19350), .ZN(n19685) );
  AOI22_X1 U21496 ( .A1(n19382), .A2(n19698), .B1(n19381), .B2(n19685), .ZN(
        n19352) );
  NAND2_X1 U21497 ( .A1(n19359), .A2(n19368), .ZN(n19687) );
  NOR2_X2 U21498 ( .A1(n21830), .A2(n19358), .ZN(n19704) );
  AOI22_X1 U21499 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19687), .B1(
        n19386), .B2(n19704), .ZN(n19351) );
  OAI211_X1 U21500 ( .C1(n19389), .C2(n19609), .A(n19352), .B(n19351), .ZN(
        P3_U2931) );
  AND2_X1 U21501 ( .A1(n21856), .A2(n19354), .ZN(n19691) );
  AOI22_X1 U21502 ( .A1(n19382), .A2(n19704), .B1(n19381), .B2(n19691), .ZN(
        n19357) );
  NOR2_X1 U21503 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19376) );
  NAND2_X1 U21504 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19376), .ZN(
        n19367) );
  NOR2_X2 U21505 ( .A1(n21825), .A2(n19367), .ZN(n19710) );
  INV_X1 U21506 ( .A(n19710), .ZN(n19702) );
  INV_X1 U21507 ( .A(n19384), .ZN(n19353) );
  AOI21_X1 U21508 ( .B1(n19696), .B2(n19702), .A(n19353), .ZN(n19364) );
  AOI22_X1 U21509 ( .A1(n19355), .A2(n19364), .B1(n19384), .B2(n19354), .ZN(
        n19693) );
  AOI22_X1 U21510 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19693), .B1(
        n19386), .B2(n19710), .ZN(n19356) );
  OAI211_X1 U21511 ( .C1(n19389), .C2(n19679), .A(n19357), .B(n19356), .ZN(
        P3_U2923) );
  INV_X1 U21512 ( .A(n19367), .ZN(n19360) );
  NAND2_X1 U21513 ( .A1(n21825), .A2(n19360), .ZN(n19620) );
  NOR2_X1 U21514 ( .A1(n19358), .A2(n19375), .ZN(n19697) );
  AOI22_X1 U21515 ( .A1(n19386), .A2(n19717), .B1(n19381), .B2(n19697), .ZN(
        n19362) );
  AOI22_X1 U21516 ( .A1(n19639), .A2(n19360), .B1(n19359), .B2(n19377), .ZN(
        n19699) );
  AOI22_X1 U21517 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19699), .B1(
        n19382), .B2(n19710), .ZN(n19361) );
  OAI211_X1 U21518 ( .C1(n19389), .C2(n19690), .A(n19362), .B(n19361), .ZN(
        P3_U2915) );
  AOI21_X1 U21519 ( .B1(n19696), .B2(n19702), .A(n21848), .ZN(n19703) );
  AOI22_X1 U21520 ( .A1(n19382), .A2(n19717), .B1(n19381), .B2(n19703), .ZN(
        n19366) );
  INV_X1 U21521 ( .A(n19376), .ZN(n19374) );
  NOR2_X2 U21522 ( .A1(n19363), .A2(n19374), .ZN(n19724) );
  NAND2_X1 U21523 ( .A1(n19620), .A2(n19715), .ZN(n19371) );
  AOI21_X1 U21524 ( .B1(n19639), .B2(n19371), .A(n19364), .ZN(n19705) );
  AOI22_X1 U21525 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19705), .B1(
        n19386), .B2(n19724), .ZN(n19365) );
  OAI211_X1 U21526 ( .C1(n19389), .C2(n19696), .A(n19366), .B(n19365), .ZN(
        P3_U2907) );
  NOR2_X1 U21527 ( .A1(n21848), .A2(n19367), .ZN(n19708) );
  AOI22_X1 U21528 ( .A1(n19382), .A2(n19724), .B1(n19381), .B2(n19708), .ZN(
        n19370) );
  NAND2_X1 U21529 ( .A1(n19376), .A2(n19368), .ZN(n19711) );
  NOR2_X2 U21530 ( .A1(n21830), .A2(n19374), .ZN(n19734) );
  AOI22_X1 U21531 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19711), .B1(
        n19386), .B2(n19734), .ZN(n19369) );
  OAI211_X1 U21532 ( .C1(n19389), .C2(n19702), .A(n19370), .B(n19369), .ZN(
        P3_U2899) );
  AND2_X1 U21533 ( .A1(n21856), .A2(n19371), .ZN(n19716) );
  AOI22_X1 U21534 ( .A1(n19382), .A2(n19734), .B1(n19381), .B2(n19716), .ZN(
        n19373) );
  INV_X1 U21535 ( .A(n19734), .ZN(n19627) );
  NAND2_X1 U21536 ( .A1(n19721), .A2(n19627), .ZN(n19383) );
  AOI22_X1 U21537 ( .A1(n19639), .A2(n19383), .B1(n19384), .B2(n19371), .ZN(
        n19718) );
  INV_X1 U21538 ( .A(n19721), .ZN(n19723) );
  AOI22_X1 U21539 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19718), .B1(
        n19723), .B2(n19386), .ZN(n19372) );
  OAI211_X1 U21540 ( .C1(n19389), .C2(n19620), .A(n19373), .B(n19372), .ZN(
        P3_U2891) );
  NOR2_X1 U21541 ( .A1(n19375), .A2(n19374), .ZN(n19722) );
  AOI22_X1 U21542 ( .A1(n19382), .A2(n19723), .B1(n19381), .B2(n19722), .ZN(
        n19380) );
  AOI22_X1 U21543 ( .A1(n19639), .A2(n19378), .B1(n19377), .B2(n19376), .ZN(
        n19725) );
  INV_X1 U21544 ( .A(n19728), .ZN(n19732) );
  AOI22_X1 U21545 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19725), .B1(
        n19386), .B2(n19732), .ZN(n19379) );
  OAI211_X1 U21546 ( .C1(n19389), .C2(n19715), .A(n19380), .B(n19379), .ZN(
        P3_U2883) );
  AND2_X1 U21547 ( .A1(n21856), .A2(n19383), .ZN(n19730) );
  AOI22_X1 U21548 ( .A1(n19382), .A2(n19732), .B1(n19381), .B2(n19730), .ZN(
        n19388) );
  AOI22_X1 U21549 ( .A1(n19639), .A2(n19385), .B1(n19384), .B2(n19383), .ZN(
        n19735) );
  AOI22_X1 U21550 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19735), .B1(
        n19652), .B2(n19386), .ZN(n19387) );
  OAI211_X1 U21551 ( .C1(n19389), .C2(n19627), .A(n19388), .B(n19387), .ZN(
        P3_U2875) );
  OAI22_X1 U21552 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n19593), .ZN(n19390) );
  INV_X1 U21553 ( .A(n19390), .ZN(U257) );
  NAND2_X1 U21554 ( .A1(n19429), .A2(n21232), .ZN(n19427) );
  AND2_X1 U21555 ( .A1(n19639), .A2(BUF2_REG_22__SCAN_IN), .ZN(n19424) );
  NOR2_X2 U21556 ( .A1(n19552), .A2(n21207), .ZN(n19422) );
  AOI22_X1 U21557 ( .A1(n19652), .A2(n19424), .B1(n19641), .B2(n19422), .ZN(
        n19393) );
  INV_X1 U21558 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n19391) );
  NOR2_X2 U21559 ( .A1(n19391), .A2(n19551), .ZN(n19423) );
  AOI22_X1 U21560 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19643), .B1(
        n19658), .B2(n19423), .ZN(n19392) );
  OAI211_X1 U21561 ( .C1(n19721), .C2(n19427), .A(n19393), .B(n19392), .ZN(
        P3_U2994) );
  AOI22_X1 U21562 ( .A1(n19658), .A2(n19424), .B1(n19646), .B2(n19422), .ZN(
        n19395) );
  AOI22_X1 U21563 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19647), .B1(
        n19663), .B2(n19423), .ZN(n19394) );
  OAI211_X1 U21564 ( .C1(n19728), .C2(n19427), .A(n19395), .B(n19394), .ZN(
        P3_U2986) );
  AOI22_X1 U21565 ( .A1(n19669), .A2(n19423), .B1(n19651), .B2(n19422), .ZN(
        n19397) );
  AOI22_X1 U21566 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19653), .B1(
        n19663), .B2(n19424), .ZN(n19396) );
  OAI211_X1 U21567 ( .C1(n19739), .C2(n19427), .A(n19397), .B(n19396), .ZN(
        P3_U2978) );
  AOI22_X1 U21568 ( .A1(n19669), .A2(n19424), .B1(n19657), .B2(n19422), .ZN(
        n19399) );
  AOI22_X1 U21569 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19659), .B1(
        n19675), .B2(n19423), .ZN(n19398) );
  OAI211_X1 U21570 ( .C1(n19556), .C2(n19427), .A(n19399), .B(n19398), .ZN(
        P3_U2970) );
  AOI22_X1 U21571 ( .A1(n19675), .A2(n19424), .B1(n19662), .B2(n19422), .ZN(
        n19401) );
  AOI22_X1 U21572 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19664), .B1(
        n19681), .B2(n19423), .ZN(n19400) );
  OAI211_X1 U21573 ( .C1(n19650), .C2(n19427), .A(n19401), .B(n19400), .ZN(
        P3_U2962) );
  AOI22_X1 U21574 ( .A1(n19686), .A2(n19423), .B1(n19668), .B2(n19422), .ZN(
        n19403) );
  AOI22_X1 U21575 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19670), .B1(
        n19681), .B2(n19424), .ZN(n19402) );
  OAI211_X1 U21576 ( .C1(n19656), .C2(n19427), .A(n19403), .B(n19402), .ZN(
        P3_U2954) );
  AOI22_X1 U21577 ( .A1(n19686), .A2(n19424), .B1(n19674), .B2(n19422), .ZN(
        n19405) );
  AOI22_X1 U21578 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19676), .B1(
        n19692), .B2(n19423), .ZN(n19404) );
  OAI211_X1 U21579 ( .C1(n19667), .C2(n19427), .A(n19405), .B(n19404), .ZN(
        P3_U2946) );
  AOI22_X1 U21580 ( .A1(n19692), .A2(n19424), .B1(n19680), .B2(n19422), .ZN(
        n19407) );
  AOI22_X1 U21581 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19682), .B1(
        n19698), .B2(n19423), .ZN(n19406) );
  OAI211_X1 U21582 ( .C1(n19673), .C2(n19427), .A(n19407), .B(n19406), .ZN(
        P3_U2938) );
  AOI22_X1 U21583 ( .A1(n19704), .A2(n19423), .B1(n19685), .B2(n19422), .ZN(
        n19409) );
  AOI22_X1 U21584 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19687), .B1(
        n19698), .B2(n19424), .ZN(n19408) );
  OAI211_X1 U21585 ( .C1(n19609), .C2(n19427), .A(n19409), .B(n19408), .ZN(
        P3_U2930) );
  AOI22_X1 U21586 ( .A1(n19704), .A2(n19424), .B1(n19691), .B2(n19422), .ZN(
        n19411) );
  AOI22_X1 U21587 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19693), .B1(
        n19710), .B2(n19423), .ZN(n19410) );
  OAI211_X1 U21588 ( .C1(n19679), .C2(n19427), .A(n19411), .B(n19410), .ZN(
        P3_U2922) );
  AOI22_X1 U21589 ( .A1(n19697), .A2(n19422), .B1(n19717), .B2(n19423), .ZN(
        n19413) );
  AOI22_X1 U21590 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19699), .B1(
        n19710), .B2(n19424), .ZN(n19412) );
  OAI211_X1 U21591 ( .C1(n19690), .C2(n19427), .A(n19413), .B(n19412), .ZN(
        P3_U2914) );
  AOI22_X1 U21592 ( .A1(n19724), .A2(n19423), .B1(n19703), .B2(n19422), .ZN(
        n19415) );
  AOI22_X1 U21593 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19705), .B1(
        n19717), .B2(n19424), .ZN(n19414) );
  OAI211_X1 U21594 ( .C1(n19696), .C2(n19427), .A(n19415), .B(n19414), .ZN(
        P3_U2906) );
  AOI22_X1 U21595 ( .A1(n19734), .A2(n19423), .B1(n19708), .B2(n19422), .ZN(
        n19417) );
  AOI22_X1 U21596 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19711), .B1(
        n19724), .B2(n19424), .ZN(n19416) );
  OAI211_X1 U21597 ( .C1(n19702), .C2(n19427), .A(n19417), .B(n19416), .ZN(
        P3_U2898) );
  AOI22_X1 U21598 ( .A1(n19723), .A2(n19423), .B1(n19716), .B2(n19422), .ZN(
        n19419) );
  AOI22_X1 U21599 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19718), .B1(
        n19734), .B2(n19424), .ZN(n19418) );
  OAI211_X1 U21600 ( .C1(n19620), .C2(n19427), .A(n19419), .B(n19418), .ZN(
        P3_U2890) );
  AOI22_X1 U21601 ( .A1(n19732), .A2(n19423), .B1(n19722), .B2(n19422), .ZN(
        n19421) );
  AOI22_X1 U21602 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19725), .B1(
        n19723), .B2(n19424), .ZN(n19420) );
  OAI211_X1 U21603 ( .C1(n19715), .C2(n19427), .A(n19421), .B(n19420), .ZN(
        P3_U2882) );
  AOI22_X1 U21604 ( .A1(n19652), .A2(n19423), .B1(n19730), .B2(n19422), .ZN(
        n19426) );
  AOI22_X1 U21605 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19735), .B1(
        n19732), .B2(n19424), .ZN(n19425) );
  OAI211_X1 U21606 ( .C1(n19627), .C2(n19427), .A(n19426), .B(n19425), .ZN(
        P3_U2874) );
  OAI22_X1 U21607 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n19593), .ZN(n19428) );
  INV_X1 U21608 ( .A(n19428), .ZN(U256) );
  NAND2_X1 U21609 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19639), .ZN(n19468) );
  NAND2_X1 U21610 ( .A1(n19639), .A2(BUF2_REG_21__SCAN_IN), .ZN(n19462) );
  INV_X1 U21611 ( .A(n19462), .ZN(n19464) );
  INV_X1 U21612 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n21211) );
  NOR2_X2 U21613 ( .A1(n19552), .A2(n21211), .ZN(n19463) );
  AOI22_X1 U21614 ( .A1(n19652), .A2(n19464), .B1(n19641), .B2(n19463), .ZN(
        n19432) );
  INV_X1 U21615 ( .A(n19429), .ZN(n19642) );
  NOR2_X2 U21616 ( .A1(n19430), .A2(n19642), .ZN(n19465) );
  AOI22_X1 U21617 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19643), .B1(
        n19723), .B2(n19465), .ZN(n19431) );
  OAI211_X1 U21618 ( .C1(n19556), .C2(n19468), .A(n19432), .B(n19431), .ZN(
        P3_U2993) );
  AOI22_X1 U21619 ( .A1(n19658), .A2(n19464), .B1(n19646), .B2(n19463), .ZN(
        n19434) );
  AOI22_X1 U21620 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19647), .B1(
        n19732), .B2(n19465), .ZN(n19433) );
  OAI211_X1 U21621 ( .C1(n19650), .C2(n19468), .A(n19434), .B(n19433), .ZN(
        P3_U2985) );
  AOI22_X1 U21622 ( .A1(n19663), .A2(n19464), .B1(n19651), .B2(n19463), .ZN(
        n19436) );
  AOI22_X1 U21623 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19653), .B1(
        n19652), .B2(n19465), .ZN(n19435) );
  OAI211_X1 U21624 ( .C1(n19656), .C2(n19468), .A(n19436), .B(n19435), .ZN(
        P3_U2977) );
  AOI22_X1 U21625 ( .A1(n19669), .A2(n19464), .B1(n19657), .B2(n19463), .ZN(
        n19438) );
  AOI22_X1 U21626 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19659), .B1(
        n19658), .B2(n19465), .ZN(n19437) );
  OAI211_X1 U21627 ( .C1(n19667), .C2(n19468), .A(n19438), .B(n19437), .ZN(
        P3_U2969) );
  INV_X1 U21628 ( .A(n19468), .ZN(n19459) );
  AOI22_X1 U21629 ( .A1(n19681), .A2(n19459), .B1(n19662), .B2(n19463), .ZN(
        n19440) );
  AOI22_X1 U21630 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19664), .B1(
        n19663), .B2(n19465), .ZN(n19439) );
  OAI211_X1 U21631 ( .C1(n19667), .C2(n19462), .A(n19440), .B(n19439), .ZN(
        P3_U2961) );
  AOI22_X1 U21632 ( .A1(n19681), .A2(n19464), .B1(n19668), .B2(n19463), .ZN(
        n19442) );
  AOI22_X1 U21633 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19670), .B1(
        n19669), .B2(n19465), .ZN(n19441) );
  OAI211_X1 U21634 ( .C1(n19609), .C2(n19468), .A(n19442), .B(n19441), .ZN(
        P3_U2953) );
  AOI22_X1 U21635 ( .A1(n19686), .A2(n19464), .B1(n19674), .B2(n19463), .ZN(
        n19444) );
  AOI22_X1 U21636 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19676), .B1(
        n19675), .B2(n19465), .ZN(n19443) );
  OAI211_X1 U21637 ( .C1(n19679), .C2(n19468), .A(n19444), .B(n19443), .ZN(
        P3_U2945) );
  AOI22_X1 U21638 ( .A1(n19698), .A2(n19459), .B1(n19680), .B2(n19463), .ZN(
        n19446) );
  AOI22_X1 U21639 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19682), .B1(
        n19681), .B2(n19465), .ZN(n19445) );
  OAI211_X1 U21640 ( .C1(n19679), .C2(n19462), .A(n19446), .B(n19445), .ZN(
        P3_U2937) );
  AOI22_X1 U21641 ( .A1(n19698), .A2(n19464), .B1(n19685), .B2(n19463), .ZN(
        n19448) );
  AOI22_X1 U21642 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19687), .B1(
        n19686), .B2(n19465), .ZN(n19447) );
  OAI211_X1 U21643 ( .C1(n19696), .C2(n19468), .A(n19448), .B(n19447), .ZN(
        P3_U2929) );
  AOI22_X1 U21644 ( .A1(n19710), .A2(n19459), .B1(n19691), .B2(n19463), .ZN(
        n19450) );
  AOI22_X1 U21645 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19693), .B1(
        n19692), .B2(n19465), .ZN(n19449) );
  OAI211_X1 U21646 ( .C1(n19696), .C2(n19462), .A(n19450), .B(n19449), .ZN(
        P3_U2921) );
  AOI22_X1 U21647 ( .A1(n19710), .A2(n19464), .B1(n19697), .B2(n19463), .ZN(
        n19452) );
  AOI22_X1 U21648 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19699), .B1(
        n19698), .B2(n19465), .ZN(n19451) );
  OAI211_X1 U21649 ( .C1(n19620), .C2(n19468), .A(n19452), .B(n19451), .ZN(
        P3_U2913) );
  AOI22_X1 U21650 ( .A1(n19724), .A2(n19459), .B1(n19703), .B2(n19463), .ZN(
        n19454) );
  AOI22_X1 U21651 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19705), .B1(
        n19704), .B2(n19465), .ZN(n19453) );
  OAI211_X1 U21652 ( .C1(n19620), .C2(n19462), .A(n19454), .B(n19453), .ZN(
        P3_U2905) );
  AOI22_X1 U21653 ( .A1(n19724), .A2(n19464), .B1(n19708), .B2(n19463), .ZN(
        n19456) );
  AOI22_X1 U21654 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19711), .B1(
        n19710), .B2(n19465), .ZN(n19455) );
  OAI211_X1 U21655 ( .C1(n19627), .C2(n19468), .A(n19456), .B(n19455), .ZN(
        P3_U2897) );
  AOI22_X1 U21656 ( .A1(n19734), .A2(n19464), .B1(n19716), .B2(n19463), .ZN(
        n19458) );
  AOI22_X1 U21657 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19718), .B1(
        n19717), .B2(n19465), .ZN(n19457) );
  OAI211_X1 U21658 ( .C1(n19721), .C2(n19468), .A(n19458), .B(n19457), .ZN(
        P3_U2889) );
  AOI22_X1 U21659 ( .A1(n19732), .A2(n19459), .B1(n19722), .B2(n19463), .ZN(
        n19461) );
  AOI22_X1 U21660 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19725), .B1(
        n19724), .B2(n19465), .ZN(n19460) );
  OAI211_X1 U21661 ( .C1(n19721), .C2(n19462), .A(n19461), .B(n19460), .ZN(
        P3_U2881) );
  AOI22_X1 U21662 ( .A1(n19732), .A2(n19464), .B1(n19730), .B2(n19463), .ZN(
        n19467) );
  AOI22_X1 U21663 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19735), .B1(
        n19734), .B2(n19465), .ZN(n19466) );
  OAI211_X1 U21664 ( .C1(n19739), .C2(n19468), .A(n19467), .B(n19466), .ZN(
        P3_U2873) );
  OAI22_X1 U21665 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n19593), .ZN(n19469) );
  INV_X1 U21666 ( .A(n19469), .ZN(U255) );
  INV_X1 U21667 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n21294) );
  NOR2_X1 U21668 ( .A1(n21294), .A2(n19551), .ZN(n19504) );
  INV_X1 U21669 ( .A(n19504), .ZN(n19500) );
  NAND2_X1 U21670 ( .A1(n19639), .A2(BUF2_REG_20__SCAN_IN), .ZN(n19508) );
  INV_X1 U21671 ( .A(n19508), .ZN(n19497) );
  NOR2_X2 U21672 ( .A1(n19552), .A2(n21216), .ZN(n19503) );
  AOI22_X1 U21673 ( .A1(n19652), .A2(n19497), .B1(n19641), .B2(n19503), .ZN(
        n19472) );
  NOR2_X2 U21674 ( .A1(n19470), .A2(n19642), .ZN(n19505) );
  AOI22_X1 U21675 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19643), .B1(
        n19723), .B2(n19505), .ZN(n19471) );
  OAI211_X1 U21676 ( .C1(n19556), .C2(n19500), .A(n19472), .B(n19471), .ZN(
        P3_U2992) );
  AOI22_X1 U21677 ( .A1(n19658), .A2(n19497), .B1(n19646), .B2(n19503), .ZN(
        n19474) );
  AOI22_X1 U21678 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19647), .B1(
        n19732), .B2(n19505), .ZN(n19473) );
  OAI211_X1 U21679 ( .C1(n19650), .C2(n19500), .A(n19474), .B(n19473), .ZN(
        P3_U2984) );
  AOI22_X1 U21680 ( .A1(n19663), .A2(n19497), .B1(n19651), .B2(n19503), .ZN(
        n19476) );
  AOI22_X1 U21681 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19653), .B1(
        n19652), .B2(n19505), .ZN(n19475) );
  OAI211_X1 U21682 ( .C1(n19656), .C2(n19500), .A(n19476), .B(n19475), .ZN(
        P3_U2976) );
  AOI22_X1 U21683 ( .A1(n19675), .A2(n19504), .B1(n19657), .B2(n19503), .ZN(
        n19478) );
  AOI22_X1 U21684 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19659), .B1(
        n19658), .B2(n19505), .ZN(n19477) );
  OAI211_X1 U21685 ( .C1(n19656), .C2(n19508), .A(n19478), .B(n19477), .ZN(
        P3_U2968) );
  AOI22_X1 U21686 ( .A1(n19681), .A2(n19504), .B1(n19662), .B2(n19503), .ZN(
        n19480) );
  AOI22_X1 U21687 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19664), .B1(
        n19663), .B2(n19505), .ZN(n19479) );
  OAI211_X1 U21688 ( .C1(n19667), .C2(n19508), .A(n19480), .B(n19479), .ZN(
        P3_U2960) );
  AOI22_X1 U21689 ( .A1(n19681), .A2(n19497), .B1(n19668), .B2(n19503), .ZN(
        n19482) );
  AOI22_X1 U21690 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19670), .B1(
        n19669), .B2(n19505), .ZN(n19481) );
  OAI211_X1 U21691 ( .C1(n19609), .C2(n19500), .A(n19482), .B(n19481), .ZN(
        P3_U2952) );
  AOI22_X1 U21692 ( .A1(n19692), .A2(n19504), .B1(n19674), .B2(n19503), .ZN(
        n19484) );
  AOI22_X1 U21693 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19676), .B1(
        n19675), .B2(n19505), .ZN(n19483) );
  OAI211_X1 U21694 ( .C1(n19609), .C2(n19508), .A(n19484), .B(n19483), .ZN(
        P3_U2944) );
  AOI22_X1 U21695 ( .A1(n19698), .A2(n19504), .B1(n19680), .B2(n19503), .ZN(
        n19486) );
  AOI22_X1 U21696 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19682), .B1(
        n19681), .B2(n19505), .ZN(n19485) );
  OAI211_X1 U21697 ( .C1(n19679), .C2(n19508), .A(n19486), .B(n19485), .ZN(
        P3_U2936) );
  AOI22_X1 U21698 ( .A1(n19698), .A2(n19497), .B1(n19685), .B2(n19503), .ZN(
        n19488) );
  AOI22_X1 U21699 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19687), .B1(
        n19686), .B2(n19505), .ZN(n19487) );
  OAI211_X1 U21700 ( .C1(n19696), .C2(n19500), .A(n19488), .B(n19487), .ZN(
        P3_U2928) );
  AOI22_X1 U21701 ( .A1(n19704), .A2(n19497), .B1(n19691), .B2(n19503), .ZN(
        n19490) );
  AOI22_X1 U21702 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19693), .B1(
        n19692), .B2(n19505), .ZN(n19489) );
  OAI211_X1 U21703 ( .C1(n19702), .C2(n19500), .A(n19490), .B(n19489), .ZN(
        P3_U2920) );
  AOI22_X1 U21704 ( .A1(n19710), .A2(n19497), .B1(n19697), .B2(n19503), .ZN(
        n19492) );
  AOI22_X1 U21705 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19699), .B1(
        n19698), .B2(n19505), .ZN(n19491) );
  OAI211_X1 U21706 ( .C1(n19620), .C2(n19500), .A(n19492), .B(n19491), .ZN(
        P3_U2912) );
  AOI22_X1 U21707 ( .A1(n19717), .A2(n19497), .B1(n19703), .B2(n19503), .ZN(
        n19494) );
  AOI22_X1 U21708 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19705), .B1(
        n19704), .B2(n19505), .ZN(n19493) );
  OAI211_X1 U21709 ( .C1(n19715), .C2(n19500), .A(n19494), .B(n19493), .ZN(
        P3_U2904) );
  AOI22_X1 U21710 ( .A1(n19734), .A2(n19504), .B1(n19708), .B2(n19503), .ZN(
        n19496) );
  AOI22_X1 U21711 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19711), .B1(
        n19710), .B2(n19505), .ZN(n19495) );
  OAI211_X1 U21712 ( .C1(n19715), .C2(n19508), .A(n19496), .B(n19495), .ZN(
        P3_U2896) );
  AOI22_X1 U21713 ( .A1(n19734), .A2(n19497), .B1(n19716), .B2(n19503), .ZN(
        n19499) );
  AOI22_X1 U21714 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19718), .B1(
        n19717), .B2(n19505), .ZN(n19498) );
  OAI211_X1 U21715 ( .C1(n19721), .C2(n19500), .A(n19499), .B(n19498), .ZN(
        P3_U2888) );
  AOI22_X1 U21716 ( .A1(n19732), .A2(n19504), .B1(n19722), .B2(n19503), .ZN(
        n19502) );
  AOI22_X1 U21717 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19725), .B1(
        n19724), .B2(n19505), .ZN(n19501) );
  OAI211_X1 U21718 ( .C1(n19721), .C2(n19508), .A(n19502), .B(n19501), .ZN(
        P3_U2880) );
  AOI22_X1 U21719 ( .A1(n19652), .A2(n19504), .B1(n19730), .B2(n19503), .ZN(
        n19507) );
  AOI22_X1 U21720 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19735), .B1(
        n19734), .B2(n19505), .ZN(n19506) );
  OAI211_X1 U21721 ( .C1(n19728), .C2(n19508), .A(n19507), .B(n19506), .ZN(
        P3_U2872) );
  OAI22_X1 U21722 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n19593), .ZN(n19509) );
  INV_X1 U21723 ( .A(n19509), .ZN(U254) );
  INV_X1 U21724 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n19510) );
  NOR2_X1 U21725 ( .A1(n19551), .A2(n19510), .ZN(n19545) );
  INV_X1 U21726 ( .A(n19545), .ZN(n19543) );
  NAND2_X1 U21727 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19639), .ZN(n19549) );
  INV_X1 U21728 ( .A(n19549), .ZN(n19540) );
  INV_X1 U21729 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n21220) );
  NOR2_X2 U21730 ( .A1(n19552), .A2(n21220), .ZN(n19544) );
  AOI22_X1 U21731 ( .A1(n19658), .A2(n19540), .B1(n19641), .B2(n19544), .ZN(
        n19513) );
  NOR2_X2 U21732 ( .A1(n19511), .A2(n19642), .ZN(n19546) );
  AOI22_X1 U21733 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19643), .B1(
        n19723), .B2(n19546), .ZN(n19512) );
  OAI211_X1 U21734 ( .C1(n19739), .C2(n19543), .A(n19513), .B(n19512), .ZN(
        P3_U2991) );
  AOI22_X1 U21735 ( .A1(n19663), .A2(n19540), .B1(n19646), .B2(n19544), .ZN(
        n19515) );
  AOI22_X1 U21736 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19647), .B1(
        n19732), .B2(n19546), .ZN(n19514) );
  OAI211_X1 U21737 ( .C1(n19556), .C2(n19543), .A(n19515), .B(n19514), .ZN(
        P3_U2983) );
  AOI22_X1 U21738 ( .A1(n19663), .A2(n19545), .B1(n19651), .B2(n19544), .ZN(
        n19517) );
  AOI22_X1 U21739 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19653), .B1(
        n19652), .B2(n19546), .ZN(n19516) );
  OAI211_X1 U21740 ( .C1(n19656), .C2(n19549), .A(n19517), .B(n19516), .ZN(
        P3_U2975) );
  AOI22_X1 U21741 ( .A1(n19675), .A2(n19540), .B1(n19657), .B2(n19544), .ZN(
        n19519) );
  AOI22_X1 U21742 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19659), .B1(
        n19658), .B2(n19546), .ZN(n19518) );
  OAI211_X1 U21743 ( .C1(n19656), .C2(n19543), .A(n19519), .B(n19518), .ZN(
        P3_U2967) );
  AOI22_X1 U21744 ( .A1(n19681), .A2(n19540), .B1(n19662), .B2(n19544), .ZN(
        n19521) );
  AOI22_X1 U21745 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19664), .B1(
        n19663), .B2(n19546), .ZN(n19520) );
  OAI211_X1 U21746 ( .C1(n19667), .C2(n19543), .A(n19521), .B(n19520), .ZN(
        P3_U2959) );
  AOI22_X1 U21747 ( .A1(n19686), .A2(n19540), .B1(n19668), .B2(n19544), .ZN(
        n19523) );
  AOI22_X1 U21748 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19670), .B1(
        n19669), .B2(n19546), .ZN(n19522) );
  OAI211_X1 U21749 ( .C1(n19673), .C2(n19543), .A(n19523), .B(n19522), .ZN(
        P3_U2951) );
  AOI22_X1 U21750 ( .A1(n19686), .A2(n19545), .B1(n19674), .B2(n19544), .ZN(
        n19525) );
  AOI22_X1 U21751 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19676), .B1(
        n19675), .B2(n19546), .ZN(n19524) );
  OAI211_X1 U21752 ( .C1(n19679), .C2(n19549), .A(n19525), .B(n19524), .ZN(
        P3_U2943) );
  AOI22_X1 U21753 ( .A1(n19692), .A2(n19545), .B1(n19680), .B2(n19544), .ZN(
        n19527) );
  AOI22_X1 U21754 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19682), .B1(
        n19681), .B2(n19546), .ZN(n19526) );
  OAI211_X1 U21755 ( .C1(n19690), .C2(n19549), .A(n19527), .B(n19526), .ZN(
        P3_U2935) );
  AOI22_X1 U21756 ( .A1(n19698), .A2(n19545), .B1(n19685), .B2(n19544), .ZN(
        n19529) );
  AOI22_X1 U21757 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19687), .B1(
        n19686), .B2(n19546), .ZN(n19528) );
  OAI211_X1 U21758 ( .C1(n19696), .C2(n19549), .A(n19529), .B(n19528), .ZN(
        P3_U2927) );
  AOI22_X1 U21759 ( .A1(n19710), .A2(n19540), .B1(n19691), .B2(n19544), .ZN(
        n19531) );
  AOI22_X1 U21760 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19693), .B1(
        n19692), .B2(n19546), .ZN(n19530) );
  OAI211_X1 U21761 ( .C1(n19696), .C2(n19543), .A(n19531), .B(n19530), .ZN(
        P3_U2919) );
  AOI22_X1 U21762 ( .A1(n19710), .A2(n19545), .B1(n19697), .B2(n19544), .ZN(
        n19533) );
  AOI22_X1 U21763 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19699), .B1(
        n19698), .B2(n19546), .ZN(n19532) );
  OAI211_X1 U21764 ( .C1(n19620), .C2(n19549), .A(n19533), .B(n19532), .ZN(
        P3_U2911) );
  AOI22_X1 U21765 ( .A1(n19724), .A2(n19540), .B1(n19703), .B2(n19544), .ZN(
        n19535) );
  AOI22_X1 U21766 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19705), .B1(
        n19704), .B2(n19546), .ZN(n19534) );
  OAI211_X1 U21767 ( .C1(n19620), .C2(n19543), .A(n19535), .B(n19534), .ZN(
        P3_U2903) );
  AOI22_X1 U21768 ( .A1(n19734), .A2(n19540), .B1(n19708), .B2(n19544), .ZN(
        n19537) );
  AOI22_X1 U21769 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19711), .B1(
        n19710), .B2(n19546), .ZN(n19536) );
  OAI211_X1 U21770 ( .C1(n19715), .C2(n19543), .A(n19537), .B(n19536), .ZN(
        P3_U2895) );
  AOI22_X1 U21771 ( .A1(n19734), .A2(n19545), .B1(n19716), .B2(n19544), .ZN(
        n19539) );
  AOI22_X1 U21772 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19718), .B1(
        n19717), .B2(n19546), .ZN(n19538) );
  OAI211_X1 U21773 ( .C1(n19721), .C2(n19549), .A(n19539), .B(n19538), .ZN(
        P3_U2887) );
  AOI22_X1 U21774 ( .A1(n19732), .A2(n19540), .B1(n19722), .B2(n19544), .ZN(
        n19542) );
  AOI22_X1 U21775 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19725), .B1(
        n19724), .B2(n19546), .ZN(n19541) );
  OAI211_X1 U21776 ( .C1(n19721), .C2(n19543), .A(n19542), .B(n19541), .ZN(
        P3_U2879) );
  AOI22_X1 U21777 ( .A1(n19732), .A2(n19545), .B1(n19730), .B2(n19544), .ZN(
        n19548) );
  AOI22_X1 U21778 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19735), .B1(
        n19734), .B2(n19546), .ZN(n19547) );
  OAI211_X1 U21779 ( .C1(n19739), .C2(n19549), .A(n19548), .B(n19547), .ZN(
        P3_U2871) );
  OAI22_X1 U21780 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n19593), .ZN(n19550) );
  INV_X1 U21781 ( .A(n19550), .ZN(U253) );
  NOR2_X1 U21782 ( .A1(n16774), .A2(n19551), .ZN(n19583) );
  NAND2_X1 U21783 ( .A1(n19639), .A2(BUF2_REG_18__SCAN_IN), .ZN(n19586) );
  INV_X1 U21784 ( .A(n19586), .ZN(n19588) );
  INV_X1 U21785 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n21228) );
  NOR2_X2 U21786 ( .A1(n19552), .A2(n21228), .ZN(n19587) );
  AOI22_X1 U21787 ( .A1(n19652), .A2(n19588), .B1(n19641), .B2(n19587), .ZN(
        n19555) );
  NOR2_X2 U21788 ( .A1(n19553), .A2(n19642), .ZN(n19589) );
  AOI22_X1 U21789 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19643), .B1(
        n19723), .B2(n19589), .ZN(n19554) );
  OAI211_X1 U21790 ( .C1(n19556), .C2(n19592), .A(n19555), .B(n19554), .ZN(
        P3_U2990) );
  AOI22_X1 U21791 ( .A1(n19658), .A2(n19588), .B1(n19646), .B2(n19587), .ZN(
        n19558) );
  AOI22_X1 U21792 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19647), .B1(
        n19732), .B2(n19589), .ZN(n19557) );
  OAI211_X1 U21793 ( .C1(n19650), .C2(n19592), .A(n19558), .B(n19557), .ZN(
        P3_U2982) );
  AOI22_X1 U21794 ( .A1(n19663), .A2(n19588), .B1(n19651), .B2(n19587), .ZN(
        n19560) );
  AOI22_X1 U21795 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19653), .B1(
        n19652), .B2(n19589), .ZN(n19559) );
  OAI211_X1 U21796 ( .C1(n19656), .C2(n19592), .A(n19560), .B(n19559), .ZN(
        P3_U2974) );
  AOI22_X1 U21797 ( .A1(n19675), .A2(n19583), .B1(n19657), .B2(n19587), .ZN(
        n19562) );
  AOI22_X1 U21798 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19659), .B1(
        n19658), .B2(n19589), .ZN(n19561) );
  OAI211_X1 U21799 ( .C1(n19656), .C2(n19586), .A(n19562), .B(n19561), .ZN(
        P3_U2966) );
  AOI22_X1 U21800 ( .A1(n19675), .A2(n19588), .B1(n19662), .B2(n19587), .ZN(
        n19564) );
  AOI22_X1 U21801 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19664), .B1(
        n19663), .B2(n19589), .ZN(n19563) );
  OAI211_X1 U21802 ( .C1(n19673), .C2(n19592), .A(n19564), .B(n19563), .ZN(
        P3_U2958) );
  AOI22_X1 U21803 ( .A1(n19681), .A2(n19588), .B1(n19668), .B2(n19587), .ZN(
        n19566) );
  AOI22_X1 U21804 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19670), .B1(
        n19669), .B2(n19589), .ZN(n19565) );
  OAI211_X1 U21805 ( .C1(n19609), .C2(n19592), .A(n19566), .B(n19565), .ZN(
        P3_U2950) );
  AOI22_X1 U21806 ( .A1(n19692), .A2(n19583), .B1(n19674), .B2(n19587), .ZN(
        n19568) );
  AOI22_X1 U21807 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19676), .B1(
        n19675), .B2(n19589), .ZN(n19567) );
  OAI211_X1 U21808 ( .C1(n19609), .C2(n19586), .A(n19568), .B(n19567), .ZN(
        P3_U2942) );
  AOI22_X1 U21809 ( .A1(n19692), .A2(n19588), .B1(n19680), .B2(n19587), .ZN(
        n19570) );
  AOI22_X1 U21810 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19682), .B1(
        n19681), .B2(n19589), .ZN(n19569) );
  OAI211_X1 U21811 ( .C1(n19690), .C2(n19592), .A(n19570), .B(n19569), .ZN(
        P3_U2934) );
  AOI22_X1 U21812 ( .A1(n19704), .A2(n19583), .B1(n19685), .B2(n19587), .ZN(
        n19572) );
  AOI22_X1 U21813 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19687), .B1(
        n19686), .B2(n19589), .ZN(n19571) );
  OAI211_X1 U21814 ( .C1(n19690), .C2(n19586), .A(n19572), .B(n19571), .ZN(
        P3_U2926) );
  AOI22_X1 U21815 ( .A1(n19710), .A2(n19583), .B1(n19691), .B2(n19587), .ZN(
        n19574) );
  AOI22_X1 U21816 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19693), .B1(
        n19692), .B2(n19589), .ZN(n19573) );
  OAI211_X1 U21817 ( .C1(n19696), .C2(n19586), .A(n19574), .B(n19573), .ZN(
        P3_U2918) );
  AOI22_X1 U21818 ( .A1(n19710), .A2(n19588), .B1(n19697), .B2(n19587), .ZN(
        n19576) );
  AOI22_X1 U21819 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19699), .B1(
        n19698), .B2(n19589), .ZN(n19575) );
  OAI211_X1 U21820 ( .C1(n19620), .C2(n19592), .A(n19576), .B(n19575), .ZN(
        P3_U2910) );
  AOI22_X1 U21821 ( .A1(n19724), .A2(n19583), .B1(n19703), .B2(n19587), .ZN(
        n19578) );
  AOI22_X1 U21822 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19705), .B1(
        n19704), .B2(n19589), .ZN(n19577) );
  OAI211_X1 U21823 ( .C1(n19620), .C2(n19586), .A(n19578), .B(n19577), .ZN(
        P3_U2902) );
  AOI22_X1 U21824 ( .A1(n19724), .A2(n19588), .B1(n19708), .B2(n19587), .ZN(
        n19580) );
  AOI22_X1 U21825 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19711), .B1(
        n19710), .B2(n19589), .ZN(n19579) );
  OAI211_X1 U21826 ( .C1(n19627), .C2(n19592), .A(n19580), .B(n19579), .ZN(
        P3_U2894) );
  AOI22_X1 U21827 ( .A1(n19734), .A2(n19588), .B1(n19716), .B2(n19587), .ZN(
        n19582) );
  AOI22_X1 U21828 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19718), .B1(
        n19717), .B2(n19589), .ZN(n19581) );
  OAI211_X1 U21829 ( .C1(n19721), .C2(n19592), .A(n19582), .B(n19581), .ZN(
        P3_U2886) );
  AOI22_X1 U21830 ( .A1(n19732), .A2(n19583), .B1(n19722), .B2(n19587), .ZN(
        n19585) );
  AOI22_X1 U21831 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19725), .B1(
        n19724), .B2(n19589), .ZN(n19584) );
  OAI211_X1 U21832 ( .C1(n19721), .C2(n19586), .A(n19585), .B(n19584), .ZN(
        P3_U2878) );
  AOI22_X1 U21833 ( .A1(n19732), .A2(n19588), .B1(n19730), .B2(n19587), .ZN(
        n19591) );
  AOI22_X1 U21834 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19735), .B1(
        n19734), .B2(n19589), .ZN(n19590) );
  OAI211_X1 U21835 ( .C1(n19739), .C2(n19592), .A(n19591), .B(n19590), .ZN(
        P3_U2870) );
  OAI22_X1 U21836 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19593), .ZN(n19594) );
  INV_X1 U21837 ( .A(n19594), .ZN(U252) );
  NAND2_X1 U21838 ( .A1(n19639), .A2(BUF2_REG_17__SCAN_IN), .ZN(n19626) );
  NAND2_X1 U21839 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19639), .ZN(n19635) );
  INV_X1 U21840 ( .A(n19635), .ZN(n19623) );
  AND2_X1 U21841 ( .A1(n19640), .A2(BUF2_REG_1__SCAN_IN), .ZN(n19630) );
  AOI22_X1 U21842 ( .A1(n19658), .A2(n19623), .B1(n19641), .B2(n19630), .ZN(
        n19596) );
  NOR2_X2 U21843 ( .A1(n20738), .A2(n19642), .ZN(n19632) );
  AOI22_X1 U21844 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19643), .B1(
        n19723), .B2(n19632), .ZN(n19595) );
  OAI211_X1 U21845 ( .C1(n19739), .C2(n19626), .A(n19596), .B(n19595), .ZN(
        P3_U2989) );
  INV_X1 U21846 ( .A(n19626), .ZN(n19631) );
  AOI22_X1 U21847 ( .A1(n19658), .A2(n19631), .B1(n19646), .B2(n19630), .ZN(
        n19598) );
  AOI22_X1 U21848 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19647), .B1(
        n19732), .B2(n19632), .ZN(n19597) );
  OAI211_X1 U21849 ( .C1(n19650), .C2(n19635), .A(n19598), .B(n19597), .ZN(
        P3_U2981) );
  AOI22_X1 U21850 ( .A1(n19663), .A2(n19631), .B1(n19651), .B2(n19630), .ZN(
        n19600) );
  AOI22_X1 U21851 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19653), .B1(
        n19652), .B2(n19632), .ZN(n19599) );
  OAI211_X1 U21852 ( .C1(n19656), .C2(n19635), .A(n19600), .B(n19599), .ZN(
        P3_U2973) );
  AOI22_X1 U21853 ( .A1(n19669), .A2(n19631), .B1(n19657), .B2(n19630), .ZN(
        n19602) );
  AOI22_X1 U21854 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19659), .B1(
        n19658), .B2(n19632), .ZN(n19601) );
  OAI211_X1 U21855 ( .C1(n19667), .C2(n19635), .A(n19602), .B(n19601), .ZN(
        P3_U2965) );
  AOI22_X1 U21856 ( .A1(n19675), .A2(n19631), .B1(n19662), .B2(n19630), .ZN(
        n19604) );
  AOI22_X1 U21857 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19664), .B1(
        n19663), .B2(n19632), .ZN(n19603) );
  OAI211_X1 U21858 ( .C1(n19673), .C2(n19635), .A(n19604), .B(n19603), .ZN(
        P3_U2957) );
  AOI22_X1 U21859 ( .A1(n19686), .A2(n19623), .B1(n19668), .B2(n19630), .ZN(
        n19606) );
  AOI22_X1 U21860 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19670), .B1(
        n19669), .B2(n19632), .ZN(n19605) );
  OAI211_X1 U21861 ( .C1(n19673), .C2(n19626), .A(n19606), .B(n19605), .ZN(
        P3_U2949) );
  AOI22_X1 U21862 ( .A1(n19692), .A2(n19623), .B1(n19674), .B2(n19630), .ZN(
        n19608) );
  AOI22_X1 U21863 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19676), .B1(
        n19675), .B2(n19632), .ZN(n19607) );
  OAI211_X1 U21864 ( .C1(n19609), .C2(n19626), .A(n19608), .B(n19607), .ZN(
        P3_U2941) );
  AOI22_X1 U21865 ( .A1(n19692), .A2(n19631), .B1(n19680), .B2(n19630), .ZN(
        n19611) );
  AOI22_X1 U21866 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19682), .B1(
        n19681), .B2(n19632), .ZN(n19610) );
  OAI211_X1 U21867 ( .C1(n19690), .C2(n19635), .A(n19611), .B(n19610), .ZN(
        P3_U2933) );
  AOI22_X1 U21868 ( .A1(n19704), .A2(n19623), .B1(n19685), .B2(n19630), .ZN(
        n19613) );
  AOI22_X1 U21869 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19687), .B1(
        n19686), .B2(n19632), .ZN(n19612) );
  OAI211_X1 U21870 ( .C1(n19690), .C2(n19626), .A(n19613), .B(n19612), .ZN(
        P3_U2925) );
  AOI22_X1 U21871 ( .A1(n19710), .A2(n19623), .B1(n19691), .B2(n19630), .ZN(
        n19615) );
  AOI22_X1 U21872 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19693), .B1(
        n19692), .B2(n19632), .ZN(n19614) );
  OAI211_X1 U21873 ( .C1(n19696), .C2(n19626), .A(n19615), .B(n19614), .ZN(
        P3_U2917) );
  AOI22_X1 U21874 ( .A1(n19710), .A2(n19631), .B1(n19697), .B2(n19630), .ZN(
        n19617) );
  AOI22_X1 U21875 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19699), .B1(
        n19698), .B2(n19632), .ZN(n19616) );
  OAI211_X1 U21876 ( .C1(n19620), .C2(n19635), .A(n19617), .B(n19616), .ZN(
        P3_U2909) );
  AOI22_X1 U21877 ( .A1(n19724), .A2(n19623), .B1(n19703), .B2(n19630), .ZN(
        n19619) );
  AOI22_X1 U21878 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19705), .B1(
        n19704), .B2(n19632), .ZN(n19618) );
  OAI211_X1 U21879 ( .C1(n19620), .C2(n19626), .A(n19619), .B(n19618), .ZN(
        P3_U2901) );
  AOI22_X1 U21880 ( .A1(n19734), .A2(n19623), .B1(n19708), .B2(n19630), .ZN(
        n19622) );
  AOI22_X1 U21881 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19711), .B1(
        n19710), .B2(n19632), .ZN(n19621) );
  OAI211_X1 U21882 ( .C1(n19715), .C2(n19626), .A(n19622), .B(n19621), .ZN(
        P3_U2893) );
  AOI22_X1 U21883 ( .A1(n19723), .A2(n19623), .B1(n19716), .B2(n19630), .ZN(
        n19625) );
  AOI22_X1 U21884 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19718), .B1(
        n19717), .B2(n19632), .ZN(n19624) );
  OAI211_X1 U21885 ( .C1(n19627), .C2(n19626), .A(n19625), .B(n19624), .ZN(
        P3_U2885) );
  AOI22_X1 U21886 ( .A1(n19723), .A2(n19631), .B1(n19722), .B2(n19630), .ZN(
        n19629) );
  AOI22_X1 U21887 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19725), .B1(
        n19724), .B2(n19632), .ZN(n19628) );
  OAI211_X1 U21888 ( .C1(n19728), .C2(n19635), .A(n19629), .B(n19628), .ZN(
        P3_U2877) );
  AOI22_X1 U21889 ( .A1(n19732), .A2(n19631), .B1(n19730), .B2(n19630), .ZN(
        n19634) );
  AOI22_X1 U21890 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19735), .B1(
        n19734), .B2(n19632), .ZN(n19633) );
  OAI211_X1 U21891 ( .C1(n19739), .C2(n19635), .A(n19634), .B(n19633), .ZN(
        P3_U2869) );
  OAI22_X1 U21892 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n19636), .ZN(n19638) );
  INV_X1 U21893 ( .A(n19638), .ZN(U251) );
  NAND2_X1 U21894 ( .A1(n19639), .A2(BUF2_REG_16__SCAN_IN), .ZN(n19714) );
  NAND2_X1 U21895 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19639), .ZN(n19738) );
  INV_X1 U21896 ( .A(n19738), .ZN(n19709) );
  AND2_X1 U21897 ( .A1(n19640), .A2(BUF2_REG_0__SCAN_IN), .ZN(n19729) );
  AOI22_X1 U21898 ( .A1(n19658), .A2(n19709), .B1(n19641), .B2(n19729), .ZN(
        n19645) );
  NOR2_X2 U21899 ( .A1(n20736), .A2(n19642), .ZN(n19733) );
  AOI22_X1 U21900 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19643), .B1(
        n19723), .B2(n19733), .ZN(n19644) );
  OAI211_X1 U21901 ( .C1(n19739), .C2(n19714), .A(n19645), .B(n19644), .ZN(
        P3_U2988) );
  INV_X1 U21902 ( .A(n19714), .ZN(n19731) );
  AOI22_X1 U21903 ( .A1(n19658), .A2(n19731), .B1(n19646), .B2(n19729), .ZN(
        n19649) );
  AOI22_X1 U21904 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19647), .B1(
        n19732), .B2(n19733), .ZN(n19648) );
  OAI211_X1 U21905 ( .C1(n19650), .C2(n19738), .A(n19649), .B(n19648), .ZN(
        P3_U2980) );
  AOI22_X1 U21906 ( .A1(n19663), .A2(n19731), .B1(n19651), .B2(n19729), .ZN(
        n19655) );
  AOI22_X1 U21907 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19653), .B1(
        n19652), .B2(n19733), .ZN(n19654) );
  OAI211_X1 U21908 ( .C1(n19656), .C2(n19738), .A(n19655), .B(n19654), .ZN(
        P3_U2972) );
  AOI22_X1 U21909 ( .A1(n19669), .A2(n19731), .B1(n19657), .B2(n19729), .ZN(
        n19661) );
  AOI22_X1 U21910 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19659), .B1(
        n19658), .B2(n19733), .ZN(n19660) );
  OAI211_X1 U21911 ( .C1(n19667), .C2(n19738), .A(n19661), .B(n19660), .ZN(
        P3_U2964) );
  AOI22_X1 U21912 ( .A1(n19681), .A2(n19709), .B1(n19662), .B2(n19729), .ZN(
        n19666) );
  AOI22_X1 U21913 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19664), .B1(
        n19663), .B2(n19733), .ZN(n19665) );
  OAI211_X1 U21914 ( .C1(n19667), .C2(n19714), .A(n19666), .B(n19665), .ZN(
        P3_U2956) );
  AOI22_X1 U21915 ( .A1(n19686), .A2(n19709), .B1(n19668), .B2(n19729), .ZN(
        n19672) );
  AOI22_X1 U21916 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19670), .B1(
        n19669), .B2(n19733), .ZN(n19671) );
  OAI211_X1 U21917 ( .C1(n19673), .C2(n19714), .A(n19672), .B(n19671), .ZN(
        P3_U2948) );
  AOI22_X1 U21918 ( .A1(n19686), .A2(n19731), .B1(n19674), .B2(n19729), .ZN(
        n19678) );
  AOI22_X1 U21919 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19676), .B1(
        n19675), .B2(n19733), .ZN(n19677) );
  OAI211_X1 U21920 ( .C1(n19679), .C2(n19738), .A(n19678), .B(n19677), .ZN(
        P3_U2940) );
  AOI22_X1 U21921 ( .A1(n19692), .A2(n19731), .B1(n19680), .B2(n19729), .ZN(
        n19684) );
  AOI22_X1 U21922 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19682), .B1(
        n19681), .B2(n19733), .ZN(n19683) );
  OAI211_X1 U21923 ( .C1(n19690), .C2(n19738), .A(n19684), .B(n19683), .ZN(
        P3_U2932) );
  AOI22_X1 U21924 ( .A1(n19704), .A2(n19709), .B1(n19685), .B2(n19729), .ZN(
        n19689) );
  AOI22_X1 U21925 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19687), .B1(
        n19686), .B2(n19733), .ZN(n19688) );
  OAI211_X1 U21926 ( .C1(n19690), .C2(n19714), .A(n19689), .B(n19688), .ZN(
        P3_U2924) );
  AOI22_X1 U21927 ( .A1(n19710), .A2(n19709), .B1(n19691), .B2(n19729), .ZN(
        n19695) );
  AOI22_X1 U21928 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19693), .B1(
        n19692), .B2(n19733), .ZN(n19694) );
  OAI211_X1 U21929 ( .C1(n19696), .C2(n19714), .A(n19695), .B(n19694), .ZN(
        P3_U2916) );
  AOI22_X1 U21930 ( .A1(n19697), .A2(n19729), .B1(n19717), .B2(n19709), .ZN(
        n19701) );
  AOI22_X1 U21931 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19699), .B1(
        n19698), .B2(n19733), .ZN(n19700) );
  OAI211_X1 U21932 ( .C1(n19702), .C2(n19714), .A(n19701), .B(n19700), .ZN(
        P3_U2908) );
  AOI22_X1 U21933 ( .A1(n19717), .A2(n19731), .B1(n19703), .B2(n19729), .ZN(
        n19707) );
  AOI22_X1 U21934 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19705), .B1(
        n19704), .B2(n19733), .ZN(n19706) );
  OAI211_X1 U21935 ( .C1(n19715), .C2(n19738), .A(n19707), .B(n19706), .ZN(
        P3_U2900) );
  AOI22_X1 U21936 ( .A1(n19734), .A2(n19709), .B1(n19708), .B2(n19729), .ZN(
        n19713) );
  AOI22_X1 U21937 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19711), .B1(
        n19710), .B2(n19733), .ZN(n19712) );
  OAI211_X1 U21938 ( .C1(n19715), .C2(n19714), .A(n19713), .B(n19712), .ZN(
        P3_U2892) );
  AOI22_X1 U21939 ( .A1(n19734), .A2(n19731), .B1(n19716), .B2(n19729), .ZN(
        n19720) );
  AOI22_X1 U21940 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19718), .B1(
        n19717), .B2(n19733), .ZN(n19719) );
  OAI211_X1 U21941 ( .C1(n19721), .C2(n19738), .A(n19720), .B(n19719), .ZN(
        P3_U2884) );
  AOI22_X1 U21942 ( .A1(n19723), .A2(n19731), .B1(n19722), .B2(n19729), .ZN(
        n19727) );
  AOI22_X1 U21943 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19725), .B1(
        n19724), .B2(n19733), .ZN(n19726) );
  OAI211_X1 U21944 ( .C1(n19728), .C2(n19738), .A(n19727), .B(n19726), .ZN(
        P3_U2876) );
  AOI22_X1 U21945 ( .A1(n19732), .A2(n19731), .B1(n19730), .B2(n19729), .ZN(
        n19737) );
  AOI22_X1 U21946 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19735), .B1(
        n19734), .B2(n19733), .ZN(n19736) );
  OAI211_X1 U21947 ( .C1(n19739), .C2(n19738), .A(n19737), .B(n19736), .ZN(
        P3_U2868) );
  AOI22_X1 U21948 ( .A1(n19158), .A2(n20067), .B1(BUF1_REG_31__SCAN_IN), .B2(
        n20064), .ZN(n19741) );
  AOI22_X1 U21949 ( .A1(n20063), .A2(BUF2_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n20060), .ZN(n19740) );
  NAND2_X1 U21950 ( .A1(n19741), .A2(n19740), .ZN(P2_U2888) );
  AOI22_X1 U21951 ( .A1(n20011), .A2(n19742), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n20060), .ZN(n19743) );
  OAI21_X1 U21952 ( .B1(n20018), .B2(n19744), .A(n19743), .ZN(P2_U2905) );
  AOI22_X1 U21953 ( .A1(n20011), .A2(n19745), .B1(P2_EAX_REG_12__SCAN_IN), 
        .B2(n20060), .ZN(n19746) );
  OAI21_X1 U21954 ( .B1(n20018), .B2(n19747), .A(n19746), .ZN(P2_U2907) );
  AOI22_X1 U21955 ( .A1(n20011), .A2(n19748), .B1(P2_EAX_REG_10__SCAN_IN), 
        .B2(n20060), .ZN(n19749) );
  OAI21_X1 U21956 ( .B1(n20018), .B2(n19750), .A(n19749), .ZN(P2_U2909) );
  OAI22_X1 U21957 ( .A1(n20667), .A2(n19764), .B1(n19753), .B2(n19765), .ZN(
        n19952) );
  INV_X1 U21958 ( .A(n19952), .ZN(n19939) );
  NAND3_X1 U21959 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19769) );
  INV_X1 U21960 ( .A(n19755), .ZN(n20248) );
  OAI21_X1 U21961 ( .B1(n19754), .B2(n20248), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19756) );
  OAI21_X1 U21962 ( .B1(n19769), .B2(n19942), .A(n19756), .ZN(n20249) );
  NOR2_X2 U21963 ( .A1(n19757), .A2(n20244), .ZN(n19957) );
  AOI22_X1 U21964 ( .A1(n20249), .A2(n19957), .B1(n20248), .B2(n19951), .ZN(
        n19767) );
  INV_X1 U21965 ( .A(n19768), .ZN(n19759) );
  OAI21_X1 U21966 ( .B1(n19759), .B2(n19844), .A(n19769), .ZN(n19763) );
  NAND2_X1 U21967 ( .A1(n19760), .A2(n19916), .ZN(n19945) );
  INV_X1 U21968 ( .A(n19945), .ZN(n19933) );
  AOI211_X1 U21969 ( .C1(n19754), .C2(n19933), .A(n20248), .B(n19932), .ZN(
        n19761) );
  NOR2_X1 U21970 ( .A1(n20244), .A2(n19761), .ZN(n19762) );
  NAND2_X1 U21971 ( .A1(n19763), .A2(n19762), .ZN(n20252) );
  NAND2_X1 U21972 ( .A1(n19768), .A2(n19881), .ZN(n20199) );
  AOI22_X1 U21973 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20252), .B1(
        n19956), .B2(n20348), .ZN(n19766) );
  OAI211_X1 U21974 ( .C1(n19939), .C2(n20261), .A(n19767), .B(n19766), .ZN(
        P2_U3175) );
  NAND2_X1 U21975 ( .A1(n19768), .A2(n19820), .ZN(n19783) );
  INV_X1 U21976 ( .A(n20267), .ZN(n20256) );
  NOR2_X1 U21977 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19769), .ZN(
        n20255) );
  AOI22_X1 U21978 ( .A1(n20256), .A2(n19952), .B1(n19951), .B2(n20255), .ZN(
        n19777) );
  NAND2_X1 U21979 ( .A1(n20267), .A2(n20261), .ZN(n19770) );
  AOI21_X1 U21980 ( .B1(n19770), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19942), 
        .ZN(n19773) );
  NAND3_X1 U21981 ( .A1(n19926), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19789) );
  NOR2_X1 U21982 ( .A1(n19927), .A2(n19789), .ZN(n20262) );
  INV_X1 U21983 ( .A(n20262), .ZN(n19780) );
  AOI21_X1 U21984 ( .B1(n11982), .B2(n19933), .A(n19902), .ZN(n19771) );
  AOI21_X1 U21985 ( .B1(n19773), .B2(n19780), .A(n19771), .ZN(n19772) );
  OAI21_X1 U21986 ( .B1(n20255), .B2(n20262), .A(n19773), .ZN(n19775) );
  OAI21_X1 U21987 ( .B1(n11982), .B2(n20255), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19774) );
  NAND2_X1 U21988 ( .A1(n19775), .A2(n19774), .ZN(n20257) );
  AOI22_X1 U21989 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20258), .B1(
        n19957), .B2(n20257), .ZN(n19776) );
  OAI211_X1 U21990 ( .C1(n19924), .C2(n20261), .A(n19777), .B(n19776), .ZN(
        P2_U3167) );
  OAI21_X1 U21991 ( .B1(n19778), .B2(n20262), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19779) );
  OAI21_X1 U21992 ( .B1(n19789), .B2(n19942), .A(n19779), .ZN(n20263) );
  AOI22_X1 U21993 ( .A1(n20263), .A2(n19957), .B1(n19951), .B2(n20262), .ZN(
        n19785) );
  OAI21_X1 U21994 ( .B1(n19783), .B2(n22292), .A(n19789), .ZN(n19782) );
  OAI211_X1 U21995 ( .C1(n11980), .C2(n19945), .A(n19780), .B(n19942), .ZN(
        n19781) );
  NAND3_X1 U21996 ( .A1(n19782), .A2(n19781), .A3(n19919), .ZN(n20264) );
  NOR2_X2 U21997 ( .A1(n19783), .A2(n19915), .ZN(n20270) );
  AOI22_X1 U21998 ( .A1(n20264), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n20270), .B2(n19952), .ZN(n19784) );
  OAI211_X1 U21999 ( .C1(n19924), .C2(n20267), .A(n19785), .B(n19784), .ZN(
        P2_U3159) );
  INV_X1 U22000 ( .A(n19786), .ZN(n19791) );
  INV_X1 U22001 ( .A(n19787), .ZN(n19788) );
  NAND2_X1 U22002 ( .A1(n19788), .A2(n19858), .ZN(n19885) );
  NOR2_X1 U22003 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19789), .ZN(
        n20268) );
  OAI21_X1 U22004 ( .B1(n11978), .B2(n20268), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19790) );
  OAI21_X1 U22005 ( .B1(n19791), .B2(n19885), .A(n19790), .ZN(n20269) );
  AOI22_X1 U22006 ( .A1(n20269), .A2(n19957), .B1(n19951), .B2(n20268), .ZN(
        n19798) );
  OAI21_X1 U22007 ( .B1(n20277), .B2(n20270), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19792) );
  OAI21_X1 U22008 ( .B1(n19885), .B2(n19809), .A(n19792), .ZN(n19796) );
  INV_X1 U22009 ( .A(n20268), .ZN(n19793) );
  OAI211_X1 U22010 ( .C1(n19794), .C2(n19945), .A(n19793), .B(n19942), .ZN(
        n19795) );
  NAND3_X1 U22011 ( .A1(n19796), .A2(n19795), .A3(n19919), .ZN(n20271) );
  AOI22_X1 U22012 ( .A1(n20271), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n20270), .B2(n19956), .ZN(n19797) );
  OAI211_X1 U22013 ( .C1(n19939), .C2(n20274), .A(n19798), .B(n19797), .ZN(
        P2_U3151) );
  NAND3_X1 U22014 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n19832), .ZN(n19807) );
  NOR2_X1 U22015 ( .A1(n19927), .A2(n19807), .ZN(n20275) );
  OAI21_X1 U22016 ( .B1(n19800), .B2(n20275), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19799) );
  OAI21_X1 U22017 ( .B1(n19807), .B2(n19942), .A(n19799), .ZN(n20276) );
  AOI22_X1 U22018 ( .A1(n20276), .A2(n19957), .B1(n19951), .B2(n20275), .ZN(
        n19806) );
  INV_X1 U22019 ( .A(n20275), .ZN(n19802) );
  NOR2_X1 U22020 ( .A1(n20275), .A2(n19800), .ZN(n19801) );
  AOI211_X1 U22021 ( .C1(n19945), .C2(n19802), .A(n20244), .B(n19801), .ZN(
        n19804) );
  OAI21_X1 U22022 ( .B1(n19880), .B2(n19898), .A(n19807), .ZN(n19803) );
  OAI21_X1 U22023 ( .B1(n19804), .B2(n19902), .A(n19803), .ZN(n20278) );
  AOI22_X1 U22024 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20278), .B1(
        n20208), .B2(n19952), .ZN(n19805) );
  OAI211_X1 U22025 ( .C1(n19924), .C2(n20274), .A(n19806), .B(n19805), .ZN(
        P2_U3143) );
  AND2_X1 U22026 ( .A1(n19820), .A2(n19915), .ZN(n19855) );
  NOR2_X1 U22027 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19807), .ZN(
        n20281) );
  AOI22_X1 U22028 ( .A1(n20288), .A2(n19952), .B1(n19951), .B2(n20281), .ZN(
        n19818) );
  OAI21_X1 U22029 ( .B1(n20288), .B2(n20208), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19808) );
  NAND2_X1 U22030 ( .A1(n19808), .A2(n19932), .ZN(n19816) );
  NOR3_X1 U22031 ( .A1(n19809), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19824) );
  INV_X1 U22032 ( .A(n19824), .ZN(n19830) );
  NOR2_X1 U22033 ( .A1(n19927), .A2(n19830), .ZN(n20287) );
  NOR2_X1 U22034 ( .A1(n20287), .A2(n20281), .ZN(n19815) );
  INV_X1 U22035 ( .A(n19815), .ZN(n19812) );
  AOI21_X1 U22036 ( .B1(n19813), .B2(n19916), .A(n20281), .ZN(n19810) );
  OAI21_X1 U22037 ( .B1(n19810), .B2(n20244), .A(n19944), .ZN(n19811) );
  OAI21_X1 U22038 ( .B1(n19813), .B2(n20281), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19814) );
  AOI22_X1 U22039 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20283), .B1(
        n19957), .B2(n20282), .ZN(n19817) );
  OAI211_X1 U22040 ( .C1(n19924), .C2(n20286), .A(n19818), .B(n19817), .ZN(
        P2_U3135) );
  AND2_X1 U22041 ( .A1(n19820), .A2(n19925), .ZN(n19865) );
  AOI22_X1 U22042 ( .A1(n20211), .A2(n19952), .B1(n19951), .B2(n20287), .ZN(
        n19829) );
  INV_X1 U22043 ( .A(n19819), .ZN(n19821) );
  NAND2_X1 U22044 ( .A1(n19820), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19867) );
  OAI21_X1 U22045 ( .B1(n19821), .B2(n19867), .A(n19932), .ZN(n19827) );
  NOR2_X1 U22046 ( .A1(n20244), .A2(n19822), .ZN(n19823) );
  OAI21_X1 U22047 ( .B1(n19827), .B2(n19824), .A(n19823), .ZN(n20290) );
  OAI21_X1 U22048 ( .B1(n19825), .B2(n20287), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19826) );
  OAI21_X1 U22049 ( .B1(n19827), .B2(n19830), .A(n19826), .ZN(n20289) );
  AOI22_X1 U22050 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20290), .B1(
        n19957), .B2(n20289), .ZN(n19828) );
  OAI211_X1 U22051 ( .C1(n19924), .C2(n20214), .A(n19829), .B(n19828), .ZN(
        P2_U3127) );
  NOR2_X1 U22052 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19830), .ZN(
        n20293) );
  AOI22_X1 U22053 ( .A1(n19956), .A2(n20211), .B1(n19951), .B2(n20293), .ZN(
        n19841) );
  NAND2_X1 U22054 ( .A1(n20298), .A2(n20219), .ZN(n19831) );
  AOI21_X1 U22055 ( .B1(n19831), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19942), 
        .ZN(n19836) );
  NOR2_X1 U22056 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19832), .ZN(
        n19883) );
  NAND2_X1 U22057 ( .A1(n19897), .A2(n19883), .ZN(n19845) );
  OAI21_X1 U22058 ( .B1(n19837), .B2(n19833), .A(n19916), .ZN(n19834) );
  AOI21_X1 U22059 ( .B1(n19836), .B2(n19845), .A(n19834), .ZN(n19835) );
  INV_X1 U22060 ( .A(n19845), .ZN(n20299) );
  OAI21_X1 U22061 ( .B1(n20299), .B2(n20293), .A(n19836), .ZN(n19839) );
  OAI21_X1 U22062 ( .B1(n19837), .B2(n20293), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19838) );
  NAND2_X1 U22063 ( .A1(n19839), .A2(n19838), .ZN(n20294) );
  AOI22_X1 U22064 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20295), .B1(
        n19957), .B2(n20294), .ZN(n19840) );
  OAI211_X1 U22065 ( .C1(n19939), .C2(n20219), .A(n19841), .B(n19840), .ZN(
        P2_U3119) );
  NAND2_X1 U22066 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19883), .ZN(
        n19850) );
  OAI21_X1 U22067 ( .B1(n19842), .B2(n20299), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19843) );
  OAI21_X1 U22068 ( .B1(n19850), .B2(n19942), .A(n19843), .ZN(n20300) );
  AOI22_X1 U22069 ( .A1(n20300), .A2(n19957), .B1(n20299), .B2(n19951), .ZN(
        n19849) );
  INV_X1 U22070 ( .A(n19866), .ZN(n19868) );
  OAI21_X1 U22071 ( .B1(n19868), .B2(n19844), .A(n19850), .ZN(n19847) );
  OAI211_X1 U22072 ( .C1(n11979), .C2(n19945), .A(n19942), .B(n19845), .ZN(
        n19846) );
  NAND3_X1 U22073 ( .A1(n19847), .A2(n19919), .A3(n19846), .ZN(n20302) );
  AOI22_X1 U22074 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20302), .B1(
        n20301), .B2(n19956), .ZN(n19848) );
  OAI211_X1 U22075 ( .C1(n19939), .C2(n20311), .A(n19849), .B(n19848), .ZN(
        P2_U3111) );
  INV_X1 U22076 ( .A(n19883), .ZN(n19854) );
  INV_X1 U22077 ( .A(n19911), .ZN(n19853) );
  NOR2_X1 U22078 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19850), .ZN(
        n20305) );
  OAI21_X1 U22079 ( .B1(n19851), .B2(n20305), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19852) );
  OAI21_X1 U22080 ( .B1(n19854), .B2(n19853), .A(n19852), .ZN(n20306) );
  AOI22_X1 U22081 ( .A1(n20306), .A2(n19957), .B1(n19951), .B2(n20305), .ZN(
        n19864) );
  INV_X1 U22082 ( .A(n20305), .ZN(n19856) );
  OAI211_X1 U22083 ( .C1(n19857), .C2(n19945), .A(n19942), .B(n19856), .ZN(
        n19862) );
  INV_X1 U22084 ( .A(n19858), .ZN(n19859) );
  NAND2_X1 U22085 ( .A1(n19859), .A2(n19883), .ZN(n19860) );
  OAI221_X1 U22086 ( .B1(n22292), .B2(n20311), .C1(n22292), .C2(n20317), .A(
        n19860), .ZN(n19861) );
  NAND3_X1 U22087 ( .A1(n19862), .A2(n19919), .A3(n19861), .ZN(n20307) );
  AOI22_X1 U22088 ( .A1(n20308), .A2(n19952), .B1(
        P2_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n20307), .ZN(n19863) );
  OAI211_X1 U22089 ( .C1(n19924), .C2(n20311), .A(n19864), .B(n19863), .ZN(
        P2_U3103) );
  NAND2_X1 U22090 ( .A1(n19866), .A2(n19865), .ZN(n19882) );
  NAND2_X1 U22091 ( .A1(n19883), .A2(n19926), .ZN(n19875) );
  NOR2_X1 U22092 ( .A1(n19927), .A2(n19875), .ZN(n20312) );
  AOI22_X1 U22093 ( .A1(n19956), .A2(n20308), .B1(n19951), .B2(n20312), .ZN(
        n19878) );
  OAI21_X1 U22094 ( .B1(n19868), .B2(n19867), .A(n19932), .ZN(n19876) );
  INV_X1 U22095 ( .A(n19875), .ZN(n19872) );
  OAI21_X1 U22096 ( .B1(n19932), .B2(n20312), .A(n19919), .ZN(n19869) );
  OAI21_X1 U22097 ( .B1(n19870), .B2(n19945), .A(n19869), .ZN(n19871) );
  OAI21_X1 U22098 ( .B1(n19876), .B2(n19872), .A(n19871), .ZN(n20314) );
  OAI21_X1 U22099 ( .B1(n19873), .B2(n20312), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19874) );
  OAI21_X1 U22100 ( .B1(n19876), .B2(n19875), .A(n19874), .ZN(n20313) );
  AOI22_X1 U22101 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20314), .B1(
        n19957), .B2(n20313), .ZN(n19877) );
  OAI211_X1 U22102 ( .C1(n19939), .C2(n19882), .A(n19878), .B(n19877), .ZN(
        P2_U3095) );
  NAND2_X1 U22103 ( .A1(n19880), .A2(n19879), .ZN(n19914) );
  NOR2_X1 U22104 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19941) );
  AND2_X1 U22105 ( .A1(n19941), .A2(n19883), .ZN(n20318) );
  AOI22_X1 U22106 ( .A1(n19956), .A2(n20319), .B1(n19951), .B2(n20318), .ZN(
        n19894) );
  OAI21_X1 U22107 ( .B1(n20326), .B2(n20319), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19884) );
  NAND2_X1 U22108 ( .A1(n19884), .A2(n19932), .ZN(n19892) );
  NOR2_X1 U22109 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19885), .ZN(
        n19888) );
  AOI21_X1 U22110 ( .B1(n19889), .B2(n19933), .A(n20318), .ZN(n19886) );
  OAI21_X1 U22111 ( .B1(n19886), .B2(n20244), .A(n19944), .ZN(n19887) );
  INV_X1 U22112 ( .A(n19888), .ZN(n19891) );
  OAI21_X1 U22113 ( .B1(n19889), .B2(n20318), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19890) );
  AOI22_X1 U22114 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20321), .B1(
        n19957), .B2(n20320), .ZN(n19893) );
  OAI211_X1 U22115 ( .C1(n19939), .C2(n20324), .A(n19894), .B(n19893), .ZN(
        P2_U3087) );
  INV_X1 U22116 ( .A(n20336), .ZN(n20228) );
  NOR2_X1 U22117 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19940) );
  AND2_X1 U22118 ( .A1(n19897), .A2(n19940), .ZN(n20325) );
  AOI22_X1 U22119 ( .A1(n20228), .A2(n19952), .B1(n19951), .B2(n20325), .ZN(
        n19909) );
  NOR2_X1 U22120 ( .A1(n19899), .A2(n19898), .ZN(n19907) );
  NAND2_X1 U22121 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19940), .ZN(
        n19910) );
  INV_X1 U22122 ( .A(n19910), .ZN(n19903) );
  AOI21_X1 U22123 ( .B1(n19904), .B2(n19933), .A(n20325), .ZN(n19900) );
  NOR2_X1 U22124 ( .A1(n20244), .A2(n19900), .ZN(n19901) );
  OAI22_X1 U22125 ( .A1(n19907), .A2(n19903), .B1(n19902), .B2(n19901), .ZN(
        n20328) );
  NAND2_X1 U22126 ( .A1(n19932), .A2(n19903), .ZN(n19906) );
  OAI21_X1 U22127 ( .B1(n19904), .B2(n20325), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19905) );
  OAI21_X1 U22128 ( .B1(n19907), .B2(n19906), .A(n19905), .ZN(n20327) );
  AOI22_X1 U22129 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20328), .B1(
        n19957), .B2(n20327), .ZN(n19908) );
  OAI211_X1 U22130 ( .C1(n19924), .C2(n20324), .A(n19909), .B(n19908), .ZN(
        P2_U3079) );
  NOR2_X1 U22131 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19910), .ZN(
        n20331) );
  OAI21_X1 U22132 ( .B1(n11969), .B2(n20331), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19912) );
  NAND2_X1 U22133 ( .A1(n19911), .A2(n19940), .ZN(n19917) );
  NAND2_X1 U22134 ( .A1(n19912), .A2(n19917), .ZN(n20332) );
  AOI22_X1 U22135 ( .A1(n20332), .A2(n19957), .B1(n19951), .B2(n20331), .ZN(
        n19923) );
  AOI211_X1 U22136 ( .C1(n20336), .C2(n20235), .A(n19942), .B(n22292), .ZN(
        n19921) );
  AOI21_X1 U22137 ( .B1(n11969), .B2(n19916), .A(n20331), .ZN(n19918) );
  OAI21_X1 U22138 ( .B1(n19918), .B2(n19932), .A(n19917), .ZN(n19920) );
  AOI22_X1 U22139 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20333), .B1(
        n20340), .B2(n19952), .ZN(n19922) );
  OAI211_X1 U22140 ( .C1(n19924), .C2(n20336), .A(n19923), .B(n19922), .ZN(
        P2_U3071) );
  NAND2_X1 U22141 ( .A1(n19929), .A2(n19925), .ZN(n20344) );
  NAND2_X1 U22142 ( .A1(n19940), .A2(n19926), .ZN(n19930) );
  NOR2_X1 U22143 ( .A1(n19927), .A2(n19930), .ZN(n20338) );
  OAI21_X1 U22144 ( .B1(n11972), .B2(n20338), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19928) );
  OAI21_X1 U22145 ( .B1(n19930), .B2(n19942), .A(n19928), .ZN(n20339) );
  AOI22_X1 U22146 ( .A1(n20339), .A2(n19957), .B1(n19951), .B2(n20338), .ZN(
        n19938) );
  INV_X1 U22147 ( .A(n19929), .ZN(n19931) );
  OAI21_X1 U22148 ( .B1(n19931), .B2(n22292), .A(n19930), .ZN(n19936) );
  NOR2_X1 U22149 ( .A1(n20244), .A2(n19934), .ZN(n19935) );
  NAND2_X1 U22150 ( .A1(n19936), .A2(n19935), .ZN(n20341) );
  AOI22_X1 U22151 ( .A1(n20341), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n19956), .B2(n20340), .ZN(n19937) );
  OAI211_X1 U22152 ( .C1(n19939), .C2(n20344), .A(n19938), .B(n19937), .ZN(
        P2_U3063) );
  NAND2_X1 U22153 ( .A1(n19941), .A2(n19940), .ZN(n19950) );
  AOI21_X1 U22154 ( .B1(n20344), .B2(n20199), .A(n22292), .ZN(n19943) );
  NOR2_X1 U22155 ( .A1(n19943), .A2(n19942), .ZN(n19953) );
  INV_X1 U22156 ( .A(n19953), .ZN(n19948) );
  INV_X1 U22157 ( .A(n11971), .ZN(n19946) );
  OAI21_X1 U22158 ( .B1(n19946), .B2(n19945), .A(n19944), .ZN(n19947) );
  OAI21_X1 U22159 ( .B1(n19948), .B2(n20248), .A(n19947), .ZN(n19949) );
  INV_X1 U22160 ( .A(n19950), .ZN(n20346) );
  AOI22_X1 U22161 ( .A1(n20348), .A2(n19952), .B1(n19951), .B2(n20346), .ZN(
        n19959) );
  OAI21_X1 U22162 ( .B1(n20248), .B2(n20346), .A(n19953), .ZN(n19955) );
  OAI21_X1 U22163 ( .B1(n11971), .B2(n20346), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19954) );
  NAND2_X1 U22164 ( .A1(n19955), .A2(n19954), .ZN(n20351) );
  AOI22_X1 U22165 ( .A1(n19957), .A2(n20351), .B1(n20353), .B2(n19956), .ZN(
        n19958) );
  OAI211_X1 U22166 ( .C1(n20357), .C2(n19960), .A(n19959), .B(n19958), .ZN(
        P2_U3055) );
  AOI22_X1 U22167 ( .A1(n20062), .A2(n19961), .B1(P2_EAX_REG_22__SCAN_IN), 
        .B2(n20060), .ZN(n19968) );
  AOI22_X1 U22168 ( .A1(n20064), .A2(BUF1_REG_22__SCAN_IN), .B1(n20063), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n19967) );
  INV_X1 U22169 ( .A(n19962), .ZN(n19965) );
  INV_X1 U22170 ( .A(n19963), .ZN(n19964) );
  AOI22_X1 U22171 ( .A1(n19965), .A2(n20068), .B1(n20067), .B2(n19964), .ZN(
        n19966) );
  NAND3_X1 U22172 ( .A1(n19968), .A2(n19967), .A3(n19966), .ZN(P2_U2897) );
  AOI22_X2 U22173 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20251), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n20250), .ZN(n20002) );
  NOR2_X2 U22174 ( .A1(n19969), .A2(n20244), .ZN(n20005) );
  NOR2_X2 U22175 ( .A1(n19970), .A2(n20154), .ZN(n20003) );
  AOI22_X1 U22176 ( .A1(n20249), .A2(n20005), .B1(n20248), .B2(n20003), .ZN(
        n19972) );
  AOI22_X1 U22177 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20251), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n20250), .ZN(n19997) );
  AOI22_X1 U22178 ( .A1(n20252), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n20196), .B2(n20004), .ZN(n19971) );
  OAI211_X1 U22179 ( .C1(n20002), .C2(n20199), .A(n19972), .B(n19971), .ZN(
        P2_U3174) );
  INV_X1 U22180 ( .A(n20002), .ZN(n20006) );
  AOI22_X1 U22181 ( .A1(n20006), .A2(n20196), .B1(n20255), .B2(n20003), .ZN(
        n19974) );
  AOI22_X1 U22182 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20258), .B1(
        n20005), .B2(n20257), .ZN(n19973) );
  OAI211_X1 U22183 ( .C1(n19997), .C2(n20267), .A(n19974), .B(n19973), .ZN(
        P2_U3166) );
  AOI22_X1 U22184 ( .A1(n20263), .A2(n20005), .B1(n20003), .B2(n20262), .ZN(
        n19976) );
  AOI22_X1 U22185 ( .A1(n20264), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n20270), .B2(n20004), .ZN(n19975) );
  OAI211_X1 U22186 ( .C1(n20002), .C2(n20267), .A(n19976), .B(n19975), .ZN(
        P2_U3158) );
  AOI22_X1 U22187 ( .A1(n20269), .A2(n20005), .B1(n20003), .B2(n20268), .ZN(
        n19978) );
  AOI22_X1 U22188 ( .A1(n20271), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n20270), .B2(n20006), .ZN(n19977) );
  OAI211_X1 U22189 ( .C1(n19997), .C2(n20274), .A(n19978), .B(n19977), .ZN(
        P2_U3150) );
  AOI22_X1 U22190 ( .A1(n20276), .A2(n20005), .B1(n20003), .B2(n20275), .ZN(
        n19980) );
  AOI22_X1 U22191 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20278), .B1(
        n20208), .B2(n20004), .ZN(n19979) );
  OAI211_X1 U22192 ( .C1(n20002), .C2(n20274), .A(n19980), .B(n19979), .ZN(
        P2_U3142) );
  AOI22_X1 U22193 ( .A1(n20004), .A2(n20288), .B1(n20281), .B2(n20003), .ZN(
        n19982) );
  AOI22_X1 U22194 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20283), .B1(
        n20005), .B2(n20282), .ZN(n19981) );
  OAI211_X1 U22195 ( .C1(n20002), .C2(n20286), .A(n19982), .B(n19981), .ZN(
        P2_U3134) );
  AOI22_X1 U22196 ( .A1(n20004), .A2(n20211), .B1(n20287), .B2(n20003), .ZN(
        n19984) );
  AOI22_X1 U22197 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20290), .B1(
        n20005), .B2(n20289), .ZN(n19983) );
  OAI211_X1 U22198 ( .C1(n20002), .C2(n20214), .A(n19984), .B(n19983), .ZN(
        P2_U3126) );
  AOI22_X1 U22199 ( .A1(n20004), .A2(n20301), .B1(n20293), .B2(n20003), .ZN(
        n19986) );
  AOI22_X1 U22200 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20295), .B1(
        n20005), .B2(n20294), .ZN(n19985) );
  OAI211_X1 U22201 ( .C1(n20002), .C2(n20298), .A(n19986), .B(n19985), .ZN(
        P2_U3118) );
  AOI22_X1 U22202 ( .A1(n20300), .A2(n20005), .B1(n20299), .B2(n20003), .ZN(
        n19988) );
  AOI22_X1 U22203 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20302), .B1(
        n20220), .B2(n20004), .ZN(n19987) );
  OAI211_X1 U22204 ( .C1(n20002), .C2(n20219), .A(n19988), .B(n19987), .ZN(
        P2_U3110) );
  AOI22_X1 U22205 ( .A1(n20306), .A2(n20005), .B1(n20003), .B2(n20305), .ZN(
        n19990) );
  AOI22_X1 U22206 ( .A1(n20004), .A2(n20308), .B1(
        P2_INSTQUEUE_REG_6__6__SCAN_IN), .B2(n20307), .ZN(n19989) );
  OAI211_X1 U22207 ( .C1(n20002), .C2(n20311), .A(n19990), .B(n19989), .ZN(
        P2_U3102) );
  AOI22_X1 U22208 ( .A1(n20004), .A2(n20319), .B1(n20003), .B2(n20312), .ZN(
        n19992) );
  AOI22_X1 U22209 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20314), .B1(
        n20005), .B2(n20313), .ZN(n19991) );
  OAI211_X1 U22210 ( .C1(n20002), .C2(n20317), .A(n19992), .B(n19991), .ZN(
        P2_U3094) );
  AOI22_X1 U22211 ( .A1(n20006), .A2(n20319), .B1(n20003), .B2(n20318), .ZN(
        n19994) );
  AOI22_X1 U22212 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20321), .B1(
        n20005), .B2(n20320), .ZN(n19993) );
  OAI211_X1 U22213 ( .C1(n19997), .C2(n20324), .A(n19994), .B(n19993), .ZN(
        P2_U3086) );
  AOI22_X1 U22214 ( .A1(n20006), .A2(n20326), .B1(n20325), .B2(n20003), .ZN(
        n19996) );
  AOI22_X1 U22215 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20328), .B1(
        n20005), .B2(n20327), .ZN(n19995) );
  OAI211_X1 U22216 ( .C1(n19997), .C2(n20336), .A(n19996), .B(n19995), .ZN(
        P2_U3078) );
  AOI22_X1 U22217 ( .A1(n20332), .A2(n20005), .B1(n20003), .B2(n20331), .ZN(
        n19999) );
  AOI22_X1 U22218 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20333), .B1(
        n20340), .B2(n20004), .ZN(n19998) );
  OAI211_X1 U22219 ( .C1(n20002), .C2(n20336), .A(n19999), .B(n19998), .ZN(
        P2_U3070) );
  AOI22_X1 U22220 ( .A1(n20339), .A2(n20005), .B1(n20003), .B2(n20338), .ZN(
        n20001) );
  AOI22_X1 U22221 ( .A1(n20341), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n20353), .B2(n20004), .ZN(n20000) );
  OAI211_X1 U22222 ( .C1(n20002), .C2(n20235), .A(n20001), .B(n20000), .ZN(
        P2_U3062) );
  AOI22_X1 U22223 ( .A1(n20004), .A2(n20348), .B1(n20346), .B2(n20003), .ZN(
        n20008) );
  AOI22_X1 U22224 ( .A1(n20353), .A2(n20006), .B1(n20351), .B2(n20005), .ZN(
        n20007) );
  OAI211_X1 U22225 ( .C1(n20357), .C2(n20009), .A(n20008), .B(n20007), .ZN(
        P2_U3054) );
  INV_X1 U22226 ( .A(n20019), .ZN(n20010) );
  AOI22_X1 U22227 ( .A1(n20011), .A2(n20010), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n20060), .ZN(n20016) );
  OR3_X1 U22228 ( .A1(n20014), .A2(n20013), .A3(n20012), .ZN(n20015) );
  OAI211_X1 U22229 ( .C1(n20018), .C2(n20017), .A(n20016), .B(n20015), .ZN(
        P2_U2914) );
  NOR2_X2 U22230 ( .A1(n20019), .A2(n20244), .ZN(n20055) );
  NOR2_X2 U22231 ( .A1(n20020), .A2(n20154), .ZN(n20053) );
  AOI22_X1 U22232 ( .A1(n20249), .A2(n20055), .B1(n20248), .B2(n20053), .ZN(
        n20022) );
  AOI22_X1 U22233 ( .A1(n20252), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n20054), .B2(n20348), .ZN(n20021) );
  OAI211_X1 U22234 ( .C1(n20045), .C2(n20261), .A(n20022), .B(n20021), .ZN(
        P2_U3173) );
  AOI22_X1 U22235 ( .A1(n20256), .A2(n20056), .B1(n20255), .B2(n20053), .ZN(
        n20024) );
  AOI22_X1 U22236 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20258), .B1(
        n20055), .B2(n20257), .ZN(n20023) );
  OAI211_X1 U22237 ( .C1(n20052), .C2(n20261), .A(n20024), .B(n20023), .ZN(
        P2_U3165) );
  AOI22_X1 U22238 ( .A1(n20263), .A2(n20055), .B1(n20053), .B2(n20262), .ZN(
        n20026) );
  AOI22_X1 U22239 ( .A1(n20264), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n20270), .B2(n20056), .ZN(n20025) );
  OAI211_X1 U22240 ( .C1(n20052), .C2(n20267), .A(n20026), .B(n20025), .ZN(
        P2_U3157) );
  AOI22_X1 U22241 ( .A1(n20269), .A2(n20055), .B1(n20053), .B2(n20268), .ZN(
        n20028) );
  AOI22_X1 U22242 ( .A1(n20271), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n20270), .B2(n20054), .ZN(n20027) );
  OAI211_X1 U22243 ( .C1(n20045), .C2(n20274), .A(n20028), .B(n20027), .ZN(
        P2_U3149) );
  AOI22_X1 U22244 ( .A1(n20276), .A2(n20055), .B1(n20053), .B2(n20275), .ZN(
        n20030) );
  AOI22_X1 U22245 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20278), .B1(
        n20277), .B2(n20054), .ZN(n20029) );
  OAI211_X1 U22246 ( .C1(n20045), .C2(n20286), .A(n20030), .B(n20029), .ZN(
        P2_U3141) );
  AOI22_X1 U22247 ( .A1(n20054), .A2(n20208), .B1(n20053), .B2(n20281), .ZN(
        n20032) );
  AOI22_X1 U22248 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20283), .B1(
        n20055), .B2(n20282), .ZN(n20031) );
  OAI211_X1 U22249 ( .C1(n20045), .C2(n20214), .A(n20032), .B(n20031), .ZN(
        P2_U3133) );
  AOI22_X1 U22250 ( .A1(n20054), .A2(n20288), .B1(n20053), .B2(n20287), .ZN(
        n20034) );
  AOI22_X1 U22251 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20290), .B1(
        n20055), .B2(n20289), .ZN(n20033) );
  OAI211_X1 U22252 ( .C1(n20045), .C2(n20298), .A(n20034), .B(n20033), .ZN(
        P2_U3125) );
  AOI22_X1 U22253 ( .A1(n20054), .A2(n20211), .B1(n20053), .B2(n20293), .ZN(
        n20036) );
  AOI22_X1 U22254 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20295), .B1(
        n20055), .B2(n20294), .ZN(n20035) );
  OAI211_X1 U22255 ( .C1(n20045), .C2(n20219), .A(n20036), .B(n20035), .ZN(
        P2_U3117) );
  AOI22_X1 U22256 ( .A1(n20300), .A2(n20055), .B1(n20299), .B2(n20053), .ZN(
        n20038) );
  AOI22_X1 U22257 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20302), .B1(
        n20301), .B2(n20054), .ZN(n20037) );
  OAI211_X1 U22258 ( .C1(n20045), .C2(n20311), .A(n20038), .B(n20037), .ZN(
        P2_U3109) );
  AOI22_X1 U22259 ( .A1(n20306), .A2(n20055), .B1(n20053), .B2(n20305), .ZN(
        n20040) );
  AOI22_X1 U22260 ( .A1(n20056), .A2(n20308), .B1(
        P2_INSTQUEUE_REG_6__5__SCAN_IN), .B2(n20307), .ZN(n20039) );
  OAI211_X1 U22261 ( .C1(n20052), .C2(n20311), .A(n20040), .B(n20039), .ZN(
        P2_U3101) );
  AOI22_X1 U22262 ( .A1(n20056), .A2(n20319), .B1(n20053), .B2(n20312), .ZN(
        n20042) );
  AOI22_X1 U22263 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20314), .B1(
        n20055), .B2(n20313), .ZN(n20041) );
  OAI211_X1 U22264 ( .C1(n20052), .C2(n20317), .A(n20042), .B(n20041), .ZN(
        P2_U3093) );
  AOI22_X1 U22265 ( .A1(n20054), .A2(n20319), .B1(n20053), .B2(n20318), .ZN(
        n20044) );
  AOI22_X1 U22266 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20321), .B1(
        n20055), .B2(n20320), .ZN(n20043) );
  OAI211_X1 U22267 ( .C1(n20045), .C2(n20324), .A(n20044), .B(n20043), .ZN(
        P2_U3085) );
  AOI22_X1 U22268 ( .A1(n20056), .A2(n20228), .B1(n20053), .B2(n20325), .ZN(
        n20047) );
  AOI22_X1 U22269 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20328), .B1(
        n20055), .B2(n20327), .ZN(n20046) );
  OAI211_X1 U22270 ( .C1(n20052), .C2(n20324), .A(n20047), .B(n20046), .ZN(
        P2_U3077) );
  AOI22_X1 U22271 ( .A1(n20332), .A2(n20055), .B1(n20053), .B2(n20331), .ZN(
        n20049) );
  AOI22_X1 U22272 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20333), .B1(
        n20340), .B2(n20056), .ZN(n20048) );
  OAI211_X1 U22273 ( .C1(n20052), .C2(n20336), .A(n20049), .B(n20048), .ZN(
        P2_U3069) );
  AOI22_X1 U22274 ( .A1(n20339), .A2(n20055), .B1(n20053), .B2(n20338), .ZN(
        n20051) );
  AOI22_X1 U22275 ( .A1(n20341), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n20353), .B2(n20056), .ZN(n20050) );
  OAI211_X1 U22276 ( .C1(n20052), .C2(n20235), .A(n20051), .B(n20050), .ZN(
        P2_U3061) );
  AOI22_X1 U22277 ( .A1(n20054), .A2(n20353), .B1(n20053), .B2(n20346), .ZN(
        n20058) );
  AOI22_X1 U22278 ( .A1(n20348), .A2(n20056), .B1(n20351), .B2(n20055), .ZN(
        n20057) );
  OAI211_X1 U22279 ( .C1(n20357), .C2(n20059), .A(n20058), .B(n20057), .ZN(
        P2_U3053) );
  AOI22_X1 U22280 ( .A1(n20062), .A2(n20061), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n20060), .ZN(n20072) );
  AOI22_X1 U22281 ( .A1(n20064), .A2(BUF1_REG_20__SCAN_IN), .B1(n20063), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n20071) );
  INV_X1 U22282 ( .A(n20065), .ZN(n20069) );
  AOI22_X1 U22283 ( .A1(n20069), .A2(n20068), .B1(n20067), .B2(n20066), .ZN(
        n20070) );
  NAND3_X1 U22284 ( .A1(n20072), .A2(n20071), .A3(n20070), .ZN(P2_U2899) );
  NOR2_X2 U22285 ( .A1(n20073), .A2(n20244), .ZN(n20108) );
  AOI22_X1 U22286 ( .A1(n20249), .A2(n20108), .B1(n20248), .B2(n11138), .ZN(
        n20075) );
  AOI22_X1 U22287 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20251), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n20250), .ZN(n20100) );
  AOI22_X1 U22288 ( .A1(n20252), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n20107), .B2(n20196), .ZN(n20074) );
  OAI211_X1 U22289 ( .C1(n20105), .C2(n20199), .A(n20075), .B(n20074), .ZN(
        P2_U3172) );
  INV_X1 U22290 ( .A(n20105), .ZN(n20109) );
  AOI22_X1 U22291 ( .A1(n20109), .A2(n20196), .B1(n20255), .B2(n11138), .ZN(
        n20077) );
  AOI22_X1 U22292 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20258), .B1(
        n20108), .B2(n20257), .ZN(n20076) );
  OAI211_X1 U22293 ( .C1(n20100), .C2(n20267), .A(n20077), .B(n20076), .ZN(
        P2_U3164) );
  AOI22_X1 U22294 ( .A1(n20263), .A2(n20108), .B1(n11138), .B2(n20262), .ZN(
        n20079) );
  AOI22_X1 U22295 ( .A1(n20264), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n20270), .B2(n20107), .ZN(n20078) );
  OAI211_X1 U22296 ( .C1(n20105), .C2(n20267), .A(n20079), .B(n20078), .ZN(
        P2_U3156) );
  AOI22_X1 U22297 ( .A1(n20269), .A2(n20108), .B1(n11138), .B2(n20268), .ZN(
        n20081) );
  AOI22_X1 U22298 ( .A1(n20271), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n20270), .B2(n20109), .ZN(n20080) );
  OAI211_X1 U22299 ( .C1(n20100), .C2(n20274), .A(n20081), .B(n20080), .ZN(
        P2_U3148) );
  AOI22_X1 U22300 ( .A1(n20276), .A2(n20108), .B1(n11138), .B2(n20275), .ZN(
        n20083) );
  AOI22_X1 U22301 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20278), .B1(
        n20277), .B2(n20109), .ZN(n20082) );
  OAI211_X1 U22302 ( .C1(n20100), .C2(n20286), .A(n20083), .B(n20082), .ZN(
        P2_U3140) );
  AOI22_X1 U22303 ( .A1(n20107), .A2(n20288), .B1(n20281), .B2(n11138), .ZN(
        n20085) );
  AOI22_X1 U22304 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20283), .B1(
        n20108), .B2(n20282), .ZN(n20084) );
  OAI211_X1 U22305 ( .C1(n20105), .C2(n20286), .A(n20085), .B(n20084), .ZN(
        P2_U3132) );
  AOI22_X1 U22306 ( .A1(n20107), .A2(n20211), .B1(n20287), .B2(n11138), .ZN(
        n20087) );
  AOI22_X1 U22307 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20290), .B1(
        n20108), .B2(n20289), .ZN(n20086) );
  OAI211_X1 U22308 ( .C1(n20105), .C2(n20214), .A(n20087), .B(n20086), .ZN(
        P2_U3124) );
  AOI22_X1 U22309 ( .A1(n20107), .A2(n20301), .B1(n20293), .B2(n11138), .ZN(
        n20089) );
  AOI22_X1 U22310 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20295), .B1(
        n20108), .B2(n20294), .ZN(n20088) );
  OAI211_X1 U22311 ( .C1(n20105), .C2(n20298), .A(n20089), .B(n20088), .ZN(
        P2_U3116) );
  AOI22_X1 U22312 ( .A1(n20300), .A2(n20108), .B1(n20299), .B2(n11138), .ZN(
        n20091) );
  AOI22_X1 U22313 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20302), .B1(
        n20220), .B2(n20107), .ZN(n20090) );
  OAI211_X1 U22314 ( .C1(n20105), .C2(n20219), .A(n20091), .B(n20090), .ZN(
        P2_U3108) );
  AOI22_X1 U22315 ( .A1(n20306), .A2(n20108), .B1(n11138), .B2(n20305), .ZN(
        n20093) );
  AOI22_X1 U22316 ( .A1(n20107), .A2(n20308), .B1(
        P2_INSTQUEUE_REG_6__4__SCAN_IN), .B2(n20307), .ZN(n20092) );
  OAI211_X1 U22317 ( .C1(n20105), .C2(n20311), .A(n20093), .B(n20092), .ZN(
        P2_U3100) );
  AOI22_X1 U22318 ( .A1(n20107), .A2(n20319), .B1(n11138), .B2(n20312), .ZN(
        n20095) );
  AOI22_X1 U22319 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20314), .B1(
        n20108), .B2(n20313), .ZN(n20094) );
  OAI211_X1 U22320 ( .C1(n20105), .C2(n20317), .A(n20095), .B(n20094), .ZN(
        P2_U3092) );
  AOI22_X1 U22321 ( .A1(n20109), .A2(n20319), .B1(n11138), .B2(n20318), .ZN(
        n20097) );
  AOI22_X1 U22322 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20321), .B1(
        n20108), .B2(n20320), .ZN(n20096) );
  OAI211_X1 U22323 ( .C1(n20100), .C2(n20324), .A(n20097), .B(n20096), .ZN(
        P2_U3084) );
  AOI22_X1 U22324 ( .A1(n20109), .A2(n20326), .B1(n20325), .B2(n11138), .ZN(
        n20099) );
  AOI22_X1 U22325 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20328), .B1(
        n20108), .B2(n20327), .ZN(n20098) );
  OAI211_X1 U22326 ( .C1(n20100), .C2(n20336), .A(n20099), .B(n20098), .ZN(
        P2_U3076) );
  AOI22_X1 U22327 ( .A1(n20332), .A2(n20108), .B1(n11138), .B2(n20331), .ZN(
        n20102) );
  AOI22_X1 U22328 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20333), .B1(
        n20340), .B2(n20107), .ZN(n20101) );
  OAI211_X1 U22329 ( .C1(n20105), .C2(n20336), .A(n20102), .B(n20101), .ZN(
        P2_U3068) );
  AOI22_X1 U22330 ( .A1(n20339), .A2(n20108), .B1(n11138), .B2(n20338), .ZN(
        n20104) );
  AOI22_X1 U22331 ( .A1(n20341), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n20353), .B2(n20107), .ZN(n20103) );
  OAI211_X1 U22332 ( .C1(n20105), .C2(n20235), .A(n20104), .B(n20103), .ZN(
        P2_U3060) );
  AOI22_X1 U22333 ( .A1(n20107), .A2(n20348), .B1(n20346), .B2(n11138), .ZN(
        n20111) );
  AOI22_X1 U22334 ( .A1(n20353), .A2(n20109), .B1(n20351), .B2(n20108), .ZN(
        n20110) );
  OAI211_X1 U22335 ( .C1(n20357), .C2(n20112), .A(n20111), .B(n20110), .ZN(
        P2_U3052) );
  NOR2_X2 U22336 ( .A1(n20113), .A2(n20244), .ZN(n20148) );
  NOR2_X2 U22337 ( .A1(n11770), .A2(n20154), .ZN(n20146) );
  AOI22_X1 U22338 ( .A1(n20249), .A2(n20148), .B1(n20248), .B2(n20146), .ZN(
        n20115) );
  AOI22_X1 U22339 ( .A1(n20252), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n20147), .B2(n20196), .ZN(n20114) );
  OAI211_X1 U22340 ( .C1(n20145), .C2(n20199), .A(n20115), .B(n20114), .ZN(
        P2_U3171) );
  AOI22_X1 U22341 ( .A1(n20149), .A2(n20196), .B1(n20255), .B2(n20146), .ZN(
        n20117) );
  AOI22_X1 U22342 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20258), .B1(
        n20148), .B2(n20257), .ZN(n20116) );
  OAI211_X1 U22343 ( .C1(n20138), .C2(n20267), .A(n20117), .B(n20116), .ZN(
        P2_U3163) );
  AOI22_X1 U22344 ( .A1(n20263), .A2(n20148), .B1(n20146), .B2(n20262), .ZN(
        n20119) );
  AOI22_X1 U22345 ( .A1(n20264), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n20270), .B2(n20147), .ZN(n20118) );
  OAI211_X1 U22346 ( .C1(n20145), .C2(n20267), .A(n20119), .B(n20118), .ZN(
        P2_U3155) );
  AOI22_X1 U22347 ( .A1(n20269), .A2(n20148), .B1(n20146), .B2(n20268), .ZN(
        n20121) );
  AOI22_X1 U22348 ( .A1(n20271), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n20270), .B2(n20149), .ZN(n20120) );
  OAI211_X1 U22349 ( .C1(n20138), .C2(n20274), .A(n20121), .B(n20120), .ZN(
        P2_U3147) );
  AOI22_X1 U22350 ( .A1(n20276), .A2(n20148), .B1(n20146), .B2(n20275), .ZN(
        n20123) );
  AOI22_X1 U22351 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20278), .B1(
        n20277), .B2(n20149), .ZN(n20122) );
  OAI211_X1 U22352 ( .C1(n20138), .C2(n20286), .A(n20123), .B(n20122), .ZN(
        P2_U3139) );
  AOI22_X1 U22353 ( .A1(n20149), .A2(n20208), .B1(n20281), .B2(n20146), .ZN(
        n20125) );
  AOI22_X1 U22354 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20283), .B1(
        n20148), .B2(n20282), .ZN(n20124) );
  OAI211_X1 U22355 ( .C1(n20138), .C2(n20214), .A(n20125), .B(n20124), .ZN(
        P2_U3131) );
  AOI22_X1 U22356 ( .A1(n20147), .A2(n20211), .B1(n20146), .B2(n20287), .ZN(
        n20127) );
  AOI22_X1 U22357 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20290), .B1(
        n20148), .B2(n20289), .ZN(n20126) );
  OAI211_X1 U22358 ( .C1(n20145), .C2(n20214), .A(n20127), .B(n20126), .ZN(
        P2_U3123) );
  AOI22_X1 U22359 ( .A1(n20149), .A2(n20211), .B1(n20146), .B2(n20293), .ZN(
        n20129) );
  AOI22_X1 U22360 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20295), .B1(
        n20148), .B2(n20294), .ZN(n20128) );
  OAI211_X1 U22361 ( .C1(n20138), .C2(n20219), .A(n20129), .B(n20128), .ZN(
        P2_U3115) );
  AOI22_X1 U22362 ( .A1(n20300), .A2(n20148), .B1(n20299), .B2(n20146), .ZN(
        n20131) );
  AOI22_X1 U22363 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20302), .B1(
        n20220), .B2(n20147), .ZN(n20130) );
  OAI211_X1 U22364 ( .C1(n20145), .C2(n20219), .A(n20131), .B(n20130), .ZN(
        P2_U3107) );
  AOI22_X1 U22365 ( .A1(n20306), .A2(n20148), .B1(n20146), .B2(n20305), .ZN(
        n20133) );
  AOI22_X1 U22366 ( .A1(n20149), .A2(n20220), .B1(
        P2_INSTQUEUE_REG_6__3__SCAN_IN), .B2(n20307), .ZN(n20132) );
  OAI211_X1 U22367 ( .C1(n20138), .C2(n20317), .A(n20133), .B(n20132), .ZN(
        P2_U3099) );
  AOI22_X1 U22368 ( .A1(n20147), .A2(n20319), .B1(n20146), .B2(n20312), .ZN(
        n20135) );
  AOI22_X1 U22369 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20314), .B1(
        n20148), .B2(n20313), .ZN(n20134) );
  OAI211_X1 U22370 ( .C1(n20145), .C2(n20317), .A(n20135), .B(n20134), .ZN(
        P2_U3091) );
  AOI22_X1 U22371 ( .A1(n20149), .A2(n20319), .B1(n20146), .B2(n20318), .ZN(
        n20137) );
  AOI22_X1 U22372 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20321), .B1(
        n20148), .B2(n20320), .ZN(n20136) );
  OAI211_X1 U22373 ( .C1(n20138), .C2(n20324), .A(n20137), .B(n20136), .ZN(
        P2_U3083) );
  AOI22_X1 U22374 ( .A1(n20147), .A2(n20228), .B1(n20325), .B2(n20146), .ZN(
        n20140) );
  AOI22_X1 U22375 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20328), .B1(
        n20148), .B2(n20327), .ZN(n20139) );
  OAI211_X1 U22376 ( .C1(n20145), .C2(n20324), .A(n20140), .B(n20139), .ZN(
        P2_U3075) );
  AOI22_X1 U22377 ( .A1(n20332), .A2(n20148), .B1(n20146), .B2(n20331), .ZN(
        n20142) );
  AOI22_X1 U22378 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20333), .B1(
        n20340), .B2(n20147), .ZN(n20141) );
  OAI211_X1 U22379 ( .C1(n20145), .C2(n20336), .A(n20142), .B(n20141), .ZN(
        P2_U3067) );
  AOI22_X1 U22380 ( .A1(n20339), .A2(n20148), .B1(n20146), .B2(n20338), .ZN(
        n20144) );
  AOI22_X1 U22381 ( .A1(n20341), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n20353), .B2(n20147), .ZN(n20143) );
  OAI211_X1 U22382 ( .C1(n20145), .C2(n20235), .A(n20144), .B(n20143), .ZN(
        P2_U3059) );
  AOI22_X1 U22383 ( .A1(n20147), .A2(n20348), .B1(n20346), .B2(n20146), .ZN(
        n20151) );
  AOI22_X1 U22384 ( .A1(n20353), .A2(n20149), .B1(n20351), .B2(n20148), .ZN(
        n20150) );
  OAI211_X1 U22385 ( .C1(n20357), .C2(n20152), .A(n20151), .B(n20150), .ZN(
        P2_U3051) );
  NOR2_X2 U22386 ( .A1(n20153), .A2(n20244), .ZN(n20190) );
  NOR2_X2 U22387 ( .A1(n20155), .A2(n20154), .ZN(n20188) );
  AOI22_X1 U22388 ( .A1(n20249), .A2(n20190), .B1(n20248), .B2(n20188), .ZN(
        n20157) );
  AOI22_X1 U22389 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20252), .B1(
        n20191), .B2(n20196), .ZN(n20156) );
  OAI211_X1 U22390 ( .C1(n20184), .C2(n20199), .A(n20157), .B(n20156), .ZN(
        P2_U3170) );
  AOI22_X1 U22391 ( .A1(n20256), .A2(n20191), .B1(n20255), .B2(n20188), .ZN(
        n20159) );
  AOI22_X1 U22392 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20258), .B1(
        n20190), .B2(n20257), .ZN(n20158) );
  OAI211_X1 U22393 ( .C1(n20184), .C2(n20261), .A(n20159), .B(n20158), .ZN(
        P2_U3162) );
  AOI22_X1 U22394 ( .A1(n20263), .A2(n20190), .B1(n20188), .B2(n20262), .ZN(
        n20161) );
  AOI22_X1 U22395 ( .A1(n20264), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n20270), .B2(n20191), .ZN(n20160) );
  OAI211_X1 U22396 ( .C1(n20184), .C2(n20267), .A(n20161), .B(n20160), .ZN(
        P2_U3154) );
  AOI22_X1 U22397 ( .A1(n20269), .A2(n20190), .B1(n20188), .B2(n20268), .ZN(
        n20163) );
  AOI22_X1 U22398 ( .A1(n20271), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n20270), .B2(n20189), .ZN(n20162) );
  OAI211_X1 U22399 ( .C1(n20187), .C2(n20274), .A(n20163), .B(n20162), .ZN(
        P2_U3146) );
  AOI22_X1 U22400 ( .A1(n20276), .A2(n20190), .B1(n20188), .B2(n20275), .ZN(
        n20165) );
  AOI22_X1 U22401 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20278), .B1(
        n20277), .B2(n20189), .ZN(n20164) );
  OAI211_X1 U22402 ( .C1(n20187), .C2(n20286), .A(n20165), .B(n20164), .ZN(
        P2_U3138) );
  AOI22_X1 U22403 ( .A1(n20191), .A2(n20288), .B1(n20188), .B2(n20281), .ZN(
        n20167) );
  AOI22_X1 U22404 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20283), .B1(
        n20190), .B2(n20282), .ZN(n20166) );
  OAI211_X1 U22405 ( .C1(n20184), .C2(n20286), .A(n20167), .B(n20166), .ZN(
        P2_U3130) );
  AOI22_X1 U22406 ( .A1(n20189), .A2(n20288), .B1(n20188), .B2(n20287), .ZN(
        n20169) );
  AOI22_X1 U22407 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20290), .B1(
        n20190), .B2(n20289), .ZN(n20168) );
  OAI211_X1 U22408 ( .C1(n20187), .C2(n20298), .A(n20169), .B(n20168), .ZN(
        P2_U3122) );
  AOI22_X1 U22409 ( .A1(n20191), .A2(n20301), .B1(n20188), .B2(n20293), .ZN(
        n20171) );
  AOI22_X1 U22410 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20295), .B1(
        n20190), .B2(n20294), .ZN(n20170) );
  OAI211_X1 U22411 ( .C1(n20184), .C2(n20298), .A(n20171), .B(n20170), .ZN(
        P2_U3114) );
  AOI22_X1 U22412 ( .A1(n20300), .A2(n20190), .B1(n20299), .B2(n20188), .ZN(
        n20173) );
  AOI22_X1 U22413 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20302), .B1(
        n20301), .B2(n20189), .ZN(n20172) );
  OAI211_X1 U22414 ( .C1(n20187), .C2(n20311), .A(n20173), .B(n20172), .ZN(
        P2_U3106) );
  AOI22_X1 U22415 ( .A1(n20306), .A2(n20190), .B1(n20188), .B2(n20305), .ZN(
        n20175) );
  AOI22_X1 U22416 ( .A1(n20189), .A2(n20220), .B1(
        P2_INSTQUEUE_REG_6__2__SCAN_IN), .B2(n20307), .ZN(n20174) );
  OAI211_X1 U22417 ( .C1(n20187), .C2(n20317), .A(n20175), .B(n20174), .ZN(
        P2_U3098) );
  AOI22_X1 U22418 ( .A1(n20191), .A2(n20319), .B1(n20188), .B2(n20312), .ZN(
        n20177) );
  AOI22_X1 U22419 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20314), .B1(
        n20190), .B2(n20313), .ZN(n20176) );
  OAI211_X1 U22420 ( .C1(n20184), .C2(n20317), .A(n20177), .B(n20176), .ZN(
        P2_U3090) );
  AOI22_X1 U22421 ( .A1(n20189), .A2(n20319), .B1(n20188), .B2(n20318), .ZN(
        n20179) );
  AOI22_X1 U22422 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20321), .B1(
        n20190), .B2(n20320), .ZN(n20178) );
  OAI211_X1 U22423 ( .C1(n20187), .C2(n20324), .A(n20179), .B(n20178), .ZN(
        P2_U3082) );
  AOI22_X1 U22424 ( .A1(n20189), .A2(n20326), .B1(n20188), .B2(n20325), .ZN(
        n20181) );
  AOI22_X1 U22425 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20328), .B1(
        n20190), .B2(n20327), .ZN(n20180) );
  OAI211_X1 U22426 ( .C1(n20187), .C2(n20336), .A(n20181), .B(n20180), .ZN(
        P2_U3074) );
  AOI22_X1 U22427 ( .A1(n20332), .A2(n20190), .B1(n20188), .B2(n20331), .ZN(
        n20183) );
  AOI22_X1 U22428 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20333), .B1(
        n20340), .B2(n20191), .ZN(n20182) );
  OAI211_X1 U22429 ( .C1(n20184), .C2(n20336), .A(n20183), .B(n20182), .ZN(
        P2_U3066) );
  AOI22_X1 U22430 ( .A1(n20339), .A2(n20190), .B1(n20188), .B2(n20338), .ZN(
        n20186) );
  AOI22_X1 U22431 ( .A1(n20341), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n20189), .B2(n20340), .ZN(n20185) );
  OAI211_X1 U22432 ( .C1(n20187), .C2(n20344), .A(n20186), .B(n20185), .ZN(
        P2_U3058) );
  AOI22_X1 U22433 ( .A1(n20189), .A2(n20353), .B1(n20188), .B2(n20346), .ZN(
        n20193) );
  AOI22_X1 U22434 ( .A1(n20348), .A2(n20191), .B1(n20351), .B2(n20190), .ZN(
        n20192) );
  OAI211_X1 U22435 ( .C1(n20357), .C2(n20194), .A(n20193), .B(n20192), .ZN(
        P2_U3050) );
  AOI22_X2 U22436 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20251), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n20250), .ZN(n20236) );
  NOR2_X2 U22437 ( .A1(n20195), .A2(n20244), .ZN(n20239) );
  AOI22_X1 U22438 ( .A1(n20249), .A2(n20239), .B1(n20248), .B2(n20237), .ZN(
        n20198) );
  AOI22_X1 U22439 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20251), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n20250), .ZN(n20227) );
  AOI22_X1 U22440 ( .A1(n20252), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n20196), .B2(n20238), .ZN(n20197) );
  OAI211_X1 U22441 ( .C1(n20236), .C2(n20199), .A(n20198), .B(n20197), .ZN(
        P2_U3169) );
  AOI22_X1 U22442 ( .A1(n20256), .A2(n20238), .B1(n20255), .B2(n20237), .ZN(
        n20201) );
  AOI22_X1 U22443 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20258), .B1(
        n20239), .B2(n20257), .ZN(n20200) );
  OAI211_X1 U22444 ( .C1(n20236), .C2(n20261), .A(n20201), .B(n20200), .ZN(
        P2_U3161) );
  AOI22_X1 U22445 ( .A1(n20263), .A2(n20239), .B1(n20237), .B2(n20262), .ZN(
        n20203) );
  AOI22_X1 U22446 ( .A1(n20264), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n20270), .B2(n20238), .ZN(n20202) );
  OAI211_X1 U22447 ( .C1(n20236), .C2(n20267), .A(n20203), .B(n20202), .ZN(
        P2_U3153) );
  AOI22_X1 U22448 ( .A1(n20269), .A2(n20239), .B1(n20237), .B2(n20268), .ZN(
        n20205) );
  INV_X1 U22449 ( .A(n20236), .ZN(n20240) );
  AOI22_X1 U22450 ( .A1(n20271), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n20270), .B2(n20240), .ZN(n20204) );
  OAI211_X1 U22451 ( .C1(n20227), .C2(n20274), .A(n20205), .B(n20204), .ZN(
        P2_U3145) );
  AOI22_X1 U22452 ( .A1(n20276), .A2(n20239), .B1(n20237), .B2(n20275), .ZN(
        n20207) );
  AOI22_X1 U22453 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20278), .B1(
        n20208), .B2(n20238), .ZN(n20206) );
  OAI211_X1 U22454 ( .C1(n20236), .C2(n20274), .A(n20207), .B(n20206), .ZN(
        P2_U3137) );
  AOI22_X1 U22455 ( .A1(n20240), .A2(n20208), .B1(n20237), .B2(n20281), .ZN(
        n20210) );
  AOI22_X1 U22456 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20283), .B1(
        n20239), .B2(n20282), .ZN(n20209) );
  OAI211_X1 U22457 ( .C1(n20227), .C2(n20214), .A(n20210), .B(n20209), .ZN(
        P2_U3129) );
  AOI22_X1 U22458 ( .A1(n20238), .A2(n20211), .B1(n20237), .B2(n20287), .ZN(
        n20213) );
  AOI22_X1 U22459 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20290), .B1(
        n20239), .B2(n20289), .ZN(n20212) );
  OAI211_X1 U22460 ( .C1(n20236), .C2(n20214), .A(n20213), .B(n20212), .ZN(
        P2_U3121) );
  AOI22_X1 U22461 ( .A1(n20238), .A2(n20301), .B1(n20237), .B2(n20293), .ZN(
        n20216) );
  AOI22_X1 U22462 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20295), .B1(
        n20239), .B2(n20294), .ZN(n20215) );
  OAI211_X1 U22463 ( .C1(n20236), .C2(n20298), .A(n20216), .B(n20215), .ZN(
        P2_U3113) );
  AOI22_X1 U22464 ( .A1(n20300), .A2(n20239), .B1(n20299), .B2(n20237), .ZN(
        n20218) );
  AOI22_X1 U22465 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20302), .B1(
        n20220), .B2(n20238), .ZN(n20217) );
  OAI211_X1 U22466 ( .C1(n20236), .C2(n20219), .A(n20218), .B(n20217), .ZN(
        P2_U3105) );
  AOI22_X1 U22467 ( .A1(n20306), .A2(n20239), .B1(n20237), .B2(n20305), .ZN(
        n20222) );
  AOI22_X1 U22468 ( .A1(n20240), .A2(n20220), .B1(
        P2_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n20307), .ZN(n20221) );
  OAI211_X1 U22469 ( .C1(n20227), .C2(n20317), .A(n20222), .B(n20221), .ZN(
        P2_U3097) );
  AOI22_X1 U22470 ( .A1(n20238), .A2(n20319), .B1(n20237), .B2(n20312), .ZN(
        n20224) );
  AOI22_X1 U22471 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20314), .B1(
        n20239), .B2(n20313), .ZN(n20223) );
  OAI211_X1 U22472 ( .C1(n20236), .C2(n20317), .A(n20224), .B(n20223), .ZN(
        P2_U3089) );
  AOI22_X1 U22473 ( .A1(n20240), .A2(n20319), .B1(n20237), .B2(n20318), .ZN(
        n20226) );
  AOI22_X1 U22474 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20321), .B1(
        n20239), .B2(n20320), .ZN(n20225) );
  OAI211_X1 U22475 ( .C1(n20227), .C2(n20324), .A(n20226), .B(n20225), .ZN(
        P2_U3081) );
  AOI22_X1 U22476 ( .A1(n20238), .A2(n20228), .B1(n20237), .B2(n20325), .ZN(
        n20230) );
  AOI22_X1 U22477 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20328), .B1(
        n20239), .B2(n20327), .ZN(n20229) );
  OAI211_X1 U22478 ( .C1(n20236), .C2(n20324), .A(n20230), .B(n20229), .ZN(
        P2_U3073) );
  AOI22_X1 U22479 ( .A1(n20332), .A2(n20239), .B1(n20237), .B2(n20331), .ZN(
        n20232) );
  AOI22_X1 U22480 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20333), .B1(
        n20340), .B2(n20238), .ZN(n20231) );
  OAI211_X1 U22481 ( .C1(n20236), .C2(n20336), .A(n20232), .B(n20231), .ZN(
        P2_U3065) );
  AOI22_X1 U22482 ( .A1(n20339), .A2(n20239), .B1(n20237), .B2(n20338), .ZN(
        n20234) );
  AOI22_X1 U22483 ( .A1(n20341), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n20353), .B2(n20238), .ZN(n20233) );
  OAI211_X1 U22484 ( .C1(n20236), .C2(n20235), .A(n20234), .B(n20233), .ZN(
        P2_U3057) );
  AOI22_X1 U22485 ( .A1(n20238), .A2(n20348), .B1(n20237), .B2(n20346), .ZN(
        n20242) );
  AOI22_X1 U22486 ( .A1(n20353), .A2(n20240), .B1(n20351), .B2(n20239), .ZN(
        n20241) );
  OAI211_X1 U22487 ( .C1(n20357), .C2(n20243), .A(n20242), .B(n20241), .ZN(
        P2_U3049) );
  NOR2_X2 U22488 ( .A1(n20245), .A2(n20244), .ZN(n20350) );
  AOI22_X1 U22489 ( .A1(n20249), .A2(n20350), .B1(n20248), .B2(n20347), .ZN(
        n20254) );
  AOI22_X1 U22490 ( .A1(n20252), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n20352), .B2(n20348), .ZN(n20253) );
  OAI211_X1 U22491 ( .C1(n20345), .C2(n20261), .A(n20254), .B(n20253), .ZN(
        P2_U3168) );
  AOI22_X1 U22492 ( .A1(n20256), .A2(n20349), .B1(n20255), .B2(n20347), .ZN(
        n20260) );
  AOI22_X1 U22493 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20258), .B1(
        n20350), .B2(n20257), .ZN(n20259) );
  OAI211_X1 U22494 ( .C1(n20337), .C2(n20261), .A(n20260), .B(n20259), .ZN(
        P2_U3160) );
  AOI22_X1 U22495 ( .A1(n20263), .A2(n20350), .B1(n20347), .B2(n20262), .ZN(
        n20266) );
  AOI22_X1 U22496 ( .A1(n20264), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n20270), .B2(n20349), .ZN(n20265) );
  OAI211_X1 U22497 ( .C1(n20337), .C2(n20267), .A(n20266), .B(n20265), .ZN(
        P2_U3152) );
  AOI22_X1 U22498 ( .A1(n20269), .A2(n20350), .B1(n20347), .B2(n20268), .ZN(
        n20273) );
  AOI22_X1 U22499 ( .A1(n20271), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n20270), .B2(n20352), .ZN(n20272) );
  OAI211_X1 U22500 ( .C1(n20345), .C2(n20274), .A(n20273), .B(n20272), .ZN(
        P2_U3144) );
  AOI22_X1 U22501 ( .A1(n20276), .A2(n20350), .B1(n20347), .B2(n20275), .ZN(
        n20280) );
  AOI22_X1 U22502 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20278), .B1(
        n20277), .B2(n20352), .ZN(n20279) );
  OAI211_X1 U22503 ( .C1(n20345), .C2(n20286), .A(n20280), .B(n20279), .ZN(
        P2_U3136) );
  AOI22_X1 U22504 ( .A1(n20349), .A2(n20288), .B1(n20347), .B2(n20281), .ZN(
        n20285) );
  AOI22_X1 U22505 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20283), .B1(
        n20350), .B2(n20282), .ZN(n20284) );
  OAI211_X1 U22506 ( .C1(n20337), .C2(n20286), .A(n20285), .B(n20284), .ZN(
        P2_U3128) );
  AOI22_X1 U22507 ( .A1(n20352), .A2(n20288), .B1(n20347), .B2(n20287), .ZN(
        n20292) );
  AOI22_X1 U22508 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20290), .B1(
        n20350), .B2(n20289), .ZN(n20291) );
  OAI211_X1 U22509 ( .C1(n20345), .C2(n20298), .A(n20292), .B(n20291), .ZN(
        P2_U3120) );
  AOI22_X1 U22510 ( .A1(n20349), .A2(n20301), .B1(n20347), .B2(n20293), .ZN(
        n20297) );
  AOI22_X1 U22511 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20295), .B1(
        n20350), .B2(n20294), .ZN(n20296) );
  OAI211_X1 U22512 ( .C1(n20337), .C2(n20298), .A(n20297), .B(n20296), .ZN(
        P2_U3112) );
  AOI22_X1 U22513 ( .A1(n20300), .A2(n20350), .B1(n20299), .B2(n20347), .ZN(
        n20304) );
  AOI22_X1 U22514 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20302), .B1(
        n20301), .B2(n20352), .ZN(n20303) );
  OAI211_X1 U22515 ( .C1(n20345), .C2(n20311), .A(n20304), .B(n20303), .ZN(
        P2_U3104) );
  AOI22_X1 U22516 ( .A1(n20306), .A2(n20350), .B1(n20347), .B2(n20305), .ZN(
        n20310) );
  AOI22_X1 U22517 ( .A1(n20349), .A2(n20308), .B1(
        P2_INSTQUEUE_REG_6__0__SCAN_IN), .B2(n20307), .ZN(n20309) );
  OAI211_X1 U22518 ( .C1(n20337), .C2(n20311), .A(n20310), .B(n20309), .ZN(
        P2_U3096) );
  AOI22_X1 U22519 ( .A1(n20349), .A2(n20319), .B1(n20347), .B2(n20312), .ZN(
        n20316) );
  AOI22_X1 U22520 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20314), .B1(
        n20350), .B2(n20313), .ZN(n20315) );
  OAI211_X1 U22521 ( .C1(n20337), .C2(n20317), .A(n20316), .B(n20315), .ZN(
        P2_U3088) );
  AOI22_X1 U22522 ( .A1(n20352), .A2(n20319), .B1(n20347), .B2(n20318), .ZN(
        n20323) );
  AOI22_X1 U22523 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20321), .B1(
        n20350), .B2(n20320), .ZN(n20322) );
  OAI211_X1 U22524 ( .C1(n20345), .C2(n20324), .A(n20323), .B(n20322), .ZN(
        P2_U3080) );
  AOI22_X1 U22525 ( .A1(n20352), .A2(n20326), .B1(n20347), .B2(n20325), .ZN(
        n20330) );
  AOI22_X1 U22526 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20328), .B1(
        n20350), .B2(n20327), .ZN(n20329) );
  OAI211_X1 U22527 ( .C1(n20345), .C2(n20336), .A(n20330), .B(n20329), .ZN(
        P2_U3072) );
  AOI22_X1 U22528 ( .A1(n20332), .A2(n20350), .B1(n20347), .B2(n20331), .ZN(
        n20335) );
  AOI22_X1 U22529 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20333), .B1(
        n20340), .B2(n20349), .ZN(n20334) );
  OAI211_X1 U22530 ( .C1(n20337), .C2(n20336), .A(n20335), .B(n20334), .ZN(
        P2_U3064) );
  AOI22_X1 U22531 ( .A1(n20339), .A2(n20350), .B1(n20347), .B2(n20338), .ZN(
        n20343) );
  AOI22_X1 U22532 ( .A1(n20341), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n20352), .B2(n20340), .ZN(n20342) );
  OAI211_X1 U22533 ( .C1(n20345), .C2(n20344), .A(n20343), .B(n20342), .ZN(
        P2_U3056) );
  AOI22_X1 U22534 ( .A1(n20349), .A2(n20348), .B1(n20347), .B2(n20346), .ZN(
        n20355) );
  AOI22_X1 U22535 ( .A1(n20353), .A2(n20352), .B1(n20351), .B2(n20350), .ZN(
        n20354) );
  OAI211_X1 U22536 ( .C1(n20357), .C2(n20356), .A(n20355), .B(n20354), .ZN(
        P2_U3048) );
  INV_X1 U22537 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n20668) );
  INV_X1 U22538 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n20358) );
  AOI222_X1 U22539 ( .A1(n20666), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n20668), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .C1(n20358), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n20359) );
  AOI22_X1 U22540 ( .A1(n20413), .A2(n20361), .B1(n20360), .B2(n20410), .ZN(
        U376) );
  INV_X2 U22541 ( .A(n20410), .ZN(n20413) );
  AOI22_X1 U22542 ( .A1(n20413), .A2(n20363), .B1(n20362), .B2(n20410), .ZN(
        U365) );
  AOI22_X1 U22543 ( .A1(n20413), .A2(n20365), .B1(n20364), .B2(n20410), .ZN(
        U354) );
  AOI22_X1 U22544 ( .A1(n20413), .A2(n20367), .B1(n20366), .B2(n20410), .ZN(
        U353) );
  AOI22_X1 U22545 ( .A1(n20413), .A2(n20369), .B1(n20368), .B2(n20410), .ZN(
        U352) );
  AOI22_X1 U22546 ( .A1(n20413), .A2(n20371), .B1(n20370), .B2(n20410), .ZN(
        U351) );
  OAI22_X1 U22547 ( .A1(n20410), .A2(P3_ADDRESS_REG_6__SCAN_IN), .B1(
        P2_ADDRESS_REG_6__SCAN_IN), .B2(n20359), .ZN(n20372) );
  INV_X1 U22548 ( .A(n20372), .ZN(U350) );
  OAI22_X1 U22549 ( .A1(n20410), .A2(P3_ADDRESS_REG_7__SCAN_IN), .B1(
        P2_ADDRESS_REG_7__SCAN_IN), .B2(n20413), .ZN(n20373) );
  INV_X1 U22550 ( .A(n20373), .ZN(U349) );
  OAI22_X1 U22551 ( .A1(n20410), .A2(P3_ADDRESS_REG_8__SCAN_IN), .B1(
        P2_ADDRESS_REG_8__SCAN_IN), .B2(n20413), .ZN(n20374) );
  INV_X1 U22552 ( .A(n20374), .ZN(U348) );
  OAI22_X1 U22553 ( .A1(n20410), .A2(P3_ADDRESS_REG_9__SCAN_IN), .B1(
        P2_ADDRESS_REG_9__SCAN_IN), .B2(n20413), .ZN(n20375) );
  INV_X1 U22554 ( .A(n20375), .ZN(U347) );
  AOI22_X1 U22555 ( .A1(n20413), .A2(n20377), .B1(n20376), .B2(n20410), .ZN(
        U375) );
  AOI22_X1 U22556 ( .A1(n20413), .A2(n20379), .B1(n20378), .B2(n20410), .ZN(
        U374) );
  AOI22_X1 U22557 ( .A1(n20413), .A2(n20381), .B1(n20380), .B2(n20410), .ZN(
        U373) );
  AOI22_X1 U22558 ( .A1(n20413), .A2(n20383), .B1(n20382), .B2(n20410), .ZN(
        U372) );
  AOI22_X1 U22559 ( .A1(n20413), .A2(n20385), .B1(n20384), .B2(n20410), .ZN(
        U371) );
  AOI22_X1 U22560 ( .A1(n20413), .A2(n20387), .B1(n20386), .B2(n20410), .ZN(
        U370) );
  OAI22_X1 U22561 ( .A1(n20410), .A2(P3_ADDRESS_REG_16__SCAN_IN), .B1(
        P2_ADDRESS_REG_16__SCAN_IN), .B2(n20413), .ZN(n20388) );
  INV_X1 U22562 ( .A(n20388), .ZN(U369) );
  OAI22_X1 U22563 ( .A1(n20410), .A2(P3_ADDRESS_REG_17__SCAN_IN), .B1(
        P2_ADDRESS_REG_17__SCAN_IN), .B2(n20359), .ZN(n20389) );
  INV_X1 U22564 ( .A(n20389), .ZN(U368) );
  AOI22_X1 U22565 ( .A1(n20413), .A2(n20391), .B1(n20390), .B2(n20410), .ZN(
        U367) );
  AOI22_X1 U22566 ( .A1(n20413), .A2(n20393), .B1(n20392), .B2(n20410), .ZN(
        U366) );
  AOI22_X1 U22567 ( .A1(n20413), .A2(n20395), .B1(n20394), .B2(n20410), .ZN(
        U364) );
  AOI22_X1 U22568 ( .A1(n20413), .A2(n20397), .B1(n20396), .B2(n20410), .ZN(
        U363) );
  AOI22_X1 U22569 ( .A1(n20413), .A2(n20399), .B1(n20398), .B2(n20410), .ZN(
        U362) );
  AOI22_X1 U22570 ( .A1(n20413), .A2(n20401), .B1(n20400), .B2(n20410), .ZN(
        U361) );
  OAI22_X1 U22571 ( .A1(n20410), .A2(P3_ADDRESS_REG_24__SCAN_IN), .B1(
        P2_ADDRESS_REG_24__SCAN_IN), .B2(n20359), .ZN(n20402) );
  INV_X1 U22572 ( .A(n20402), .ZN(U360) );
  OAI22_X1 U22573 ( .A1(n20410), .A2(P3_ADDRESS_REG_25__SCAN_IN), .B1(
        P2_ADDRESS_REG_25__SCAN_IN), .B2(n20359), .ZN(n20403) );
  INV_X1 U22574 ( .A(n20403), .ZN(U359) );
  AOI22_X1 U22575 ( .A1(n20413), .A2(n20405), .B1(n20404), .B2(n20410), .ZN(
        U358) );
  AOI22_X1 U22576 ( .A1(n20413), .A2(n20407), .B1(n20406), .B2(n20410), .ZN(
        U357) );
  AOI22_X1 U22577 ( .A1(n20413), .A2(n20409), .B1(n20408), .B2(n20410), .ZN(
        U356) );
  AOI22_X1 U22578 ( .A1(n20413), .A2(n20412), .B1(n20411), .B2(n20410), .ZN(
        U355) );
  AOI22_X1 U22579 ( .A1(n21877), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n20429), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20415) );
  OAI21_X1 U22580 ( .B1(n20416), .B2(n20437), .A(n20415), .ZN(P1_U2936) );
  AOI22_X1 U22581 ( .A1(n20425), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n20429), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20417) );
  OAI21_X1 U22582 ( .B1(n13333), .B2(n20437), .A(n20417), .ZN(P1_U2935) );
  AOI22_X1 U22583 ( .A1(n20425), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n20429), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20418) );
  OAI21_X1 U22584 ( .B1(n13327), .B2(n20437), .A(n20418), .ZN(P1_U2934) );
  AOI22_X1 U22585 ( .A1(n20425), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n20429), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20419) );
  OAI21_X1 U22586 ( .B1(n13322), .B2(n20437), .A(n20419), .ZN(P1_U2933) );
  AOI22_X1 U22587 ( .A1(n20425), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n20429), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20420) );
  OAI21_X1 U22588 ( .B1(n20421), .B2(n20437), .A(n20420), .ZN(P1_U2932) );
  AOI22_X1 U22589 ( .A1(n20425), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n20429), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20422) );
  OAI21_X1 U22590 ( .B1(n15426), .B2(n20437), .A(n20422), .ZN(P1_U2931) );
  AOI22_X1 U22591 ( .A1(n20425), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n20429), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20423) );
  OAI21_X1 U22592 ( .B1(n13370), .B2(n20437), .A(n20423), .ZN(P1_U2930) );
  AOI22_X1 U22593 ( .A1(n21877), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n20429), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20424) );
  OAI21_X1 U22594 ( .B1(n13316), .B2(n20437), .A(n20424), .ZN(P1_U2929) );
  AOI22_X1 U22595 ( .A1(n20425), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n20429), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20426) );
  OAI21_X1 U22596 ( .B1(n20427), .B2(n20437), .A(n20426), .ZN(P1_U2928) );
  AOI22_X1 U22597 ( .A1(n21877), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n20429), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20428) );
  OAI21_X1 U22598 ( .B1(n15902), .B2(n20437), .A(n20428), .ZN(P1_U2927) );
  AOI22_X1 U22599 ( .A1(n21877), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n20429), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20430) );
  OAI21_X1 U22600 ( .B1(n15904), .B2(n20437), .A(n20430), .ZN(P1_U2926) );
  AOI22_X1 U22601 ( .A1(n21877), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n20429), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20431) );
  OAI21_X1 U22602 ( .B1(n15924), .B2(n20437), .A(n20431), .ZN(P1_U2925) );
  AOI22_X1 U22603 ( .A1(n21877), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n20429), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20432) );
  OAI21_X1 U22604 ( .B1(n15932), .B2(n20437), .A(n20432), .ZN(P1_U2924) );
  AOI22_X1 U22605 ( .A1(n21877), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n20429), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20433) );
  OAI21_X1 U22606 ( .B1(n16266), .B2(n20437), .A(n20433), .ZN(P1_U2923) );
  AOI22_X1 U22607 ( .A1(n21877), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n20429), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20434) );
  OAI21_X1 U22608 ( .B1(n20435), .B2(n20437), .A(n20434), .ZN(P1_U2922) );
  AOI22_X1 U22609 ( .A1(n21877), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n20429), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20436) );
  OAI21_X1 U22610 ( .B1(n16263), .B2(n20437), .A(n20436), .ZN(P1_U2921) );
  INV_X2 U22611 ( .A(n22682), .ZN(n20472) );
  NOR2_X1 U22612 ( .A1(n20472), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20474) );
  INV_X1 U22613 ( .A(n20474), .ZN(n20466) );
  OR2_X1 U22614 ( .A1(n22312), .A2(n20472), .ZN(n20463) );
  INV_X2 U22615 ( .A(n20463), .ZN(n20469) );
  AOI222_X1 U22616 ( .A1(n20470), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n20472), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n20469), .ZN(n20438) );
  INV_X1 U22617 ( .A(n20438), .ZN(P1_U3197) );
  AOI222_X1 U22618 ( .A1(n20469), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n20472), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n20470), .ZN(n20439) );
  INV_X1 U22619 ( .A(n20439), .ZN(P1_U3198) );
  AOI222_X1 U22620 ( .A1(n20469), .A2(P1_REIP_REG_3__SCAN_IN), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n20472), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20474), .ZN(n20440) );
  INV_X1 U22621 ( .A(n20440), .ZN(P1_U3199) );
  AOI222_X1 U22622 ( .A1(n20469), .A2(P1_REIP_REG_4__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20472), .C1(P1_REIP_REG_5__SCAN_IN), 
        .C2(n20470), .ZN(n20441) );
  INV_X1 U22623 ( .A(n20441), .ZN(P1_U3200) );
  AOI222_X1 U22624 ( .A1(n20469), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20472), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n20474), .ZN(n20442) );
  INV_X1 U22625 ( .A(n20442), .ZN(P1_U3201) );
  AOI222_X1 U22626 ( .A1(n20469), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20472), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n20470), .ZN(n20443) );
  INV_X1 U22627 ( .A(n20443), .ZN(P1_U3202) );
  AOI222_X1 U22628 ( .A1(n20469), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n20472), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20470), .ZN(n20444) );
  INV_X1 U22629 ( .A(n20444), .ZN(P1_U3203) );
  AOI222_X1 U22630 ( .A1(n20469), .A2(P1_REIP_REG_8__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n20472), .C1(P1_REIP_REG_9__SCAN_IN), 
        .C2(n20470), .ZN(n20445) );
  INV_X1 U22631 ( .A(n20445), .ZN(P1_U3204) );
  AOI222_X1 U22632 ( .A1(n20469), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20472), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20470), .ZN(n20446) );
  INV_X1 U22633 ( .A(n20446), .ZN(P1_U3205) );
  AOI222_X1 U22634 ( .A1(n20469), .A2(P1_REIP_REG_10__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20472), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n20470), .ZN(n20447) );
  INV_X1 U22635 ( .A(n20447), .ZN(P1_U3206) );
  AOI222_X1 U22636 ( .A1(n20474), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20472), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n20469), .ZN(n20448) );
  INV_X1 U22637 ( .A(n20448), .ZN(P1_U3207) );
  AOI222_X1 U22638 ( .A1(n20469), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20472), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n20470), .ZN(n20449) );
  INV_X1 U22639 ( .A(n20449), .ZN(P1_U3208) );
  AOI222_X1 U22640 ( .A1(n20469), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n20472), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20470), .ZN(n20450) );
  INV_X1 U22641 ( .A(n20450), .ZN(P1_U3209) );
  AOI222_X1 U22642 ( .A1(n20469), .A2(P1_REIP_REG_14__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n20472), .C1(P1_REIP_REG_15__SCAN_IN), 
        .C2(n20470), .ZN(n20451) );
  INV_X1 U22643 ( .A(n20451), .ZN(P1_U3210) );
  AOI222_X1 U22644 ( .A1(n20474), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20472), .C1(P1_REIP_REG_15__SCAN_IN), 
        .C2(n20469), .ZN(n20452) );
  INV_X1 U22645 ( .A(n20452), .ZN(P1_U3211) );
  AOI222_X1 U22646 ( .A1(n20469), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n20472), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n20470), .ZN(n20453) );
  INV_X1 U22647 ( .A(n20453), .ZN(P1_U3212) );
  AOI222_X1 U22648 ( .A1(n20469), .A2(P1_REIP_REG_17__SCAN_IN), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n20472), .C1(P1_REIP_REG_18__SCAN_IN), 
        .C2(n20470), .ZN(n20454) );
  INV_X1 U22649 ( .A(n20454), .ZN(P1_U3213) );
  AOI222_X1 U22650 ( .A1(n20469), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n20472), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20470), .ZN(n20455) );
  INV_X1 U22651 ( .A(n20455), .ZN(P1_U3214) );
  AOI222_X1 U22652 ( .A1(n20474), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n20472), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20469), .ZN(n20456) );
  INV_X1 U22653 ( .A(n20456), .ZN(P1_U3215) );
  AOI222_X1 U22654 ( .A1(n20469), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n20472), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n20470), .ZN(n20457) );
  INV_X1 U22655 ( .A(n20457), .ZN(P1_U3216) );
  AOI222_X1 U22656 ( .A1(n20474), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20472), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n20469), .ZN(n20458) );
  INV_X1 U22657 ( .A(n20458), .ZN(P1_U3217) );
  AOI222_X1 U22658 ( .A1(n20469), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n20472), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n20470), .ZN(n20459) );
  INV_X1 U22659 ( .A(n20459), .ZN(P1_U3218) );
  AOI222_X1 U22660 ( .A1(n20474), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n20472), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n20469), .ZN(n20460) );
  INV_X1 U22661 ( .A(n20460), .ZN(P1_U3219) );
  AOI222_X1 U22662 ( .A1(n20469), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20472), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20474), .ZN(n20461) );
  INV_X1 U22663 ( .A(n20461), .ZN(P1_U3220) );
  AOI22_X1 U22664 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n20470), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20472), .ZN(n20462) );
  OAI21_X1 U22665 ( .B1(n20464), .B2(n20463), .A(n20462), .ZN(P1_U3221) );
  AOI22_X1 U22666 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n20469), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20472), .ZN(n20465) );
  OAI21_X1 U22667 ( .B1(n20467), .B2(n20466), .A(n20465), .ZN(P1_U3222) );
  AOI222_X1 U22668 ( .A1(n20474), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20472), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20469), .ZN(n20468) );
  INV_X1 U22669 ( .A(n20468), .ZN(P1_U3223) );
  AOI222_X1 U22670 ( .A1(n20470), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20472), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20469), .ZN(n20471) );
  INV_X1 U22671 ( .A(n20471), .ZN(P1_U3224) );
  AOI222_X1 U22672 ( .A1(n20469), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20472), .C1(P1_REIP_REG_30__SCAN_IN), 
        .C2(n20474), .ZN(n20473) );
  INV_X1 U22673 ( .A(n20473), .ZN(P1_U3225) );
  AOI222_X1 U22674 ( .A1(n20469), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20472), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20474), .ZN(n20475) );
  INV_X1 U22675 ( .A(n20475), .ZN(P1_U3226) );
  OAI22_X1 U22676 ( .A1(n20472), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n22682), .ZN(n20476) );
  INV_X1 U22677 ( .A(n20476), .ZN(P1_U3458) );
  AOI221_X1 U22678 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(P1_REIP_REG_1__SCAN_IN), 
        .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(P1_REIP_REG_1__SCAN_IN), .A(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20487) );
  NOR4_X1 U22679 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20480) );
  NOR4_X1 U22680 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20479) );
  NOR4_X1 U22681 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n20478) );
  NOR4_X1 U22682 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n20477) );
  NAND4_X1 U22683 ( .A1(n20480), .A2(n20479), .A3(n20478), .A4(n20477), .ZN(
        n20486) );
  NOR4_X1 U22684 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n20484) );
  AOI211_X1 U22685 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_31__SCAN_IN), .B(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n20483) );
  NOR4_X1 U22686 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n20482) );
  NOR4_X1 U22687 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n20481) );
  NAND4_X1 U22688 ( .A1(n20484), .A2(n20483), .A3(n20482), .A4(n20481), .ZN(
        n20485) );
  NOR2_X1 U22689 ( .A1(n20486), .A2(n20485), .ZN(n20500) );
  INV_X1 U22690 ( .A(n20500), .ZN(n20497) );
  MUX2_X1 U22691 ( .A(n20487), .B(P1_BYTEENABLE_REG_3__SCAN_IN), .S(n20497), 
        .Z(P1_U2808) );
  OAI22_X1 U22692 ( .A1(n20472), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n22682), .ZN(n20488) );
  INV_X1 U22693 ( .A(n20488), .ZN(P1_U3459) );
  AOI211_X1 U22694 ( .C1(P1_REIP_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_REIP_REG_1__SCAN_IN), .B(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20489) );
  AOI21_X1 U22695 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20489), .ZN(n20491) );
  AOI22_X1 U22696 ( .A1(n20500), .A2(n20491), .B1(n20490), .B2(n20497), .ZN(
        P1_U3481) );
  OAI22_X1 U22697 ( .A1(n20472), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n22682), .ZN(n20492) );
  INV_X1 U22698 ( .A(n20492), .ZN(P1_U3460) );
  NOR3_X1 U22699 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20493) );
  NOR2_X1 U22700 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(n20493), .ZN(n20495) );
  AOI22_X1 U22701 ( .A1(n20500), .A2(n20495), .B1(n20494), .B2(n20497), .ZN(
        P1_U2807) );
  OAI22_X1 U22702 ( .A1(n20472), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n22682), .ZN(n20496) );
  INV_X1 U22703 ( .A(n20496), .ZN(P1_U3461) );
  NOR2_X1 U22704 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n20499) );
  INV_X1 U22705 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20498) );
  AOI22_X1 U22706 ( .A1(n20500), .A2(n20499), .B1(n20498), .B2(n20497), .ZN(
        P1_U3482) );
  INV_X1 U22707 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n20502) );
  XNOR2_X1 U22708 ( .A(n11203), .B(n11274), .ZN(n22105) );
  AOI22_X1 U22709 ( .A1(n22112), .A2(n13916), .B1(n20528), .B2(n22105), .ZN(
        n20501) );
  OAI21_X1 U22710 ( .B1(n20524), .B2(n20502), .A(n20501), .ZN(P1_U2866) );
  INV_X1 U22711 ( .A(n20503), .ZN(n20585) );
  AOI22_X1 U22712 ( .A1(n20585), .A2(n13916), .B1(n20528), .B2(n22026), .ZN(
        n20504) );
  OAI21_X1 U22713 ( .B1(n20524), .B2(n20505), .A(n20504), .ZN(P1_U2855) );
  INV_X1 U22714 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n22160) );
  NOR2_X1 U22715 ( .A1(n20507), .A2(n20506), .ZN(n20508) );
  OR2_X1 U22716 ( .A1(n20509), .A2(n20508), .ZN(n22010) );
  OAI22_X1 U22717 ( .A1(n20569), .A2(n16189), .B1(n20510), .B2(n22010), .ZN(
        n20511) );
  INV_X1 U22718 ( .A(n20511), .ZN(n20512) );
  OAI21_X1 U22719 ( .B1(n20524), .B2(n22160), .A(n20512), .ZN(P1_U2857) );
  INV_X1 U22720 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n20515) );
  OAI22_X1 U22721 ( .A1(n22247), .A2(n16189), .B1(n22245), .B2(n20510), .ZN(
        n20513) );
  INV_X1 U22722 ( .A(n20513), .ZN(n20514) );
  OAI21_X1 U22723 ( .B1(n20524), .B2(n20515), .A(n20514), .ZN(P1_U2849) );
  NOR2_X1 U22724 ( .A1(n22214), .A2(n20510), .ZN(n20516) );
  AOI21_X1 U22725 ( .B1(n22216), .B2(n13916), .A(n20516), .ZN(n20517) );
  OAI21_X1 U22726 ( .B1(n20524), .B2(n20518), .A(n20517), .ZN(P1_U2851) );
  INV_X1 U22727 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n22194) );
  AND2_X1 U22728 ( .A1(n20520), .A2(n20519), .ZN(n20521) );
  NOR2_X1 U22729 ( .A1(n20522), .A2(n20521), .ZN(n22198) );
  AOI22_X1 U22730 ( .A1(n22200), .A2(n13916), .B1(n22198), .B2(n20528), .ZN(
        n20523) );
  OAI21_X1 U22731 ( .B1(n20524), .B2(n22194), .A(n20523), .ZN(P1_U2853) );
  INV_X1 U22732 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20530) );
  NAND2_X1 U22733 ( .A1(n20526), .A2(n20525), .ZN(n20527) );
  AND2_X1 U22734 ( .A1(n11203), .A2(n20527), .ZN(n22091) );
  AOI22_X1 U22735 ( .A1(n22100), .A2(n13916), .B1(n20528), .B2(n22091), .ZN(
        n20529) );
  OAI21_X1 U22736 ( .B1(n20524), .B2(n20530), .A(n20529), .ZN(P1_U2867) );
  AOI22_X1 U22737 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n22052), .B1(
        P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n20588), .ZN(n20537) );
  OAI21_X1 U22738 ( .B1(n20533), .B2(n20532), .A(n20531), .ZN(n20534) );
  INV_X1 U22739 ( .A(n20534), .ZN(n21928) );
  AOI22_X1 U22740 ( .A1(n21928), .A2(n20591), .B1(n20555), .B2(n20535), .ZN(
        n20536) );
  OAI211_X1 U22741 ( .C1(n20594), .C2(n22090), .A(n20537), .B(n20536), .ZN(
        P1_U2995) );
  AOI22_X1 U22742 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n22052), .B1(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n20588), .ZN(n20543) );
  OAI21_X1 U22743 ( .B1(n20540), .B2(n20539), .A(n20538), .ZN(n20541) );
  INV_X1 U22744 ( .A(n20541), .ZN(n21952) );
  AOI22_X1 U22745 ( .A1(n21952), .A2(n20591), .B1(n20555), .B2(n22100), .ZN(
        n20542) );
  OAI211_X1 U22746 ( .C1(n20594), .C2(n22103), .A(n20543), .B(n20542), .ZN(
        P1_U2994) );
  AOI22_X1 U22747 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n22052), .B1(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n20588), .ZN(n20549) );
  OAI21_X1 U22748 ( .B1(n20546), .B2(n20545), .A(n20544), .ZN(n20547) );
  INV_X1 U22749 ( .A(n20547), .ZN(n21946) );
  AOI22_X1 U22750 ( .A1(n21946), .A2(n20591), .B1(n20555), .B2(n22112), .ZN(
        n20548) );
  OAI211_X1 U22751 ( .C1(n20594), .C2(n22114), .A(n20549), .B(n20548), .ZN(
        P1_U2993) );
  AOI22_X1 U22752 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n22052), .B1(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n20588), .ZN(n20557) );
  OAI21_X1 U22753 ( .B1(n20552), .B2(n20551), .A(n20550), .ZN(n20553) );
  INV_X1 U22754 ( .A(n20553), .ZN(n21961) );
  AOI22_X1 U22755 ( .A1(n21961), .A2(n20591), .B1(n20555), .B2(n20554), .ZN(
        n20556) );
  OAI211_X1 U22756 ( .C1(n20594), .C2(n22126), .A(n20557), .B(n20556), .ZN(
        P1_U2992) );
  AOI21_X1 U22757 ( .B1(n20560), .B2(n20559), .A(n20558), .ZN(n20563) );
  INV_X1 U22758 ( .A(n20561), .ZN(n20562) );
  NOR2_X1 U22759 ( .A1(n20563), .A2(n20562), .ZN(n21995) );
  AOI22_X1 U22760 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(n22052), .B1(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n20588), .ZN(n20566) );
  INV_X1 U22761 ( .A(n22159), .ZN(n20564) );
  AOI22_X1 U22762 ( .A1(n20584), .A2(n22156), .B1(n20555), .B2(n20564), .ZN(
        n20565) );
  OAI211_X1 U22763 ( .C1(n21995), .C2(n22268), .A(n20566), .B(n20565), .ZN(
        P1_U2987) );
  XNOR2_X1 U22764 ( .A(n11452), .B(n22015), .ZN(n20567) );
  XNOR2_X1 U22765 ( .A(n20568), .B(n20567), .ZN(n22018) );
  AOI22_X1 U22766 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n22052), .B1(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n20588), .ZN(n20571) );
  INV_X1 U22767 ( .A(n20569), .ZN(n22165) );
  AOI22_X1 U22768 ( .A1(n22165), .A2(n20555), .B1(n20584), .B2(n22164), .ZN(
        n20570) );
  OAI211_X1 U22769 ( .C1(n22268), .C2(n22018), .A(n20571), .B(n20570), .ZN(
        P1_U2984) );
  INV_X1 U22770 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n20582) );
  INV_X1 U22771 ( .A(n16375), .ZN(n20575) );
  INV_X1 U22772 ( .A(n20572), .ZN(n20573) );
  AOI21_X1 U22773 ( .B1(n20575), .B2(n20574), .A(n20573), .ZN(n20577) );
  INV_X1 U22774 ( .A(n20577), .ZN(n20576) );
  INV_X1 U22775 ( .A(n22028), .ZN(n22038) );
  NOR2_X1 U22776 ( .A1(n20576), .A2(n22038), .ZN(n20580) );
  NOR2_X1 U22777 ( .A1(n20577), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n20579) );
  MUX2_X1 U22778 ( .A(n20580), .B(n20579), .S(n20578), .Z(n20581) );
  XOR2_X1 U22779 ( .A(n20582), .B(n20581), .Z(n22032) );
  AOI22_X1 U22780 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n22052), .B1(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n20588), .ZN(n20587) );
  AOI22_X1 U22781 ( .A1(n20585), .A2(n20555), .B1(n20584), .B2(n20583), .ZN(
        n20586) );
  OAI211_X1 U22782 ( .C1(n22032), .C2(n22268), .A(n20587), .B(n20586), .ZN(
        P1_U2982) );
  AOI22_X1 U22783 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n22052), .B1(
        P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n20588), .ZN(n20593) );
  XNOR2_X1 U22784 ( .A(n11452), .B(n22045), .ZN(n20589) );
  XNOR2_X1 U22785 ( .A(n20590), .B(n20589), .ZN(n22042) );
  AOI22_X1 U22786 ( .A1(n22200), .A2(n20555), .B1(n20591), .B2(n22042), .ZN(
        n20592) );
  OAI211_X1 U22787 ( .C1(n20594), .C2(n22195), .A(n20593), .B(n20592), .ZN(
        P1_U2980) );
  INV_X1 U22788 ( .A(n20595), .ZN(n20596) );
  OAI21_X1 U22789 ( .B1(n20596), .B2(n22283), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20597) );
  OAI21_X1 U22790 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20598), .A(n20597), 
        .ZN(P1_U2803) );
  OAI21_X1 U22791 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n22312), .A(n14846), 
        .ZN(n20599) );
  AOI22_X1 U22792 ( .A1(n22682), .A2(P1_CODEFETCH_REG_SCAN_IN), .B1(n20600), 
        .B2(n20599), .ZN(P1_U2804) );
  INV_X1 U22793 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n20603) );
  AOI22_X1 U22794 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(n20663), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n20662), .ZN(n20602) );
  OAI21_X1 U22795 ( .B1(n20603), .B2(n20648), .A(n20602), .ZN(U247) );
  INV_X1 U22796 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n20605) );
  AOI22_X1 U22797 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(n20663), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n20662), .ZN(n20604) );
  OAI21_X1 U22798 ( .B1(n20605), .B2(n20648), .A(n20604), .ZN(U246) );
  INV_X1 U22799 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n20607) );
  AOI22_X1 U22800 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(n20663), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n20662), .ZN(n20606) );
  OAI21_X1 U22801 ( .B1(n20607), .B2(n20648), .A(n20606), .ZN(U245) );
  INV_X1 U22802 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n20609) );
  AOI22_X1 U22803 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(n20663), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n20662), .ZN(n20608) );
  OAI21_X1 U22804 ( .B1(n20609), .B2(n20648), .A(n20608), .ZN(U244) );
  AOI22_X1 U22805 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n20663), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n20662), .ZN(n20610) );
  OAI21_X1 U22806 ( .B1(n20611), .B2(n20648), .A(n20610), .ZN(U243) );
  AOI22_X1 U22807 ( .A1(P2_DATAO_REG_5__SCAN_IN), .A2(n20663), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n20662), .ZN(n20612) );
  OAI21_X1 U22808 ( .B1(n20613), .B2(n20648), .A(n20612), .ZN(U242) );
  AOI22_X1 U22809 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(n20663), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n20662), .ZN(n20614) );
  OAI21_X1 U22810 ( .B1(n20615), .B2(n20648), .A(n20614), .ZN(U241) );
  INV_X1 U22811 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n20617) );
  AOI22_X1 U22812 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(n20663), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n20662), .ZN(n20616) );
  OAI21_X1 U22813 ( .B1(n20617), .B2(n20648), .A(n20616), .ZN(U240) );
  AOI22_X1 U22814 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(n20663), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n20662), .ZN(n20618) );
  OAI21_X1 U22815 ( .B1(n20619), .B2(n20648), .A(n20618), .ZN(U239) );
  AOI22_X1 U22816 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(n20663), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n20662), .ZN(n20620) );
  OAI21_X1 U22817 ( .B1(n14720), .B2(n20648), .A(n20620), .ZN(U238) );
  AOI22_X1 U22818 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(n20663), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n20662), .ZN(n20621) );
  OAI21_X1 U22819 ( .B1(n20622), .B2(n20648), .A(n20621), .ZN(U237) );
  INV_X1 U22820 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n20624) );
  AOI22_X1 U22821 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(n20663), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n20662), .ZN(n20623) );
  OAI21_X1 U22822 ( .B1(n20624), .B2(n20648), .A(n20623), .ZN(U236) );
  AOI22_X1 U22823 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(n20663), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n20662), .ZN(n20625) );
  OAI21_X1 U22824 ( .B1(n20626), .B2(n20648), .A(n20625), .ZN(U235) );
  INV_X1 U22825 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n20628) );
  AOI22_X1 U22826 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(n20663), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n20662), .ZN(n20627) );
  OAI21_X1 U22827 ( .B1(n20628), .B2(n20648), .A(n20627), .ZN(U234) );
  AOI22_X1 U22828 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(n20663), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n20662), .ZN(n20629) );
  OAI21_X1 U22829 ( .B1(n20630), .B2(n20648), .A(n20629), .ZN(U233) );
  AOI22_X1 U22830 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(n20663), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n20662), .ZN(n20631) );
  OAI21_X1 U22831 ( .B1(n20632), .B2(n20648), .A(n20631), .ZN(U232) );
  AOI22_X1 U22832 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n20663), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n20662), .ZN(n20633) );
  OAI21_X1 U22833 ( .B1(n20634), .B2(n20648), .A(n20633), .ZN(U231) );
  AOI22_X1 U22834 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n20663), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n20662), .ZN(n20635) );
  OAI21_X1 U22835 ( .B1(n20636), .B2(n20648), .A(n20635), .ZN(U230) );
  AOI22_X1 U22836 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n20663), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n20662), .ZN(n20637) );
  OAI21_X1 U22837 ( .B1(n20638), .B2(n20648), .A(n20637), .ZN(U229) );
  AOI22_X1 U22838 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n20663), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n20662), .ZN(n20639) );
  OAI21_X1 U22839 ( .B1(n20640), .B2(n20648), .A(n20639), .ZN(U228) );
  AOI22_X1 U22840 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n20663), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n20662), .ZN(n20641) );
  OAI21_X1 U22841 ( .B1(n20642), .B2(n20648), .A(n20641), .ZN(U227) );
  AOI22_X1 U22842 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n20663), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n20662), .ZN(n20643) );
  OAI21_X1 U22843 ( .B1(n20644), .B2(n20648), .A(n20643), .ZN(U226) );
  AOI22_X1 U22844 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n20663), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n20662), .ZN(n20645) );
  OAI21_X1 U22845 ( .B1(n20646), .B2(n20648), .A(n20645), .ZN(U225) );
  AOI22_X1 U22846 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n20663), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n20662), .ZN(n20647) );
  OAI21_X1 U22847 ( .B1(n20649), .B2(n20648), .A(n20647), .ZN(U224) );
  AOI22_X1 U22848 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n20663), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n20662), .ZN(n20650) );
  OAI21_X1 U22849 ( .B1(n20651), .B2(n20648), .A(n20650), .ZN(U223) );
  AOI22_X1 U22850 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n20663), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n20662), .ZN(n20652) );
  OAI21_X1 U22851 ( .B1(n20653), .B2(n20648), .A(n20652), .ZN(U222) );
  AOI22_X1 U22852 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n20663), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n20662), .ZN(n20654) );
  OAI21_X1 U22853 ( .B1(n20655), .B2(n20648), .A(n20654), .ZN(U221) );
  AOI22_X1 U22854 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n20663), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n20662), .ZN(n20656) );
  OAI21_X1 U22855 ( .B1(n20657), .B2(n20648), .A(n20656), .ZN(U220) );
  AOI22_X1 U22856 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n20663), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n20662), .ZN(n20658) );
  OAI21_X1 U22857 ( .B1(n20659), .B2(n20648), .A(n20658), .ZN(U219) );
  AOI22_X1 U22858 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n20663), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n20662), .ZN(n20660) );
  OAI21_X1 U22859 ( .B1(n20661), .B2(n20648), .A(n20660), .ZN(U218) );
  AOI22_X1 U22860 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n20663), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n20662), .ZN(n20664) );
  OAI21_X1 U22861 ( .B1(n20665), .B2(n20648), .A(n20664), .ZN(U217) );
  OAI222_X1 U22862 ( .A1(U214), .A2(n20668), .B1(n20648), .B2(n20667), .C1(
        U212), .C2(n20666), .ZN(U216) );
  AOI22_X1 U22863 ( .A1(n22682), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20669), 
        .B2(n20472), .ZN(P1_U3483) );
  AOI21_X1 U22864 ( .B1(n22296), .B2(n20738), .A(n20735), .ZN(n20670) );
  OAI211_X1 U22865 ( .C1(n20671), .C2(n20670), .A(n22352), .B(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n20672) );
  INV_X1 U22866 ( .A(n20672), .ZN(n20673) );
  OAI21_X1 U22867 ( .B1(n20673), .B2(n21862), .A(n21863), .ZN(n20678) );
  INV_X1 U22868 ( .A(n20674), .ZN(n20675) );
  AOI22_X1 U22869 ( .A1(n21805), .A2(n22352), .B1(n20675), .B2(n21868), .ZN(
        n20676) );
  NAND2_X1 U22870 ( .A1(n20676), .A2(n20745), .ZN(n20677) );
  MUX2_X1 U22871 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .B(n20678), .S(n20677), 
        .Z(P3_U3296) );
  AND3_X2 U22872 ( .A1(n20682), .A2(n20681), .A3(n22352), .ZN(n20732) );
  AOI22_X1 U22873 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20732), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n20728), .ZN(n20684) );
  OAI21_X1 U22874 ( .B1(n20685), .B2(n20734), .A(n20684), .ZN(P3_U2768) );
  AOI22_X1 U22875 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20732), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n20728), .ZN(n20686) );
  OAI21_X1 U22876 ( .B1(n20687), .B2(n20734), .A(n20686), .ZN(P3_U2769) );
  AOI22_X1 U22877 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20732), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n20728), .ZN(n20688) );
  OAI21_X1 U22878 ( .B1(n21255), .B2(n20734), .A(n20688), .ZN(P3_U2770) );
  AOI22_X1 U22879 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20732), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n20728), .ZN(n20689) );
  OAI21_X1 U22880 ( .B1(n21229), .B2(n20734), .A(n20689), .ZN(P3_U2771) );
  AOI22_X1 U22881 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20732), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n20728), .ZN(n20690) );
  OAI21_X1 U22882 ( .B1(n21242), .B2(n20734), .A(n20690), .ZN(P3_U2772) );
  AOI22_X1 U22883 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20732), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n20728), .ZN(n20691) );
  OAI21_X1 U22884 ( .B1(n21236), .B2(n20734), .A(n20691), .ZN(P3_U2773) );
  AOI22_X1 U22885 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20732), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n20728), .ZN(n20692) );
  OAI21_X1 U22886 ( .B1(n21265), .B2(n20734), .A(n20692), .ZN(P3_U2774) );
  AOI22_X1 U22887 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20732), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n20728), .ZN(n20693) );
  OAI21_X1 U22888 ( .B1(n20694), .B2(n20734), .A(n20693), .ZN(P3_U2775) );
  AOI22_X1 U22889 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20732), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n20728), .ZN(n20695) );
  OAI21_X1 U22890 ( .B1(n20696), .B2(n20734), .A(n20695), .ZN(P3_U2776) );
  AOI22_X1 U22891 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20732), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n20728), .ZN(n20697) );
  OAI21_X1 U22892 ( .B1(n20698), .B2(n20734), .A(n20697), .ZN(P3_U2777) );
  AOI22_X1 U22893 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20732), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n20728), .ZN(n20699) );
  OAI21_X1 U22894 ( .B1(n21274), .B2(n20734), .A(n20699), .ZN(P3_U2778) );
  AOI22_X1 U22895 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20732), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n20728), .ZN(n20700) );
  OAI21_X1 U22896 ( .B1(n20701), .B2(n20734), .A(n20700), .ZN(P3_U2779) );
  AOI22_X1 U22897 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20732), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n20728), .ZN(n20702) );
  OAI21_X1 U22898 ( .B1(n21290), .B2(n20734), .A(n20702), .ZN(P3_U2780) );
  AOI22_X1 U22899 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20732), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n20728), .ZN(n20703) );
  OAI21_X1 U22900 ( .B1(n20704), .B2(n20734), .A(n20703), .ZN(P3_U2781) );
  AOI22_X1 U22901 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20732), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n20728), .ZN(n20705) );
  OAI21_X1 U22902 ( .B1(n20706), .B2(n20734), .A(n20705), .ZN(P3_U2782) );
  AOI22_X1 U22903 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20732), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n20728), .ZN(n20707) );
  OAI21_X1 U22904 ( .B1(n21198), .B2(n20734), .A(n20707), .ZN(P3_U2783) );
  AOI22_X1 U22905 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20732), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n20728), .ZN(n20708) );
  OAI21_X1 U22906 ( .B1(n20709), .B2(n20734), .A(n20708), .ZN(P3_U2784) );
  AOI22_X1 U22907 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20732), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n20728), .ZN(n20710) );
  OAI21_X1 U22908 ( .B1(n21222), .B2(n20734), .A(n20710), .ZN(P3_U2785) );
  AOI22_X1 U22909 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20732), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n20731), .ZN(n20711) );
  OAI21_X1 U22910 ( .B1(n20712), .B2(n20734), .A(n20711), .ZN(P3_U2786) );
  AOI22_X1 U22911 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20732), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n20731), .ZN(n20713) );
  OAI21_X1 U22912 ( .B1(n21199), .B2(n20734), .A(n20713), .ZN(P3_U2787) );
  AOI22_X1 U22913 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20732), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n20731), .ZN(n20714) );
  OAI21_X1 U22914 ( .B1(n20715), .B2(n20734), .A(n20714), .ZN(P3_U2788) );
  AOI22_X1 U22915 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20732), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n20731), .ZN(n20716) );
  OAI21_X1 U22916 ( .B1(n21200), .B2(n20734), .A(n20716), .ZN(P3_U2789) );
  AOI22_X1 U22917 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20732), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n20731), .ZN(n20717) );
  OAI21_X1 U22918 ( .B1(n20718), .B2(n20734), .A(n20717), .ZN(P3_U2790) );
  AOI22_X1 U22919 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20732), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n20728), .ZN(n20719) );
  OAI21_X1 U22920 ( .B1(n21330), .B2(n20734), .A(n20719), .ZN(P3_U2791) );
  AOI22_X1 U22921 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20732), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n20731), .ZN(n20720) );
  OAI21_X1 U22922 ( .B1(n21190), .B2(n20734), .A(n20720), .ZN(P3_U2792) );
  AOI22_X1 U22923 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20732), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n20731), .ZN(n20721) );
  OAI21_X1 U22924 ( .B1(n20722), .B2(n20734), .A(n20721), .ZN(P3_U2793) );
  AOI22_X1 U22925 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20732), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n20731), .ZN(n20723) );
  OAI21_X1 U22926 ( .B1(n21179), .B2(n20734), .A(n20723), .ZN(P3_U2794) );
  AOI22_X1 U22927 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20732), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n20731), .ZN(n20724) );
  OAI21_X1 U22928 ( .B1(n20725), .B2(n20734), .A(n20724), .ZN(P3_U2795) );
  AOI22_X1 U22929 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20732), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n20731), .ZN(n20726) );
  OAI21_X1 U22930 ( .B1(n20727), .B2(n20734), .A(n20726), .ZN(P3_U2796) );
  AOI22_X1 U22931 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20732), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n20728), .ZN(n20729) );
  OAI21_X1 U22932 ( .B1(n20730), .B2(n20734), .A(n20729), .ZN(P3_U2797) );
  AOI22_X1 U22933 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n20732), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n20731), .ZN(n20733) );
  OAI21_X1 U22934 ( .B1(n21325), .B2(n20734), .A(n20733), .ZN(P3_U2798) );
  AOI211_X1 U22935 ( .C1(n20738), .C2(n20735), .A(n22341), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n20737) );
  INV_X1 U22936 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n20739) );
  INV_X1 U22937 ( .A(n20737), .ZN(n21847) );
  OAI211_X2 U22938 ( .C1(n20739), .C2(n20738), .A(n21847), .B(n20742), .ZN(
        n21132) );
  NAND2_X1 U22939 ( .A1(n22352), .A2(n22296), .ZN(n20740) );
  AOI22_X1 U22940 ( .A1(n21161), .A2(P3_EBX_REG_1__SCAN_IN), .B1(n21160), .B2(
        n20743), .ZN(n20751) );
  INV_X1 U22941 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n21156) );
  AND4_X1 U22942 ( .A1(n21862), .A2(n20744), .A3(n22296), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n20970) );
  NOR2_X1 U22943 ( .A1(n21128), .A2(n21851), .ZN(n20847) );
  INV_X1 U22944 ( .A(n20847), .ZN(n21143) );
  NOR2_X1 U22945 ( .A1(n21774), .A2(n20970), .ZN(n20746) );
  OAI211_X1 U22946 ( .C1(n21156), .C2(n21143), .A(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B(n21146), .ZN(n20749) );
  AOI21_X1 U22947 ( .B1(n20817), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n21851), .ZN(n20901) );
  NAND2_X1 U22948 ( .A1(n20747), .A2(n21360), .ZN(n21352) );
  OAI22_X1 U22949 ( .A1(n21077), .A2(n21429), .B1(n21352), .B2(n21164), .ZN(
        n20748) );
  AOI221_X1 U22950 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20749), .C1(
        n20901), .C2(n20749), .A(n20748), .ZN(n20750) );
  OAI211_X1 U22951 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(n21076), .A(n20751), .B(
        n20750), .ZN(P3_U2670) );
  AOI21_X1 U22952 ( .B1(n20755), .B2(n21429), .A(n21076), .ZN(n20752) );
  NAND2_X1 U22953 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .ZN(n20766) );
  AOI22_X1 U22954 ( .A1(n21161), .A2(P3_EBX_REG_2__SCAN_IN), .B1(n20752), .B2(
        n20766), .ZN(n20763) );
  NAND2_X1 U22955 ( .A1(n21371), .A2(n21360), .ZN(n21385) );
  AND2_X1 U22956 ( .A1(n21380), .A2(n21385), .ZN(n21366) );
  NOR3_X1 U22957 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .ZN(n20773) );
  OAI21_X1 U22958 ( .B1(n20754), .B2(n20753), .A(n21160), .ZN(n20756) );
  OAI22_X1 U22959 ( .A1(n20773), .A2(n20756), .B1(n20755), .B2(n21077), .ZN(
        n20761) );
  NOR2_X1 U22960 ( .A1(n20757), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n20887) );
  OAI22_X1 U22961 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20767), .B1(
        n20887), .B2(n20758), .ZN(n20759) );
  AOI221_X1 U22962 ( .B1(n20817), .B2(n20759), .C1(n20933), .C2(n20758), .A(
        n21851), .ZN(n20760) );
  AOI211_X1 U22963 ( .C1(n21366), .C2(n20781), .A(n20761), .B(n20760), .ZN(
        n20762) );
  OAI211_X1 U22964 ( .C1(n20764), .C2(n21146), .A(n20763), .B(n20762), .ZN(
        P3_U2669) );
  INV_X1 U22965 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n20776) );
  NOR2_X1 U22966 ( .A1(n21440), .A2(n20766), .ZN(n20792) );
  OAI21_X1 U22967 ( .B1(n21076), .B2(n20792), .A(n21077), .ZN(n20765) );
  INV_X1 U22968 ( .A(n20765), .ZN(n20791) );
  AOI221_X1 U22969 ( .B1(n21076), .B2(n21440), .C1(n20766), .C2(n21440), .A(
        n20791), .ZN(n20772) );
  AOI21_X1 U22970 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n21380), .A(
        n11175), .ZN(n21391) );
  OAI21_X1 U22971 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20767), .A(
        n20817), .ZN(n20768) );
  XNOR2_X1 U22972 ( .A(n20769), .B(n20768), .ZN(n20770) );
  OAI22_X1 U22973 ( .A1(n21391), .A2(n21164), .B1(n21851), .B2(n20770), .ZN(
        n20771) );
  AOI211_X1 U22974 ( .C1(n21127), .C2(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n20772), .B(n20771), .ZN(n20775) );
  NAND2_X1 U22975 ( .A1(n20773), .A2(n20776), .ZN(n20780) );
  OAI211_X1 U22976 ( .C1(n20773), .C2(n20776), .A(n21160), .B(n20780), .ZN(
        n20774) );
  OAI211_X1 U22977 ( .C1(n20776), .C2(n21132), .A(n20775), .B(n20774), .ZN(
        P3_U2668) );
  AOI221_X1 U22978 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20817), .C1(
        n20777), .C2(n20817), .A(n21851), .ZN(n20778) );
  AOI22_X1 U22979 ( .A1(n21161), .A2(P3_EBX_REG_4__SCAN_IN), .B1(n20779), .B2(
        n20778), .ZN(n20789) );
  NOR2_X1 U22980 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n20780), .ZN(n20799) );
  AOI211_X1 U22981 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n20780), .A(n20799), .B(
        n21135), .ZN(n20787) );
  NAND3_X1 U22982 ( .A1(n21075), .A2(n20792), .A3(n20790), .ZN(n20785) );
  OAI21_X1 U22983 ( .B1(n11147), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n20781), .ZN(n20784) );
  INV_X1 U22984 ( .A(n20887), .ZN(n20794) );
  OAI211_X1 U22985 ( .C1(n20795), .C2(n20794), .A(n20847), .B(n20782), .ZN(
        n20783) );
  NAND4_X1 U22986 ( .A1(n11142), .A2(n20785), .A3(n20784), .A4(n20783), .ZN(
        n20786) );
  AOI211_X1 U22987 ( .C1(n21127), .C2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20787), .B(n20786), .ZN(n20788) );
  OAI211_X1 U22988 ( .C1(n20791), .C2(n20790), .A(n20789), .B(n20788), .ZN(
        P3_U2667) );
  NAND2_X1 U22989 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n20792), .ZN(n20806) );
  NOR2_X1 U22990 ( .A1(n21464), .A2(n20806), .ZN(n20821) );
  OR2_X1 U22991 ( .A1(n21076), .A2(n20821), .ZN(n20805) );
  OAI21_X1 U22992 ( .B1(n20821), .B2(n21076), .A(n21077), .ZN(n20823) );
  OAI22_X1 U22993 ( .A1(n20793), .A2(n21146), .B1(n21132), .B2(n20798), .ZN(
        n20803) );
  OAI21_X1 U22994 ( .B1(n20795), .B2(n20794), .A(n20817), .ZN(n20796) );
  XOR2_X1 U22995 ( .A(n20797), .B(n20796), .Z(n20801) );
  NAND2_X1 U22996 ( .A1(n20799), .A2(n20798), .ZN(n20807) );
  OAI211_X1 U22997 ( .C1(n20799), .C2(n20798), .A(n21160), .B(n20807), .ZN(
        n20800) );
  OAI211_X1 U22998 ( .C1(n20801), .C2(n21851), .A(n11142), .B(n20800), .ZN(
        n20802) );
  AOI211_X1 U22999 ( .C1(P3_REIP_REG_5__SCAN_IN), .C2(n20823), .A(n20803), .B(
        n20802), .ZN(n20804) );
  OAI21_X1 U23000 ( .B1(n20806), .B2(n20805), .A(n20804), .ZN(P3_U2666) );
  AOI211_X1 U23001 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n20807), .A(n20826), .B(
        n21135), .ZN(n20808) );
  AOI21_X1 U23002 ( .B1(n21127), .B2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n20808), .ZN(n20815) );
  OAI21_X1 U23003 ( .B1(n20809), .B2(n21128), .A(n20901), .ZN(n20811) );
  OAI211_X1 U23004 ( .C1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n20818), .A(
        n20847), .B(n20812), .ZN(n20810) );
  NAND3_X1 U23005 ( .A1(n21075), .A2(n20821), .A3(n21476), .ZN(n20822) );
  OAI211_X1 U23006 ( .C1(n20812), .C2(n20811), .A(n20810), .B(n20822), .ZN(
        n20813) );
  AOI211_X1 U23007 ( .C1(P3_REIP_REG_6__SCAN_IN), .C2(n20823), .A(n21774), .B(
        n20813), .ZN(n20814) );
  OAI211_X1 U23008 ( .C1(n21132), .C2(n20816), .A(n20815), .B(n20814), .ZN(
        P3_U2665) );
  OAI21_X1 U23009 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20818), .A(
        n20817), .ZN(n20819) );
  XNOR2_X1 U23010 ( .A(n20820), .B(n20819), .ZN(n20833) );
  NAND2_X1 U23011 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n20821), .ZN(n20838) );
  NOR3_X1 U23012 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n21076), .A3(n20838), .ZN(
        n20831) );
  INV_X1 U23013 ( .A(n20822), .ZN(n20824) );
  OAI21_X1 U23014 ( .B1(n20824), .B2(n20823), .A(P3_REIP_REG_7__SCAN_IN), .ZN(
        n20828) );
  NAND2_X1 U23015 ( .A1(n20826), .A2(n20825), .ZN(n20837) );
  OAI211_X1 U23016 ( .C1(n20826), .C2(n20825), .A(n21160), .B(n20837), .ZN(
        n20827) );
  OAI211_X1 U23017 ( .C1(n21146), .C2(n20829), .A(n20828), .B(n20827), .ZN(
        n20830) );
  AOI211_X1 U23018 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n21161), .A(n20831), .B(
        n20830), .ZN(n20832) );
  OAI211_X1 U23019 ( .C1(n21851), .C2(n20833), .A(n20832), .B(n11142), .ZN(
        P3_U2664) );
  AOI21_X1 U23020 ( .B1(n20834), .B2(n20887), .A(n21128), .ZN(n20835) );
  XNOR2_X1 U23021 ( .A(n20836), .B(n20835), .ZN(n20846) );
  AOI211_X1 U23022 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n20837), .A(n20855), .B(
        n21135), .ZN(n20844) );
  NOR2_X1 U23023 ( .A1(n20839), .A2(n20838), .ZN(n20840) );
  AOI21_X1 U23024 ( .B1(n21075), .B2(n20840), .A(P3_REIP_REG_8__SCAN_IN), .ZN(
        n20842) );
  NAND2_X1 U23025 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n20840), .ZN(n20859) );
  INV_X1 U23026 ( .A(n21077), .ZN(n21157) );
  AOI21_X1 U23027 ( .B1(n20859), .B2(n21075), .A(n21157), .ZN(n20861) );
  OAI22_X1 U23028 ( .A1(n20842), .A2(n20861), .B1(n20841), .B2(n21146), .ZN(
        n20843) );
  AOI211_X1 U23029 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n21161), .A(n20844), .B(
        n20843), .ZN(n20845) );
  OAI211_X1 U23030 ( .C1(n21851), .C2(n20846), .A(n20845), .B(n11142), .ZN(
        P3_U2663) );
  AOI22_X1 U23031 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n21127), .B1(
        n21161), .B2(P3_EBX_REG_9__SCAN_IN), .ZN(n20858) );
  INV_X1 U23032 ( .A(n20861), .ZN(n20853) );
  INV_X1 U23033 ( .A(n20850), .ZN(n20851) );
  OAI21_X1 U23034 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20863), .A(
        n20847), .ZN(n20866) );
  OAI21_X1 U23035 ( .B1(n20848), .B2(n20933), .A(n20901), .ZN(n20849) );
  OAI221_X1 U23036 ( .B1(n20851), .B2(n20866), .C1(n20850), .C2(n20849), .A(
        n11142), .ZN(n20852) );
  AOI21_X1 U23037 ( .B1(P3_REIP_REG_9__SCAN_IN), .B2(n20853), .A(n20852), .ZN(
        n20857) );
  OR3_X1 U23038 ( .A1(n21076), .A2(n20859), .A3(P3_REIP_REG_9__SCAN_IN), .ZN(
        n20860) );
  INV_X1 U23039 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n20854) );
  NAND2_X1 U23040 ( .A1(n20855), .A2(n20854), .ZN(n20862) );
  OAI211_X1 U23041 ( .C1(n20855), .C2(n20854), .A(n21160), .B(n20862), .ZN(
        n20856) );
  NAND4_X1 U23042 ( .A1(n20858), .A2(n20857), .A3(n20860), .A4(n20856), .ZN(
        P3_U2662) );
  NAND2_X1 U23043 ( .A1(n21075), .A2(n20886), .ZN(n20873) );
  AOI22_X1 U23044 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n21127), .B1(
        n21161), .B2(P3_EBX_REG_10__SCAN_IN), .ZN(n20872) );
  NAND2_X1 U23045 ( .A1(n20861), .A2(n20860), .ZN(n20870) );
  AOI211_X1 U23046 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n20862), .A(n20882), .B(
        n21135), .ZN(n20869) );
  NOR2_X1 U23047 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20863), .ZN(
        n20864) );
  OAI211_X1 U23048 ( .C1(n20864), .C2(n21128), .A(n20970), .B(n20867), .ZN(
        n20865) );
  OAI211_X1 U23049 ( .C1(n20867), .C2(n20866), .A(n11142), .B(n20865), .ZN(
        n20868) );
  AOI211_X1 U23050 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(n20870), .A(n20869), 
        .B(n20868), .ZN(n20871) );
  OAI211_X1 U23051 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(n20873), .A(n20872), 
        .B(n20871), .ZN(P3_U2661) );
  AOI22_X1 U23052 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n21127), .B1(
        n21161), .B2(P3_EBX_REG_11__SCAN_IN), .ZN(n20885) );
  AOI21_X1 U23053 ( .B1(n20874), .B2(n21156), .A(n20933), .ZN(n20876) );
  XNOR2_X1 U23054 ( .A(n20876), .B(n20875), .ZN(n20880) );
  NAND3_X1 U23055 ( .A1(n21075), .A2(P3_REIP_REG_10__SCAN_IN), .A3(n20886), 
        .ZN(n20877) );
  NAND3_X1 U23056 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_11__SCAN_IN), 
        .A3(n20886), .ZN(n20918) );
  AOI21_X1 U23057 ( .B1(n21075), .B2(n20918), .A(n21157), .ZN(n20913) );
  AOI21_X1 U23058 ( .B1(n20878), .B2(n20877), .A(n20913), .ZN(n20879) );
  AOI211_X1 U23059 ( .C1(n20970), .C2(n20880), .A(n21774), .B(n20879), .ZN(
        n20884) );
  INV_X1 U23060 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n20881) );
  NAND2_X1 U23061 ( .A1(n20882), .A2(n20881), .ZN(n20891) );
  OAI211_X1 U23062 ( .C1(n20882), .C2(n20881), .A(n21160), .B(n20891), .ZN(
        n20883) );
  NAND3_X1 U23063 ( .A1(n20885), .A2(n20884), .A3(n20883), .ZN(P3_U2660) );
  NAND4_X1 U23064 ( .A1(n21075), .A2(P3_REIP_REG_10__SCAN_IN), .A3(
        P3_REIP_REG_11__SCAN_IN), .A4(n20886), .ZN(n20921) );
  AND2_X1 U23065 ( .A1(n18399), .A2(n20887), .ZN(n20899) );
  NOR2_X1 U23066 ( .A1(n20899), .A2(n21128), .ZN(n20889) );
  OAI21_X1 U23067 ( .B1(n20890), .B2(n20889), .A(n20970), .ZN(n20888) );
  AOI21_X1 U23068 ( .B1(n20890), .B2(n20889), .A(n20888), .ZN(n20896) );
  AOI211_X1 U23069 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n20891), .A(n20904), .B(
        n21135), .ZN(n20895) );
  OAI22_X1 U23070 ( .A1(n20893), .A2(n21146), .B1(n21132), .B2(n20892), .ZN(
        n20894) );
  NOR4_X1 U23071 ( .A1(n21774), .A2(n20896), .A3(n20895), .A4(n20894), .ZN(
        n20897) );
  OAI221_X1 U23072 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n20921), .C1(n20898), 
        .C2(n20913), .A(n20897), .ZN(P3_U2659) );
  AOI22_X1 U23073 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n21127), .B1(
        n21161), .B2(P3_EBX_REG_13__SCAN_IN), .ZN(n20912) );
  AOI21_X1 U23074 ( .B1(n20914), .B2(n20898), .A(n20921), .ZN(n20910) );
  NAND2_X1 U23075 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(P3_REIP_REG_12__SCAN_IN), 
        .ZN(n20922) );
  AOI21_X1 U23076 ( .B1(n20900), .B2(n20899), .A(n20933), .ZN(n20915) );
  NAND2_X1 U23077 ( .A1(n20970), .A2(n20915), .ZN(n20907) );
  OAI211_X1 U23078 ( .C1(n20902), .C2(n20933), .A(n20908), .B(n20901), .ZN(
        n20906) );
  INV_X1 U23079 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n20903) );
  NAND2_X1 U23080 ( .A1(n20904), .A2(n20903), .ZN(n20917) );
  OAI211_X1 U23081 ( .C1(n20904), .C2(n20903), .A(n21160), .B(n20917), .ZN(
        n20905) );
  OAI211_X1 U23082 ( .C1(n20908), .C2(n20907), .A(n20906), .B(n20905), .ZN(
        n20909) );
  AOI211_X1 U23083 ( .C1(n20910), .C2(n20922), .A(n21774), .B(n20909), .ZN(
        n20911) );
  OAI211_X1 U23084 ( .C1(n20914), .C2(n20913), .A(n20912), .B(n20911), .ZN(
        P3_U2658) );
  XNOR2_X1 U23085 ( .A(n20916), .B(n20915), .ZN(n20928) );
  AOI211_X1 U23086 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n20917), .A(n20931), .B(
        n21135), .ZN(n20926) );
  NOR3_X1 U23087 ( .A1(n20919), .A2(n20918), .A3(n20922), .ZN(n20958) );
  OAI21_X1 U23088 ( .B1(n21076), .B2(n20958), .A(n21077), .ZN(n20920) );
  INV_X1 U23089 ( .A(n20920), .ZN(n20944) );
  NOR2_X1 U23090 ( .A1(n20922), .A2(n20921), .ZN(n20929) );
  NOR2_X1 U23091 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n20929), .ZN(n20924) );
  OAI22_X1 U23092 ( .A1(n20944), .A2(n20924), .B1(n20923), .B2(n21146), .ZN(
        n20925) );
  AOI211_X1 U23093 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n21161), .A(n20926), .B(
        n20925), .ZN(n20927) );
  OAI211_X1 U23094 ( .C1(n21851), .C2(n20928), .A(n20927), .B(n11142), .ZN(
        P3_U2657) );
  NAND2_X1 U23095 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n20929), .ZN(n20946) );
  AOI22_X1 U23096 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n21127), .B1(
        n21161), .B2(P3_EBX_REG_15__SCAN_IN), .ZN(n20939) );
  NAND2_X1 U23097 ( .A1(n20931), .A2(n20930), .ZN(n20942) );
  OAI211_X1 U23098 ( .C1(n20931), .C2(n20930), .A(n21160), .B(n20942), .ZN(
        n20938) );
  NOR2_X1 U23099 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20932), .ZN(
        n20949) );
  INV_X1 U23100 ( .A(n20936), .ZN(n20965) );
  OAI221_X1 U23101 ( .B1(n20936), .B2(n20935), .C1(n20965), .C2(n20934), .A(
        n20970), .ZN(n20937) );
  AND4_X1 U23102 ( .A1(n20939), .A2(n11142), .A3(n20938), .A4(n20937), .ZN(
        n20940) );
  OAI221_X1 U23103 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n20946), .C1(n20941), 
        .C2(n20944), .A(n20940), .ZN(P3_U2656) );
  AOI211_X1 U23104 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n20942), .A(n20957), .B(
        n21135), .ZN(n20948) );
  XNOR2_X1 U23105 ( .A(P3_REIP_REG_16__SCAN_IN), .B(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n20945) );
  OAI22_X1 U23106 ( .A1(n20946), .A2(n20945), .B1(n20944), .B2(n20943), .ZN(
        n20947) );
  AOI211_X1 U23107 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n21161), .A(n20948), .B(
        n20947), .ZN(n20954) );
  AOI21_X1 U23108 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n20949), .A(
        n21128), .ZN(n20950) );
  XNOR2_X1 U23109 ( .A(n20951), .B(n20950), .ZN(n20952) );
  AOI21_X1 U23110 ( .B1(n20952), .B2(n20970), .A(n21774), .ZN(n20953) );
  OAI211_X1 U23111 ( .C1(n21146), .C2(n20955), .A(n20954), .B(n20953), .ZN(
        P3_U2655) );
  INV_X1 U23112 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n20961) );
  OAI21_X1 U23113 ( .B1(n20961), .B2(n20957), .A(n21160), .ZN(n20956) );
  INV_X1 U23114 ( .A(n20956), .ZN(n20964) );
  NAND2_X1 U23115 ( .A1(n20957), .A2(n20961), .ZN(n20977) );
  NAND3_X1 U23116 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .A3(n20958), .ZN(n20959) );
  NOR2_X1 U23117 ( .A1(n20960), .A2(n20959), .ZN(n20980) );
  AOI211_X1 U23118 ( .C1(n20960), .C2(n20959), .A(n20980), .B(n21076), .ZN(
        n20963) );
  OAI22_X1 U23119 ( .A1(n21132), .A2(n20961), .B1(n21077), .B2(n20960), .ZN(
        n20962) );
  AOI211_X1 U23120 ( .C1(n20964), .C2(n20977), .A(n20963), .B(n20962), .ZN(
        n20972) );
  OAI21_X1 U23121 ( .B1(n20966), .B2(n20933), .A(n20965), .ZN(n20967) );
  NOR2_X1 U23122 ( .A1(n20968), .A2(n20967), .ZN(n20974) );
  AOI21_X1 U23123 ( .B1(n20968), .B2(n20967), .A(n20974), .ZN(n20969) );
  AOI21_X1 U23124 ( .B1(n20970), .B2(n20969), .A(n21774), .ZN(n20971) );
  OAI211_X1 U23125 ( .C1(n21146), .C2(n20973), .A(n20972), .B(n20971), .ZN(
        P3_U2654) );
  AOI21_X1 U23126 ( .B1(n21161), .B2(P3_EBX_REG_18__SCAN_IN), .A(n21774), .ZN(
        n20983) );
  NOR2_X1 U23127 ( .A1(n20974), .A2(n21128), .ZN(n20975) );
  NOR2_X1 U23128 ( .A1(n20976), .A2(n20975), .ZN(n20984) );
  AOI211_X1 U23129 ( .C1(n20976), .C2(n20975), .A(n20984), .B(n21851), .ZN(
        n20979) );
  AOI211_X1 U23130 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n20977), .A(n20993), .B(
        n21135), .ZN(n20978) );
  AOI211_X1 U23131 ( .C1(n21127), .C2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n20979), .B(n20978), .ZN(n20982) );
  NAND2_X1 U23132 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n20980), .ZN(n20997) );
  INV_X1 U23133 ( .A(n20997), .ZN(n20987) );
  OAI21_X1 U23134 ( .B1(n20987), .B2(n21076), .A(n21077), .ZN(n20991) );
  OAI221_X1 U23135 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n21075), .C1(
        P3_REIP_REG_18__SCAN_IN), .C2(n20980), .A(n20991), .ZN(n20981) );
  NAND3_X1 U23136 ( .A1(n20983), .A2(n20982), .A3(n20981), .ZN(P3_U2653) );
  NOR2_X1 U23137 ( .A1(n20985), .A2(n20986), .ZN(n21001) );
  AOI211_X1 U23138 ( .C1(n20986), .C2(n20985), .A(n21001), .B(n21851), .ZN(
        n20990) );
  NAND3_X1 U23139 ( .A1(n21075), .A2(n20987), .A3(n20998), .ZN(n20988) );
  OAI211_X1 U23140 ( .C1(n21132), .C2(n20992), .A(n11142), .B(n20988), .ZN(
        n20989) );
  AOI211_X1 U23141 ( .C1(n20991), .C2(P3_REIP_REG_19__SCAN_IN), .A(n20990), 
        .B(n20989), .ZN(n20995) );
  NAND2_X1 U23142 ( .A1(n20993), .A2(n20992), .ZN(n21004) );
  OAI211_X1 U23143 ( .C1(n20993), .C2(n20992), .A(n21160), .B(n21004), .ZN(
        n20994) );
  OAI211_X1 U23144 ( .C1(n21146), .C2(n20996), .A(n20995), .B(n20994), .ZN(
        P3_U2652) );
  NOR2_X1 U23145 ( .A1(n20998), .A2(n20997), .ZN(n21000) );
  NAND2_X1 U23146 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n21000), .ZN(n21035) );
  INV_X1 U23147 ( .A(n21035), .ZN(n21014) );
  OAI21_X1 U23148 ( .B1(n21076), .B2(n21014), .A(n21077), .ZN(n21017) );
  INV_X1 U23149 ( .A(n21017), .ZN(n21034) );
  NOR2_X1 U23150 ( .A1(n21014), .A2(n21076), .ZN(n20999) );
  AOI22_X1 U23151 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n21127), .B1(
        n21000), .B2(n20999), .ZN(n21008) );
  NOR2_X1 U23152 ( .A1(n21001), .A2(n21128), .ZN(n21002) );
  NOR2_X1 U23153 ( .A1(n21003), .A2(n21002), .ZN(n21010) );
  AOI211_X1 U23154 ( .C1(n21003), .C2(n21002), .A(n21010), .B(n21851), .ZN(
        n21006) );
  AOI211_X1 U23155 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n21004), .A(n21019), .B(
        n21135), .ZN(n21005) );
  AOI211_X1 U23156 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n21161), .A(n21006), .B(
        n21005), .ZN(n21007) );
  OAI211_X1 U23157 ( .C1(n21034), .C2(n21009), .A(n21008), .B(n21007), .ZN(
        P3_U2651) );
  INV_X1 U23158 ( .A(n21011), .ZN(n21012) );
  NOR2_X1 U23159 ( .A1(n21013), .A2(n21012), .ZN(n21025) );
  AOI211_X1 U23160 ( .C1(n21013), .C2(n21012), .A(n21025), .B(n21851), .ZN(
        n21016) );
  NAND2_X1 U23161 ( .A1(n21075), .A2(n21014), .ZN(n21037) );
  OAI22_X1 U23162 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n21037), .B1(n21132), 
        .B2(n21018), .ZN(n21015) );
  AOI211_X1 U23163 ( .C1(P3_REIP_REG_21__SCAN_IN), .C2(n21017), .A(n21016), 
        .B(n21015), .ZN(n21021) );
  NAND2_X1 U23164 ( .A1(n21019), .A2(n21018), .ZN(n21024) );
  OAI211_X1 U23165 ( .C1(n21019), .C2(n21018), .A(n21160), .B(n21024), .ZN(
        n21020) );
  OAI211_X1 U23166 ( .C1(n21146), .C2(n21022), .A(n21021), .B(n21020), .ZN(
        P3_U2650) );
  AOI22_X1 U23167 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n21127), .B1(
        n21161), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n21032) );
  AOI21_X1 U23168 ( .B1(n21033), .B2(n21023), .A(n21037), .ZN(n21030) );
  NAND2_X1 U23169 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .ZN(n21038) );
  AOI211_X1 U23170 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n21024), .A(n21046), .B(
        n21135), .ZN(n21029) );
  AOI211_X1 U23171 ( .C1(n21027), .C2(n21026), .A(n11265), .B(n21851), .ZN(
        n21028) );
  AOI211_X1 U23172 ( .C1(n21030), .C2(n21038), .A(n21029), .B(n21028), .ZN(
        n21031) );
  OAI211_X1 U23173 ( .C1(n21034), .C2(n21033), .A(n21032), .B(n21031), .ZN(
        P3_U2649) );
  NOR3_X1 U23174 ( .A1(n21036), .A2(n21035), .A3(n21038), .ZN(n21063) );
  OAI21_X1 U23175 ( .B1(n21063), .B2(n21076), .A(n21077), .ZN(n21059) );
  OAI21_X1 U23176 ( .B1(n21038), .B2(n21037), .A(n21036), .ZN(n21044) );
  AOI211_X1 U23177 ( .C1(n21040), .C2(n21039), .A(n21051), .B(n21851), .ZN(
        n21043) );
  OAI22_X1 U23178 ( .A1(n21041), .A2(n21146), .B1(n21132), .B2(n21045), .ZN(
        n21042) );
  AOI211_X1 U23179 ( .C1(n21059), .C2(n21044), .A(n21043), .B(n21042), .ZN(
        n21048) );
  NAND2_X1 U23180 ( .A1(n21046), .A2(n21045), .ZN(n21050) );
  OAI211_X1 U23181 ( .C1(n21046), .C2(n21045), .A(n21160), .B(n21050), .ZN(
        n21047) );
  NAND2_X1 U23182 ( .A1(n21048), .A2(n21047), .ZN(P3_U2648) );
  NOR2_X1 U23183 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n21076), .ZN(n21049) );
  AOI22_X1 U23184 ( .A1(n21161), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n21063), 
        .B2(n21049), .ZN(n21057) );
  AOI211_X1 U23185 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n21050), .A(n21069), .B(
        n21135), .ZN(n21055) );
  NOR2_X1 U23186 ( .A1(n21051), .A2(n21128), .ZN(n21052) );
  NOR2_X1 U23187 ( .A1(n21052), .A2(n21053), .ZN(n21060) );
  AOI211_X1 U23188 ( .C1(n21053), .C2(n21052), .A(n21060), .B(n21851), .ZN(
        n21054) );
  AOI211_X1 U23189 ( .C1(n21059), .C2(P3_REIP_REG_24__SCAN_IN), .A(n21055), 
        .B(n21054), .ZN(n21056) );
  OAI211_X1 U23190 ( .C1(n21058), .C2(n21146), .A(n21057), .B(n21056), .ZN(
        P3_U2647) );
  AOI21_X1 U23191 ( .B1(n21075), .B2(n21702), .A(n21059), .ZN(n21072) );
  AOI211_X1 U23192 ( .C1(n21062), .C2(n21061), .A(n21081), .B(n21851), .ZN(
        n21067) );
  NAND2_X1 U23193 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n21063), .ZN(n21073) );
  NOR3_X1 U23194 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n21076), .A3(n21073), 
        .ZN(n21066) );
  OAI22_X1 U23195 ( .A1(n21064), .A2(n21146), .B1(n21132), .B2(n21068), .ZN(
        n21065) );
  NOR3_X1 U23196 ( .A1(n21067), .A2(n21066), .A3(n21065), .ZN(n21071) );
  NAND2_X1 U23197 ( .A1(n21069), .A2(n21068), .ZN(n21079) );
  OAI211_X1 U23198 ( .C1(n21069), .C2(n21068), .A(n21160), .B(n21079), .ZN(
        n21070) );
  OAI211_X1 U23199 ( .C1(n21072), .C2(n21074), .A(n21071), .B(n21070), .ZN(
        P3_U2646) );
  AOI22_X1 U23200 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n21127), .B1(
        n21161), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n21088) );
  NOR2_X1 U23201 ( .A1(n21074), .A2(n21073), .ZN(n21078) );
  NAND2_X1 U23202 ( .A1(n21077), .A2(n21076), .ZN(n21159) );
  NAND3_X1 U23203 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n21078), .A3(n21077), 
        .ZN(n21111) );
  AND2_X1 U23204 ( .A1(n21159), .A2(n21111), .ZN(n21107) );
  OAI21_X1 U23205 ( .B1(P3_REIP_REG_26__SCAN_IN), .B2(n21089), .A(n21107), 
        .ZN(n21087) );
  AOI211_X1 U23206 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n21079), .A(n21097), .B(
        n21135), .ZN(n21085) );
  INV_X1 U23207 ( .A(n21080), .ZN(n21083) );
  AOI211_X1 U23208 ( .C1(n21083), .C2(n21082), .A(n21090), .B(n21851), .ZN(
        n21084) );
  NOR2_X1 U23209 ( .A1(n21085), .A2(n21084), .ZN(n21086) );
  NAND3_X1 U23210 ( .A1(n21088), .A2(n21087), .A3(n21086), .ZN(P3_U2645) );
  NAND2_X1 U23211 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n21089), .ZN(n21125) );
  NOR2_X1 U23212 ( .A1(n21090), .A2(n21128), .ZN(n21091) );
  NOR2_X1 U23213 ( .A1(n21091), .A2(n21092), .ZN(n21102) );
  AOI211_X1 U23214 ( .C1(n21092), .C2(n21091), .A(n21102), .B(n21851), .ZN(
        n21095) );
  INV_X1 U23215 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n21096) );
  OAI22_X1 U23216 ( .A1(n21093), .A2(n21146), .B1(n21132), .B2(n21096), .ZN(
        n21094) );
  AOI211_X1 U23217 ( .C1(n21107), .C2(P3_REIP_REG_27__SCAN_IN), .A(n21095), 
        .B(n21094), .ZN(n21099) );
  NAND2_X1 U23218 ( .A1(n21097), .A2(n21096), .ZN(n21100) );
  OAI211_X1 U23219 ( .C1(n21097), .C2(n21096), .A(n21160), .B(n21100), .ZN(
        n21098) );
  OAI211_X1 U23220 ( .C1(P3_REIP_REG_27__SCAN_IN), .C2(n21125), .A(n21099), 
        .B(n21098), .ZN(P3_U2644) );
  NAND2_X1 U23221 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n21115) );
  OAI21_X1 U23222 ( .B1(P3_REIP_REG_28__SCAN_IN), .B2(P3_REIP_REG_27__SCAN_IN), 
        .A(n21115), .ZN(n21110) );
  AOI22_X1 U23223 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n21127), .B1(
        n21161), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n21109) );
  NOR2_X1 U23224 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n21100), .ZN(n21113) );
  AOI211_X1 U23225 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n21100), .A(n21113), .B(
        n21135), .ZN(n21106) );
  INV_X1 U23226 ( .A(n21101), .ZN(n21104) );
  AOI211_X1 U23227 ( .C1(n21104), .C2(n21103), .A(n21116), .B(n21851), .ZN(
        n21105) );
  AOI211_X1 U23228 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n21107), .A(n21106), 
        .B(n21105), .ZN(n21108) );
  OAI211_X1 U23229 ( .C1(n21125), .C2(n21110), .A(n21109), .B(n21108), .ZN(
        P3_U2643) );
  NAND3_X1 U23230 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n21126) );
  OAI21_X1 U23231 ( .B1(n21126), .B2(n21111), .A(n21159), .ZN(n21148) );
  AOI22_X1 U23232 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n21127), .B1(
        n21161), .B2(P3_EBX_REG_29__SCAN_IN), .ZN(n21123) );
  INV_X1 U23233 ( .A(n21113), .ZN(n21114) );
  NAND2_X1 U23234 ( .A1(n21113), .A2(n21112), .ZN(n21134) );
  NAND2_X1 U23235 ( .A1(n21160), .A2(n21134), .ZN(n21133) );
  AOI21_X1 U23236 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n21114), .A(n21133), .ZN(
        n21121) );
  NOR3_X1 U23237 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n21115), .A3(n21125), 
        .ZN(n21120) );
  AOI211_X1 U23238 ( .C1(n21118), .C2(n21117), .A(n21129), .B(n21851), .ZN(
        n21119) );
  NOR3_X1 U23239 ( .A1(n21121), .A2(n21120), .A3(n21119), .ZN(n21122) );
  OAI211_X1 U23240 ( .C1(n21124), .C2(n21148), .A(n21123), .B(n21122), .ZN(
        P3_U2642) );
  NOR2_X1 U23241 ( .A1(n21126), .A2(n21125), .ZN(n21151) );
  AOI22_X1 U23242 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n21127), .B1(
        n21151), .B2(n21152), .ZN(n21142) );
  INV_X1 U23243 ( .A(n21130), .ZN(n21145) );
  XNOR2_X1 U23244 ( .A(n21144), .B(n21145), .ZN(n21139) );
  INV_X1 U23245 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n21131) );
  INV_X1 U23246 ( .A(n21140), .ZN(n21141) );
  OAI211_X1 U23247 ( .C1(n21152), .C2(n21148), .A(n21142), .B(n21141), .ZN(
        P3_U2641) );
  NOR3_X1 U23248 ( .A1(n21145), .A2(n21144), .A3(n21143), .ZN(n21150) );
  OAI22_X1 U23249 ( .A1(n21153), .A2(n21148), .B1(n21147), .B2(n21146), .ZN(
        n21149) );
  AOI211_X1 U23250 ( .C1(n21161), .C2(P3_EBX_REG_31__SCAN_IN), .A(n21150), .B(
        n21149), .ZN(n21155) );
  OAI221_X1 U23251 ( .B1(P3_REIP_REG_31__SCAN_IN), .B2(P3_REIP_REG_30__SCAN_IN), .C1(n21153), .C2(n21152), .A(n21151), .ZN(n21154) );
  OAI211_X1 U23252 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n11646), .A(n21155), .B(
        n21154), .ZN(P3_U2640) );
  NOR3_X1 U23253 ( .A1(n21390), .A2(n21157), .A3(n21156), .ZN(n21158) );
  AOI21_X1 U23254 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(n21159), .A(n21158), .ZN(
        n21163) );
  OAI21_X1 U23255 ( .B1(n21161), .B2(n21160), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n21162) );
  OAI211_X1 U23256 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n21164), .A(
        n21163), .B(n21162), .ZN(P3_U2671) );
  NAND4_X1 U23257 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_5__SCAN_IN), 
        .A3(P3_EAX_REG_6__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n21168) );
  NAND4_X1 U23258 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(P3_EAX_REG_3__SCAN_IN), 
        .A3(P3_EAX_REG_4__SCAN_IN), .A4(n21169), .ZN(n21332) );
  NOR2_X1 U23259 ( .A1(n21267), .A2(n21332), .ZN(n21331) );
  NAND2_X1 U23260 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n21331), .ZN(n21189) );
  NAND2_X1 U23261 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n21194), .ZN(n21186) );
  NAND2_X1 U23262 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n21183), .ZN(n21175) );
  NAND2_X1 U23263 ( .A1(n21175), .A2(P3_EAX_REG_13__SCAN_IN), .ZN(n21174) );
  AOI22_X1 U23264 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n21345), .B1(n21338), .B2(
        n21172), .ZN(n21173) );
  OAI221_X1 U23265 ( .B1(n21175), .B2(P3_EAX_REG_13__SCAN_IN), .C1(n21174), 
        .C2(n21324), .A(n21173), .ZN(P3_U2722) );
  INV_X1 U23266 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n21178) );
  INV_X1 U23267 ( .A(n21175), .ZN(n21318) );
  AOI21_X1 U23268 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n21333), .A(n21183), .ZN(
        n21177) );
  OAI222_X1 U23269 ( .A1(n21227), .A2(n21178), .B1(n21318), .B2(n21177), .C1(
        n21349), .C2(n21176), .ZN(P3_U2723) );
  INV_X1 U23270 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n21184) );
  OAI21_X1 U23271 ( .B1(n21179), .B2(n21324), .A(n21186), .ZN(n21180) );
  INV_X1 U23272 ( .A(n21180), .ZN(n21182) );
  OAI222_X1 U23273 ( .A1(n21227), .A2(n21184), .B1(n21183), .B2(n21182), .C1(
        n21349), .C2(n21181), .ZN(P3_U2724) );
  AOI22_X1 U23274 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n21345), .B1(n21338), .B2(
        n21185), .ZN(n21188) );
  OAI211_X1 U23275 ( .C1(P3_EAX_REG_10__SCAN_IN), .C2(n21194), .A(n21333), .B(
        n21186), .ZN(n21187) );
  NAND2_X1 U23276 ( .A1(n21188), .A2(n21187), .ZN(P3_U2725) );
  INV_X1 U23277 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n21195) );
  OAI21_X1 U23278 ( .B1(n21190), .B2(n21324), .A(n21189), .ZN(n21191) );
  INV_X1 U23279 ( .A(n21191), .ZN(n21193) );
  OAI222_X1 U23280 ( .A1(n21227), .A2(n21195), .B1(n21194), .B2(n21193), .C1(
        n21349), .C2(n21192), .ZN(P3_U2726) );
  NAND2_X1 U23281 ( .A1(n21197), .A2(n21196), .ZN(n21339) );
  NOR2_X1 U23282 ( .A1(n21198), .A2(n21339), .ZN(n21341) );
  NAND2_X1 U23283 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n21341), .ZN(n21221) );
  NAND2_X1 U23284 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n21226), .ZN(n21212) );
  NOR2_X1 U23285 ( .A1(n21199), .A2(n21212), .ZN(n21215) );
  NAND2_X1 U23286 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n21215), .ZN(n21203) );
  NOR2_X1 U23287 ( .A1(n21200), .A2(n21203), .ZN(n21206) );
  AOI21_X1 U23288 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n21333), .A(n21206), .ZN(
        n21201) );
  OAI222_X1 U23289 ( .A1(n21202), .A2(n21227), .B1(n21331), .B2(n21201), .C1(
        n21349), .C2(n21653), .ZN(P3_U2728) );
  INV_X1 U23290 ( .A(n21203), .ZN(n21210) );
  AOI21_X1 U23291 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n21333), .A(n21210), .ZN(
        n21205) );
  OAI222_X1 U23292 ( .A1(n21207), .A2(n21227), .B1(n21206), .B2(n21205), .C1(
        n21349), .C2(n21204), .ZN(P3_U2729) );
  AOI21_X1 U23293 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n21333), .A(n21215), .ZN(
        n21209) );
  OAI222_X1 U23294 ( .A1(n21211), .A2(n21227), .B1(n21210), .B2(n21209), .C1(
        n21349), .C2(n21208), .ZN(P3_U2730) );
  INV_X1 U23295 ( .A(n21212), .ZN(n21219) );
  AOI21_X1 U23296 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n21333), .A(n21219), .ZN(
        n21214) );
  OAI222_X1 U23297 ( .A1(n21216), .A2(n21227), .B1(n21215), .B2(n21214), .C1(
        n21349), .C2(n21213), .ZN(P3_U2731) );
  AOI21_X1 U23298 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n21333), .A(n21226), .ZN(
        n21218) );
  OAI222_X1 U23299 ( .A1(n21220), .A2(n21227), .B1(n21219), .B2(n21218), .C1(
        n21349), .C2(n21217), .ZN(P3_U2732) );
  OAI21_X1 U23300 ( .B1(n21222), .B2(n21324), .A(n21221), .ZN(n21223) );
  INV_X1 U23301 ( .A(n21223), .ZN(n21225) );
  OAI222_X1 U23302 ( .A1(n21228), .A2(n21227), .B1(n21226), .B2(n21225), .C1(
        n21349), .C2(n21224), .ZN(P3_U2733) );
  NOR2_X1 U23303 ( .A1(n21242), .A2(n21229), .ZN(n21243) );
  NAND4_X1 U23304 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_14__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(P3_EAX_REG_13__SCAN_IN), .ZN(n21230)
         );
  NAND2_X1 U23305 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n21261), .ZN(n21260) );
  NAND2_X1 U23306 ( .A1(n21243), .A2(n21254), .ZN(n21238) );
  NAND2_X1 U23307 ( .A1(n21333), .A2(n21238), .ZN(n21245) );
  NOR2_X2 U23308 ( .A1(n21231), .A2(n21333), .ZN(n21313) );
  NAND2_X1 U23309 ( .A1(n21232), .A2(n21324), .ZN(n21306) );
  OAI22_X1 U23310 ( .A1(n21233), .A2(n21349), .B1(n16811), .B2(n21306), .ZN(
        n21234) );
  AOI21_X1 U23311 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n21313), .A(n21234), .ZN(
        n21235) );
  OAI221_X1 U23312 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n21238), .C1(n21236), 
        .C2(n21245), .A(n21235), .ZN(P3_U2714) );
  AOI22_X1 U23313 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n21312), .B1(n21338), .B2(
        n21237), .ZN(n21241) );
  NAND2_X1 U23314 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n21254), .ZN(n21250) );
  INV_X1 U23315 ( .A(n21250), .ZN(n21239) );
  AOI22_X1 U23316 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n21313), .B1(n21239), .B2(
        n21238), .ZN(n21240) );
  OAI211_X1 U23317 ( .C1(n21242), .C2(n21245), .A(n21241), .B(n21240), .ZN(
        P3_U2715) );
  NAND4_X1 U23318 ( .A1(n21243), .A2(P3_EAX_REG_18__SCAN_IN), .A3(
        P3_EAX_REG_17__SCAN_IN), .A4(P3_EAX_REG_21__SCAN_IN), .ZN(n21266) );
  NAND2_X1 U23319 ( .A1(n21261), .A2(n21265), .ZN(n21249) );
  AOI22_X1 U23320 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n21312), .B1(n21338), .B2(
        n21244), .ZN(n21248) );
  OAI21_X1 U23321 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n21339), .A(n21245), .ZN(
        n21246) );
  AOI22_X1 U23322 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n21313), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n21246), .ZN(n21247) );
  OAI211_X1 U23323 ( .C1(n21266), .C2(n21249), .A(n21248), .B(n21247), .ZN(
        P3_U2713) );
  AOI22_X1 U23324 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n21313), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n21312), .ZN(n21252) );
  OAI211_X1 U23325 ( .C1(n21254), .C2(P3_EAX_REG_19__SCAN_IN), .A(n21333), .B(
        n21250), .ZN(n21251) );
  OAI211_X1 U23326 ( .C1(n21253), .C2(n21349), .A(n21252), .B(n21251), .ZN(
        P3_U2716) );
  AOI22_X1 U23327 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n21313), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n21312), .ZN(n21258) );
  AOI211_X1 U23328 ( .C1(n21255), .C2(n21260), .A(n21254), .B(n21324), .ZN(
        n21256) );
  INV_X1 U23329 ( .A(n21256), .ZN(n21257) );
  OAI211_X1 U23330 ( .C1(n21259), .C2(n21349), .A(n21258), .B(n21257), .ZN(
        P3_U2717) );
  AOI22_X1 U23331 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n21313), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n21312), .ZN(n21263) );
  OAI211_X1 U23332 ( .C1(n21261), .C2(P3_EAX_REG_17__SCAN_IN), .A(n21333), .B(
        n21260), .ZN(n21262) );
  OAI211_X1 U23333 ( .C1(n21264), .C2(n21349), .A(n21263), .B(n21262), .ZN(
        P3_U2718) );
  AOI22_X1 U23334 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n21313), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n21312), .ZN(n21270) );
  NAND2_X1 U23335 ( .A1(n21308), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n21307) );
  NAND2_X1 U23336 ( .A1(n21302), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n21301) );
  OAI211_X1 U23337 ( .C1(n21268), .C2(P3_EAX_REG_25__SCAN_IN), .A(n21333), .B(
        n21273), .ZN(n21269) );
  OAI211_X1 U23338 ( .C1(n21271), .C2(n21349), .A(n21270), .B(n21269), .ZN(
        P3_U2710) );
  AOI22_X1 U23339 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n21313), .B1(n21338), .B2(
        n21272), .ZN(n21277) );
  AOI211_X1 U23340 ( .C1(n21274), .C2(n21273), .A(n21296), .B(n21324), .ZN(
        n21275) );
  INV_X1 U23341 ( .A(n21275), .ZN(n21276) );
  OAI211_X1 U23342 ( .C1(n21306), .C2(n16774), .A(n21277), .B(n21276), .ZN(
        P3_U2709) );
  NAND2_X1 U23343 ( .A1(n21281), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n21280) );
  NAND2_X1 U23344 ( .A1(n21280), .A2(P3_EAX_REG_31__SCAN_IN), .ZN(n21279) );
  NAND2_X1 U23345 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n21312), .ZN(n21278) );
  OAI221_X1 U23346 ( .B1(n21280), .B2(P3_EAX_REG_31__SCAN_IN), .C1(n21279), 
        .C2(n21324), .A(n21278), .ZN(P3_U2704) );
  AOI22_X1 U23347 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n21313), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n21312), .ZN(n21283) );
  OAI211_X1 U23348 ( .C1(n21281), .C2(P3_EAX_REG_30__SCAN_IN), .A(n21333), .B(
        n21280), .ZN(n21282) );
  OAI211_X1 U23349 ( .C1(n21284), .C2(n21349), .A(n21283), .B(n21282), .ZN(
        P3_U2705) );
  AOI22_X1 U23350 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n21313), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n21312), .ZN(n21287) );
  OAI211_X1 U23351 ( .C1(n11227), .C2(P3_EAX_REG_29__SCAN_IN), .A(n21333), .B(
        n21285), .ZN(n21286) );
  OAI211_X1 U23352 ( .C1(n21288), .C2(n21349), .A(n21287), .B(n21286), .ZN(
        P3_U2706) );
  AOI22_X1 U23353 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n21313), .B1(n21338), .B2(
        n21289), .ZN(n21293) );
  AOI211_X1 U23354 ( .C1(n21290), .C2(n21295), .A(n11227), .B(n21324), .ZN(
        n21291) );
  INV_X1 U23355 ( .A(n21291), .ZN(n21292) );
  OAI211_X1 U23356 ( .C1(n21306), .C2(n21294), .A(n21293), .B(n21292), .ZN(
        P3_U2707) );
  AOI22_X1 U23357 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n21313), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n21312), .ZN(n21298) );
  OAI211_X1 U23358 ( .C1(n21296), .C2(P3_EAX_REG_27__SCAN_IN), .A(n21333), .B(
        n21295), .ZN(n21297) );
  OAI211_X1 U23359 ( .C1(n21299), .C2(n21349), .A(n21298), .B(n21297), .ZN(
        P3_U2708) );
  INV_X1 U23360 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n21305) );
  AOI22_X1 U23361 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n21313), .B1(n21338), .B2(
        n21300), .ZN(n21304) );
  OAI211_X1 U23362 ( .C1(n21302), .C2(P3_EAX_REG_24__SCAN_IN), .A(n21333), .B(
        n21301), .ZN(n21303) );
  OAI211_X1 U23363 ( .C1(n21306), .C2(n21305), .A(n21304), .B(n21303), .ZN(
        P3_U2711) );
  AOI22_X1 U23364 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n21313), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n21312), .ZN(n21310) );
  OAI211_X1 U23365 ( .C1(n21308), .C2(P3_EAX_REG_23__SCAN_IN), .A(n21333), .B(
        n21307), .ZN(n21309) );
  OAI211_X1 U23366 ( .C1(n21311), .C2(n21349), .A(n21310), .B(n21309), .ZN(
        P3_U2712) );
  AOI22_X1 U23367 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n21313), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n21312), .ZN(n21316) );
  OAI211_X1 U23368 ( .C1(n21323), .C2(P3_EAX_REG_16__SCAN_IN), .A(n21333), .B(
        n21314), .ZN(n21315) );
  OAI211_X1 U23369 ( .C1(n21317), .C2(n21349), .A(n21316), .B(n21315), .ZN(
        P3_U2719) );
  NAND2_X1 U23370 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n21318), .ZN(n21322) );
  AOI22_X1 U23371 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n21345), .B1(n21338), .B2(
        n21319), .ZN(n21321) );
  NAND3_X1 U23372 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n21333), .A3(n21326), 
        .ZN(n21320) );
  OAI211_X1 U23373 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n21322), .A(n21321), .B(
        n21320), .ZN(P3_U2721) );
  AOI211_X1 U23374 ( .C1(n21326), .C2(n21325), .A(n21324), .B(n21323), .ZN(
        n21327) );
  AOI21_X1 U23375 ( .B1(n21345), .B2(BUF2_REG_15__SCAN_IN), .A(n21327), .ZN(
        n21328) );
  OAI21_X1 U23376 ( .B1(n21329), .B2(n21349), .A(n21328), .ZN(P3_U2720) );
  AOI22_X1 U23377 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n21345), .B1(n21331), .B2(
        n21330), .ZN(n21335) );
  NAND3_X1 U23378 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n21333), .A3(n21332), .ZN(
        n21334) );
  OAI211_X1 U23379 ( .C1(n21336), .C2(n21349), .A(n21335), .B(n21334), .ZN(
        P3_U2727) );
  AOI22_X1 U23380 ( .A1(n21345), .A2(BUF2_REG_1__SCAN_IN), .B1(n21338), .B2(
        n21337), .ZN(n21343) );
  NOR2_X1 U23381 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n21339), .ZN(n21346) );
  OAI22_X1 U23382 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n21341), .B1(n21346), .B2(
        n21340), .ZN(n21342) );
  NAND2_X1 U23383 ( .A1(n21343), .A2(n21342), .ZN(P3_U2734) );
  AOI22_X1 U23384 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n21345), .B1(
        P3_EAX_REG_0__SCAN_IN), .B2(n21344), .ZN(n21348) );
  INV_X1 U23385 ( .A(n21346), .ZN(n21347) );
  OAI211_X1 U23386 ( .C1(n21350), .C2(n21349), .A(n21348), .B(n21347), .ZN(
        P3_U2735) );
  INV_X1 U23387 ( .A(n21393), .ZN(n21372) );
  AOI21_X1 U23388 ( .B1(n21576), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n21776), .ZN(n21381) );
  OAI22_X1 U23389 ( .A1(n21351), .A2(n21352), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n21381), .ZN(n21829) );
  INV_X1 U23390 ( .A(n21352), .ZN(n21355) );
  OAI22_X1 U23391 ( .A1(n21443), .A2(n21353), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21365) );
  NOR2_X1 U23392 ( .A1(n21354), .A2(n21508), .ZN(n21369) );
  AOI222_X1 U23393 ( .A1(n21829), .A2(n21390), .B1(n21367), .B2(n21355), .C1(
        n21365), .C2(n21369), .ZN(n21356) );
  AOI22_X1 U23394 ( .A1(n21372), .A2(n21382), .B1(n21356), .B2(n21393), .ZN(
        P3_U3289) );
  INV_X1 U23395 ( .A(n21377), .ZN(n21361) );
  OAI22_X1 U23396 ( .A1(n21359), .A2(n21358), .B1(n21373), .B2(n21357), .ZN(
        n21379) );
  OAI211_X1 U23397 ( .C1(n21361), .C2(n21379), .A(n21360), .B(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n21364) );
  AOI211_X1 U23398 ( .C1(n21371), .C2(n21382), .A(n21381), .B(n21376), .ZN(
        n21362) );
  INV_X1 U23399 ( .A(n21362), .ZN(n21363) );
  OAI211_X1 U23400 ( .C1(n21812), .C2(n21366), .A(n21364), .B(n21363), .ZN(
        n21823) );
  INV_X1 U23401 ( .A(n21365), .ZN(n21368) );
  AOI222_X1 U23402 ( .A1(n21823), .A2(n21390), .B1(n21369), .B2(n21368), .C1(
        n21367), .C2(n21366), .ZN(n21370) );
  AOI22_X1 U23403 ( .A1(n21372), .A2(n21371), .B1(n21370), .B2(n21393), .ZN(
        P3_U3288) );
  NOR2_X1 U23404 ( .A1(n21374), .A2(n21373), .ZN(n21375) );
  OAI22_X1 U23405 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21377), .B1(
        n21376), .B2(n21375), .ZN(n21378) );
  AOI21_X1 U23406 ( .B1(n21380), .B2(n21379), .A(n21378), .ZN(n21389) );
  OR3_X1 U23407 ( .A1(n21383), .A2(n21382), .A3(n21381), .ZN(n21387) );
  INV_X1 U23408 ( .A(n21385), .ZN(n21384) );
  OAI221_X1 U23409 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n21385), 
        .C1(n21388), .C2(n21384), .A(n21736), .ZN(n21386) );
  OAI211_X1 U23410 ( .C1(n21389), .C2(n21388), .A(n21387), .B(n21386), .ZN(
        n21821) );
  NAND2_X1 U23411 ( .A1(n21821), .A2(n21390), .ZN(n21395) );
  OAI21_X1 U23412 ( .B1(n21864), .B2(n21391), .A(n21393), .ZN(n21392) );
  OAI21_X1 U23413 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n21393), .A(
        n21392), .ZN(n21394) );
  OAI21_X1 U23414 ( .B1(n21396), .B2(n21395), .A(n21394), .ZN(P3_U3285) );
  OAI22_X1 U23415 ( .A1(n21397), .A2(n21811), .B1(n21731), .B2(n21509), .ZN(
        n21506) );
  NAND2_X1 U23416 ( .A1(n21725), .A2(n21506), .ZN(n21574) );
  AOI221_X1 U23417 ( .B1(n21399), .B2(n21574), .C1(n21727), .C2(n21574), .A(
        n21398), .ZN(n21400) );
  OAI211_X1 U23418 ( .C1(n21401), .C2(n21400), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B(n21793), .ZN(n21723) );
  AOI22_X1 U23419 ( .A1(n14606), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n21801), 
        .B2(n21402), .ZN(n21414) );
  OAI221_X1 U23420 ( .B1(n21790), .B2(n21403), .C1(n21790), .C2(n21556), .A(
        n21793), .ZN(n21703) );
  INV_X1 U23421 ( .A(n21735), .ZN(n21406) );
  OAI21_X1 U23422 ( .B1(n21727), .B2(n21404), .A(n21776), .ZN(n21405) );
  OAI221_X1 U23423 ( .B1(n21812), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), 
        .C1(n21812), .C2(n21406), .A(n21405), .ZN(n21704) );
  OAI22_X1 U23424 ( .A1(n21795), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n21411), .B2(n21812), .ZN(n21410) );
  OAI22_X1 U23425 ( .A1(n21408), .A2(n21811), .B1(n21407), .B2(n21731), .ZN(
        n21409) );
  NOR3_X1 U23426 ( .A1(n21704), .A2(n21410), .A3(n21409), .ZN(n21578) );
  OAI21_X1 U23427 ( .B1(n21790), .B2(n21411), .A(n21578), .ZN(n21412) );
  OAI211_X1 U23428 ( .C1(n21703), .C2(n21412), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n11142), .ZN(n21413) );
  OAI211_X1 U23429 ( .C1(n21415), .C2(n21723), .A(n21414), .B(n21413), .ZN(
        P3_U2841) );
  NAND2_X1 U23430 ( .A1(n21793), .A2(n21656), .ZN(n21592) );
  NOR2_X1 U23431 ( .A1(n11142), .A2(n21416), .ZN(n21418) );
  NAND2_X1 U23432 ( .A1(n21508), .A2(n21625), .ZN(n21423) );
  AOI221_X1 U23433 ( .B1(n21795), .B2(n21423), .C1(n21508), .C2(n21423), .A(
        n21693), .ZN(n21417) );
  AOI211_X1 U23434 ( .C1(n21744), .C2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n21418), .B(n21417), .ZN(n21419) );
  OAI221_X1 U23435 ( .B1(n21421), .B2(n21592), .C1(n21420), .C2(n21489), .A(
        n21419), .ZN(P3_U2862) );
  AOI22_X1 U23436 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21744), .B1(
        n21606), .B2(n21422), .ZN(n21428) );
  AOI211_X1 U23437 ( .C1(n21795), .C2(n21508), .A(n21756), .B(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21426) );
  OAI22_X1 U23438 ( .A1(n21457), .A2(n21424), .B1(n21443), .B2(n21423), .ZN(
        n21425) );
  OAI21_X1 U23439 ( .B1(n21426), .B2(n21425), .A(n21793), .ZN(n21427) );
  OAI211_X1 U23440 ( .C1(n21429), .C2(n11142), .A(n21428), .B(n21427), .ZN(
        P3_U2861) );
  NAND2_X1 U23441 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21445), .ZN(
        n21435) );
  NOR2_X1 U23442 ( .A1(n21776), .A2(n21576), .ZN(n21789) );
  INV_X1 U23443 ( .A(n21789), .ZN(n21617) );
  NOR2_X1 U23444 ( .A1(n21790), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n21728) );
  AOI21_X1 U23445 ( .B1(n21443), .B2(n21617), .A(n21728), .ZN(n21434) );
  NAND2_X1 U23446 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21430) );
  OAI21_X1 U23447 ( .B1(n21430), .B2(n21444), .A(n21446), .ZN(n21432) );
  AOI22_X1 U23448 ( .A1(n21736), .A2(n21432), .B1(n21656), .B2(n21431), .ZN(
        n21433) );
  OAI221_X1 U23449 ( .B1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n21435), .C1(
        n21444), .C2(n21434), .A(n21433), .ZN(n21436) );
  AOI22_X1 U23450 ( .A1(n21739), .A2(n21436), .B1(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n21744), .ZN(n21438) );
  OAI211_X1 U23451 ( .C1(n21439), .C2(n21489), .A(n21438), .B(n21437), .ZN(
        P3_U2860) );
  OAI22_X1 U23452 ( .A1(n11142), .A2(n21440), .B1(n21447), .B2(n21680), .ZN(
        n21441) );
  AOI21_X1 U23453 ( .B1(n21606), .B2(n21442), .A(n21441), .ZN(n21452) );
  NOR2_X1 U23454 ( .A1(n21444), .A2(n21443), .ZN(n21450) );
  AOI22_X1 U23455 ( .A1(n21736), .A2(n21446), .B1(n21445), .B2(n21450), .ZN(
        n21481) );
  INV_X1 U23456 ( .A(n21481), .ZN(n21465) );
  AOI211_X1 U23457 ( .C1(n21736), .C2(n21448), .A(n21728), .B(n21447), .ZN(
        n21449) );
  OAI21_X1 U23458 ( .B1(n21789), .B2(n21450), .A(n21449), .ZN(n21454) );
  OAI211_X1 U23459 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n21465), .A(
        n21793), .B(n21454), .ZN(n21451) );
  OAI211_X1 U23460 ( .C1(n21453), .C2(n21489), .A(n21452), .B(n21451), .ZN(
        P3_U2859) );
  NAND3_X1 U23461 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n21604), .A3(
        n21454), .ZN(n21456) );
  NAND3_X1 U23462 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n21463), .A3(
        n21465), .ZN(n21455) );
  OAI211_X1 U23463 ( .C1(n21458), .C2(n21457), .A(n21456), .B(n21455), .ZN(
        n21460) );
  AOI22_X1 U23464 ( .A1(n21739), .A2(n21460), .B1(n21606), .B2(n21459), .ZN(
        n21462) );
  OAI211_X1 U23465 ( .C1(n21680), .C2(n21463), .A(n21462), .B(n21461), .ZN(
        P3_U2858) );
  NOR2_X1 U23466 ( .A1(n11142), .A2(n21464), .ZN(n21472) );
  NAND4_X1 U23467 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n21739), .A3(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A4(n21465), .ZN(n21469) );
  INV_X1 U23468 ( .A(n21466), .ZN(n21785) );
  OAI21_X1 U23469 ( .B1(n21728), .B2(n21785), .A(n21617), .ZN(n21467) );
  OAI21_X1 U23470 ( .B1(n21468), .B2(n21812), .A(n21467), .ZN(n21485) );
  AOI21_X1 U23471 ( .B1(n21793), .B2(n21485), .A(n21744), .ZN(n21477) );
  AOI21_X1 U23472 ( .B1(n21470), .B2(n21469), .A(n21477), .ZN(n21471) );
  AOI211_X1 U23473 ( .C1(n21606), .C2(n21473), .A(n21472), .B(n21471), .ZN(
        n21474) );
  OAI21_X1 U23474 ( .B1(n21489), .B2(n21475), .A(n21474), .ZN(P3_U2857) );
  OAI22_X1 U23475 ( .A1(n21477), .A2(n21787), .B1(n11142), .B2(n21476), .ZN(
        n21478) );
  AOI21_X1 U23476 ( .B1(n21606), .B2(n21479), .A(n21478), .ZN(n21483) );
  NOR2_X1 U23477 ( .A1(n21481), .A2(n21480), .ZN(n21504) );
  NAND3_X1 U23478 ( .A1(n21793), .A2(n21504), .A3(n21787), .ZN(n21482) );
  OAI211_X1 U23479 ( .C1(n21484), .C2(n21489), .A(n21483), .B(n21482), .ZN(
        P3_U2856) );
  NAND2_X1 U23480 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21504), .ZN(
        n21486) );
  AOI211_X1 U23481 ( .C1(n21604), .C2(n21787), .A(n21786), .B(n21485), .ZN(
        n21499) );
  AOI211_X1 U23482 ( .C1(n21786), .C2(n21486), .A(n21499), .B(n21693), .ZN(
        n21491) );
  OAI22_X1 U23483 ( .A1(n21489), .A2(n21488), .B1(n21592), .B2(n21487), .ZN(
        n21490) );
  NOR2_X1 U23484 ( .A1(n21491), .A2(n21490), .ZN(n21493) );
  NAND2_X1 U23485 ( .A1(n21774), .A2(P3_REIP_REG_7__SCAN_IN), .ZN(n21492) );
  OAI211_X1 U23486 ( .C1(n21680), .C2(n21786), .A(n21493), .B(n21492), .ZN(
        P3_U2855) );
  NAND2_X1 U23487 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21604), .ZN(
        n21498) );
  INV_X1 U23488 ( .A(n21731), .ZN(n21601) );
  AOI22_X1 U23489 ( .A1(n21601), .A2(n21503), .B1(n21656), .B2(n21494), .ZN(
        n21497) );
  NAND4_X1 U23490 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n21504), .A4(n21495), .ZN(
        n21496) );
  OAI211_X1 U23491 ( .C1(n21499), .C2(n21498), .A(n21497), .B(n21496), .ZN(
        n21500) );
  AOI22_X1 U23492 ( .A1(n21739), .A2(n21500), .B1(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n21744), .ZN(n21502) );
  OAI211_X1 U23493 ( .C1(n21770), .C2(n21503), .A(n21502), .B(n21501), .ZN(
        P3_U2854) );
  NAND2_X1 U23494 ( .A1(n21505), .A2(n21504), .ZN(n21562) );
  INV_X1 U23495 ( .A(n21562), .ZN(n21507) );
  OAI21_X1 U23496 ( .B1(n21507), .B2(n21506), .A(n21739), .ZN(n21783) );
  NOR2_X1 U23497 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n21783), .ZN(
        n21516) );
  NAND2_X1 U23498 ( .A1(n21731), .A2(n21811), .ZN(n21734) );
  NOR2_X1 U23499 ( .A1(n21508), .A2(n21775), .ZN(n21788) );
  AOI21_X1 U23500 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n21788), .A(
        n21790), .ZN(n21512) );
  NAND2_X1 U23501 ( .A1(n21601), .A2(n21509), .ZN(n21511) );
  NAND2_X1 U23502 ( .A1(n21736), .A2(n21510), .ZN(n21526) );
  OAI211_X1 U23503 ( .C1(n11416), .C2(n21811), .A(n21511), .B(n21526), .ZN(
        n21797) );
  AOI211_X1 U23504 ( .C1(n21513), .C2(n21734), .A(n21512), .B(n21797), .ZN(
        n21777) );
  NOR2_X1 U23505 ( .A1(n21532), .A2(n21812), .ZN(n21524) );
  AOI21_X1 U23506 ( .B1(n21517), .B2(n21540), .A(n21795), .ZN(n21527) );
  AOI211_X1 U23507 ( .C1(n21576), .C2(n21772), .A(n21524), .B(n21527), .ZN(
        n21514) );
  OAI221_X1 U23508 ( .B1(n21693), .B2(n21777), .C1(n21693), .C2(n21514), .A(
        n21680), .ZN(n21515) );
  AOI22_X1 U23509 ( .A1(n21517), .A2(n21516), .B1(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n21515), .ZN(n21520) );
  INV_X1 U23510 ( .A(n21518), .ZN(n21519) );
  OAI211_X1 U23511 ( .C1(n21521), .C2(n21770), .A(n21520), .B(n21519), .ZN(
        P3_U2851) );
  NAND2_X1 U23512 ( .A1(n21522), .A2(n21788), .ZN(n21539) );
  OAI211_X1 U23513 ( .C1(n21795), .C2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n21790), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21531) );
  INV_X1 U23514 ( .A(n21523), .ZN(n21530) );
  INV_X1 U23515 ( .A(n21524), .ZN(n21525) );
  NAND2_X1 U23516 ( .A1(n21526), .A2(n21525), .ZN(n21542) );
  AOI211_X1 U23517 ( .C1(n21656), .C2(n21528), .A(n21527), .B(n21542), .ZN(
        n21529) );
  OAI21_X1 U23518 ( .B1(n21530), .B2(n21731), .A(n21529), .ZN(n21767) );
  AOI21_X1 U23519 ( .B1(n21539), .B2(n21531), .A(n21767), .ZN(n21537) );
  INV_X1 U23520 ( .A(n21783), .ZN(n21799) );
  AOI22_X1 U23521 ( .A1(n21793), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n21799), .B2(n21532), .ZN(n21536) );
  AOI22_X1 U23522 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n21744), .B1(
        n21801), .B2(n21533), .ZN(n21535) );
  OAI211_X1 U23523 ( .C1(n21537), .C2(n21536), .A(n21535), .B(n21534), .ZN(
        P3_U2850) );
  NOR3_X1 U23524 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n21538), .A3(
        n21562), .ZN(n21547) );
  AOI22_X1 U23525 ( .A1(n21736), .A2(n21762), .B1(n21576), .B2(n21539), .ZN(
        n21765) );
  AOI21_X1 U23526 ( .B1(n21541), .B2(n21540), .A(n21795), .ZN(n21560) );
  AOI211_X1 U23527 ( .C1(n21625), .C2(n21543), .A(n21560), .B(n21542), .ZN(
        n21545) );
  AOI21_X1 U23528 ( .B1(n21765), .B2(n21545), .A(n21544), .ZN(n21546) );
  AOI211_X1 U23529 ( .C1(n21601), .C2(n21548), .A(n21547), .B(n21546), .ZN(
        n21554) );
  OAI22_X1 U23530 ( .A1(n21550), .A2(n21770), .B1(n21592), .B2(n21549), .ZN(
        n21551) );
  AOI211_X1 U23531 ( .C1(n21744), .C2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n21552), .B(n21551), .ZN(n21553) );
  OAI21_X1 U23532 ( .B1(n21554), .B2(n21693), .A(n21553), .ZN(P3_U2848) );
  AND2_X1 U23533 ( .A1(n21567), .A2(n21601), .ZN(n21566) );
  NOR3_X1 U23534 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21811), .A3(
        n21555), .ZN(n21564) );
  AOI21_X1 U23535 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n21790), .A(
        n21556), .ZN(n21559) );
  OAI22_X1 U23536 ( .A1(n21795), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n21557), .B2(n21812), .ZN(n21558) );
  NOR3_X1 U23537 ( .A1(n21560), .A2(n21559), .A3(n21558), .ZN(n21755) );
  NOR3_X1 U23538 ( .A1(n21755), .A2(n21562), .A3(n21561), .ZN(n21563) );
  AOI211_X1 U23539 ( .C1(n21566), .C2(n21565), .A(n21564), .B(n21563), .ZN(
        n21572) );
  AOI22_X1 U23540 ( .A1(n21601), .A2(n21567), .B1(n21656), .B2(n11422), .ZN(
        n21754) );
  OAI221_X1 U23541 ( .B1(n21693), .B2(n21755), .C1(n21693), .C2(n21754), .A(
        n21680), .ZN(n21569) );
  AOI22_X1 U23542 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21569), .B1(
        n21801), .B2(n21568), .ZN(n21571) );
  OAI211_X1 U23543 ( .C1(n21572), .C2(n21693), .A(n21571), .B(n21570), .ZN(
        P3_U2847) );
  AOI22_X1 U23544 ( .A1(n21774), .A2(P3_REIP_REG_22__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n21744), .ZN(n21581) );
  OAI21_X1 U23545 ( .B1(n21574), .B2(n21573), .A(n21633), .ZN(n21678) );
  NOR2_X1 U23546 ( .A1(n21736), .A2(n21776), .ZN(n21779) );
  NAND2_X1 U23547 ( .A1(n21576), .A2(n21575), .ZN(n21577) );
  OAI211_X1 U23548 ( .C1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n21779), .A(
        n21578), .B(n21577), .ZN(n21579) );
  OAI221_X1 U23549 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n21678), 
        .C1(n21679), .C2(n21579), .A(n21739), .ZN(n21580) );
  OAI211_X1 U23550 ( .C1(n21582), .C2(n21770), .A(n21581), .B(n21580), .ZN(
        P3_U2840) );
  AND2_X1 U23551 ( .A1(n21583), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n21584) );
  INV_X1 U23552 ( .A(n21728), .ZN(n21616) );
  AOI21_X1 U23553 ( .B1(n21584), .B2(n21616), .A(n21789), .ZN(n21685) );
  AOI21_X1 U23554 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n21585), .A(
        n21812), .ZN(n21687) );
  NOR3_X1 U23555 ( .A1(n21685), .A2(n21687), .A3(n21586), .ZN(n21587) );
  OAI21_X1 U23556 ( .B1(n21756), .B2(n21587), .A(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21603) );
  OAI21_X1 U23557 ( .B1(n21633), .B2(n21588), .A(n21598), .ZN(n21589) );
  AOI22_X1 U23558 ( .A1(n21601), .A2(n21590), .B1(n21603), .B2(n21589), .ZN(
        n21593) );
  OAI22_X1 U23559 ( .A1(n21593), .A2(n21693), .B1(n21592), .B2(n21591), .ZN(
        n21594) );
  AOI21_X1 U23560 ( .B1(n21801), .B2(n21595), .A(n21594), .ZN(n21597) );
  NAND2_X1 U23561 ( .A1(n21774), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n21596) );
  OAI211_X1 U23562 ( .C1(n21680), .C2(n21598), .A(n21597), .B(n21596), .ZN(
        P3_U2837) );
  NAND4_X1 U23563 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n21600), .A3(
        n21678), .A4(n21599), .ZN(n21612) );
  NAND2_X1 U23564 ( .A1(n21601), .A2(n21631), .ZN(n21614) );
  INV_X1 U23565 ( .A(n21614), .ZN(n21602) );
  AOI21_X1 U23566 ( .B1(n21604), .B2(n21603), .A(n21602), .ZN(n21607) );
  NAND2_X1 U23567 ( .A1(n21606), .A2(n21605), .ZN(n21619) );
  OAI211_X1 U23568 ( .C1(n21607), .C2(n21693), .A(n21619), .B(n21680), .ZN(
        n21609) );
  AOI22_X1 U23569 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n21609), .B1(
        n21801), .B2(n21608), .ZN(n21611) );
  OAI211_X1 U23570 ( .C1(n21693), .C2(n21612), .A(n21611), .B(n21610), .ZN(
        P3_U2836) );
  NAND2_X1 U23571 ( .A1(n21613), .A2(n21678), .ZN(n21666) );
  NAND4_X1 U23572 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n21616), .A3(
        n21615), .A4(n21614), .ZN(n21618) );
  OAI221_X1 U23573 ( .B1(n21618), .B2(n21617), .C1(n21618), .C2(n21657), .A(
        n21739), .ZN(n21620) );
  AOI22_X1 U23574 ( .A1(n21666), .A2(n21665), .B1(n21620), .B2(n21619), .ZN(
        n21621) );
  AOI21_X1 U23575 ( .B1(n21801), .B2(n21622), .A(n21621), .ZN(n21624) );
  OAI211_X1 U23576 ( .C1(n21680), .C2(n21665), .A(n21624), .B(n21623), .ZN(
        P3_U2835) );
  INV_X1 U23577 ( .A(n21625), .ZN(n21717) );
  OAI22_X1 U23578 ( .A1(n21627), .A2(n21731), .B1(n21626), .B2(n21811), .ZN(
        n21647) );
  AOI21_X1 U23579 ( .B1(n21736), .B2(n21665), .A(n21647), .ZN(n21628) );
  OAI211_X1 U23580 ( .C1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n21717), .A(
        n21629), .B(n21628), .ZN(n21630) );
  AOI21_X1 U23581 ( .B1(n21793), .B2(n21630), .A(n21744), .ZN(n21642) );
  OAI22_X1 U23582 ( .A1(n21633), .A2(n21632), .B1(n21731), .B2(n21631), .ZN(
        n21634) );
  AOI21_X1 U23583 ( .B1(n21656), .B2(n21635), .A(n21634), .ZN(n21645) );
  NOR3_X1 U23584 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n21645), .A3(
        n21636), .ZN(n21638) );
  AOI22_X1 U23585 ( .A1(n21739), .A2(n21638), .B1(n21801), .B2(n21637), .ZN(
        n21640) );
  NAND2_X1 U23586 ( .A1(n21774), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n21639) );
  OAI211_X1 U23587 ( .C1(n21642), .C2(n21641), .A(n21640), .B(n21639), .ZN(
        P3_U2833) );
  AOI22_X1 U23588 ( .A1(n21774), .A2(P3_REIP_REG_30__SCAN_IN), .B1(n21744), 
        .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21650) );
  OAI21_X1 U23589 ( .B1(n21645), .B2(n21644), .A(n21643), .ZN(n21646) );
  OAI211_X1 U23590 ( .C1(n21648), .C2(n21647), .A(n21793), .B(n21646), .ZN(
        n21649) );
  OAI211_X1 U23591 ( .C1(n21651), .C2(n21770), .A(n21650), .B(n21649), .ZN(
        P3_U2832) );
  INV_X1 U23592 ( .A(n21657), .ZN(n21658) );
  OAI22_X1 U23593 ( .A1(n21795), .A2(n21658), .B1(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n21779), .ZN(n21659) );
  NOR3_X1 U23594 ( .A1(n21744), .A2(n21660), .A3(n21659), .ZN(n21663) );
  OR2_X1 U23595 ( .A1(n21661), .A2(n21731), .ZN(n21662) );
  NAND3_X1 U23596 ( .A1(n21664), .A2(n21663), .A3(n21662), .ZN(n21672) );
  OAI22_X1 U23597 ( .A1(n21668), .A2(n21667), .B1(n21666), .B2(n21665), .ZN(
        n21669) );
  NAND2_X1 U23598 ( .A1(n21669), .A2(n21793), .ZN(n21670) );
  NAND2_X1 U23599 ( .A1(n21672), .A2(n21671), .ZN(n21677) );
  OR3_X1 U23600 ( .A1(n21674), .A2(n21770), .A3(n21673), .ZN(n21675) );
  OAI221_X1 U23601 ( .B1(n21774), .B2(n21677), .C1(n11142), .C2(n21676), .A(
        n21675), .ZN(P3_U2834) );
  INV_X1 U23602 ( .A(n21678), .ZN(n21694) );
  NOR2_X1 U23603 ( .A1(n21694), .A2(n21679), .ZN(n21681) );
  AOI21_X1 U23604 ( .B1(n21681), .B2(n21680), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21691) );
  OAI22_X1 U23605 ( .A1(n21683), .A2(n21811), .B1(n21682), .B2(n21731), .ZN(
        n21684) );
  NOR3_X1 U23606 ( .A1(n21744), .A2(n21685), .A3(n21684), .ZN(n21697) );
  NAND2_X1 U23607 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n21697), .ZN(
        n21686) );
  OAI21_X1 U23608 ( .B1(n21687), .B2(n21686), .A(n11142), .ZN(n21695) );
  AOI21_X1 U23609 ( .B1(n21689), .B2(n21801), .A(n21688), .ZN(n21690) );
  OAI21_X1 U23610 ( .B1(n21691), .B2(n21695), .A(n21690), .ZN(P3_U2839) );
  NOR4_X1 U23611 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n21694), .A3(
        n21693), .A4(n21692), .ZN(n21699) );
  AOI211_X1 U23612 ( .C1(n21756), .C2(n21697), .A(n21696), .B(n21695), .ZN(
        n21698) );
  AOI211_X1 U23613 ( .C1(n21801), .C2(n21700), .A(n21699), .B(n21698), .ZN(
        n21701) );
  OAI21_X1 U23614 ( .B1(n11142), .B2(n21702), .A(n21701), .ZN(P3_U2838) );
  INV_X1 U23615 ( .A(n21703), .ZN(n21710) );
  INV_X1 U23616 ( .A(n21704), .ZN(n21709) );
  OAI22_X1 U23617 ( .A1(n21706), .A2(n21731), .B1(n21705), .B2(n21811), .ZN(
        n21707) );
  INV_X1 U23618 ( .A(n21707), .ZN(n21708) );
  NAND3_X1 U23619 ( .A1(n21710), .A2(n21709), .A3(n21708), .ZN(n21711) );
  NAND2_X1 U23620 ( .A1(n11142), .A2(n21711), .ZN(n21715) );
  AOI22_X1 U23621 ( .A1(n14606), .A2(P3_REIP_REG_19__SCAN_IN), .B1(n21801), 
        .B2(n21712), .ZN(n21713) );
  OAI221_X1 U23622 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n21723), 
        .C1(n21714), .C2(n21715), .A(n21713), .ZN(P3_U2843) );
  NAND2_X1 U23623 ( .A1(n21714), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n21716) );
  OAI21_X1 U23624 ( .B1(n21717), .B2(n21716), .A(n21715), .ZN(n21720) );
  INV_X1 U23625 ( .A(n21718), .ZN(n21719) );
  AOI22_X1 U23626 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n21720), .B1(
        n21801), .B2(n21719), .ZN(n21722) );
  OAI211_X1 U23627 ( .C1(n21724), .C2(n21723), .A(n21722), .B(n21721), .ZN(
        P3_U2842) );
  AOI22_X1 U23628 ( .A1(n21774), .A2(P3_REIP_REG_18__SCAN_IN), .B1(n21753), 
        .B2(n21726), .ZN(n21742) );
  NOR3_X1 U23629 ( .A1(n21728), .A2(n21727), .A3(n21752), .ZN(n21738) );
  OAI211_X1 U23630 ( .C1(n21732), .C2(n21731), .A(n21730), .B(n21729), .ZN(
        n21733) );
  AOI22_X1 U23631 ( .A1(n21736), .A2(n21735), .B1(n21734), .B2(n21733), .ZN(
        n21737) );
  OAI21_X1 U23632 ( .B1(n21789), .B2(n21738), .A(n21737), .ZN(n21745) );
  OAI21_X1 U23633 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n21789), .A(
        n21739), .ZN(n21740) );
  OAI211_X1 U23634 ( .C1(n21745), .C2(n21740), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B(n11142), .ZN(n21741) );
  OAI211_X1 U23635 ( .C1(n21743), .C2(n21770), .A(n21742), .B(n21741), .ZN(
        P3_U2844) );
  AOI21_X1 U23636 ( .B1(n21793), .B2(n21745), .A(n21744), .ZN(n21751) );
  AOI22_X1 U23637 ( .A1(n21801), .A2(n21747), .B1(n21753), .B2(n21746), .ZN(
        n21749) );
  OAI211_X1 U23638 ( .C1(n21751), .C2(n21750), .A(n21749), .B(n21748), .ZN(
        P3_U2845) );
  AOI22_X1 U23639 ( .A1(n21774), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n21753), 
        .B2(n21752), .ZN(n21759) );
  OAI211_X1 U23640 ( .C1(n21756), .C2(n21755), .A(n21793), .B(n21754), .ZN(
        n21757) );
  NAND3_X1 U23641 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n11142), .A3(
        n21757), .ZN(n21758) );
  OAI211_X1 U23642 ( .C1(n21770), .C2(n21760), .A(n21759), .B(n21758), .ZN(
        P3_U2846) );
  AOI22_X1 U23643 ( .A1(n21774), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n21799), 
        .B2(n21761), .ZN(n21769) );
  OAI21_X1 U23644 ( .B1(n21763), .B2(n21762), .A(n21776), .ZN(n21764) );
  NAND3_X1 U23645 ( .A1(n21793), .A2(n21765), .A3(n21764), .ZN(n21766) );
  OAI211_X1 U23646 ( .C1(n21767), .C2(n21766), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n11142), .ZN(n21768) );
  OAI211_X1 U23647 ( .C1(n21771), .C2(n21770), .A(n21769), .B(n21768), .ZN(
        P3_U2849) );
  NAND2_X1 U23648 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n21772), .ZN(
        n21784) );
  AOI22_X1 U23649 ( .A1(n21774), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n21801), 
        .B2(n21773), .ZN(n21782) );
  AOI21_X1 U23650 ( .B1(n21776), .B2(n21775), .A(n21798), .ZN(n21778) );
  OAI211_X1 U23651 ( .C1(n21779), .C2(n21778), .A(n21793), .B(n21777), .ZN(
        n21780) );
  NAND3_X1 U23652 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n11142), .A3(
        n21780), .ZN(n21781) );
  OAI211_X1 U23653 ( .C1(n21784), .C2(n21783), .A(n21782), .B(n21781), .ZN(
        P3_U2852) );
  NOR3_X1 U23654 ( .A1(n21787), .A2(n21786), .A3(n21785), .ZN(n21794) );
  AOI211_X1 U23655 ( .C1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n21790), .A(
        n21789), .B(n21788), .ZN(n21791) );
  INV_X1 U23656 ( .A(n21791), .ZN(n21792) );
  OAI211_X1 U23657 ( .C1(n21795), .C2(n21794), .A(n21793), .B(n21792), .ZN(
        n21796) );
  OAI21_X1 U23658 ( .B1(n21797), .B2(n21796), .A(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21804) );
  AOI22_X1 U23659 ( .A1(n21801), .A2(n21800), .B1(n21799), .B2(n21798), .ZN(
        n21802) );
  OAI221_X1 U23660 ( .B1(n21774), .B2(n21804), .C1(n11142), .C2(n21803), .A(
        n21802), .ZN(P3_U2853) );
  NAND2_X1 U23661 ( .A1(n22341), .A2(n21805), .ZN(n21861) );
  INV_X1 U23662 ( .A(n21806), .ZN(n21850) );
  AOI22_X1 U23663 ( .A1(n21809), .A2(n21808), .B1(n21817), .B2(n21807), .ZN(
        n21810) );
  OAI221_X1 U23664 ( .B1(n21813), .B2(n21812), .C1(n21813), .C2(n21811), .A(
        n21810), .ZN(n21870) );
  INV_X1 U23665 ( .A(n21814), .ZN(n21815) );
  NOR3_X1 U23666 ( .A1(n21817), .A2(n21816), .A3(n21815), .ZN(n21869) );
  OAI21_X1 U23667 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(P3_MORE_REG_SCAN_IN), .A(
        n21869), .ZN(n21819) );
  OAI211_X1 U23668 ( .C1(n21826), .C2(n21820), .A(n21819), .B(n21818), .ZN(
        n21843) );
  INV_X1 U23669 ( .A(n21826), .ZN(n21822) );
  AOI22_X1 U23670 ( .A1(n21822), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n21821), .B2(n21826), .ZN(n21841) );
  OAI22_X1 U23671 ( .A1(n21826), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n21823), .B2(n21822), .ZN(n21824) );
  INV_X1 U23672 ( .A(n21824), .ZN(n21836) );
  NOR3_X1 U23673 ( .A1(n21828), .A2(n21825), .A3(n21827), .ZN(n21832) );
  OAI221_X1 U23674 ( .B1(n21829), .B2(n21828), .C1(n21829), .C2(n21827), .A(
        n21826), .ZN(n21831) );
  OAI21_X1 U23675 ( .B1(n21832), .B2(n21831), .A(n21830), .ZN(n21835) );
  AND2_X1 U23676 ( .A1(n21836), .A2(n21835), .ZN(n21833) );
  OAI221_X1 U23677 ( .B1(n21836), .B2(n21835), .C1(n21834), .C2(n21833), .A(
        n21838), .ZN(n21840) );
  AOI21_X1 U23678 ( .B1(n21838), .B2(n21837), .A(n21836), .ZN(n21839) );
  AOI222_X1 U23679 ( .A1(n21841), .A2(n21840), .B1(n21841), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n21840), .C2(n21839), .ZN(
        n21842) );
  NOR4_X1 U23680 ( .A1(n21844), .A2(n21870), .A3(n21843), .A4(n21842), .ZN(
        n21867) );
  OAI211_X1 U23681 ( .C1(n21847), .C2(n21846), .A(n21845), .B(n21867), .ZN(
        n21854) );
  OAI21_X1 U23682 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n22352), .A(n21854), 
        .ZN(n21859) );
  OR3_X1 U23683 ( .A1(n21848), .A2(n21857), .A3(n21859), .ZN(n21849) );
  NAND4_X1 U23684 ( .A1(n21851), .A2(n21861), .A3(n21850), .A4(n21849), .ZN(
        P3_U2997) );
  OAI211_X1 U23685 ( .C1(n21855), .C2(n21854), .A(n21853), .B(n21852), .ZN(
        P3_U3282) );
  NOR2_X1 U23686 ( .A1(n21857), .A2(n21856), .ZN(n21858) );
  AOI221_X1 U23687 ( .B1(n21860), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n21859), 
        .C2(P3_STATE2_REG_0__SCAN_IN), .A(n21858), .ZN(n21866) );
  OAI211_X1 U23688 ( .C1(n21864), .C2(n21863), .A(n21862), .B(n21861), .ZN(
        n21865) );
  OAI211_X1 U23689 ( .C1(n21867), .C2(n21868), .A(n21866), .B(n21865), .ZN(
        P3_U2996) );
  NOR2_X1 U23690 ( .A1(n21869), .A2(n21868), .ZN(n21873) );
  MUX2_X1 U23691 ( .A(P3_MORE_REG_SCAN_IN), .B(n21870), .S(n21873), .Z(
        P3_U3295) );
  OAI21_X1 U23692 ( .B1(n21873), .B2(n21872), .A(n21871), .ZN(P3_U2637) );
  AOI211_X1 U23693 ( .C1(n21877), .C2(n21876), .A(n21875), .B(n21874), .ZN(
        n21885) );
  INV_X1 U23694 ( .A(n21878), .ZN(n21881) );
  INV_X1 U23695 ( .A(n21879), .ZN(n21880) );
  OAI211_X1 U23696 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n21881), .A(n21880), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n21882) );
  AOI21_X1 U23697 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n21882), .A(n22278), 
        .ZN(n21884) );
  NAND2_X1 U23698 ( .A1(n21885), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n21883) );
  OAI21_X1 U23699 ( .B1(n21885), .B2(n21884), .A(n21883), .ZN(P1_U3485) );
  NOR2_X1 U23700 ( .A1(n21886), .A2(n21907), .ZN(n22006) );
  AOI21_X1 U23701 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n21887), .A(
        n21892), .ZN(n21891) );
  OAI21_X1 U23702 ( .B1(n21889), .B2(n21888), .A(n22062), .ZN(n21890) );
  NOR3_X1 U23703 ( .A1(n22006), .A2(n21891), .A3(n21890), .ZN(n21898) );
  AOI221_X1 U23704 ( .B1(n22014), .B2(n21899), .C1(n21892), .C2(n21899), .A(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n21893) );
  AOI21_X1 U23705 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n22052), .A(n21893), 
        .ZN(n21897) );
  AOI22_X1 U23706 ( .A1(n22056), .A2(n21895), .B1(n22053), .B2(n21894), .ZN(
        n21896) );
  OAI211_X1 U23707 ( .C1(n21898), .C2(n21901), .A(n21897), .B(n21896), .ZN(
        P1_U3018) );
  OAI21_X1 U23708 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n21899), .A(
        n21898), .ZN(n21900) );
  AOI22_X1 U23709 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n22052), .B1(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n21900), .ZN(n21905) );
  NOR4_X1 U23710 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n21901), .A3(
        n16414), .A4(n16401), .ZN(n21902) );
  AOI22_X1 U23711 ( .A1(n22053), .A2(n21903), .B1(n21902), .B2(n21999), .ZN(
        n21904) );
  OAI211_X1 U23712 ( .C1(n22033), .C2(n21906), .A(n21905), .B(n21904), .ZN(
        P1_U3017) );
  NOR2_X1 U23713 ( .A1(n21907), .A2(n21924), .ZN(n21921) );
  AOI21_X1 U23714 ( .B1(n22052), .B2(P1_REIP_REG_2__SCAN_IN), .A(n21921), .ZN(
        n21918) );
  NOR2_X1 U23715 ( .A1(n21908), .A2(n22064), .ZN(n21910) );
  AOI22_X1 U23716 ( .A1(n21910), .A2(n22007), .B1(n22064), .B2(n21909), .ZN(
        n21911) );
  NAND2_X1 U23717 ( .A1(n21911), .A2(n22002), .ZN(n21912) );
  NAND2_X1 U23718 ( .A1(n21912), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n21914) );
  OR3_X1 U23719 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n22064), .A3(
        n22012), .ZN(n21913) );
  OAI211_X1 U23720 ( .C1(n21915), .C2(n22031), .A(n21914), .B(n21913), .ZN(
        n21916) );
  INV_X1 U23721 ( .A(n21916), .ZN(n21917) );
  OAI211_X1 U23722 ( .C1(n22033), .C2(n21919), .A(n21918), .B(n21917), .ZN(
        P1_U3029) );
  INV_X1 U23723 ( .A(n21923), .ZN(n21920) );
  OAI21_X1 U23724 ( .B1(n22004), .B2(n21920), .A(n22002), .ZN(n21957) );
  NOR2_X1 U23725 ( .A1(n21921), .A2(n21957), .ZN(n21938) );
  OAI22_X1 U23726 ( .A1(n22077), .A2(n22033), .B1(n22049), .B2(n21922), .ZN(
        n21927) );
  NOR2_X1 U23727 ( .A1(n21923), .A2(n22012), .ZN(n21944) );
  AND2_X1 U23728 ( .A1(n22007), .A2(n21924), .ZN(n21925) );
  AOI211_X1 U23729 ( .C1(n21930), .C2(n21937), .A(n21956), .B(n21942), .ZN(
        n21926) );
  AOI211_X1 U23730 ( .C1(n21928), .C2(n22053), .A(n21927), .B(n21926), .ZN(
        n21929) );
  OAI21_X1 U23731 ( .B1(n21938), .B2(n21930), .A(n21929), .ZN(P1_U3027) );
  AOI22_X1 U23732 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n22052), .B1(n22056), 
        .B2(n21931), .ZN(n21936) );
  INV_X1 U23733 ( .A(n21932), .ZN(n21934) );
  AOI22_X1 U23734 ( .A1(n21934), .A2(n22053), .B1(n21937), .B2(n21933), .ZN(
        n21935) );
  OAI211_X1 U23735 ( .C1(n21938), .C2(n21937), .A(n21936), .B(n21935), .ZN(
        P1_U3028) );
  NAND2_X1 U23736 ( .A1(n21939), .A2(n21942), .ZN(n21955) );
  INV_X1 U23737 ( .A(n21955), .ZN(n21943) );
  AOI21_X1 U23738 ( .B1(n22007), .B2(n21940), .A(n21957), .ZN(n21941) );
  OAI21_X1 U23739 ( .B1(n22004), .B2(n21942), .A(n21941), .ZN(n21951) );
  AOI21_X1 U23740 ( .B1(n21944), .B2(n21943), .A(n21951), .ZN(n21950) );
  AOI22_X1 U23741 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n22052), .B1(n22056), 
        .B2(n22105), .ZN(n21948) );
  NOR2_X1 U23742 ( .A1(n21956), .A2(n21945), .ZN(n21962) );
  AOI22_X1 U23743 ( .A1(n21946), .A2(n22053), .B1(n21962), .B2(n21949), .ZN(
        n21947) );
  OAI211_X1 U23744 ( .C1(n21950), .C2(n21949), .A(n21948), .B(n21947), .ZN(
        P1_U3025) );
  AOI22_X1 U23745 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n22052), .B1(n22056), 
        .B2(n22091), .ZN(n21954) );
  AOI22_X1 U23746 ( .A1(n21952), .A2(n22053), .B1(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n21951), .ZN(n21953) );
  OAI211_X1 U23747 ( .C1(n21956), .C2(n21955), .A(n21954), .B(n21953), .ZN(
        P1_U3026) );
  INV_X1 U23748 ( .A(n22002), .ZN(n21959) );
  OAI22_X1 U23749 ( .A1(n22051), .A2(n21959), .B1(n21958), .B2(n21957), .ZN(
        n21967) );
  AOI222_X1 U23750 ( .A1(n21961), .A2(n22053), .B1(n22056), .B2(n21960), .C1(
        n22052), .C2(P1_REIP_REG_7__SCAN_IN), .ZN(n21963) );
  NAND2_X1 U23751 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21962), .ZN(
        n21979) );
  OR2_X1 U23752 ( .A1(n21979), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n21968) );
  OAI211_X1 U23753 ( .C1(n21965), .C2(n21967), .A(n21963), .B(n21968), .ZN(
        P1_U3024) );
  INV_X1 U23754 ( .A(n21964), .ZN(n21971) );
  NOR3_X1 U23755 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21965), .A3(
        n21979), .ZN(n21970) );
  AOI21_X1 U23756 ( .B1(n21968), .B2(n21967), .A(n21966), .ZN(n21969) );
  AOI211_X1 U23757 ( .C1(n21971), .C2(n22053), .A(n21970), .B(n21969), .ZN(
        n21973) );
  NAND2_X1 U23758 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n22052), .ZN(n21972) );
  OAI211_X1 U23759 ( .C1(n22033), .C2(n22129), .A(n21973), .B(n21972), .ZN(
        P1_U3023) );
  OAI21_X1 U23760 ( .B1(n22004), .B2(n21974), .A(n22002), .ZN(n21975) );
  AOI21_X1 U23761 ( .B1(n22007), .B2(n21976), .A(n21975), .ZN(n21994) );
  INV_X1 U23762 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21984) );
  AOI22_X1 U23763 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n22052), .B1(n22056), 
        .B2(n21977), .ZN(n21983) );
  INV_X1 U23764 ( .A(n21978), .ZN(n21981) );
  NOR2_X1 U23765 ( .A1(n21980), .A2(n21979), .ZN(n21990) );
  AOI22_X1 U23766 ( .A1(n21981), .A2(n22053), .B1(n21990), .B2(n21984), .ZN(
        n21982) );
  OAI211_X1 U23767 ( .C1(n21994), .C2(n21984), .A(n21983), .B(n21982), .ZN(
        P1_U3022) );
  NOR2_X1 U23768 ( .A1(n21985), .A2(n22033), .ZN(n21986) );
  AOI211_X1 U23769 ( .C1(n21988), .C2(n22053), .A(n21987), .B(n21986), .ZN(
        n21992) );
  OAI211_X1 U23770 ( .C1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n21990), .B(n21989), .ZN(
        n21991) );
  OAI211_X1 U23771 ( .C1(n21994), .C2(n21993), .A(n21992), .B(n21991), .ZN(
        P1_U3021) );
  NOR2_X1 U23772 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n22012), .ZN(
        n21998) );
  OAI22_X1 U23773 ( .A1(n21995), .A2(n22031), .B1(n22033), .B2(n22149), .ZN(
        n21996) );
  AOI221_X1 U23774 ( .B1(n21998), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), 
        .C1(n21997), .C2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n21996), .ZN(
        n22001) );
  NAND3_X1 U23775 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16401), .A3(
        n21999), .ZN(n22000) );
  OAI211_X1 U23776 ( .C1(n22049), .C2(n22151), .A(n22001), .B(n22000), .ZN(
        P1_U3019) );
  NOR2_X1 U23777 ( .A1(n22011), .A2(n22014), .ZN(n22003) );
  OAI21_X1 U23778 ( .B1(n22004), .B2(n22003), .A(n22002), .ZN(n22005) );
  AOI211_X1 U23779 ( .C1(n22007), .C2(n22011), .A(n22006), .B(n22005), .ZN(
        n22035) );
  OAI22_X1 U23780 ( .A1(n22008), .A2(n22049), .B1(n22015), .B2(n22035), .ZN(
        n22009) );
  INV_X1 U23781 ( .A(n22009), .ZN(n22017) );
  INV_X1 U23782 ( .A(n22010), .ZN(n22163) );
  AOI221_X1 U23783 ( .B1(n22014), .B2(n22013), .C1(n22012), .C2(n22013), .A(
        n22011), .ZN(n22039) );
  AOI22_X1 U23784 ( .A1(n22163), .A2(n22056), .B1(n22015), .B2(n22039), .ZN(
        n22016) );
  OAI211_X1 U23785 ( .C1(n22031), .C2(n22018), .A(n22017), .B(n22016), .ZN(
        P1_U3016) );
  INV_X1 U23786 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n22187) );
  OAI21_X1 U23787 ( .B1(n22023), .B2(n22019), .A(n22035), .ZN(n22027) );
  OAI22_X1 U23788 ( .A1(n22020), .A2(n22031), .B1(n22033), .B2(n22193), .ZN(
        n22021) );
  AOI21_X1 U23789 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n22027), .A(
        n22021), .ZN(n22025) );
  NAND3_X1 U23790 ( .A1(n22023), .A2(n22022), .A3(n22039), .ZN(n22024) );
  OAI211_X1 U23791 ( .C1(n22049), .C2(n22187), .A(n22025), .B(n22024), .ZN(
        P1_U3013) );
  AOI22_X1 U23792 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n22052), .B1(n22056), 
        .B2(n22026), .ZN(n22030) );
  OAI221_X1 U23793 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n22028), 
        .C1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n22039), .A(n22027), .ZN(
        n22029) );
  OAI211_X1 U23794 ( .C1(n22032), .C2(n22031), .A(n22030), .B(n22029), .ZN(
        P1_U3014) );
  OAI22_X1 U23795 ( .A1(n22035), .A2(n22034), .B1(n22033), .B2(n22183), .ZN(
        n22036) );
  AOI21_X1 U23796 ( .B1(n22053), .B2(n22037), .A(n22036), .ZN(n22041) );
  OAI211_X1 U23797 ( .C1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A(n22039), .B(n22038), .ZN(
        n22040) );
  OAI211_X1 U23798 ( .C1(n22049), .C2(n22176), .A(n22041), .B(n22040), .ZN(
        P1_U3015) );
  INV_X1 U23799 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n22203) );
  AOI22_X1 U23800 ( .A1(n22042), .A2(n22053), .B1(n22056), .B2(n22198), .ZN(
        n22048) );
  OAI22_X1 U23801 ( .A1(n22045), .A2(n22044), .B1(n22043), .B2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n22046) );
  INV_X1 U23802 ( .A(n22046), .ZN(n22047) );
  OAI211_X1 U23803 ( .C1(n22049), .C2(n22203), .A(n22048), .B(n22047), .ZN(
        P1_U3012) );
  NAND3_X1 U23804 ( .A1(n22064), .A2(n22051), .A3(n22050), .ZN(n22060) );
  NAND2_X1 U23805 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(n22052), .ZN(n22059) );
  NAND3_X1 U23806 ( .A1(n15071), .A2(n22054), .A3(n22053), .ZN(n22058) );
  NAND2_X1 U23807 ( .A1(n22056), .A2(n22055), .ZN(n22057) );
  AND4_X1 U23808 ( .A1(n22060), .A2(n22059), .A3(n22058), .A4(n22057), .ZN(
        n22061) );
  OAI221_X1 U23809 ( .B1(n22064), .B2(n22063), .C1(n22064), .C2(n22062), .A(
        n22061), .ZN(P1_U3030) );
  INV_X1 U23810 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n22066) );
  AOI22_X1 U23811 ( .A1(n22427), .A2(n22074), .B1(n22235), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n22065) );
  OAI21_X1 U23812 ( .B1(n22104), .B2(n22066), .A(n22065), .ZN(n22067) );
  AOI21_X1 U23813 ( .B1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n22244), .A(
        n22067), .ZN(n22068) );
  OAI21_X1 U23814 ( .B1(n22085), .B2(n22069), .A(n22068), .ZN(n22070) );
  AOI21_X1 U23815 ( .B1(n22260), .B2(n22071), .A(n22070), .ZN(n22073) );
  OR2_X1 U23816 ( .A1(n22220), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n22072) );
  OAI211_X1 U23817 ( .C1(n22267), .C2(n15028), .A(n22073), .B(n22072), .ZN(
        P1_U2839) );
  AOI22_X1 U23818 ( .A1(n22075), .A2(n22074), .B1(n22235), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n22076) );
  OAI21_X1 U23819 ( .B1(n22267), .B2(n22077), .A(n22076), .ZN(n22078) );
  AOI211_X1 U23820 ( .C1(n22244), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n22197), .B(n22078), .ZN(n22089) );
  INV_X1 U23821 ( .A(n22096), .ZN(n22079) );
  NAND2_X1 U23822 ( .A1(n22236), .A2(n22079), .ZN(n22080) );
  NAND2_X1 U23823 ( .A1(n22104), .A2(n22080), .ZN(n22098) );
  INV_X1 U23824 ( .A(n22098), .ZN(n22084) );
  INV_X1 U23825 ( .A(n22081), .ZN(n22082) );
  AOI21_X1 U23826 ( .B1(n22236), .B2(n22082), .A(P1_REIP_REG_4__SCAN_IN), .ZN(
        n22083) );
  OAI22_X1 U23827 ( .A1(n22086), .A2(n22085), .B1(n22084), .B2(n22083), .ZN(
        n22087) );
  INV_X1 U23828 ( .A(n22087), .ZN(n22088) );
  OAI211_X1 U23829 ( .C1(n22090), .C2(n22251), .A(n22089), .B(n22088), .ZN(
        P1_U2836) );
  NOR2_X1 U23830 ( .A1(n22220), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n22097) );
  INV_X1 U23831 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n22094) );
  AOI22_X1 U23832 ( .A1(n22091), .A2(n22199), .B1(n22235), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n22093) );
  OAI211_X1 U23833 ( .C1(n22256), .C2(n22094), .A(n22093), .B(n22092), .ZN(
        n22095) );
  AOI21_X1 U23834 ( .B1(n22097), .B2(n22096), .A(n22095), .ZN(n22102) );
  AOI22_X1 U23835 ( .A1(n22100), .A2(n22099), .B1(P1_REIP_REG_5__SCAN_IN), 
        .B2(n22098), .ZN(n22101) );
  OAI211_X1 U23836 ( .C1(n22103), .C2(n22251), .A(n22102), .B(n22101), .ZN(
        P1_U2835) );
  INV_X1 U23837 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n22110) );
  OAI21_X1 U23838 ( .B1(n22116), .B2(n22220), .A(n22104), .ZN(n22124) );
  AOI22_X1 U23839 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n22124), .B1(n22199), 
        .B2(n22105), .ZN(n22109) );
  NOR3_X1 U23840 ( .A1(n22220), .A2(n22116), .A3(n22106), .ZN(n22107) );
  AOI211_X1 U23841 ( .C1(n22235), .C2(P1_EBX_REG_6__SCAN_IN), .A(n22107), .B(
        n22197), .ZN(n22108) );
  OAI211_X1 U23842 ( .C1(n22110), .C2(n22256), .A(n22109), .B(n22108), .ZN(
        n22111) );
  AOI21_X1 U23843 ( .B1(n22112), .B2(n22262), .A(n22111), .ZN(n22113) );
  OAI21_X1 U23844 ( .B1(n22114), .B2(n22251), .A(n22113), .ZN(P1_U2834) );
  NAND2_X1 U23845 ( .A1(n22235), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n22118) );
  INV_X1 U23846 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n22115) );
  NAND3_X1 U23847 ( .A1(n22236), .A2(n22116), .A3(n22115), .ZN(n22117) );
  OAI211_X1 U23848 ( .C1(n22119), .C2(n22267), .A(n22118), .B(n22117), .ZN(
        n22120) );
  AOI211_X1 U23849 ( .C1(n22244), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n22120), .B(n22197), .ZN(n22121) );
  OAI21_X1 U23850 ( .B1(n22122), .B2(n22246), .A(n22121), .ZN(n22123) );
  AOI21_X1 U23851 ( .B1(P1_REIP_REG_7__SCAN_IN), .B2(n22124), .A(n22123), .ZN(
        n22125) );
  OAI21_X1 U23852 ( .B1(n22126), .B2(n22251), .A(n22125), .ZN(P1_U2833) );
  NOR2_X1 U23853 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n22127), .ZN(n22137) );
  OAI22_X1 U23854 ( .A1(n22129), .A2(n22267), .B1(n22254), .B2(n22128), .ZN(
        n22130) );
  AOI211_X1 U23855 ( .C1(n22244), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n22197), .B(n22130), .ZN(n22135) );
  INV_X1 U23856 ( .A(n22131), .ZN(n22132) );
  AOI22_X1 U23857 ( .A1(n22133), .A2(n22262), .B1(n22132), .B2(n22260), .ZN(
        n22134) );
  OAI211_X1 U23858 ( .C1(n22137), .C2(n22136), .A(n22135), .B(n22134), .ZN(
        P1_U2832) );
  OAI22_X1 U23859 ( .A1(n22256), .A2(n22139), .B1(n22254), .B2(n22138), .ZN(
        n22140) );
  AOI211_X1 U23860 ( .C1(P1_REIP_REG_11__SCAN_IN), .C2(n22141), .A(n22197), 
        .B(n22140), .ZN(n22146) );
  OAI22_X1 U23861 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n22152), .B1(n22142), 
        .B2(n22267), .ZN(n22143) );
  AOI21_X1 U23862 ( .B1(n22262), .B2(n22144), .A(n22143), .ZN(n22145) );
  OAI211_X1 U23863 ( .C1(n22147), .C2(n22251), .A(n22146), .B(n22145), .ZN(
        P1_U2829) );
  OAI22_X1 U23864 ( .A1(n22149), .A2(n22267), .B1(n22254), .B2(n22148), .ZN(
        n22150) );
  AOI211_X1 U23865 ( .C1(n22244), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n22197), .B(n22150), .ZN(n22158) );
  OAI21_X1 U23866 ( .B1(n22153), .B2(n22152), .A(n22151), .ZN(n22154) );
  AOI22_X1 U23867 ( .A1(n22156), .A2(n22260), .B1(n22155), .B2(n22154), .ZN(
        n22157) );
  OAI211_X1 U23868 ( .C1(n22246), .C2(n22159), .A(n22158), .B(n22157), .ZN(
        P1_U2828) );
  OAI22_X1 U23869 ( .A1(n22256), .A2(n22161), .B1(n22254), .B2(n22160), .ZN(
        n22162) );
  AOI211_X1 U23870 ( .C1(n22163), .C2(n22199), .A(n22197), .B(n22162), .ZN(
        n22170) );
  AOI22_X1 U23871 ( .A1(n22165), .A2(n22262), .B1(n22260), .B2(n22164), .ZN(
        n22169) );
  NAND2_X1 U23872 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n22167), .ZN(n22175) );
  OAI211_X1 U23873 ( .C1(n22167), .C2(P1_REIP_REG_15__SCAN_IN), .A(n22166), 
        .B(n22175), .ZN(n22168) );
  NAND3_X1 U23874 ( .A1(n22170), .A2(n22169), .A3(n22168), .ZN(P1_U2825) );
  OAI22_X1 U23875 ( .A1(n22256), .A2(n22172), .B1(n22171), .B2(n22254), .ZN(
        n22173) );
  AOI211_X1 U23876 ( .C1(n22260), .C2(n22174), .A(n22197), .B(n22173), .ZN(
        n22182) );
  OAI21_X1 U23877 ( .B1(n22177), .B2(n22176), .A(n22175), .ZN(n22178) );
  AOI22_X1 U23878 ( .A1(n22180), .A2(n22262), .B1(n22179), .B2(n22178), .ZN(
        n22181) );
  OAI211_X1 U23879 ( .C1(n22267), .C2(n22183), .A(n22182), .B(n22181), .ZN(
        P1_U2824) );
  OAI22_X1 U23880 ( .A1(n22185), .A2(n22256), .B1(n22251), .B2(n22184), .ZN(
        n22186) );
  AOI211_X1 U23881 ( .C1(P1_EBX_REG_18__SCAN_IN), .C2(n22235), .A(n22197), .B(
        n22186), .ZN(n22189) );
  AND2_X1 U23882 ( .A1(n22187), .A2(n22204), .ZN(n22201) );
  INV_X1 U23883 ( .A(n22201), .ZN(n22188) );
  OAI211_X1 U23884 ( .C1(n22190), .C2(n22246), .A(n22189), .B(n22188), .ZN(
        n22191) );
  AOI21_X1 U23885 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(n22202), .A(n22191), 
        .ZN(n22192) );
  OAI21_X1 U23886 ( .B1(n22267), .B2(n22193), .A(n22192), .ZN(P1_U2822) );
  OAI22_X1 U23887 ( .A1(n22251), .A2(n22195), .B1(n22254), .B2(n22194), .ZN(
        n22196) );
  AOI211_X1 U23888 ( .C1(n22244), .C2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n22197), .B(n22196), .ZN(n22208) );
  AOI22_X1 U23889 ( .A1(n22200), .A2(n22262), .B1(n22199), .B2(n22198), .ZN(
        n22207) );
  OAI21_X1 U23890 ( .B1(n22202), .B2(n22201), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n22206) );
  NAND3_X1 U23891 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n22204), .A3(n22203), 
        .ZN(n22205) );
  NAND4_X1 U23892 ( .A1(n22208), .A2(n22207), .A3(n22206), .A4(n22205), .ZN(
        P1_U2821) );
  NOR2_X1 U23893 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n22220), .ZN(n22209) );
  AOI22_X1 U23894 ( .A1(n22210), .A2(n22209), .B1(n22235), .B2(
        P1_EBX_REG_21__SCAN_IN), .ZN(n22211) );
  OAI21_X1 U23895 ( .B1(n22256), .B2(n22212), .A(n22211), .ZN(n22213) );
  AOI21_X1 U23896 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n22222), .A(n22213), 
        .ZN(n22218) );
  NOR2_X1 U23897 ( .A1(n22214), .A2(n22267), .ZN(n22215) );
  AOI21_X1 U23898 ( .B1(n22216), .B2(n22262), .A(n22215), .ZN(n22217) );
  OAI211_X1 U23899 ( .C1(n22219), .C2(n22251), .A(n22218), .B(n22217), .ZN(
        P1_U2819) );
  NOR3_X1 U23900 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n22221), .A3(n22220), 
        .ZN(n22228) );
  AOI21_X1 U23901 ( .B1(n22236), .B2(n22223), .A(n22222), .ZN(n22226) );
  OAI22_X1 U23902 ( .A1(n22226), .A2(n22225), .B1(n22254), .B2(n22224), .ZN(
        n22227) );
  AOI211_X1 U23903 ( .C1(n22244), .C2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n22228), .B(n22227), .ZN(n22233) );
  OAI22_X1 U23904 ( .A1(n22230), .A2(n22246), .B1(n22229), .B2(n22251), .ZN(
        n22231) );
  INV_X1 U23905 ( .A(n22231), .ZN(n22232) );
  OAI211_X1 U23906 ( .C1(n22267), .C2(n22234), .A(n22233), .B(n22232), .ZN(
        P1_U2818) );
  NAND2_X1 U23907 ( .A1(n22235), .A2(P1_EBX_REG_23__SCAN_IN), .ZN(n22240) );
  NAND3_X1 U23908 ( .A1(n22238), .A2(n22237), .A3(n22236), .ZN(n22239) );
  OAI211_X1 U23909 ( .C1(n22242), .C2(n22241), .A(n22240), .B(n22239), .ZN(
        n22243) );
  AOI21_X1 U23910 ( .B1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n22244), .A(
        n22243), .ZN(n22250) );
  OAI22_X1 U23911 ( .A1(n22247), .A2(n22246), .B1(n22245), .B2(n22267), .ZN(
        n22248) );
  INV_X1 U23912 ( .A(n22248), .ZN(n22249) );
  OAI211_X1 U23913 ( .C1(n22252), .C2(n22251), .A(n22250), .B(n22249), .ZN(
        P1_U2817) );
  INV_X1 U23914 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n22255) );
  OAI22_X1 U23915 ( .A1(n22256), .A2(n22255), .B1(n22254), .B2(n22253), .ZN(
        n22257) );
  AOI221_X1 U23916 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n22259), .C1(n22258), 
        .C2(n22259), .A(n22257), .ZN(n22265) );
  AOI22_X1 U23917 ( .A1(n22263), .A2(n22262), .B1(n22261), .B2(n22260), .ZN(
        n22264) );
  OAI211_X1 U23918 ( .C1(n22267), .C2(n22266), .A(n22265), .B(n22264), .ZN(
        P1_U2816) );
  OAI21_X1 U23919 ( .B1(n22270), .B2(n22269), .A(n22268), .ZN(P1_U2806) );
  NAND2_X1 U23920 ( .A1(n22272), .A2(n22271), .ZN(P1_U3163) );
  OAI22_X1 U23921 ( .A1(n22275), .A2(n22435), .B1(n22274), .B2(n22273), .ZN(
        P1_U3466) );
  AOI21_X1 U23922 ( .B1(n22278), .B2(n22277), .A(n22276), .ZN(n22279) );
  OAI22_X1 U23923 ( .A1(n22281), .A2(n22280), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n22279), .ZN(n22282) );
  OAI21_X1 U23924 ( .B1(n22284), .B2(n22283), .A(n22282), .ZN(P1_U3161) );
  OAI21_X1 U23925 ( .B1(n22287), .B2(n22286), .A(n22285), .ZN(P1_U2805) );
  AOI21_X1 U23926 ( .B1(n22289), .B2(P1_DATAWIDTH_REG_1__SCAN_IN), .A(n22288), 
        .ZN(n22290) );
  INV_X1 U23927 ( .A(n22290), .ZN(P1_U3465) );
  INV_X1 U23928 ( .A(n22291), .ZN(n22293) );
  OAI21_X1 U23929 ( .B1(n22295), .B2(n22292), .A(n22293), .ZN(P2_U2818) );
  OAI21_X1 U23930 ( .B1(n22295), .B2(n22294), .A(n22293), .ZN(P2_U3592) );
  OAI21_X1 U23931 ( .B1(n22299), .B2(n22296), .A(n22297), .ZN(P3_U2636) );
  INV_X1 U23932 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n22298) );
  OAI21_X1 U23933 ( .B1(n22299), .B2(n22298), .A(n22297), .ZN(P3_U3281) );
  NAND2_X1 U23934 ( .A1(HOLD), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n22344) );
  INV_X1 U23935 ( .A(n22344), .ZN(n22300) );
  INV_X1 U23936 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n22343) );
  AOI211_X1 U23937 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(HOLD), .A(n22300), .B(
        n22343), .ZN(n22302) );
  AOI21_X1 U23938 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n22341), .A(n22345), 
        .ZN(n22356) );
  AOI21_X1 U23939 ( .B1(NA), .B2(n22346), .A(n22301), .ZN(n22349) );
  OAI22_X1 U23940 ( .A1(n22303), .A2(n22302), .B1(n22356), .B2(n22349), .ZN(
        P3_U3029) );
  NAND2_X1 U23941 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n22305), .ZN(n22316) );
  AOI22_X1 U23942 ( .A1(NA), .A2(n22311), .B1(P1_STATE_REG_0__SCAN_IN), .B2(
        n22316), .ZN(n22309) );
  INV_X1 U23943 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n22307) );
  INV_X1 U23944 ( .A(HOLD), .ZN(n22339) );
  INV_X1 U23945 ( .A(NA), .ZN(n22350) );
  AOI21_X1 U23946 ( .B1(n22305), .B2(n22350), .A(n22304), .ZN(n22306) );
  OAI21_X1 U23947 ( .B1(n22339), .B2(n22312), .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n22317) );
  INV_X1 U23948 ( .A(n22317), .ZN(n22313) );
  OAI33_X1 U23949 ( .A1(n22316), .A2(NA), .A3(n22307), .B1(n22339), .B2(n22306), .B3(n22313), .ZN(n22308) );
  AOI22_X1 U23950 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n22309), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(n22308), .ZN(n22310) );
  INV_X1 U23951 ( .A(n22310), .ZN(P1_U3196) );
  NOR2_X1 U23952 ( .A1(n22339), .A2(n22311), .ZN(n22318) );
  AOI22_X1 U23953 ( .A1(n22313), .A2(P1_STATE_REG_0__SCAN_IN), .B1(n22318), 
        .B2(n22312), .ZN(n22315) );
  NAND3_X1 U23954 ( .A1(n22315), .A2(n22314), .A3(n22316), .ZN(P1_U3195) );
  AND2_X1 U23955 ( .A1(n22316), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n22320) );
  AOI211_X1 U23956 ( .C1(NA), .C2(n14846), .A(n22318), .B(n22317), .ZN(n22319)
         );
  OAI22_X1 U23957 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n22320), .B1(n22682), 
        .B2(n22319), .ZN(P1_U3194) );
  NOR2_X1 U23958 ( .A1(n17987), .A2(n22339), .ZN(n22325) );
  NAND2_X1 U23959 ( .A1(n22321), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n22334) );
  NAND2_X1 U23960 ( .A1(n22334), .A2(P2_STATE_REG_0__SCAN_IN), .ZN(n22333) );
  INV_X1 U23961 ( .A(n22322), .ZN(n22323) );
  OAI21_X1 U23962 ( .B1(n22323), .B2(n22350), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n22338) );
  AOI22_X1 U23963 ( .A1(n22325), .A2(n22324), .B1(n22333), .B2(n22338), .ZN(
        n22326) );
  OAI21_X1 U23964 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(n22327), .A(n22326), .ZN(P2_U3209) );
  OAI211_X1 U23965 ( .C1(n22328), .C2(n22339), .A(P2_STATE_REG_0__SCAN_IN), 
        .B(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n22331) );
  NAND2_X1 U23966 ( .A1(n22329), .A2(HOLD), .ZN(n22330) );
  NAND4_X1 U23967 ( .A1(n22332), .A2(n22331), .A3(n22334), .A4(n22330), .ZN(
        P2_U3210) );
  INV_X1 U23968 ( .A(n22333), .ZN(n22337) );
  OAI22_X1 U23969 ( .A1(NA), .A2(n22334), .B1(P2_STATE_REG_1__SCAN_IN), .B2(
        P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n22335) );
  OAI211_X1 U23970 ( .C1(HOLD), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n22335), .ZN(n22336) );
  OAI221_X1 U23971 ( .B1(n22338), .B2(n22337), .C1(n22338), .C2(n22339), .A(
        n22336), .ZN(P2_U3211) );
  AOI21_X1 U23972 ( .B1(n22339), .B2(n22343), .A(n22345), .ZN(n22342) );
  AOI211_X1 U23973 ( .C1(n22342), .C2(n22344), .A(n22341), .B(n22340), .ZN(
        n22348) );
  NOR2_X1 U23974 ( .A1(n22345), .A2(n22343), .ZN(n22351) );
  AOI22_X1 U23975 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n22345), .B1(n22351), 
        .B2(n22344), .ZN(n22347) );
  AOI22_X1 U23976 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n22348), .B1(n22347), 
        .B2(n22346), .ZN(P3_U3030) );
  AOI21_X1 U23977 ( .B1(n22351), .B2(n22350), .A(n22349), .ZN(n22355) );
  AOI221_X1 U23978 ( .B1(NA), .B2(P3_STATE_REG_1__SCAN_IN), .C1(n22352), .C2(
        P3_STATE_REG_1__SCAN_IN), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n22353) );
  OAI211_X1 U23979 ( .C1(P3_STATE_REG_2__SCAN_IN), .C2(n22353), .A(HOLD), .B(
        P3_STATE_REG_0__SCAN_IN), .ZN(n22354) );
  OAI21_X1 U23980 ( .B1(n22356), .B2(n22355), .A(n22354), .ZN(P3_U3031) );
  INV_X1 U23981 ( .A(n22615), .ZN(n22676) );
  NOR2_X1 U23982 ( .A1(n22676), .A2(n22424), .ZN(n22357) );
  NOR2_X1 U23983 ( .A1(n22424), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n22425) );
  AOI21_X1 U23984 ( .B1(n22366), .B2(n22357), .A(n22425), .ZN(n22365) );
  INV_X1 U23985 ( .A(n22365), .ZN(n22359) );
  NOR2_X1 U23986 ( .A1(n22382), .A2(n22427), .ZN(n22364) );
  NAND2_X1 U23987 ( .A1(n22415), .A2(n22360), .ZN(n22614) );
  OAI22_X1 U23988 ( .A1(n22615), .A2(n22401), .B1(n22614), .B2(n22400), .ZN(
        n22361) );
  INV_X1 U23989 ( .A(n22361), .ZN(n22368) );
  AOI22_X1 U23990 ( .A1(n22362), .A2(P1_STATE2_REG_2__SCAN_IN), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n22614), .ZN(n22363) );
  OAI211_X1 U23991 ( .C1(n22365), .C2(n22364), .A(n22419), .B(n22363), .ZN(
        n22618) );
  INV_X1 U23992 ( .A(n22366), .ZN(n22617) );
  AOI22_X1 U23993 ( .A1(n22618), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n22617), .B2(n22434), .ZN(n22367) );
  OAI211_X1 U23994 ( .C1(n22621), .C2(n22445), .A(n22368), .B(n22367), .ZN(
        P1_U3033) );
  NOR2_X1 U23995 ( .A1(n22633), .A2(n22424), .ZN(n22371) );
  AOI21_X1 U23996 ( .B1(n22371), .B2(n22623), .A(n22425), .ZN(n22378) );
  INV_X1 U23997 ( .A(n22378), .ZN(n22373) );
  NOR2_X1 U23998 ( .A1(n22382), .A2(n14969), .ZN(n22377) );
  NOR3_X1 U23999 ( .A1(n22374), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n22388) );
  NAND2_X1 U24000 ( .A1(n22415), .A2(n22388), .ZN(n22622) );
  OAI22_X1 U24001 ( .A1(n22623), .A2(n22401), .B1(n22622), .B2(n22400), .ZN(
        n22375) );
  INV_X1 U24002 ( .A(n22375), .ZN(n22380) );
  NOR2_X1 U24003 ( .A1(n11636), .A2(n15575), .ZN(n22403) );
  AOI21_X1 U24004 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22622), .A(n22403), 
        .ZN(n22376) );
  OAI211_X1 U24005 ( .C1(n22378), .C2(n22377), .A(n22419), .B(n22376), .ZN(
        n22625) );
  AOI22_X1 U24006 ( .A1(n22625), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n22633), .B2(n22434), .ZN(n22379) );
  OAI211_X1 U24007 ( .C1(n22628), .C2(n22445), .A(n22380), .B(n22379), .ZN(
        P1_U3049) );
  OR2_X1 U24008 ( .A1(n22382), .A2(n22381), .ZN(n22384) );
  INV_X1 U24009 ( .A(n22388), .ZN(n22383) );
  OR2_X1 U24010 ( .A1(n22415), .A2(n22383), .ZN(n22629) );
  NAND2_X1 U24011 ( .A1(n22384), .A2(n22629), .ZN(n22391) );
  OAI22_X1 U24012 ( .A1(n22592), .A2(n22401), .B1(n22629), .B2(n22400), .ZN(
        n22385) );
  INV_X1 U24013 ( .A(n22385), .ZN(n22394) );
  INV_X1 U24014 ( .A(n22386), .ZN(n22392) );
  OAI21_X1 U24015 ( .B1(n15786), .B2(n22388), .A(n22387), .ZN(n22389) );
  INV_X1 U24016 ( .A(n22389), .ZN(n22390) );
  AOI22_X1 U24017 ( .A1(n22634), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n22594), .B2(n22434), .ZN(n22393) );
  OAI211_X1 U24018 ( .C1(n22637), .C2(n22445), .A(n22394), .B(n22393), .ZN(
        P1_U3057) );
  NOR2_X1 U24019 ( .A1(n22642), .A2(n22424), .ZN(n22395) );
  AOI21_X1 U24020 ( .B1(n22395), .B2(n22640), .A(n22425), .ZN(n22406) );
  INV_X1 U24021 ( .A(n22406), .ZN(n22397) );
  AND2_X1 U24022 ( .A1(n22396), .A2(n22427), .ZN(n22405) );
  INV_X1 U24023 ( .A(n22398), .ZN(n22399) );
  NOR2_X1 U24024 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22399), .ZN(
        n22597) );
  INV_X1 U24025 ( .A(n22597), .ZN(n22638) );
  OAI22_X1 U24026 ( .A1(n22640), .A2(n22401), .B1(n22638), .B2(n22400), .ZN(
        n22402) );
  INV_X1 U24027 ( .A(n22402), .ZN(n22408) );
  AOI21_X1 U24028 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22638), .A(n22403), 
        .ZN(n22404) );
  OAI211_X1 U24029 ( .C1(n22406), .C2(n22405), .A(n22439), .B(n22404), .ZN(
        n22643) );
  AOI22_X1 U24030 ( .A1(n22643), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n22642), .B2(n22434), .ZN(n22407) );
  OAI211_X1 U24031 ( .C1(n22646), .C2(n22445), .A(n22408), .B(n22407), .ZN(
        P1_U3081) );
  NOR2_X1 U24032 ( .A1(n22654), .A2(n22424), .ZN(n22409) );
  AOI21_X1 U24033 ( .B1(n22409), .B2(n22604), .A(n22425), .ZN(n22421) );
  INV_X1 U24034 ( .A(n22421), .ZN(n22413) );
  AND2_X1 U24035 ( .A1(n22410), .A2(n22427), .ZN(n22420) );
  NAND2_X1 U24036 ( .A1(n22415), .A2(n22414), .ZN(n22602) );
  INV_X1 U24037 ( .A(n22602), .ZN(n22653) );
  AOI22_X1 U24038 ( .A1(n22654), .A2(n22434), .B1(n22653), .B2(n22433), .ZN(
        n22423) );
  INV_X1 U24039 ( .A(n22416), .ZN(n22417) );
  AOI21_X1 U24040 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22602), .A(n22417), 
        .ZN(n22418) );
  OAI211_X1 U24041 ( .C1(n22421), .C2(n22420), .A(n22419), .B(n22418), .ZN(
        n22656) );
  INV_X1 U24042 ( .A(n22604), .ZN(n22655) );
  AOI22_X1 U24043 ( .A1(n22656), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n22655), .B2(n22442), .ZN(n22422) );
  OAI211_X1 U24044 ( .C1(n22659), .C2(n22445), .A(n22423), .B(n22422), .ZN(
        P1_U3113) );
  NOR3_X1 U24045 ( .A1(n22663), .A2(n22661), .A3(n22424), .ZN(n22426) );
  NOR2_X1 U24046 ( .A1(n22426), .A2(n22425), .ZN(n22441) );
  INV_X1 U24047 ( .A(n22441), .ZN(n22431) );
  NOR2_X1 U24048 ( .A1(n22428), .A2(n22427), .ZN(n22440) );
  NOR2_X1 U24049 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22432), .ZN(
        n22660) );
  AOI22_X1 U24050 ( .A1(n22661), .A2(n22434), .B1(n22660), .B2(n22433), .ZN(
        n22444) );
  NOR2_X1 U24051 ( .A1(n22435), .A2(n22660), .ZN(n22436) );
  AOI21_X1 U24052 ( .B1(n22437), .B2(P1_STATE2_REG_2__SCAN_IN), .A(n22436), 
        .ZN(n22438) );
  OAI211_X1 U24053 ( .C1(n22441), .C2(n22440), .A(n22439), .B(n22438), .ZN(
        n22664) );
  AOI22_X1 U24054 ( .A1(n22664), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n22663), .B2(n22442), .ZN(n22443) );
  OAI211_X1 U24055 ( .C1(n22668), .C2(n22445), .A(n22444), .B(n22443), .ZN(
        P1_U3129) );
  OAI22_X1 U24056 ( .A1(n22615), .A2(n22460), .B1(n22614), .B2(n22459), .ZN(
        n22446) );
  INV_X1 U24057 ( .A(n22446), .ZN(n22448) );
  AOI22_X1 U24058 ( .A1(n22618), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n22617), .B2(n22465), .ZN(n22447) );
  OAI211_X1 U24059 ( .C1(n22621), .C2(n22469), .A(n22448), .B(n22447), .ZN(
        P1_U3034) );
  OAI22_X1 U24060 ( .A1(n22623), .A2(n22460), .B1(n22622), .B2(n22459), .ZN(
        n22449) );
  INV_X1 U24061 ( .A(n22449), .ZN(n22451) );
  AOI22_X1 U24062 ( .A1(n22625), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n22633), .B2(n22465), .ZN(n22450) );
  OAI211_X1 U24063 ( .C1(n22628), .C2(n22469), .A(n22451), .B(n22450), .ZN(
        P1_U3050) );
  OAI22_X1 U24064 ( .A1(n22631), .A2(n22452), .B1(n22459), .B2(n22629), .ZN(
        n22453) );
  INV_X1 U24065 ( .A(n22453), .ZN(n22455) );
  AOI22_X1 U24066 ( .A1(n22634), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n22633), .B2(n22466), .ZN(n22454) );
  OAI211_X1 U24067 ( .C1(n22637), .C2(n22469), .A(n22455), .B(n22454), .ZN(
        P1_U3058) );
  OAI22_X1 U24068 ( .A1(n22640), .A2(n22460), .B1(n22638), .B2(n22459), .ZN(
        n22456) );
  INV_X1 U24069 ( .A(n22456), .ZN(n22458) );
  AOI22_X1 U24070 ( .A1(n22643), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n22642), .B2(n22465), .ZN(n22457) );
  OAI211_X1 U24071 ( .C1(n22646), .C2(n22469), .A(n22458), .B(n22457), .ZN(
        P1_U3082) );
  OAI22_X1 U24072 ( .A1(n22604), .A2(n22460), .B1(n22602), .B2(n22459), .ZN(
        n22461) );
  INV_X1 U24073 ( .A(n22461), .ZN(n22463) );
  AOI22_X1 U24074 ( .A1(n22656), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n22654), .B2(n22465), .ZN(n22462) );
  OAI211_X1 U24075 ( .C1(n22659), .C2(n22469), .A(n22463), .B(n22462), .ZN(
        P1_U3114) );
  AOI22_X1 U24076 ( .A1(n22661), .A2(n22465), .B1(n22660), .B2(n22464), .ZN(
        n22468) );
  AOI22_X1 U24077 ( .A1(n22664), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n22663), .B2(n22466), .ZN(n22467) );
  OAI211_X1 U24078 ( .C1(n22668), .C2(n22469), .A(n22468), .B(n22467), .ZN(
        P1_U3130) );
  OAI22_X1 U24079 ( .A1(n22615), .A2(n22483), .B1(n22614), .B2(n22482), .ZN(
        n22470) );
  INV_X1 U24080 ( .A(n22470), .ZN(n22472) );
  AOI22_X1 U24081 ( .A1(n22618), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n22617), .B2(n22488), .ZN(n22471) );
  OAI211_X1 U24082 ( .C1(n22621), .C2(n22492), .A(n22472), .B(n22471), .ZN(
        P1_U3035) );
  OAI22_X1 U24083 ( .A1(n22623), .A2(n22483), .B1(n22622), .B2(n22482), .ZN(
        n22473) );
  INV_X1 U24084 ( .A(n22473), .ZN(n22475) );
  AOI22_X1 U24085 ( .A1(n22625), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n22633), .B2(n22488), .ZN(n22474) );
  OAI211_X1 U24086 ( .C1(n22628), .C2(n22492), .A(n22475), .B(n22474), .ZN(
        P1_U3051) );
  OAI22_X1 U24087 ( .A1(n22631), .A2(n22476), .B1(n22482), .B2(n22629), .ZN(
        n22477) );
  INV_X1 U24088 ( .A(n22477), .ZN(n22479) );
  AOI22_X1 U24089 ( .A1(n22634), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n22633), .B2(n22489), .ZN(n22478) );
  OAI211_X1 U24090 ( .C1(n22637), .C2(n22492), .A(n22479), .B(n22478), .ZN(
        P1_U3059) );
  AOI22_X1 U24091 ( .A1(n22642), .A2(n22488), .B1(n22597), .B2(n22487), .ZN(
        n22481) );
  INV_X1 U24092 ( .A(n22640), .ZN(n22598) );
  AOI22_X1 U24093 ( .A1(n22643), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n22598), .B2(n22489), .ZN(n22480) );
  OAI211_X1 U24094 ( .C1(n22646), .C2(n22492), .A(n22481), .B(n22480), .ZN(
        P1_U3083) );
  OAI22_X1 U24095 ( .A1(n22604), .A2(n22483), .B1(n22602), .B2(n22482), .ZN(
        n22484) );
  INV_X1 U24096 ( .A(n22484), .ZN(n22486) );
  AOI22_X1 U24097 ( .A1(n22656), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n22654), .B2(n22488), .ZN(n22485) );
  OAI211_X1 U24098 ( .C1(n22659), .C2(n22492), .A(n22486), .B(n22485), .ZN(
        P1_U3115) );
  AOI22_X1 U24099 ( .A1(n22661), .A2(n22488), .B1(n22660), .B2(n22487), .ZN(
        n22491) );
  AOI22_X1 U24100 ( .A1(n22664), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n22663), .B2(n22489), .ZN(n22490) );
  OAI211_X1 U24101 ( .C1(n22668), .C2(n22492), .A(n22491), .B(n22490), .ZN(
        P1_U3131) );
  OAI22_X1 U24102 ( .A1(n22615), .A2(n22507), .B1(n22614), .B2(n22506), .ZN(
        n22493) );
  INV_X1 U24103 ( .A(n22493), .ZN(n22495) );
  AOI22_X1 U24104 ( .A1(n22618), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n22617), .B2(n22512), .ZN(n22494) );
  OAI211_X1 U24105 ( .C1(n22621), .C2(n22516), .A(n22495), .B(n22494), .ZN(
        P1_U3036) );
  OAI22_X1 U24106 ( .A1(n22592), .A2(n22499), .B1(n22622), .B2(n22506), .ZN(
        n22496) );
  INV_X1 U24107 ( .A(n22496), .ZN(n22498) );
  AOI22_X1 U24108 ( .A1(n22625), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n22589), .B2(n22513), .ZN(n22497) );
  OAI211_X1 U24109 ( .C1(n22628), .C2(n22516), .A(n22498), .B(n22497), .ZN(
        P1_U3052) );
  OAI22_X1 U24110 ( .A1(n22631), .A2(n22499), .B1(n22506), .B2(n22629), .ZN(
        n22500) );
  INV_X1 U24111 ( .A(n22500), .ZN(n22502) );
  AOI22_X1 U24112 ( .A1(n22634), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n22633), .B2(n22513), .ZN(n22501) );
  OAI211_X1 U24113 ( .C1(n22637), .C2(n22516), .A(n22502), .B(n22501), .ZN(
        P1_U3060) );
  OAI22_X1 U24114 ( .A1(n22640), .A2(n22507), .B1(n22638), .B2(n22506), .ZN(
        n22503) );
  INV_X1 U24115 ( .A(n22503), .ZN(n22505) );
  AOI22_X1 U24116 ( .A1(n22643), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n22642), .B2(n22512), .ZN(n22504) );
  OAI211_X1 U24117 ( .C1(n22646), .C2(n22516), .A(n22505), .B(n22504), .ZN(
        P1_U3084) );
  OAI22_X1 U24118 ( .A1(n22604), .A2(n22507), .B1(n22602), .B2(n22506), .ZN(
        n22508) );
  INV_X1 U24119 ( .A(n22508), .ZN(n22510) );
  AOI22_X1 U24120 ( .A1(n22656), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n22654), .B2(n22512), .ZN(n22509) );
  OAI211_X1 U24121 ( .C1(n22659), .C2(n22516), .A(n22510), .B(n22509), .ZN(
        P1_U3116) );
  AOI22_X1 U24122 ( .A1(n22661), .A2(n22512), .B1(n22660), .B2(n22511), .ZN(
        n22515) );
  AOI22_X1 U24123 ( .A1(n22664), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n22663), .B2(n22513), .ZN(n22514) );
  OAI211_X1 U24124 ( .C1(n22668), .C2(n22516), .A(n22515), .B(n22514), .ZN(
        P1_U3132) );
  OAI22_X1 U24125 ( .A1(n22615), .A2(n22536), .B1(n22614), .B2(n22535), .ZN(
        n22517) );
  INV_X1 U24126 ( .A(n22517), .ZN(n22519) );
  AOI22_X1 U24127 ( .A1(n22618), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n22547), .B2(n22617), .ZN(n22518) );
  OAI211_X1 U24128 ( .C1(n22621), .C2(n22550), .A(n22519), .B(n22518), .ZN(
        P1_U3037) );
  OAI22_X1 U24129 ( .A1(n22592), .A2(n22560), .B1(n22535), .B2(n22622), .ZN(
        n22520) );
  INV_X1 U24130 ( .A(n22520), .ZN(n22522) );
  AOI22_X1 U24131 ( .A1(n22625), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n22589), .B2(n22555), .ZN(n22521) );
  OAI211_X1 U24132 ( .C1(n22628), .C2(n22550), .A(n22522), .B(n22521), .ZN(
        P1_U3053) );
  OAI22_X1 U24133 ( .A1(n22631), .A2(n22560), .B1(n22535), .B2(n22629), .ZN(
        n22523) );
  INV_X1 U24134 ( .A(n22523), .ZN(n22525) );
  AOI22_X1 U24135 ( .A1(n22634), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n22633), .B2(n22555), .ZN(n22524) );
  OAI211_X1 U24136 ( .C1(n22637), .C2(n22550), .A(n22525), .B(n22524), .ZN(
        P1_U3061) );
  AOI22_X1 U24137 ( .A1(n22642), .A2(n22547), .B1(n22554), .B2(n22597), .ZN(
        n22527) );
  AOI22_X1 U24138 ( .A1(n22643), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n22598), .B2(n22555), .ZN(n22526) );
  OAI211_X1 U24139 ( .C1(n22646), .C2(n22550), .A(n22527), .B(n22526), .ZN(
        P1_U3085) );
  INV_X1 U24140 ( .A(n22528), .ZN(n22530) );
  AOI22_X1 U24141 ( .A1(n22530), .A2(n22552), .B1(n22554), .B2(n22529), .ZN(
        n22534) );
  AOI22_X1 U24142 ( .A1(n22532), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n22531), .B2(n22555), .ZN(n22533) );
  OAI211_X1 U24143 ( .C1(n22560), .C2(n22652), .A(n22534), .B(n22533), .ZN(
        P1_U3101) );
  OAI22_X1 U24144 ( .A1(n22604), .A2(n22536), .B1(n22602), .B2(n22535), .ZN(
        n22537) );
  INV_X1 U24145 ( .A(n22537), .ZN(n22539) );
  AOI22_X1 U24146 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n22656), .B1(
        n22654), .B2(n22547), .ZN(n22538) );
  OAI211_X1 U24147 ( .C1(n22659), .C2(n22550), .A(n22539), .B(n22538), .ZN(
        P1_U3117) );
  INV_X1 U24148 ( .A(n22540), .ZN(n22542) );
  AOI22_X1 U24149 ( .A1(n22552), .A2(n22542), .B1(n22554), .B2(n22541), .ZN(
        n22545) );
  AOI22_X1 U24150 ( .A1(n22543), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n22654), .B2(n22555), .ZN(n22544) );
  OAI211_X1 U24151 ( .C1(n22560), .C2(n22546), .A(n22545), .B(n22544), .ZN(
        P1_U3125) );
  AOI22_X1 U24152 ( .A1(n22661), .A2(n22547), .B1(n22554), .B2(n22660), .ZN(
        n22549) );
  AOI22_X1 U24153 ( .A1(n22664), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n22663), .B2(n22555), .ZN(n22548) );
  OAI211_X1 U24154 ( .C1(n22668), .C2(n22550), .A(n22549), .B(n22548), .ZN(
        P1_U3133) );
  AOI22_X1 U24155 ( .A1(n22554), .A2(n22553), .B1(n22552), .B2(n22551), .ZN(
        n22559) );
  AOI22_X1 U24156 ( .A1(n22557), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n22556), .B2(n22555), .ZN(n22558) );
  OAI211_X1 U24157 ( .C1(n22560), .C2(n22680), .A(n22559), .B(n22558), .ZN(
        P1_U3149) );
  OAI22_X1 U24158 ( .A1(n22615), .A2(n22574), .B1(n22614), .B2(n22573), .ZN(
        n22561) );
  INV_X1 U24159 ( .A(n22561), .ZN(n22563) );
  AOI22_X1 U24160 ( .A1(n22618), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n22617), .B2(n22579), .ZN(n22562) );
  OAI211_X1 U24161 ( .C1(n22621), .C2(n22583), .A(n22563), .B(n22562), .ZN(
        P1_U3038) );
  OAI22_X1 U24162 ( .A1(n22623), .A2(n22574), .B1(n22622), .B2(n22573), .ZN(
        n22564) );
  INV_X1 U24163 ( .A(n22564), .ZN(n22566) );
  AOI22_X1 U24164 ( .A1(n22625), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n22633), .B2(n22579), .ZN(n22565) );
  OAI211_X1 U24165 ( .C1(n22628), .C2(n22583), .A(n22566), .B(n22565), .ZN(
        P1_U3054) );
  OAI22_X1 U24166 ( .A1(n22631), .A2(n22567), .B1(n22573), .B2(n22629), .ZN(
        n22568) );
  INV_X1 U24167 ( .A(n22568), .ZN(n22570) );
  AOI22_X1 U24168 ( .A1(n22634), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n22633), .B2(n22580), .ZN(n22569) );
  OAI211_X1 U24169 ( .C1(n22637), .C2(n22583), .A(n22570), .B(n22569), .ZN(
        P1_U3062) );
  AOI22_X1 U24170 ( .A1(n22642), .A2(n22579), .B1(n22597), .B2(n22578), .ZN(
        n22572) );
  AOI22_X1 U24171 ( .A1(n22643), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n22598), .B2(n22580), .ZN(n22571) );
  OAI211_X1 U24172 ( .C1(n22646), .C2(n22583), .A(n22572), .B(n22571), .ZN(
        P1_U3086) );
  OAI22_X1 U24173 ( .A1(n22604), .A2(n22574), .B1(n22602), .B2(n22573), .ZN(
        n22575) );
  INV_X1 U24174 ( .A(n22575), .ZN(n22577) );
  AOI22_X1 U24175 ( .A1(n22656), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n22654), .B2(n22579), .ZN(n22576) );
  OAI211_X1 U24176 ( .C1(n22659), .C2(n22583), .A(n22577), .B(n22576), .ZN(
        P1_U3118) );
  AOI22_X1 U24177 ( .A1(n22661), .A2(n22579), .B1(n22660), .B2(n22578), .ZN(
        n22582) );
  AOI22_X1 U24178 ( .A1(n22664), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n22663), .B2(n22580), .ZN(n22581) );
  OAI211_X1 U24179 ( .C1(n22668), .C2(n22583), .A(n22582), .B(n22581), .ZN(
        P1_U3134) );
  OAI22_X1 U24180 ( .A1(n22615), .A2(n22603), .B1(n22614), .B2(n22601), .ZN(
        n22584) );
  INV_X1 U24181 ( .A(n22584), .ZN(n22586) );
  AOI22_X1 U24182 ( .A1(n22618), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n22617), .B2(n22609), .ZN(n22585) );
  OAI211_X1 U24183 ( .C1(n22621), .C2(n22613), .A(n22586), .B(n22585), .ZN(
        P1_U3039) );
  OAI22_X1 U24184 ( .A1(n22592), .A2(n22587), .B1(n22622), .B2(n22601), .ZN(
        n22588) );
  INV_X1 U24185 ( .A(n22588), .ZN(n22591) );
  AOI22_X1 U24186 ( .A1(n22625), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n22589), .B2(n22610), .ZN(n22590) );
  OAI211_X1 U24187 ( .C1(n22628), .C2(n22613), .A(n22591), .B(n22590), .ZN(
        P1_U3055) );
  OAI22_X1 U24188 ( .A1(n22592), .A2(n22603), .B1(n22629), .B2(n22601), .ZN(
        n22593) );
  INV_X1 U24189 ( .A(n22593), .ZN(n22596) );
  AOI22_X1 U24190 ( .A1(n22634), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n22594), .B2(n22609), .ZN(n22595) );
  OAI211_X1 U24191 ( .C1(n22637), .C2(n22613), .A(n22596), .B(n22595), .ZN(
        P1_U3063) );
  AOI22_X1 U24192 ( .A1(n22642), .A2(n22609), .B1(n22597), .B2(n22608), .ZN(
        n22600) );
  AOI22_X1 U24193 ( .A1(n22643), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n22598), .B2(n22610), .ZN(n22599) );
  OAI211_X1 U24194 ( .C1(n22646), .C2(n22613), .A(n22600), .B(n22599), .ZN(
        P1_U3087) );
  OAI22_X1 U24195 ( .A1(n22604), .A2(n22603), .B1(n22602), .B2(n22601), .ZN(
        n22605) );
  INV_X1 U24196 ( .A(n22605), .ZN(n22607) );
  AOI22_X1 U24197 ( .A1(n22656), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n22654), .B2(n22609), .ZN(n22606) );
  OAI211_X1 U24198 ( .C1(n22659), .C2(n22613), .A(n22607), .B(n22606), .ZN(
        P1_U3119) );
  AOI22_X1 U24199 ( .A1(n22661), .A2(n22609), .B1(n22660), .B2(n22608), .ZN(
        n22612) );
  AOI22_X1 U24200 ( .A1(n22664), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n22663), .B2(n22610), .ZN(n22611) );
  OAI211_X1 U24201 ( .C1(n22668), .C2(n22613), .A(n22612), .B(n22611), .ZN(
        P1_U3135) );
  OAI22_X1 U24202 ( .A1(n22615), .A2(n22681), .B1(n22639), .B2(n22614), .ZN(
        n22616) );
  INV_X1 U24203 ( .A(n22616), .ZN(n22620) );
  AOI22_X1 U24204 ( .A1(n22618), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n22617), .B2(n22675), .ZN(n22619) );
  OAI211_X1 U24205 ( .C1(n22621), .C2(n22667), .A(n22620), .B(n22619), .ZN(
        P1_U3040) );
  OAI22_X1 U24206 ( .A1(n22623), .A2(n22681), .B1(n22639), .B2(n22622), .ZN(
        n22624) );
  INV_X1 U24207 ( .A(n22624), .ZN(n22627) );
  AOI22_X1 U24208 ( .A1(n22625), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n22633), .B2(n22675), .ZN(n22626) );
  OAI211_X1 U24209 ( .C1(n22628), .C2(n22667), .A(n22627), .B(n22626), .ZN(
        P1_U3056) );
  OAI22_X1 U24210 ( .A1(n22631), .A2(n22630), .B1(n22639), .B2(n22629), .ZN(
        n22632) );
  INV_X1 U24211 ( .A(n22632), .ZN(n22636) );
  AOI22_X1 U24212 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n22634), .B1(
        n22633), .B2(n22662), .ZN(n22635) );
  OAI211_X1 U24213 ( .C1(n22637), .C2(n22667), .A(n22636), .B(n22635), .ZN(
        P1_U3064) );
  OAI22_X1 U24214 ( .A1(n22640), .A2(n22681), .B1(n22639), .B2(n22638), .ZN(
        n22641) );
  INV_X1 U24215 ( .A(n22641), .ZN(n22645) );
  AOI22_X1 U24216 ( .A1(n22643), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n22642), .B2(n22675), .ZN(n22644) );
  OAI211_X1 U24217 ( .C1(n22646), .C2(n22667), .A(n22645), .B(n22644), .ZN(
        P1_U3088) );
  AOI22_X1 U24218 ( .A1(n22674), .A2(n22648), .B1(n22671), .B2(n22647), .ZN(
        n22651) );
  AOI22_X1 U24219 ( .A1(n22655), .A2(n22675), .B1(n22649), .B2(
        P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n22650) );
  OAI211_X1 U24220 ( .C1(n22681), .C2(n22652), .A(n22651), .B(n22650), .ZN(
        P1_U3112) );
  AOI22_X1 U24221 ( .A1(n22654), .A2(n22675), .B1(n22653), .B2(n22671), .ZN(
        n22658) );
  AOI22_X1 U24222 ( .A1(n22656), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n22662), .B2(n22655), .ZN(n22657) );
  OAI211_X1 U24223 ( .C1(n22659), .C2(n22667), .A(n22658), .B(n22657), .ZN(
        P1_U3120) );
  AOI22_X1 U24224 ( .A1(n22661), .A2(n22675), .B1(n22660), .B2(n22671), .ZN(
        n22666) );
  AOI22_X1 U24225 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n22664), .B1(
        n22663), .B2(n22662), .ZN(n22665) );
  OAI211_X1 U24226 ( .C1(n22668), .C2(n22667), .A(n22666), .B(n22665), .ZN(
        P1_U3136) );
  INV_X1 U24227 ( .A(n22669), .ZN(n22673) );
  INV_X1 U24228 ( .A(n22670), .ZN(n22672) );
  AOI22_X1 U24229 ( .A1(n22674), .A2(n22673), .B1(n22672), .B2(n22671), .ZN(
        n22679) );
  AOI22_X1 U24230 ( .A1(n22677), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n22676), .B2(n22675), .ZN(n22678) );
  OAI211_X1 U24231 ( .C1(n22681), .C2(n22680), .A(n22679), .B(n22678), .ZN(
        P1_U3160) );
  OAI22_X1 U24232 ( .A1(n20472), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(n22682), .ZN(n22683) );
  INV_X1 U24233 ( .A(n22683), .ZN(P1_U3486) );
  AND2_X1 U11861 ( .A1(n11771), .A2(n11785), .ZN(n19168) );
  OR2_X1 U12956 ( .A1(n11872), .A2(n11876), .ZN(n19857) );
  INV_X1 U11246 ( .A(n21756), .ZN(n21604) );
  CLKBUF_X1 U11245 ( .A(n13136), .Z(n13731) );
  AND2_X1 U11263 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12849) );
  NAND2_X1 U11280 ( .A1(n21388), .A2(n21371), .ZN(n14308) );
  CLKBUF_X1 U11287 ( .A(n12950), .Z(n13911) );
  CLKBUF_X1 U11288 ( .A(n14372), .Z(n18348) );
  NAND4_X1 U11292 ( .A1(n12944), .A2(n12943), .A3(n12942), .A4(n12941), .ZN(
        n12963) );
  CLKBUF_X1 U11304 ( .A(n12973), .Z(n16592) );
  NAND2_X1 U11308 ( .A1(n11739), .A2(n11738), .ZN(n11760) );
  CLKBUF_X1 U11310 ( .A(n11812), .Z(n12706) );
  INV_X1 U11353 ( .A(n11785), .ZN(n20247) );
  CLKBUF_X1 U11359 ( .A(n11769), .Z(n20155) );
  CLKBUF_X1 U11574 ( .A(n13337), .Z(n13338) );
  CLKBUF_X1 U12420 ( .A(n17928), .Z(n17948) );
  CLKBUF_X1 U12591 ( .A(n12761), .Z(n11154) );
  INV_X1 U12629 ( .A(n21656), .ZN(n21811) );
  OR2_X1 U12641 ( .A1(n11762), .A2(n20154), .ZN(n22684) );
  XOR2_X1 U13470 ( .A(n16850), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .Z(
        n22685) );
endmodule

