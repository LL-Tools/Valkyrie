

module b15_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD, 
        READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN, 
        M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN, 
        STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN, 
        W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, DATAI_29_,
         DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
         DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
         DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
         DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
         DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N,
         BS16_N, READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN,
         CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN,
         REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN,
         FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073;

  NAND2_X1 U34610 ( .A1(n4671), .A2(n4670), .ZN(n4669) );
  CLKBUF_X3 U34620 ( .A(n4448), .Z(n3431) );
  CLKBUF_X2 U34630 ( .A(n4383), .Z(n4301) );
  BUF_X2 U34640 ( .A(n3697), .Z(n4405) );
  CLKBUF_X2 U34650 ( .A(n4000), .Z(n3429) );
  CLKBUF_X2 U3466 ( .A(n3700), .Z(n3428) );
  CLKBUF_X2 U3467 ( .A(n3696), .Z(n3430) );
  CLKBUF_X2 U34680 ( .A(n3545), .Z(n4407) );
  CLKBUF_X1 U34690 ( .A(n4388), .Z(n4308) );
  AND2_X1 U34700 ( .A1(n4781), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4749) );
  NOR2_X1 U34740 ( .A1(n4549), .A2(n4548), .ZN(n4550) );
  OR2_X1 U3475 ( .A1(n3519), .A2(n3518), .ZN(n3586) );
  AND2_X1 U3476 ( .A1(n4458), .A2(n4457), .ZN(n4823) );
  INV_X1 U3477 ( .A(n6395), .ZN(n6354) );
  INV_X1 U3479 ( .A(n6375), .ZN(n6390) );
  XNOR2_X1 U3480 ( .A(n4553), .B(n4552), .ZN(n5653) );
  INV_X1 U3481 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4781) );
  OR2_X2 U3482 ( .A1(n3802), .A2(n4933), .ZN(n4990) );
  AND2_X4 U3483 ( .A1(n4749), .A2(n4799), .ZN(n3691) );
  AND2_X4 U3484 ( .A1(n4799), .A2(n3451), .ZN(n3544) );
  AND2_X2 U3485 ( .A1(n4807), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3452)
         );
  NAND2_X2 U3486 ( .A1(n3724), .A2(n3723), .ZN(n4598) );
  AND2_X2 U3487 ( .A1(n3714), .A2(n3713), .ZN(n6585) );
  XNOR2_X1 U3488 ( .A(n3876), .B(n3875), .ZN(n5652) );
  NOR2_X1 U3489 ( .A1(n5209), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3872)
         );
  CLKBUF_X1 U3490 ( .A(n5271), .Z(n5290) );
  CLKBUF_X1 U3491 ( .A(n5300), .Z(n5316) );
  CLKBUF_X1 U3492 ( .A(n5330), .Z(n5344) );
  OAI21_X1 U3493 ( .B1(n5234), .B2(n6224), .A(n5233), .ZN(n5235) );
  NAND2_X1 U3494 ( .A1(n5185), .A2(n4551), .ZN(n4553) );
  AND2_X1 U3495 ( .A1(n4990), .A2(n4992), .ZN(n3822) );
  AND2_X1 U3496 ( .A1(n4952), .A2(n4951), .ZN(n4953) );
  NOR2_X1 U3497 ( .A1(n5474), .A2(n5404), .ZN(n4509) );
  CLKBUF_X1 U3498 ( .A(n4789), .Z(n6574) );
  CLKBUF_X1 U3499 ( .A(n4886), .Z(n6518) );
  NAND2_X2 U3500 ( .A1(n6086), .A2(n5494), .ZN(n5489) );
  BUF_X2 U3502 ( .A(n4689), .Z(n4735) );
  NAND2_X2 U3503 ( .A1(n4615), .A2(n6691), .ZN(n4738) );
  AND2_X2 U3504 ( .A1(n6397), .A2(n4434), .ZN(n6119) );
  NAND2_X1 U3505 ( .A1(n4476), .A2(n4475), .ZN(n4979) );
  NAND2_X1 U3506 ( .A1(n3961), .A2(n3959), .ZN(n3679) );
  CLKBUF_X1 U3507 ( .A(n3683), .Z(n3725) );
  NOR2_X1 U3508 ( .A1(n3816), .A2(n3817), .ZN(n3814) );
  MUX2_X1 U3509 ( .A(n3667), .B(n3666), .S(n3665), .Z(n6634) );
  NAND2_X1 U3510 ( .A1(n3886), .A2(n3608), .ZN(n3918) );
  AND2_X1 U3511 ( .A1(n4831), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3886) );
  CLKBUF_X1 U3512 ( .A(n3598), .Z(n3934) );
  NAND2_X1 U3513 ( .A1(n6908), .A2(n3598), .ZN(n4681) );
  INV_X1 U3514 ( .A(n3598), .ZN(n6864) );
  NAND4_X2 U3515 ( .A1(n3487), .A2(n3486), .A3(n3485), .A4(n3484), .ZN(n3598)
         );
  OR2_X2 U3516 ( .A1(n3563), .A2(n3562), .ZN(n4444) );
  INV_X2 U3517 ( .A(n3586), .ZN(n6780) );
  INV_X1 U3518 ( .A(n6732), .ZN(n4839) );
  AND4_X1 U3519 ( .A1(n3475), .A2(n3474), .A3(n3473), .A4(n3472), .ZN(n3486)
         );
  AND4_X1 U3520 ( .A1(n3496), .A2(n3495), .A3(n3494), .A4(n3493), .ZN(n3507)
         );
  OR2_X2 U3521 ( .A1(n3467), .A2(n3466), .ZN(n5494) );
  AND4_X1 U3522 ( .A1(n3549), .A2(n3548), .A3(n3547), .A4(n3546), .ZN(n3550)
         );
  AND4_X1 U3523 ( .A1(n3456), .A2(n3455), .A3(n3454), .A4(n3453), .ZN(n3457)
         );
  AND4_X1 U3524 ( .A1(n3483), .A2(n3482), .A3(n3481), .A4(n3480), .ZN(n3484)
         );
  AND4_X1 U3525 ( .A1(n3471), .A2(n3470), .A3(n3469), .A4(n3468), .ZN(n3487)
         );
  AND4_X1 U3526 ( .A1(n3479), .A2(n3478), .A3(n3477), .A4(n3476), .ZN(n3485)
         );
  BUF_X2 U3527 ( .A(n4307), .Z(n4412) );
  INV_X2 U3528 ( .A(n4793), .ZN(n3427) );
  BUF_X2 U3529 ( .A(n3638), .Z(n4371) );
  BUF_X2 U3531 ( .A(n3691), .Z(n3627) );
  BUF_X2 U3532 ( .A(n3698), .Z(n4413) );
  BUF_X2 U3533 ( .A(n3543), .Z(n4342) );
  INV_X2 U3534 ( .A(n6474), .ZN(n6471) );
  AND2_X2 U3535 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4790) );
  NOR2_X4 U3536 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3451) );
  NAND2_X1 U3537 ( .A1(n3815), .A2(n3814), .ZN(n3838) );
  INV_X1 U3538 ( .A(n3818), .ZN(n3815) );
  BUF_X4 U3539 ( .A(n4443), .Z(n4831) );
  NOR2_X4 U3540 ( .A1(n5325), .A2(n5303), .ZN(n5302) );
  NAND2_X1 U3541 ( .A1(n4543), .A2(n3431), .ZN(n5184) );
  NAND2_X2 U3542 ( .A1(n3868), .A2(n3436), .ZN(n5539) );
  AND2_X4 U3543 ( .A1(n4750), .A2(n4798), .ZN(n3699) );
  NAND2_X1 U3544 ( .A1(n3582), .A2(n3581), .ZN(n3936) );
  AND2_X1 U3545 ( .A1(n3571), .A2(n3570), .ZN(n3593) );
  OR2_X1 U3546 ( .A1(n3633), .A2(n3632), .ZN(n3840) );
  NOR2_X1 U3547 ( .A1(n5491), .A2(n4831), .ZN(n4649) );
  AOI21_X1 U3548 ( .B1(n3658), .B2(n3665), .A(n3836), .ZN(n3677) );
  INV_X1 U3549 ( .A(n3882), .ZN(n4673) );
  NAND3_X1 U3550 ( .A1(n3529), .A2(n4673), .A3(n6780), .ZN(n4744) );
  NAND2_X1 U3551 ( .A1(n4843), .A2(n6449), .ZN(n4858) );
  AND2_X1 U3552 ( .A1(n3587), .A2(n4745), .ZN(n3606) );
  NAND2_X1 U3553 ( .A1(n6822), .A2(n3598), .ZN(n3937) );
  NAND2_X1 U3554 ( .A1(n5149), .A2(n4087), .ZN(n4100) );
  NAND2_X1 U3555 ( .A1(n5113), .A2(n5148), .ZN(n4091) );
  XNOR2_X1 U3556 ( .A(n3838), .B(n3828), .ZN(n3999) );
  INV_X1 U3557 ( .A(n6110), .ZN(n3854) );
  OR2_X1 U3558 ( .A1(n3648), .A2(n3647), .ZN(n3716) );
  NAND3_X1 U3559 ( .A1(n3595), .A2(n3594), .A3(n3593), .ZN(n3680) );
  NOR2_X1 U3560 ( .A1(n3675), .A2(n3674), .ZN(n3676) );
  NAND2_X1 U3561 ( .A1(n3708), .A2(n3707), .ZN(n3711) );
  OR2_X1 U3562 ( .A1(n4766), .A2(n4765), .ZN(n4772) );
  OR2_X1 U3563 ( .A1(n6633), .A2(n6632), .ZN(n6649) );
  NAND4_X2 U3564 ( .A1(n3553), .A2(n3552), .A3(n3551), .A4(n3550), .ZN(n4443)
         );
  AND4_X1 U3565 ( .A1(n3542), .A2(n3541), .A3(n3540), .A4(n3539), .ZN(n3551)
         );
  AND4_X1 U3566 ( .A1(n3534), .A2(n3533), .A3(n3532), .A4(n3531), .ZN(n3553)
         );
  NAND4_X1 U3567 ( .A1(n3508), .A2(n3507), .A3(n3506), .A4(n3505), .ZN(n3564)
         );
  AND4_X1 U3568 ( .A1(n3500), .A2(n3499), .A3(n3498), .A4(n3497), .ZN(n3506)
         );
  AND4_X1 U3569 ( .A1(n3492), .A2(n3491), .A3(n3490), .A4(n3489), .ZN(n3508)
         );
  AND4_X1 U3570 ( .A1(n3504), .A2(n3503), .A3(n3502), .A4(n3501), .ZN(n3505)
         );
  OR2_X1 U3571 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4425) );
  AND2_X2 U3572 ( .A1(n3530), .A2(n3529), .ZN(n4613) );
  NAND2_X1 U3573 ( .A1(n4300), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4321)
         );
  INV_X1 U3574 ( .A(n4299), .ZN(n4300) );
  INV_X1 U3575 ( .A(n4576), .ZN(n5198) );
  AND2_X1 U3576 ( .A1(n4474), .A2(n4473), .ZN(n4977) );
  OR2_X1 U3577 ( .A1(n4766), .A2(n4614), .ZN(n4679) );
  NOR2_X1 U3578 ( .A1(n4604), .A2(n4820), .ZN(n3978) );
  INV_X1 U3579 ( .A(n4819), .ZN(n3977) );
  NAND2_X1 U3580 ( .A1(n5288), .A2(n5281), .ZN(n5280) );
  NAND2_X1 U3581 ( .A1(n5280), .A2(n4645), .ZN(n5185) );
  NAND2_X1 U3582 ( .A1(n5531), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5208) );
  OR2_X1 U3583 ( .A1(n5737), .A2(n6230), .ZN(n5619) );
  AND2_X1 U3584 ( .A1(n5737), .A2(n6230), .ZN(n5620) );
  NAND2_X1 U3585 ( .A1(n5154), .A2(n5095), .ZN(n5180) );
  INV_X1 U3586 ( .A(n4744), .ZN(n3568) );
  NAND2_X1 U3587 ( .A1(n3933), .A2(n3932), .ZN(n5262) );
  OR2_X1 U3588 ( .A1(n3929), .A2(n3928), .ZN(n3933) );
  AND2_X1 U3589 ( .A1(n6440), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3939) );
  CLKBUF_X1 U3590 ( .A(n3750), .Z(n6147) );
  OR2_X1 U3591 ( .A1(n6119), .A2(n4437), .ZN(n6125) );
  OR2_X1 U3592 ( .A1(n3766), .A2(n3765), .ZN(n3791) );
  INV_X1 U3593 ( .A(n3877), .ZN(n4664) );
  OR2_X1 U3594 ( .A1(n3619), .A2(n3618), .ZN(n3715) );
  OR2_X1 U3595 ( .A1(n3608), .A2(n6491), .ZN(n3689) );
  NAND2_X1 U3596 ( .A1(n3878), .A2(n4681), .ZN(n3591) );
  OR2_X1 U3597 ( .A1(n4263), .A2(n5375), .ZN(n5376) );
  AND2_X1 U3598 ( .A1(n4776), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4422) );
  NOR2_X2 U3599 ( .A1(n5035), .A2(n5034), .ZN(n5033) );
  AND2_X1 U3600 ( .A1(n5619), .A2(n3861), .ZN(n3862) );
  INV_X1 U3601 ( .A(n4547), .ZN(n4524) );
  NAND2_X1 U3602 ( .A1(n3834), .A2(n3833), .ZN(n3844) );
  NAND2_X1 U3603 ( .A1(n4447), .A2(n4446), .ZN(n4451) );
  NAND2_X1 U3604 ( .A1(n4654), .A2(n3607), .ZN(n3959) );
  AND3_X1 U3605 ( .A1(n3606), .A2(n3605), .A3(n3604), .ZN(n3607) );
  NAND2_X1 U3606 ( .A1(n3596), .A2(n3680), .ZN(n3681) );
  XNOR2_X1 U3607 ( .A(n4598), .B(n6610), .ZN(n4789) );
  INV_X2 U3608 ( .A(n3918), .ZN(n3878) );
  OR2_X1 U3609 ( .A1(n3937), .A2(n4448), .ZN(n4745) );
  INV_X1 U3610 ( .A(n4613), .ZN(n4746) );
  INV_X1 U3611 ( .A(n6518), .ZN(n6583) );
  OAI21_X1 U3612 ( .B1(n6445), .B2(n6438), .A(n5248), .ZN(n6490) );
  AND2_X1 U3613 ( .A1(n4887), .A2(n6551), .ZN(n6575) );
  AND2_X1 U3614 ( .A1(n3664), .A2(n3654), .ZN(n3666) );
  NOR2_X1 U3615 ( .A1(n3937), .A2(n3565), .ZN(n3566) );
  XNOR2_X1 U3616 ( .A(n3681), .B(n3679), .ZN(n4741) );
  NAND2_X1 U3617 ( .A1(n5178), .A2(n4100), .ZN(n5357) );
  NAND2_X1 U3618 ( .A1(n5357), .A2(n5482), .ZN(n5481) );
  AND2_X1 U3619 ( .A1(n4322), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4323)
         );
  NAND2_X1 U3620 ( .A1(n4323), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4359)
         );
  NAND2_X1 U3621 ( .A1(n4282), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4299)
         );
  NAND2_X1 U3622 ( .A1(n4178), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4177)
         );
  NOR2_X1 U3623 ( .A1(n4214), .A2(n5613), .ZN(n4211) );
  NAND2_X1 U3624 ( .A1(n4211), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4210)
         );
  AND2_X1 U3625 ( .A1(n5470), .A2(n5469), .ZN(n5467) );
  AND2_X1 U3626 ( .A1(n4247), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4229)
         );
  NOR2_X1 U3627 ( .A1(n4093), .A2(n5164), .ZN(n4094) );
  NAND2_X1 U3628 ( .A1(n4094), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4265)
         );
  OAI21_X1 U3629 ( .B1(n4091), .B2(n4090), .A(n4089), .ZN(n4092) );
  NAND2_X1 U3630 ( .A1(n4099), .A2(n4098), .ZN(n5178) );
  INV_X1 U3631 ( .A(n5175), .ZN(n4098) );
  INV_X1 U3632 ( .A(n5176), .ZN(n4099) );
  NOR2_X1 U3633 ( .A1(n4045), .A2(n5119), .ZN(n4058) );
  NAND2_X1 U3634 ( .A1(n3995), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4015)
         );
  NOR2_X1 U3635 ( .A1(n3988), .A2(n6292), .ZN(n3995) );
  NAND2_X1 U3636 ( .A1(n3994), .A2(n3993), .ZN(n4974) );
  NAND2_X1 U3637 ( .A1(n3987), .A2(n4274), .ZN(n3994) );
  NAND2_X1 U3638 ( .A1(n4953), .A2(n4974), .ZN(n5003) );
  INV_X1 U3639 ( .A(n3980), .ZN(n3981) );
  NAND2_X1 U3640 ( .A1(n3981), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3988)
         );
  INV_X1 U3641 ( .A(n3945), .ZN(n3946) );
  AND3_X1 U3642 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A3(PHYADDRPOINTER_REG_3__SCAN_IN), 
        .ZN(n3948) );
  NAND2_X1 U3643 ( .A1(n4643), .A2(n4642), .ZN(n4784) );
  CLKBUF_X1 U3644 ( .A(n5565), .Z(n5566) );
  NAND2_X1 U3645 ( .A1(n5566), .A2(n5604), .ZN(n5735) );
  NOR2_X1 U3647 ( .A1(n3434), .A2(n3854), .ZN(n3855) );
  INV_X1 U3648 ( .A(n5181), .ZN(n4498) );
  INV_X1 U3649 ( .A(n5180), .ZN(n4499) );
  INV_X1 U3650 ( .A(n5126), .ZN(n4490) );
  INV_X1 U3651 ( .A(n4976), .ZN(n4476) );
  OR2_X1 U3652 ( .A1(n4858), .A2(n5258), .ZN(n6179) );
  OR2_X1 U3653 ( .A1(n4637), .A2(n5763), .ZN(n4875) );
  XNOR2_X1 U3654 ( .A(n3678), .B(n3677), .ZN(n4886) );
  AND2_X2 U3655 ( .A1(n4753), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4750)
         );
  INV_X1 U3656 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4753) );
  NAND3_X1 U3657 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6491), .A3(n6490), .ZN(
        n6966) );
  NOR2_X1 U3658 ( .A1(n6561), .A2(n6584), .ZN(n6496) );
  INV_X1 U3659 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5057) );
  INV_X1 U3660 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6292) );
  OR2_X1 U3661 ( .A1(n6150), .A2(n4564), .ZN(n6283) );
  NAND2_X1 U3662 ( .A1(n5198), .A2(n4580), .ZN(n6301) );
  CLKBUF_X1 U3663 ( .A(n4741), .Z(n4742) );
  AND2_X1 U3664 ( .A1(n6283), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6370) );
  INV_X1 U3665 ( .A(n6334), .ZN(n6389) );
  INV_X1 U3666 ( .A(n5479), .ZN(n6082) );
  AND2_X1 U3667 ( .A1(n4668), .A2(n6449), .ZN(n6086) );
  NAND2_X1 U3668 ( .A1(n6086), .A2(n6965), .ZN(n5479) );
  AND2_X1 U3669 ( .A1(n5520), .A2(n5495), .ZN(n6687) );
  NAND2_X1 U3670 ( .A1(n4680), .A2(n4679), .ZN(n5520) );
  INV_X1 U3671 ( .A(n4679), .ZN(n4736) );
  OR2_X1 U3672 ( .A1(n4567), .A2(n4566), .ZN(n4568) );
  AND2_X1 U3673 ( .A1(n5458), .A2(n5457), .ZN(n6479) );
  XOR2_X1 U3674 ( .A(n5188), .B(n5187), .Z(n5234) );
  OAI21_X1 U3675 ( .B1(n5280), .B2(n5186), .A(n5185), .ZN(n5187) );
  XNOR2_X1 U3676 ( .A(n5214), .B(n5229), .ZN(n5242) );
  NAND2_X1 U3677 ( .A1(n5213), .A2(n3438), .ZN(n5214) );
  AND2_X1 U3678 ( .A1(n5208), .A2(n5207), .ZN(n5213) );
  BUF_X1 U3679 ( .A(n5539), .Z(n5541) );
  OR2_X1 U3680 ( .A1(n5721), .A2(n5226), .ZN(n5703) );
  CLKBUF_X1 U3681 ( .A(n5622), .Z(n5623) );
  INV_X1 U3682 ( .A(n6215), .ZN(n6233) );
  OR2_X1 U3683 ( .A1(n4858), .A2(n4857), .ZN(n6224) );
  INV_X1 U3684 ( .A(n6225), .ZN(n6244) );
  INV_X1 U3685 ( .A(n6585), .ZN(n6537) );
  OR2_X1 U3686 ( .A1(n3744), .A2(n6560), .ZN(n3745) );
  OR2_X1 U3687 ( .A1(n5262), .A2(n6678), .ZN(n5248) );
  INV_X1 U3688 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6404) );
  INV_X1 U3689 ( .A(n7036), .ZN(n7039) );
  AND2_X1 U3690 ( .A1(n6597), .A2(n6634), .ZN(n7031) );
  OR2_X1 U3691 ( .A1(n6526), .A2(n6634), .ZN(n6924) );
  INV_X1 U3692 ( .A(n6984), .ZN(n6913) );
  INV_X1 U3693 ( .A(n6869), .ZN(n6975) );
  INV_X1 U3694 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6440) );
  OR2_X1 U3695 ( .A1(n5243), .A2(n6862), .ZN(n4440) );
  NAND2_X1 U3696 ( .A1(n5652), .A2(n6121), .ZN(n4441) );
  INV_X2 U3697 ( .A(n3851), .ZN(n5748) );
  NAND2_X2 U3698 ( .A1(n3838), .A2(n3837), .ZN(n3851) );
  INV_X1 U3699 ( .A(n4455), .ZN(n4670) );
  INV_X2 U3700 ( .A(n4670), .ZN(n4518) );
  NAND2_X1 U3701 ( .A1(n6908), .A2(n5494), .ZN(n4662) );
  NOR3_X2 U3702 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6667), .ZN(n7063) );
  INV_X1 U3703 ( .A(n6369), .ZN(n6382) );
  NOR2_X4 U3704 ( .A1(n4576), .A2(n4572), .ZN(n6369) );
  XNOR2_X1 U3705 ( .A(n5272), .B(n5190), .ZN(n5243) );
  NAND2_X1 U3706 ( .A1(n5737), .A2(n3858), .ZN(n3433) );
  AND2_X1 U3707 ( .A1(n5737), .A2(n5215), .ZN(n3434) );
  NOR2_X1 U3708 ( .A1(n6574), .A2(n6573), .ZN(n3435) );
  NAND2_X1 U3709 ( .A1(n5737), .A2(n5693), .ZN(n3436) );
  NAND2_X1 U3710 ( .A1(n4451), .A2(n4450), .ZN(n4456) );
  INV_X1 U3711 ( .A(n4644), .ZN(n3581) );
  NOR2_X1 U3712 ( .A1(n6604), .A2(n6632), .ZN(n3437) );
  AND2_X1 U3713 ( .A1(n5212), .A2(n5211), .ZN(n3438) );
  AND2_X1 U3714 ( .A1(n6112), .A2(n6108), .ZN(n3439) );
  OR2_X1 U3715 ( .A1(n5653), .A2(n6389), .ZN(n3440) );
  INV_X4 U3716 ( .A(n5748), .ZN(n5737) );
  AND4_X1 U3717 ( .A1(n3450), .A2(n3449), .A3(n3448), .A4(n3447), .ZN(n3441)
         );
  AND3_X1 U3718 ( .A1(n3527), .A2(n3526), .A3(n3525), .ZN(n3442) );
  AND3_X1 U3719 ( .A1(n3645), .A2(n3644), .A3(n3643), .ZN(n3443) );
  NAND2_X1 U3720 ( .A1(n6864), .A2(n6732), .ZN(n3575) );
  AND4_X1 U3721 ( .A1(n3524), .A2(n3523), .A3(n3522), .A4(n3521), .ZN(n3444)
         );
  AND2_X2 U3722 ( .A1(n5033), .A2(n4028), .ZN(n3445) );
  INV_X1 U3723 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3875) );
  NAND2_X1 U3724 ( .A1(n3744), .A2(n6560), .ZN(n3756) );
  INV_X1 U3725 ( .A(n5491), .ZN(n3567) );
  NAND2_X1 U3726 ( .A1(n6491), .A2(n6490), .ZN(n6963) );
  OAI21_X1 U3727 ( .B1(n3937), .B2(n6732), .A(n3575), .ZN(n3576) );
  AND2_X1 U3728 ( .A1(n3882), .A2(n3883), .ZN(n3903) );
  NOR2_X1 U3729 ( .A1(n4837), .A2(n6458), .ZN(n3583) );
  OAI21_X1 U3730 ( .B1(n4681), .B2(n3608), .A(n3585), .ZN(n4646) );
  INV_X1 U3731 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4445) );
  NOR2_X1 U3732 ( .A1(n3595), .A2(n3573), .ZN(n3574) );
  NAND2_X1 U3733 ( .A1(n4662), .A2(n3488), .ZN(n3585) );
  BUF_X1 U3734 ( .A(n3513), .Z(n3690) );
  INV_X1 U3735 ( .A(n4281), .ZN(n4282) );
  OR2_X1 U3736 ( .A1(n3812), .A2(n3811), .ZN(n3830) );
  OR2_X1 U3737 ( .A1(n3788), .A2(n3787), .ZN(n3794) );
  OR2_X1 U3738 ( .A1(n3706), .A2(n3705), .ZN(n3746) );
  NAND2_X1 U3740 ( .A1(n6691), .A2(n6492), .ZN(n3882) );
  OR2_X1 U3741 ( .A1(n4831), .A2(n6491), .ZN(n3688) );
  NAND2_X1 U3742 ( .A1(n3878), .A2(n3877), .ZN(n3927) );
  AND2_X1 U3743 ( .A1(n4360), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4361)
         );
  OR2_X1 U3744 ( .A1(n5494), .A2(n6657), .ZN(n4399) );
  AND2_X1 U3745 ( .A1(n5580), .A2(n3862), .ZN(n5565) );
  AND2_X1 U3746 ( .A1(n5024), .A2(n3845), .ZN(n3848) );
  NAND2_X1 U3747 ( .A1(n3568), .A2(n3567), .ZN(n4854) );
  AND3_X1 U3748 ( .A1(n3637), .A2(n3636), .A3(n3635), .ZN(n3673) );
  OR2_X1 U3749 ( .A1(n3741), .A2(n3740), .ZN(n3771) );
  INV_X1 U3750 ( .A(n3575), .ZN(n3529) );
  AND2_X1 U3751 ( .A1(n4588), .A2(n5203), .ZN(n4589) );
  INV_X1 U3752 ( .A(n4177), .ZN(n4125) );
  INV_X1 U3753 ( .A(n5116), .ZN(n4489) );
  NAND2_X1 U3754 ( .A1(n4670), .A2(n4448), .ZN(n4539) );
  NAND2_X1 U3755 ( .A1(n3689), .A2(n3688), .ZN(n3931) );
  NAND2_X1 U3756 ( .A1(n4361), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4428)
         );
  AND2_X1 U3757 ( .A1(n4279), .A2(n5482), .ZN(n4280) );
  INV_X1 U3758 ( .A(n4422), .ZN(n4380) );
  NOR2_X1 U3759 ( .A1(n4265), .A2(n6337), .ZN(n4247) );
  AOI21_X1 U3760 ( .B1(n3999), .B2(n4274), .A(n3998), .ZN(n5002) );
  INV_X1 U3761 ( .A(n3940), .ZN(n3947) );
  OR2_X1 U3762 ( .A1(n5230), .A2(n5237), .ZN(n5231) );
  NAND2_X1 U3763 ( .A1(n4499), .A2(n4498), .ZN(n5484) );
  INV_X1 U3764 ( .A(n4977), .ZN(n4475) );
  INV_X1 U3765 ( .A(n4938), .ZN(n4469) );
  NAND2_X1 U3766 ( .A1(n3687), .A2(n3686), .ZN(n3723) );
  AND2_X1 U3767 ( .A1(n4772), .A2(n4771), .ZN(n4842) );
  NAND2_X1 U3768 ( .A1(n3731), .A2(n3730), .ZN(n6610) );
  INV_X1 U3769 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6621) );
  NAND2_X1 U3770 ( .A1(n4789), .A2(n6491), .ZN(n3743) );
  AOI21_X1 U3771 ( .B1(n3652), .B2(n3716), .A(n3651), .ZN(n3664) );
  NOR2_X1 U3772 ( .A1(n4590), .A2(n4589), .ZN(n4591) );
  AND2_X1 U3773 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n4125), .ZN(n4141)
         );
  NOR2_X1 U3774 ( .A1(n4015), .A2(n5057), .ZN(n4029) );
  NAND2_X1 U3775 ( .A1(n3948), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3980)
         );
  NAND2_X1 U3776 ( .A1(n6283), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4576) );
  INV_X1 U3777 ( .A(n4550), .ZN(n4551) );
  NAND2_X1 U3778 ( .A1(n4490), .A2(n4489), .ZN(n5153) );
  NOR2_X1 U3779 ( .A1(n5315), .A2(n5317), .ZN(n5300) );
  OR2_X1 U3780 ( .A1(n5262), .A2(READY_N), .ZN(n4766) );
  OR2_X1 U3781 ( .A1(n4428), .A2(n5276), .ZN(n4567) );
  NAND2_X1 U3782 ( .A1(n5357), .A2(n4280), .ZN(n5361) );
  NAND2_X1 U3783 ( .A1(n4229), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4214)
         );
  AND2_X1 U3784 ( .A1(n3978), .A2(n3977), .ZN(n4952) );
  NOR2_X1 U3785 ( .A1(n5232), .A2(n5231), .ZN(n5233) );
  AND2_X1 U3786 ( .A1(n5530), .A2(n3870), .ZN(n5522) );
  NOR2_X2 U3787 ( .A1(n5486), .A2(n5415), .ZN(n5472) );
  NOR2_X1 U3788 ( .A1(n6164), .A2(n6162), .ZN(n6215) );
  AND2_X1 U3789 ( .A1(n4488), .A2(n4487), .ZN(n5116) );
  NOR2_X2 U3790 ( .A1(n4979), .A2(n4980), .ZN(n5027) );
  NAND2_X1 U3791 ( .A1(n4470), .A2(n4469), .ZN(n4976) );
  NAND2_X1 U3792 ( .A1(n3775), .A2(n3774), .ZN(n3778) );
  OR2_X1 U3793 ( .A1(n4858), .A2(n4890), .ZN(n5765) );
  AND2_X1 U3794 ( .A1(n4773), .A2(n4842), .ZN(n6410) );
  OR2_X1 U3795 ( .A1(n4887), .A2(n6551), .ZN(n6665) );
  INV_X1 U3796 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6647) );
  NAND2_X1 U3797 ( .A1(n3743), .A2(n3742), .ZN(n6560) );
  INV_X1 U3798 ( .A(n4425), .ZN(n4562) );
  NAND2_X1 U3799 ( .A1(n4613), .A2(n4831), .ZN(n5263) );
  OAI21_X1 U3800 ( .B1(n5243), .B2(n6390), .A(n4591), .ZN(n4592) );
  NAND2_X1 U3801 ( .A1(n4141), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4281)
         );
  AND2_X1 U3802 ( .A1(n6283), .A2(n4569), .ZN(n6375) );
  INV_X1 U3803 ( .A(n6370), .ZN(n6384) );
  AND2_X1 U3804 ( .A1(n6254), .A2(n4670), .ZN(n6334) );
  AND2_X2 U3805 ( .A1(n5302), .A2(n5286), .ZN(n5288) );
  NAND2_X1 U3806 ( .A1(n5025), .A2(n5127), .ZN(n5126) );
  CLKBUF_X1 U3807 ( .A(n4594), .Z(n4939) );
  INV_X1 U3808 ( .A(n5520), .ZN(n6686) );
  NOR2_X1 U3809 ( .A1(n5481), .A2(n5413), .ZN(n5470) );
  INV_X1 U3810 ( .A(n4443), .ZN(n6492) );
  XNOR2_X1 U3811 ( .A(n5194), .B(n5193), .ZN(n5490) );
  INV_X1 U3812 ( .A(n6120), .ZN(n6482) );
  NOR2_X1 U3813 ( .A1(n4210), .A2(n5605), .ZN(n4178) );
  INV_X1 U3814 ( .A(n4091), .ZN(n5149) );
  INV_X1 U3815 ( .A(n6125), .ZN(n6104) );
  INV_X1 U3816 ( .A(n6397), .ZN(n6121) );
  NOR2_X1 U3817 ( .A1(n5765), .A2(n5093), .ZN(n6162) );
  XNOR2_X1 U3818 ( .A(n3844), .B(n3835), .ZN(n5019) );
  CLKBUF_X1 U3819 ( .A(n4933), .Z(n4937) );
  INV_X1 U3820 ( .A(n6224), .ZN(n6243) );
  INV_X1 U3821 ( .A(n6179), .ZN(n5089) );
  INV_X1 U3822 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4807) );
  INV_X1 U3823 ( .A(n6956), .ZN(n7067) );
  INV_X1 U3824 ( .A(n6649), .ZN(n6646) );
  INV_X1 U3825 ( .A(n6947), .ZN(n7051) );
  AND3_X1 U3826 ( .A1(n6585), .A2(n6584), .A3(n6583), .ZN(n6597) );
  AND2_X1 U3827 ( .A1(n6571), .A2(n6645), .ZN(n7018) );
  INV_X1 U3828 ( .A(n7023), .ZN(n7012) );
  INV_X1 U3829 ( .A(n7016), .ZN(n7004) );
  INV_X1 U3830 ( .A(n6924), .ZN(n6998) );
  INV_X1 U3831 ( .A(n6916), .ZN(n6987) );
  AND2_X1 U3832 ( .A1(n6432), .A2(n6431), .ZN(n6443) );
  OR3_X1 U3833 ( .A1(n5262), .A2(n5263), .A3(n6428), .ZN(n4612) );
  NAND2_X1 U3834 ( .A1(n4612), .A2(n4610), .ZN(n6150) );
  INV_X1 U3835 ( .A(n4592), .ZN(n4593) );
  NAND2_X1 U3836 ( .A1(n6283), .A2(n4573), .ZN(n6395) );
  OR2_X1 U3837 ( .A1(n5452), .A2(n5451), .ZN(n6120) );
  INV_X1 U3838 ( .A(n5587), .ZN(n5513) );
  OR2_X1 U3839 ( .A1(n5414), .A2(n5470), .ZN(n5637) );
  NOR2_X1 U3840 ( .A1(n6152), .A2(n4623), .ZN(n5777) );
  OR3_X1 U3841 ( .A1(n5262), .A2(n4621), .A3(n4620), .ZN(n6007) );
  AOI21_X1 U3842 ( .B1(n5490), .B2(n6969), .A(n5240), .ZN(n5241) );
  OR2_X1 U3843 ( .A1(n5436), .A2(n5435), .ZN(n6391) );
  OAI21_X1 U3844 ( .B1(n5467), .B2(n5403), .A(n5456), .ZN(n5618) );
  OR2_X1 U3845 ( .A1(n6419), .A2(n6428), .ZN(n6397) );
  INV_X1 U3846 ( .A(n5235), .ZN(n5236) );
  OR2_X1 U3847 ( .A1(n4858), .A2(n4849), .ZN(n6225) );
  NAND2_X1 U3848 ( .A1(n6646), .A2(n6634), .ZN(n7062) );
  NAND2_X1 U3849 ( .A1(n3437), .A2(n6645), .ZN(n6947) );
  NAND2_X1 U3850 ( .A1(n3437), .A2(n6634), .ZN(n7048) );
  INV_X1 U3851 ( .A(n7018), .ZN(n7029) );
  OR2_X1 U3852 ( .A1(n6550), .A2(n6634), .ZN(n7016) );
  OR2_X1 U3853 ( .A1(n6550), .A2(n6645), .ZN(n7009) );
  OR2_X1 U3854 ( .A1(n6526), .A2(n6645), .ZN(n6996) );
  NAND2_X1 U3855 ( .A1(n6510), .A2(n6645), .ZN(n6916) );
  NAND2_X1 U3856 ( .A1(n6496), .A2(n6634), .ZN(n7072) );
  INV_X1 U3857 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6491) );
  INV_X1 U3858 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3446) );
  AND2_X2 U3859 ( .A1(n3446), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4791)
         );
  AND2_X2 U3860 ( .A1(n4791), .A2(n4750), .ZN(n3513) );
  BUF_X2 U3861 ( .A(n3513), .Z(n4307) );
  NOR2_X4 U3862 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4799) );
  AND2_X4 U3863 ( .A1(n4750), .A2(n4799), .ZN(n4366) );
  AOI22_X1 U3864 ( .A1(n4307), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4366), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3450) );
  AND2_X2 U3865 ( .A1(n3452), .A2(n4790), .ZN(n3609) );
  AND2_X2 U3866 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4798) );
  AOI22_X1 U3867 ( .A1(n3609), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3699), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3449) );
  AND2_X2 U3868 ( .A1(n3452), .A2(n4750), .ZN(n3696) );
  AOI22_X1 U3869 ( .A1(n3696), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3448) );
  AND2_X2 U3870 ( .A1(n4791), .A2(n4790), .ZN(n3543) );
  AND2_X2 U3871 ( .A1(n3451), .A2(n4798), .ZN(n3545) );
  AOI22_X1 U3872 ( .A1(n3543), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3447) );
  AND2_X2 U3873 ( .A1(n4749), .A2(n4798), .ZN(n4000) );
  AOI22_X1 U3874 ( .A1(n4000), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3691), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3456) );
  AND2_X2 U3875 ( .A1(n4749), .A2(n3452), .ZN(n3697) );
  AND2_X2 U3876 ( .A1(n4791), .A2(n3451), .ZN(n3698) );
  AOI22_X1 U3877 ( .A1(n3697), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3698), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3455) );
  AND2_X2 U3878 ( .A1(n3452), .A2(n3451), .ZN(n3700) );
  AND2_X4 U3879 ( .A1(n4799), .A2(n4790), .ZN(n4388) );
  AOI22_X1 U3880 ( .A1(n3700), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3454) );
  AND2_X2 U3881 ( .A1(n4749), .A2(n4791), .ZN(n3638) );
  AND2_X4 U3882 ( .A1(n4798), .A2(n4790), .ZN(n4383) );
  AOI22_X1 U3883 ( .A1(n3638), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3453) );
  AND2_X2 U3884 ( .A1(n3441), .A2(n3457), .ZN(n6908) );
  AOI22_X1 U3885 ( .A1(n4000), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3691), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3461) );
  AOI22_X1 U3886 ( .A1(n3700), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3698), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3460) );
  AOI22_X1 U3887 ( .A1(n3543), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3459) );
  AOI22_X1 U3888 ( .A1(n3638), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3458) );
  NAND4_X1 U3889 ( .A1(n3461), .A2(n3460), .A3(n3459), .A4(n3458), .ZN(n3467)
         );
  AOI22_X1 U3890 ( .A1(n3513), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4366), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3465) );
  AOI22_X1 U3891 ( .A1(n3609), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3699), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3464) );
  AOI22_X1 U3892 ( .A1(n3696), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3463) );
  AOI22_X1 U3893 ( .A1(n3697), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3462) );
  NAND4_X1 U3894 ( .A1(n3465), .A2(n3464), .A3(n3463), .A4(n3462), .ZN(n3466)
         );
  NAND2_X1 U3895 ( .A1(n4000), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3471)
         );
  NAND2_X1 U3896 ( .A1(n3691), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3470) );
  NAND2_X1 U3897 ( .A1(n3697), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3469) );
  NAND2_X1 U3898 ( .A1(n3700), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3468) );
  NAND2_X1 U3899 ( .A1(n3609), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3475) );
  NAND2_X1 U3900 ( .A1(n3690), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3474) );
  NAND2_X1 U3901 ( .A1(n3696), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3473) );
  NAND2_X1 U3902 ( .A1(n3543), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3472)
         );
  NAND2_X1 U3903 ( .A1(n3699), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3479)
         );
  NAND2_X1 U3904 ( .A1(n4366), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3478) );
  NAND2_X1 U3905 ( .A1(n3544), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3477) );
  NAND2_X1 U3906 ( .A1(n3545), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3476)
         );
  NAND2_X1 U3907 ( .A1(n3638), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3483)
         );
  NAND2_X1 U3908 ( .A1(n3698), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3482) );
  NAND2_X1 U3909 ( .A1(n4388), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3481) );
  NAND2_X1 U3910 ( .A1(n4383), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3480)
         );
  NAND2_X1 U3911 ( .A1(n3598), .A2(n5494), .ZN(n3488) );
  NAND2_X1 U3912 ( .A1(n3696), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3492) );
  NAND2_X1 U3913 ( .A1(n3543), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3491)
         );
  NAND2_X1 U3914 ( .A1(n3544), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3490) );
  NAND2_X1 U3915 ( .A1(n3545), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3489)
         );
  NAND2_X1 U3916 ( .A1(n3690), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3496) );
  NAND2_X1 U3917 ( .A1(n4366), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3495) );
  NAND2_X1 U3918 ( .A1(n3609), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3494) );
  NAND2_X1 U3919 ( .A1(n3699), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3493)
         );
  NAND2_X1 U3920 ( .A1(n3638), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3500)
         );
  NAND2_X1 U3921 ( .A1(n3700), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3499) );
  NAND2_X1 U3922 ( .A1(n4388), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3498) );
  NAND2_X1 U3923 ( .A1(n4383), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3497)
         );
  NAND2_X1 U3924 ( .A1(n4000), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3504)
         );
  NAND2_X1 U3925 ( .A1(n3691), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3503) );
  NAND2_X1 U3926 ( .A1(n3697), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3502) );
  NAND2_X1 U3927 ( .A1(n3698), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3501) );
  NAND2_X1 U3928 ( .A1(n4681), .A2(n3608), .ZN(n3520) );
  AOI22_X1 U3929 ( .A1(n3609), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4366), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3512) );
  AOI22_X1 U3930 ( .A1(n3700), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3698), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3511) );
  AOI22_X1 U3931 ( .A1(n3691), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3510) );
  AOI22_X1 U3932 ( .A1(n3543), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3509) );
  NAND4_X1 U3933 ( .A1(n3512), .A2(n3511), .A3(n3510), .A4(n3509), .ZN(n3519)
         );
  AOI22_X1 U3934 ( .A1(n4000), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3696), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3517) );
  AOI22_X1 U3935 ( .A1(n3513), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3699), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3516) );
  AOI22_X1 U3936 ( .A1(n3697), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3515) );
  AOI22_X1 U3937 ( .A1(n3638), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3514) );
  NAND4_X1 U3938 ( .A1(n3517), .A2(n3516), .A3(n3515), .A4(n3514), .ZN(n3518)
         );
  NAND3_X1 U3939 ( .A1(n3585), .A2(n3520), .A3(n4656), .ZN(n3600) );
  INV_X1 U3940 ( .A(n3600), .ZN(n3530) );
  AOI22_X1 U3941 ( .A1(n4000), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3691), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3524) );
  AOI22_X1 U3942 ( .A1(n3697), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3698), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3523) );
  AOI22_X1 U3943 ( .A1(n3700), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3522) );
  AOI22_X1 U3944 ( .A1(n3638), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3521) );
  AOI22_X1 U3945 ( .A1(n3543), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3527) );
  AOI22_X1 U3946 ( .A1(n3696), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3526) );
  AOI22_X1 U3947 ( .A1(n3609), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3699), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3525) );
  AOI22_X1 U3948 ( .A1(n4307), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4366), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3528) );
  AND3_X2 U3949 ( .A1(n3444), .A2(n3442), .A3(n3528), .ZN(n6732) );
  NAND2_X1 U3950 ( .A1(n4000), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3534)
         );
  NAND2_X1 U3951 ( .A1(n3691), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3533) );
  NAND2_X1 U3952 ( .A1(n3697), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3532) );
  NAND2_X1 U3953 ( .A1(n3698), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3531) );
  NAND2_X1 U3954 ( .A1(n3690), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3538) );
  NAND2_X1 U3955 ( .A1(n4366), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3537) );
  NAND2_X1 U3956 ( .A1(n3609), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3536) );
  NAND2_X1 U3957 ( .A1(n3699), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3535)
         );
  AND4_X2 U3958 ( .A1(n3538), .A2(n3537), .A3(n3536), .A4(n3535), .ZN(n3552)
         );
  NAND2_X1 U3959 ( .A1(n3638), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3542)
         );
  NAND2_X1 U3960 ( .A1(n3700), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3541) );
  NAND2_X1 U3961 ( .A1(n4388), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3540) );
  NAND2_X1 U3962 ( .A1(n4383), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3539)
         );
  NAND2_X1 U3963 ( .A1(n3696), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3549) );
  NAND2_X1 U3964 ( .A1(n3543), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3548)
         );
  NAND2_X1 U3965 ( .A1(n3544), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3547) );
  NAND2_X1 U3966 ( .A1(n3545), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3546)
         );
  AOI22_X1 U3967 ( .A1(n4000), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3700), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3557) );
  AOI22_X1 U3968 ( .A1(n4366), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3543), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3556) );
  AOI22_X1 U3969 ( .A1(n3691), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3555) );
  AOI22_X1 U3970 ( .A1(n3696), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3554) );
  NAND4_X1 U3971 ( .A1(n3557), .A2(n3556), .A3(n3555), .A4(n3554), .ZN(n3563)
         );
  AOI22_X1 U3972 ( .A1(n3690), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3609), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3561) );
  AOI22_X1 U3973 ( .A1(n3699), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3698), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3560) );
  AOI22_X1 U3974 ( .A1(n3697), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3559) );
  AOI22_X1 U3975 ( .A1(n3638), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3558) );
  NAND4_X1 U3976 ( .A1(n3561), .A2(n3560), .A3(n3559), .A4(n3558), .ZN(n3562)
         );
  INV_X1 U3977 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6140) );
  XNOR2_X1 U3978 ( .A(n6140), .B(STATE_REG_2__SCAN_IN), .ZN(n6458) );
  INV_X2 U3979 ( .A(n3564), .ZN(n6822) );
  NAND2_X1 U3980 ( .A1(n6780), .A2(n4839), .ZN(n3565) );
  INV_X2 U3981 ( .A(n6908), .ZN(n3941) );
  NAND2_X2 U3982 ( .A1(n3941), .A2(n5494), .ZN(n5491) );
  NAND2_X1 U3983 ( .A1(n3566), .A2(n4649), .ZN(n5264) );
  OR2_X2 U3984 ( .A1(n5264), .A2(n4837), .ZN(n4901) );
  INV_X2 U3985 ( .A(n4444), .ZN(n6691) );
  OAI211_X1 U3986 ( .C1(n5263), .C2(n3583), .A(n4901), .B(n4854), .ZN(n3569)
         );
  NAND2_X1 U3987 ( .A1(n3569), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3595) );
  NOR2_X1 U3988 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6434) );
  NAND2_X1 U3989 ( .A1(n6434), .A2(n6491), .ZN(n4433) );
  NAND2_X1 U3990 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6620) );
  OAI21_X1 U3991 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n6620), .ZN(n6606) );
  OR2_X1 U3992 ( .A1(n4433), .A2(n6606), .ZN(n3571) );
  INV_X1 U3993 ( .A(n3939), .ZN(n3728) );
  NAND2_X1 U3994 ( .A1(n3728), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3570) );
  INV_X1 U3995 ( .A(n3593), .ZN(n3572) );
  NOR2_X1 U3996 ( .A1(n3572), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3573)
         );
  INV_X1 U3997 ( .A(n3574), .ZN(n3596) );
  NAND2_X1 U3998 ( .A1(n3576), .A2(n3567), .ZN(n3578) );
  INV_X1 U3999 ( .A(n4662), .ZN(n3577) );
  NAND3_X1 U4000 ( .A1(n3577), .A2(n3608), .A3(n6732), .ZN(n4665) );
  NAND2_X1 U4001 ( .A1(n3578), .A2(n4665), .ZN(n3579) );
  AOI21_X1 U4002 ( .B1(n4681), .B2(n4656), .A(n4444), .ZN(n3603) );
  NAND2_X1 U4003 ( .A1(n3579), .A2(n3603), .ZN(n3580) );
  NAND2_X1 U4004 ( .A1(n3580), .A2(n6492), .ZN(n3599) );
  INV_X1 U4005 ( .A(n4646), .ZN(n3582) );
  NAND2_X1 U4006 ( .A1(n6732), .A2(n4656), .ZN(n4644) );
  INV_X1 U4007 ( .A(n3936), .ZN(n3589) );
  INV_X1 U4008 ( .A(n3583), .ZN(n3584) );
  NAND2_X1 U4009 ( .A1(n3584), .A2(n6864), .ZN(n3588) );
  NAND2_X1 U4010 ( .A1(n3585), .A2(n6822), .ZN(n4650) );
  NAND2_X1 U4011 ( .A1(n6691), .A2(n4443), .ZN(n3659) );
  INV_X1 U4012 ( .A(n3659), .ZN(n3750) );
  NAND2_X1 U4013 ( .A1(n4650), .A2(n3750), .ZN(n3587) );
  NAND2_X2 U4014 ( .A1(n3586), .A2(n4444), .ZN(n4448) );
  NAND4_X1 U4015 ( .A1(n3599), .A2(n3589), .A3(n3588), .A4(n3606), .ZN(n3590)
         );
  NAND2_X1 U4016 ( .A1(n3590), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3592) );
  NAND2_X1 U4017 ( .A1(n3592), .A2(n3591), .ZN(n3683) );
  NAND2_X1 U4018 ( .A1(n3683), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3594) );
  NAND2_X1 U4019 ( .A1(n3683), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3597) );
  MUX2_X1 U4020 ( .A(n3939), .B(n4433), .S(n6647), .Z(n3653) );
  NAND2_X1 U4021 ( .A1(n3597), .A2(n3653), .ZN(n3961) );
  AND2_X2 U4022 ( .A1(n4837), .A2(n3934), .ZN(n3877) );
  NOR2_X1 U4023 ( .A1(n4664), .A2(n3608), .ZN(n4660) );
  OR2_X1 U4024 ( .A1(n3599), .A2(n4660), .ZN(n4654) );
  NAND2_X1 U4025 ( .A1(n6434), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3601) );
  AOI21_X1 U4026 ( .B1(n3600), .B2(n4837), .A(n3601), .ZN(n3605) );
  OAI21_X1 U4027 ( .B1(n4665), .B2(n4656), .A(n6492), .ZN(n3602) );
  OAI21_X1 U4028 ( .B1(n3603), .B2(n4839), .A(n3602), .ZN(n3604) );
  INV_X1 U4029 ( .A(n3689), .ZN(n3620) );
  INV_X1 U4030 ( .A(n3609), .ZN(n4793) );
  AOI22_X1 U4031 ( .A1(n4412), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3427), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3613) );
  AOI22_X1 U4032 ( .A1(n3429), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3627), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3612) );
  AOI22_X1 U4033 ( .A1(n4405), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3611) );
  AOI22_X1 U4034 ( .A1(n3622), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3610) );
  NAND4_X1 U4035 ( .A1(n3613), .A2(n3612), .A3(n3611), .A4(n3610), .ZN(n3619)
         );
  AOI22_X1 U4036 ( .A1(n4366), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4342), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3617) );
  AOI22_X1 U4037 ( .A1(n3430), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3616) );
  AOI22_X1 U4038 ( .A1(n4413), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3615) );
  AOI22_X1 U4039 ( .A1(n4371), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4301), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3614) );
  NAND4_X1 U4040 ( .A1(n3617), .A2(n3616), .A3(n3615), .A4(n3614), .ZN(n3618)
         );
  NAND2_X1 U4041 ( .A1(n3620), .A2(n3715), .ZN(n3621) );
  OAI21_X2 U4042 ( .B1(n4741), .B2(STATE2_REG_0__SCAN_IN), .A(n3621), .ZN(
        n3675) );
  NAND2_X1 U4043 ( .A1(n3878), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3637) );
  BUF_X1 U4044 ( .A(n4366), .Z(n4306) );
  AOI22_X1 U4045 ( .A1(n4307), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3626) );
  AOI22_X1 U4046 ( .A1(n3427), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3622), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3625) );
  AOI22_X1 U4047 ( .A1(n3430), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3624) );
  AOI22_X1 U4048 ( .A1(n4342), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3623) );
  NAND4_X1 U4049 ( .A1(n3626), .A2(n3625), .A3(n3624), .A4(n3623), .ZN(n3633)
         );
  AOI22_X1 U4050 ( .A1(n3429), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3627), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3631) );
  AOI22_X1 U4051 ( .A1(n4405), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3630) );
  AOI22_X1 U4052 ( .A1(n3428), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3629) );
  AOI22_X1 U4053 ( .A1(n4371), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4301), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3628) );
  NAND4_X1 U4054 ( .A1(n3631), .A2(n3630), .A3(n3629), .A4(n3628), .ZN(n3632)
         );
  NOR2_X1 U4055 ( .A1(n3689), .A2(n3840), .ZN(n3652) );
  INV_X1 U4056 ( .A(n3652), .ZN(n3636) );
  INV_X1 U4057 ( .A(n3688), .ZN(n3634) );
  NAND2_X1 U4058 ( .A1(n3634), .A2(n3715), .ZN(n3635) );
  XNOR2_X2 U4059 ( .A(n3675), .B(n3673), .ZN(n3678) );
  AOI22_X1 U4060 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n4405), .B1(n3429), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3642) );
  AOI22_X1 U4061 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n3638), .B1(n3428), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3641) );
  AOI22_X1 U4062 ( .A1(n3430), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3622), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3640) );
  AOI22_X1 U4063 ( .A1(n3627), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3639) );
  NAND4_X1 U4064 ( .A1(n3642), .A2(n3641), .A3(n3640), .A4(n3639), .ZN(n3648)
         );
  AOI22_X1 U4065 ( .A1(n4412), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4366), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3646) );
  AOI22_X1 U4066 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4413), .B1(n4407), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3645) );
  AOI22_X1 U4067 ( .A1(n3427), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4342), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3644) );
  AOI22_X1 U4068 ( .A1(n4388), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4301), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3643) );
  NAND2_X1 U4069 ( .A1(n3646), .A2(n3443), .ZN(n3647) );
  INV_X1 U4070 ( .A(n3716), .ZN(n3650) );
  INV_X1 U4071 ( .A(n3840), .ZN(n3649) );
  NOR2_X1 U4072 ( .A1(n3649), .A2(n3689), .ZN(n3836) );
  AND2_X1 U4073 ( .A1(n3650), .A2(n3836), .ZN(n3651) );
  NAND2_X1 U4074 ( .A1(n3653), .A2(n6491), .ZN(n3654) );
  INV_X1 U4075 ( .A(n3666), .ZN(n3658) );
  INV_X1 U4076 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3657) );
  AOI21_X1 U4077 ( .B1(n6822), .B2(n3840), .A(n6491), .ZN(n3656) );
  NAND2_X1 U4078 ( .A1(n6492), .A2(n3716), .ZN(n3655) );
  OAI211_X1 U4079 ( .C1(n3918), .C2(n3657), .A(n3656), .B(n3655), .ZN(n3665)
         );
  NAND2_X1 U4080 ( .A1(n4886), .A2(n3877), .ZN(n3663) );
  XNOR2_X1 U4081 ( .A(n3716), .B(n3715), .ZN(n3660) );
  OAI211_X1 U4082 ( .C1(n3660), .C2(n3659), .A(n3581), .B(n3934), .ZN(n3661)
         );
  INV_X1 U4083 ( .A(n3661), .ZN(n3662) );
  NAND2_X1 U4084 ( .A1(n3663), .A2(n3662), .ZN(n4877) );
  INV_X1 U4085 ( .A(n3664), .ZN(n3667) );
  NAND2_X1 U4086 ( .A1(n6492), .A2(n4656), .ZN(n4658) );
  OAI21_X1 U4087 ( .B1(n3659), .B2(n3716), .A(n4658), .ZN(n3668) );
  AOI21_X1 U4088 ( .B1(n6634), .B2(n3877), .A(n3668), .ZN(n4637) );
  INV_X1 U4089 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5763) );
  INV_X1 U4090 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3669) );
  NAND2_X1 U4091 ( .A1(n4875), .A2(n3669), .ZN(n3670) );
  NAND2_X1 U4092 ( .A1(n4877), .A2(n3670), .ZN(n3672) );
  INV_X1 U4093 ( .A(n4875), .ZN(n4636) );
  NAND2_X1 U4094 ( .A1(n4636), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3671)
         );
  NAND2_X1 U4095 ( .A1(n3672), .A2(n3671), .ZN(n3719) );
  NAND2_X1 U4096 ( .A1(n3719), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6092)
         );
  INV_X1 U4097 ( .A(n3673), .ZN(n3674) );
  AOI21_X2 U4098 ( .B1(n3678), .B2(n3677), .A(n3676), .ZN(n3712) );
  INV_X1 U4099 ( .A(n3712), .ZN(n3710) );
  INV_X1 U4100 ( .A(n3679), .ZN(n3682) );
  OAI21_X2 U4101 ( .B1(n3682), .B2(n3681), .A(n3680), .ZN(n3722) );
  NAND2_X1 U4102 ( .A1(n3725), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3687) );
  INV_X1 U4103 ( .A(n6620), .ZN(n3684) );
  NAND2_X1 U4104 ( .A1(n3684), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6489) );
  NAND2_X1 U4105 ( .A1(n6620), .A2(n6619), .ZN(n3685) );
  AND2_X1 U4106 ( .A1(n6489), .A2(n3685), .ZN(n6502) );
  INV_X1 U4107 ( .A(n4433), .ZN(n3729) );
  AOI22_X1 U4108 ( .A1(n6502), .A2(n3729), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3728), .ZN(n3686) );
  XNOR2_X2 U4109 ( .A(n3722), .B(n3723), .ZN(n4887) );
  NAND2_X1 U4110 ( .A1(n4887), .A2(n6491), .ZN(n3708) );
  AOI22_X1 U4111 ( .A1(n3690), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3695) );
  AOI22_X1 U4112 ( .A1(n3427), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4342), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3694) );
  AOI22_X1 U4113 ( .A1(n3627), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3693) );
  AOI22_X1 U4114 ( .A1(n4371), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3692) );
  NAND4_X1 U4115 ( .A1(n3695), .A2(n3694), .A3(n3693), .A4(n3692), .ZN(n3706)
         );
  AOI22_X1 U4116 ( .A1(n3429), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3430), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3704) );
  AOI22_X1 U4117 ( .A1(n4405), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3703) );
  AOI22_X1 U4118 ( .A1(n3622), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3702) );
  AOI22_X1 U4119 ( .A1(n3428), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4301), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3701) );
  NAND4_X1 U4120 ( .A1(n3704), .A2(n3703), .A3(n3702), .A4(n3701), .ZN(n3705)
         );
  AOI22_X1 U4121 ( .A1(n3878), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3931), 
        .B2(n3746), .ZN(n3707) );
  INV_X1 U4122 ( .A(n3711), .ZN(n3709) );
  NAND2_X1 U4123 ( .A1(n3710), .A2(n3709), .ZN(n3714) );
  AND2_X2 U4124 ( .A1(n3712), .A2(n3711), .ZN(n3744) );
  INV_X1 U4125 ( .A(n3744), .ZN(n3713) );
  NAND2_X1 U4126 ( .A1(n3716), .A2(n3715), .ZN(n3748) );
  XNOR2_X1 U4127 ( .A(n3748), .B(n3746), .ZN(n3717) );
  OAI21_X1 U4128 ( .B1(n3717), .B2(n3659), .A(n4658), .ZN(n3718) );
  AOI21_X1 U4129 ( .B1(n6585), .B2(n3877), .A(n3718), .ZN(n6095) );
  NAND2_X1 U4130 ( .A1(n6092), .A2(n6095), .ZN(n3720) );
  OR2_X1 U4131 ( .A1(n3719), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6093)
         );
  NAND2_X1 U4132 ( .A1(n3720), .A2(n6093), .ZN(n3754) );
  INV_X1 U4133 ( .A(n3754), .ZN(n3721) );
  NAND2_X1 U4134 ( .A1(n3721), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4865)
         );
  INV_X1 U4135 ( .A(n3722), .ZN(n3724) );
  NAND2_X1 U4136 ( .A1(n3725), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3731) );
  INV_X1 U4137 ( .A(n6489), .ZN(n3726) );
  INV_X1 U4138 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6499) );
  NAND2_X1 U4139 ( .A1(n3726), .A2(n6499), .ZN(n6572) );
  NAND2_X1 U4140 ( .A1(n6489), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3727) );
  NAND2_X1 U4141 ( .A1(n6572), .A2(n3727), .ZN(n6605) );
  AOI22_X1 U4142 ( .A1(n6605), .A2(n3729), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3728), .ZN(n3730) );
  AOI22_X1 U4143 ( .A1(n4412), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3735) );
  AOI22_X1 U4144 ( .A1(n3427), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3622), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3734) );
  AOI22_X1 U4145 ( .A1(n3430), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3733) );
  AOI22_X1 U4146 ( .A1(n4342), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3732) );
  NAND4_X1 U4147 ( .A1(n3735), .A2(n3734), .A3(n3733), .A4(n3732), .ZN(n3741)
         );
  AOI22_X1 U4148 ( .A1(n3429), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3627), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3739) );
  AOI22_X1 U4149 ( .A1(n4405), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3738) );
  AOI22_X1 U4150 ( .A1(n3428), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3737) );
  AOI22_X1 U4151 ( .A1(n4371), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4301), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3736) );
  NAND4_X1 U4152 ( .A1(n3739), .A2(n3738), .A3(n3737), .A4(n3736), .ZN(n3740)
         );
  AOI22_X1 U4153 ( .A1(n3878), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3931), 
        .B2(n3771), .ZN(n3742) );
  AND2_X2 U4154 ( .A1(n3756), .A2(n3745), .ZN(n6632) );
  NAND2_X1 U4155 ( .A1(n6632), .A2(n3877), .ZN(n3753) );
  INV_X1 U4156 ( .A(n3746), .ZN(n3747) );
  NAND2_X1 U4157 ( .A1(n3748), .A2(n3747), .ZN(n3772) );
  INV_X1 U4158 ( .A(n3771), .ZN(n3749) );
  XNOR2_X1 U4159 ( .A(n3772), .B(n3749), .ZN(n3751) );
  NAND2_X1 U4160 ( .A1(n3751), .A2(n6147), .ZN(n3752) );
  AND2_X1 U4161 ( .A1(n3753), .A2(n3752), .ZN(n4866) );
  NAND2_X1 U4162 ( .A1(n4865), .A2(n4866), .ZN(n3755) );
  NAND2_X1 U4163 ( .A1(n3754), .A2(n4868), .ZN(n4864) );
  NAND2_X1 U4164 ( .A1(n3755), .A2(n4864), .ZN(n4830) );
  INV_X1 U4165 ( .A(n4830), .ZN(n3777) );
  INV_X1 U4166 ( .A(n3756), .ZN(n3768) );
  AOI22_X1 U4167 ( .A1(n3427), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4342), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3760) );
  AOI22_X1 U4168 ( .A1(n3429), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3627), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3759) );
  AOI22_X1 U4169 ( .A1(n4371), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3758) );
  AOI22_X1 U4170 ( .A1(n3430), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3757) );
  NAND4_X1 U4171 ( .A1(n3760), .A2(n3759), .A3(n3758), .A4(n3757), .ZN(n3766)
         );
  AOI22_X1 U4172 ( .A1(n4405), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3764) );
  AOI22_X1 U4173 ( .A1(n4412), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3763) );
  AOI22_X1 U4174 ( .A1(n3622), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3762) );
  AOI22_X1 U4175 ( .A1(n4388), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4301), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3761) );
  NAND4_X1 U4176 ( .A1(n3764), .A2(n3763), .A3(n3762), .A4(n3761), .ZN(n3765)
         );
  AOI22_X1 U4177 ( .A1(n3878), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3931), 
        .B2(n3791), .ZN(n3769) );
  INV_X1 U4178 ( .A(n3769), .ZN(n3767) );
  NAND2_X2 U4179 ( .A1(n3768), .A2(n3767), .ZN(n3818) );
  NAND2_X1 U4180 ( .A1(n3756), .A2(n3769), .ZN(n3770) );
  NAND2_X1 U4181 ( .A1(n3818), .A2(n3770), .ZN(n3940) );
  OR2_X1 U4182 ( .A1(n3940), .A2(n4664), .ZN(n3775) );
  NAND2_X1 U4183 ( .A1(n3772), .A2(n3771), .ZN(n3793) );
  XNOR2_X1 U4184 ( .A(n3793), .B(n3791), .ZN(n3773) );
  NAND2_X1 U4185 ( .A1(n3773), .A2(n6147), .ZN(n3774) );
  XNOR2_X1 U4186 ( .A(n3778), .B(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4829)
         );
  INV_X1 U4187 ( .A(n4829), .ZN(n3776) );
  NAND2_X1 U4188 ( .A1(n3777), .A2(n3776), .ZN(n4935) );
  NAND2_X1 U4189 ( .A1(n3778), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4934)
         );
  INV_X1 U4190 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3790) );
  AOI22_X1 U4191 ( .A1(n4412), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3782) );
  AOI22_X1 U4192 ( .A1(n3427), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3622), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3781) );
  AOI22_X1 U4193 ( .A1(n3430), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3780) );
  AOI22_X1 U4194 ( .A1(n4342), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3779) );
  NAND4_X1 U4195 ( .A1(n3782), .A2(n3781), .A3(n3780), .A4(n3779), .ZN(n3788)
         );
  AOI22_X1 U4196 ( .A1(n3429), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3627), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3786) );
  AOI22_X1 U4197 ( .A1(n4405), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3785) );
  AOI22_X1 U4198 ( .A1(n3428), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3784) );
  AOI22_X1 U4199 ( .A1(n4371), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4301), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3783) );
  NAND4_X1 U4200 ( .A1(n3786), .A2(n3785), .A3(n3784), .A4(n3783), .ZN(n3787)
         );
  NAND2_X1 U4201 ( .A1(n3931), .A2(n3794), .ZN(n3789) );
  OAI21_X1 U4202 ( .B1(n3918), .B2(n3790), .A(n3789), .ZN(n3813) );
  XNOR2_X1 U4203 ( .A(n3818), .B(n3813), .ZN(n3979) );
  NAND2_X1 U4204 ( .A1(n3979), .A2(n3877), .ZN(n3797) );
  INV_X1 U4205 ( .A(n3791), .ZN(n3792) );
  NOR2_X1 U4206 ( .A1(n3793), .A2(n3792), .ZN(n3795) );
  NAND2_X1 U4207 ( .A1(n3795), .A2(n3794), .ZN(n3829) );
  OAI211_X1 U4208 ( .C1(n3795), .C2(n3794), .A(n3829), .B(n6147), .ZN(n3796)
         );
  NAND2_X1 U4209 ( .A1(n3797), .A2(n3796), .ZN(n3801) );
  NAND2_X1 U4210 ( .A1(n3801), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3799)
         );
  AND2_X1 U4211 ( .A1(n4934), .A2(n3799), .ZN(n3798) );
  NAND2_X1 U4212 ( .A1(n4935), .A2(n3798), .ZN(n4989) );
  INV_X1 U4213 ( .A(n3799), .ZN(n3802) );
  INV_X1 U4214 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3800) );
  XNOR2_X1 U4215 ( .A(n3801), .B(n3800), .ZN(n4933) );
  AOI22_X1 U4216 ( .A1(n4412), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4217 ( .A1(n3627), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3430), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4218 ( .A1(n3622), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4342), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3804) );
  AOI22_X1 U4219 ( .A1(n4405), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3803) );
  NAND4_X1 U4220 ( .A1(n3806), .A2(n3805), .A3(n3804), .A4(n3803), .ZN(n3812)
         );
  AOI22_X1 U4221 ( .A1(n3428), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4222 ( .A1(n3429), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4223 ( .A1(n3427), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3808) );
  AOI22_X1 U4224 ( .A1(n4371), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4301), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3807) );
  NAND4_X1 U4225 ( .A1(n3810), .A2(n3809), .A3(n3808), .A4(n3807), .ZN(n3811)
         );
  AOI22_X1 U4226 ( .A1(n3878), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3931), 
        .B2(n3830), .ZN(n3816) );
  INV_X1 U4227 ( .A(n3813), .ZN(n3817) );
  OAI21_X1 U4228 ( .B1(n3818), .B2(n3817), .A(n3816), .ZN(n3987) );
  NAND3_X1 U4229 ( .A1(n3838), .A2(n3877), .A3(n3987), .ZN(n3821) );
  XNOR2_X1 U4230 ( .A(n3829), .B(n3830), .ZN(n3819) );
  NAND2_X1 U4231 ( .A1(n3819), .A2(n6147), .ZN(n3820) );
  NAND2_X1 U4232 ( .A1(n3821), .A2(n3820), .ZN(n3823) );
  INV_X1 U4233 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4471) );
  XNOR2_X1 U4234 ( .A(n3823), .B(n4471), .ZN(n4992) );
  NAND2_X1 U4235 ( .A1(n4989), .A2(n3822), .ZN(n3825) );
  NAND2_X1 U4236 ( .A1(n3823), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3824)
         );
  NAND2_X2 U4237 ( .A1(n3825), .A2(n3824), .ZN(n5020) );
  INV_X1 U4238 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3827) );
  NAND2_X1 U4239 ( .A1(n3931), .A2(n3840), .ZN(n3826) );
  OAI21_X1 U4240 ( .B1(n3918), .B2(n3827), .A(n3826), .ZN(n3828) );
  NAND2_X1 U4241 ( .A1(n3999), .A2(n3877), .ZN(n3834) );
  INV_X1 U4242 ( .A(n3829), .ZN(n3831) );
  NAND2_X1 U4243 ( .A1(n3831), .A2(n3830), .ZN(n3839) );
  XNOR2_X1 U4244 ( .A(n3839), .B(n3840), .ZN(n3832) );
  NAND2_X1 U4245 ( .A1(n3832), .A2(n6147), .ZN(n3833) );
  INV_X1 U4246 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3835) );
  AND2_X1 U4247 ( .A1(n3836), .A2(n3877), .ZN(n3837) );
  INV_X1 U4248 ( .A(n3839), .ZN(n3841) );
  NAND3_X1 U4249 ( .A1(n3841), .A2(n6147), .A3(n3840), .ZN(n3842) );
  NAND2_X1 U4250 ( .A1(n3851), .A2(n3842), .ZN(n3846) );
  INV_X1 U4251 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4478) );
  XNOR2_X1 U4252 ( .A(n3846), .B(n4478), .ZN(n5024) );
  AND2_X1 U4253 ( .A1(n5019), .A2(n5024), .ZN(n3843) );
  NAND2_X1 U4254 ( .A1(n5020), .A2(n3843), .ZN(n3850) );
  NAND2_X1 U4255 ( .A1(n3844), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n5021)
         );
  INV_X1 U4256 ( .A(n5021), .ZN(n3845) );
  AND2_X1 U4257 ( .A1(n3846), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3847)
         );
  NOR2_X1 U4258 ( .A1(n3848), .A2(n3847), .ZN(n3849) );
  NAND2_X1 U4259 ( .A1(n3850), .A2(n3849), .ZN(n5102) );
  XNOR2_X1 U4260 ( .A(n5737), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5103)
         );
  NAND2_X1 U4261 ( .A1(n5102), .A2(n5103), .ZN(n5076) );
  INV_X1 U4262 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6189) );
  OR2_X1 U4263 ( .A1(n5737), .A2(n6189), .ZN(n5075) );
  XNOR2_X1 U4264 ( .A(n3851), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6112)
         );
  INV_X1 U4265 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4485) );
  OR2_X1 U4266 ( .A1(n3851), .A2(n4485), .ZN(n6100) );
  INV_X1 U4267 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3853) );
  OR2_X1 U4268 ( .A1(n3851), .A2(n3853), .ZN(n6099) );
  AND2_X1 U4269 ( .A1(n6100), .A2(n6099), .ZN(n5077) );
  INV_X1 U4270 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6161) );
  OR2_X1 U4271 ( .A1(n3851), .A2(n6161), .ZN(n5080) );
  AND2_X1 U4272 ( .A1(n5077), .A2(n5080), .ZN(n6108) );
  AND2_X1 U4273 ( .A1(n5075), .A2(n3439), .ZN(n3852) );
  NAND2_X1 U4274 ( .A1(n5076), .A2(n3852), .ZN(n3856) );
  INV_X1 U4275 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5215) );
  NAND2_X1 U4276 ( .A1(n3851), .A2(n3853), .ZN(n6098) );
  NAND2_X1 U4277 ( .A1(n5737), .A2(n6161), .ZN(n5079) );
  AND2_X1 U4278 ( .A1(n6098), .A2(n5079), .ZN(n6110) );
  NAND2_X1 U4279 ( .A1(n5737), .A2(n4485), .ZN(n5131) );
  NAND3_X1 U4280 ( .A1(n3856), .A2(n3855), .A3(n5131), .ZN(n5646) );
  INV_X1 U4281 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5644) );
  AND2_X1 U4282 ( .A1(n5737), .A2(n5644), .ZN(n3857) );
  OAI22_X2 U4283 ( .A1(n5646), .A2(n3857), .B1(n5737), .B2(n5644), .ZN(n5636)
         );
  INV_X1 U4284 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6222) );
  NOR2_X1 U4285 ( .A1(n5737), .A2(n6222), .ZN(n5632) );
  NAND2_X1 U4286 ( .A1(n5737), .A2(n6222), .ZN(n5633) );
  OAI21_X1 U4287 ( .B1(n5636), .B2(n5632), .A(n5633), .ZN(n5622) );
  INV_X1 U4288 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6230) );
  OR2_X2 U4289 ( .A1(n5622), .A2(n5620), .ZN(n5611) );
  INV_X1 U4290 ( .A(n5611), .ZN(n3859) );
  AND2_X1 U4291 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5219) );
  INV_X1 U4292 ( .A(n5219), .ZN(n3858) );
  NAND2_X1 U4293 ( .A1(n3859), .A2(n3433), .ZN(n5580) );
  NOR2_X1 U4294 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3860) );
  OR2_X1 U4295 ( .A1(n5737), .A2(n3860), .ZN(n3861) );
  NOR2_X1 U4296 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5739) );
  NOR2_X1 U4297 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5712) );
  NOR2_X1 U4298 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5567) );
  NAND3_X1 U4299 ( .A1(n5739), .A2(n5712), .A3(n5567), .ZN(n3863) );
  NAND2_X1 U4300 ( .A1(n5748), .A2(n3863), .ZN(n3864) );
  NAND2_X1 U4301 ( .A1(n5565), .A2(n3864), .ZN(n3866) );
  AND2_X1 U4302 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5740) );
  AND2_X1 U4303 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5216) );
  NAND2_X1 U4304 ( .A1(n5740), .A2(n5216), .ZN(n5579) );
  NAND2_X1 U4305 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5226) );
  OAI21_X1 U4306 ( .B1(n5579), .B2(n5226), .A(n3851), .ZN(n3865) );
  NAND2_X1 U4307 ( .A1(n3866), .A2(n3865), .ZN(n5558) );
  XNOR2_X1 U4308 ( .A(n3851), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5557)
         );
  NAND2_X1 U4309 ( .A1(n5558), .A2(n5557), .ZN(n5556) );
  INV_X1 U4310 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5706) );
  NAND2_X1 U4311 ( .A1(n5737), .A2(n5706), .ZN(n3867) );
  NAND2_X1 U4312 ( .A1(n5556), .A2(n3867), .ZN(n5550) );
  INV_X1 U4313 ( .A(n5550), .ZN(n3868) );
  INV_X1 U4314 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5693) );
  AND2_X1 U4315 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5675) );
  NAND2_X1 U4316 ( .A1(n5675), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5654) );
  AND2_X1 U4317 ( .A1(n5737), .A2(n5654), .ZN(n3871) );
  NOR2_X1 U4318 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3869) );
  OR2_X1 U4319 ( .A1(n5737), .A2(n3869), .ZN(n5530) );
  INV_X1 U4320 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5676) );
  OR2_X1 U4321 ( .A1(n5737), .A2(n5676), .ZN(n3870) );
  OAI21_X2 U4322 ( .B1(n5539), .B2(n3871), .A(n5522), .ZN(n5209) );
  INV_X1 U4323 ( .A(n3872), .ZN(n3874) );
  NAND2_X1 U4324 ( .A1(n5209), .A2(n5737), .ZN(n3873) );
  OAI21_X2 U4325 ( .B1(n3874), .B2(n5737), .A(n3873), .ZN(n3876) );
  XNOR2_X1 U4326 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3898) );
  NAND2_X1 U4327 ( .A1(n6647), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3884) );
  INV_X1 U4328 ( .A(n3884), .ZN(n3897) );
  XNOR2_X1 U4329 ( .A(n3898), .B(n3897), .ZN(n4555) );
  OR2_X1 U4330 ( .A1(n4555), .A2(n6491), .ZN(n3879) );
  NAND2_X1 U4331 ( .A1(n3927), .A2(n3879), .ZN(n3894) );
  INV_X1 U4332 ( .A(n4555), .ZN(n3881) );
  NAND2_X1 U4333 ( .A1(n3931), .A2(n4837), .ZN(n3880) );
  OAI211_X1 U4334 ( .C1(n3918), .C2(n3881), .A(n3934), .B(n3880), .ZN(n3893)
         );
  NAND2_X1 U4335 ( .A1(n6691), .A2(n3934), .ZN(n3883) );
  OAI21_X1 U4336 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6647), .A(n3884), 
        .ZN(n3889) );
  INV_X1 U4337 ( .A(n3889), .ZN(n3885) );
  NAND2_X1 U4338 ( .A1(n3937), .A2(n3885), .ZN(n3887) );
  NAND2_X1 U4339 ( .A1(n3887), .A2(n3886), .ZN(n3888) );
  NAND2_X1 U4340 ( .A1(n3903), .A2(n3888), .ZN(n3892) );
  INV_X1 U4341 ( .A(n3931), .ZN(n3890) );
  OAI21_X1 U4342 ( .B1(n3890), .B2(n3889), .A(n3927), .ZN(n3891) );
  OAI211_X1 U4343 ( .C1(n3894), .C2(n3893), .A(n3892), .B(n3891), .ZN(n3896)
         );
  NAND2_X1 U4344 ( .A1(n3894), .A2(n3893), .ZN(n3895) );
  NAND2_X1 U4345 ( .A1(n3896), .A2(n3895), .ZN(n3906) );
  NAND2_X1 U4346 ( .A1(n3898), .A2(n3897), .ZN(n3900) );
  NAND2_X1 U4347 ( .A1(n6621), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3899) );
  NAND2_X1 U4348 ( .A1(n3900), .A2(n3899), .ZN(n3908) );
  MUX2_X1 U4349 ( .A(n6619), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n3907) );
  XNOR2_X1 U4350 ( .A(n3908), .B(n3907), .ZN(n4554) );
  INV_X1 U4351 ( .A(n4554), .ZN(n3901) );
  NAND2_X1 U4352 ( .A1(n3931), .A2(n3901), .ZN(n3902) );
  OAI211_X1 U4353 ( .C1(n3901), .C2(n3918), .A(n3903), .B(n3902), .ZN(n3905)
         );
  NOR2_X1 U4354 ( .A1(n3903), .A2(n3902), .ZN(n3904) );
  AOI21_X1 U4355 ( .B1(n3906), .B2(n3905), .A(n3904), .ZN(n3913) );
  NAND2_X1 U4356 ( .A1(n3908), .A2(n3907), .ZN(n3910) );
  NAND2_X1 U4357 ( .A1(n6619), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3909) );
  NAND2_X1 U4358 ( .A1(n3910), .A2(n3909), .ZN(n3916) );
  MUX2_X1 U4359 ( .A(n6499), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n3915) );
  XNOR2_X1 U4360 ( .A(n3916), .B(n3915), .ZN(n4556) );
  AND2_X1 U4361 ( .A1(n3918), .A2(n4556), .ZN(n3912) );
  INV_X1 U4362 ( .A(n4556), .ZN(n3911) );
  OAI22_X1 U4363 ( .A1(n3913), .A2(n3912), .B1(n3911), .B2(n3927), .ZN(n3921)
         );
  NOR2_X1 U4364 ( .A1(n4807), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3914)
         );
  AOI21_X1 U4365 ( .B1(n3916), .B2(n3915), .A(n3914), .ZN(n3922) );
  AND2_X1 U4366 ( .A1(n6404), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n3923)
         );
  NAND2_X1 U4367 ( .A1(n3922), .A2(n3923), .ZN(n4559) );
  INV_X1 U4368 ( .A(n4559), .ZN(n3917) );
  NAND2_X1 U4369 ( .A1(n3918), .A2(n3917), .ZN(n3920) );
  OAI22_X1 U4370 ( .A1(n3927), .A2(n4559), .B1(STATE2_REG_0__SCAN_IN), .B2(
        n6404), .ZN(n3919) );
  AOI21_X1 U4371 ( .B1(n3921), .B2(n3920), .A(n3919), .ZN(n3929) );
  INV_X1 U4372 ( .A(n3922), .ZN(n3926) );
  INV_X1 U4373 ( .A(n3923), .ZN(n3925) );
  NOR2_X1 U4374 ( .A1(n6404), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n3924)
         );
  AOI21_X1 U4375 ( .B1(n3926), .B2(n3925), .A(n3924), .ZN(n4558) );
  NOR2_X1 U4376 ( .A1(n3927), .A2(n4558), .ZN(n3928) );
  INV_X1 U4377 ( .A(n4558), .ZN(n3930) );
  NAND2_X1 U4378 ( .A1(n3931), .A2(n3930), .ZN(n3932) );
  AOI21_X1 U4379 ( .B1(n3577), .B2(n3934), .A(n4831), .ZN(n3935) );
  NOR2_X1 U4380 ( .A1(n3936), .A2(n3935), .ZN(n4769) );
  INV_X1 U4381 ( .A(n3937), .ZN(n3938) );
  NAND2_X1 U4382 ( .A1(n4769), .A2(n3938), .ZN(n4844) );
  OR2_X1 U4383 ( .A1(n5262), .A2(n4844), .ZN(n6419) );
  AND2_X1 U4384 ( .A1(n3939), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6449) );
  INV_X1 U4385 ( .A(n6449), .ZN(n6428) );
  INV_X2 U4386 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6657) );
  NOR2_X2 U4387 ( .A1(n3941), .A2(n6657), .ZN(n4274) );
  OAI21_X1 U4388 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n3948), .A(n3980), 
        .ZN(n4959) );
  NAND2_X1 U4389 ( .A1(n3567), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3954) );
  INV_X1 U4390 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6670) );
  OAI21_X1 U4391 ( .B1(n6670), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6657), 
        .ZN(n3943) );
  NAND2_X1 U4392 ( .A1(n4427), .A2(EAX_REG_4__SCAN_IN), .ZN(n3942) );
  OAI211_X1 U4393 ( .C1(n3954), .C2(n6404), .A(n3943), .B(n3942), .ZN(n3944)
         );
  OAI21_X1 U4394 ( .B1(n4425), .B2(n4959), .A(n3944), .ZN(n3945) );
  AOI21_X1 U4395 ( .B1(n3947), .B2(n4274), .A(n3946), .ZN(n4604) );
  NAND2_X1 U4396 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3967) );
  INV_X1 U4397 ( .A(n3967), .ZN(n3950) );
  INV_X1 U4398 ( .A(n3948), .ZN(n3949) );
  OAI21_X1 U4399 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3950), .A(n3949), 
        .ZN(n5062) );
  AND2_X1 U4400 ( .A1(n6657), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5191) );
  AOI22_X1 U4401 ( .A1(n4562), .A2(n5062), .B1(n5191), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3952) );
  NAND2_X1 U4402 ( .A1(n4427), .A2(EAX_REG_3__SCAN_IN), .ZN(n3951) );
  OAI211_X1 U4403 ( .C1(n3954), .C2(n4807), .A(n3952), .B(n3951), .ZN(n3953)
         );
  AOI21_X1 U4404 ( .B1(n6632), .B2(n4274), .A(n3953), .ZN(n4820) );
  NAND2_X1 U4405 ( .A1(n4886), .A2(n4274), .ZN(n3958) );
  AOI22_X1 U4406 ( .A1(n4427), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6657), .ZN(n3956) );
  INV_X1 U4407 ( .A(n3954), .ZN(n3966) );
  NAND2_X1 U4408 ( .A1(n3966), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3955) );
  AND2_X1 U4409 ( .A1(n3956), .A2(n3955), .ZN(n3957) );
  NAND2_X1 U4410 ( .A1(n3958), .A2(n3957), .ZN(n4643) );
  INV_X2 U4411 ( .A(n6634), .ZN(n6645) );
  AOI21_X1 U4412 ( .B1(n6645), .B2(n3577), .A(n6657), .ZN(n4635) );
  INV_X1 U4413 ( .A(n3959), .ZN(n3960) );
  XNOR2_X1 U4414 ( .A(n3961), .B(n3960), .ZN(n6529) );
  NAND2_X1 U4415 ( .A1(n6529), .A2(n4274), .ZN(n3965) );
  AOI22_X1 U4416 ( .A1(n4427), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6657), .ZN(n3963) );
  NAND2_X1 U4417 ( .A1(n3966), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3962) );
  AND2_X1 U4418 ( .A1(n3963), .A2(n3962), .ZN(n3964) );
  NAND2_X1 U4419 ( .A1(n3965), .A2(n3964), .ZN(n4634) );
  MUX2_X1 U4420 ( .A(n4562), .B(n4635), .S(n4634), .Z(n4642) );
  INV_X1 U4421 ( .A(n4784), .ZN(n3973) );
  NAND2_X1 U4422 ( .A1(n3966), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3971) );
  INV_X2 U4423 ( .A(n4399), .ZN(n4427) );
  INV_X1 U4424 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6269) );
  INV_X1 U4425 ( .A(n5191), .ZN(n4283) );
  OAI21_X1 U4426 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3967), .ZN(n6275) );
  NAND2_X1 U4427 ( .A1(n4562), .A2(n6275), .ZN(n3968) );
  OAI21_X1 U4428 ( .B1(n6269), .B2(n4283), .A(n3968), .ZN(n3969) );
  AOI21_X1 U4429 ( .B1(n4427), .B2(EAX_REG_2__SCAN_IN), .A(n3969), .ZN(n3970)
         );
  AND2_X1 U4430 ( .A1(n3971), .A2(n3970), .ZN(n4785) );
  INV_X1 U4431 ( .A(n4785), .ZN(n3972) );
  NAND2_X1 U4432 ( .A1(n3973), .A2(n3972), .ZN(n3974) );
  AOI21_X1 U4433 ( .B1(n6585), .B2(n4274), .A(n5191), .ZN(n4786) );
  NAND2_X1 U4434 ( .A1(n3974), .A2(n4786), .ZN(n3976) );
  NAND2_X1 U4435 ( .A1(n4784), .A2(n4785), .ZN(n3975) );
  NAND2_X1 U4436 ( .A1(n3976), .A2(n3975), .ZN(n4819) );
  NAND2_X1 U4437 ( .A1(n3979), .A2(n4274), .ZN(n3986) );
  INV_X1 U4438 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3983) );
  OAI21_X1 U4439 ( .B1(PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n3981), .A(n3988), 
        .ZN(n6276) );
  NAND2_X1 U4440 ( .A1(n4562), .A2(n6276), .ZN(n3982) );
  OAI21_X1 U4441 ( .B1(n3983), .B2(n4283), .A(n3982), .ZN(n3984) );
  AOI21_X1 U4442 ( .B1(n4427), .B2(EAX_REG_5__SCAN_IN), .A(n3984), .ZN(n3985)
         );
  NAND2_X1 U4443 ( .A1(n3986), .A2(n3985), .ZN(n4951) );
  INV_X1 U4444 ( .A(n3988), .ZN(n3990) );
  INV_X1 U4445 ( .A(n3995), .ZN(n3989) );
  OAI21_X1 U4446 ( .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n3990), .A(n3989), 
        .ZN(n6293) );
  NAND2_X1 U4447 ( .A1(n4562), .A2(n6293), .ZN(n3991) );
  OAI21_X1 U4448 ( .B1(n6292), .B2(n4283), .A(n3991), .ZN(n3992) );
  AOI21_X1 U4449 ( .B1(n4427), .B2(EAX_REG_6__SCAN_IN), .A(n3992), .ZN(n3993)
         );
  INV_X1 U4450 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3997) );
  OAI21_X1 U4451 ( .B1(PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n3995), .A(n4015), 
        .ZN(n6303) );
  AOI22_X1 U4452 ( .A1(n4562), .A2(n6303), .B1(n5191), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3996) );
  OAI21_X1 U4453 ( .B1(n4399), .B2(n3997), .A(n3996), .ZN(n3998) );
  OR2_X2 U4454 ( .A1(n5003), .A2(n5002), .ZN(n5035) );
  AOI22_X1 U4455 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n3427), .B1(n4306), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4004) );
  AOI22_X1 U4456 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n3429), .B1(n4413), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4003) );
  AOI22_X1 U4457 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4342), .B1(n4407), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4002) );
  AOI22_X1 U4458 ( .A1(n4388), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4301), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4001) );
  NAND4_X1 U4459 ( .A1(n4004), .A2(n4003), .A3(n4002), .A4(n4001), .ZN(n4010)
         );
  AOI22_X1 U4460 ( .A1(n3627), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4405), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U4461 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n4371), .B1(n3428), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4007) );
  AOI22_X1 U4462 ( .A1(n4412), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3622), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4006) );
  AOI22_X1 U4463 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n3430), .B1(n4406), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4005) );
  NAND4_X1 U4464 ( .A1(n4008), .A2(n4007), .A3(n4006), .A4(n4005), .ZN(n4009)
         );
  OAI21_X1 U4465 ( .B1(n4010), .B2(n4009), .A(n4274), .ZN(n4014) );
  INV_X1 U4466 ( .A(n4015), .ZN(n4011) );
  XNOR2_X1 U4467 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n4011), .ZN(n5051) );
  AOI22_X1 U4468 ( .A1(n4562), .A2(n5051), .B1(n5191), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4013) );
  NAND2_X1 U4469 ( .A1(n4427), .A2(EAX_REG_8__SCAN_IN), .ZN(n4012) );
  AND3_X1 U4470 ( .A1(n4014), .A2(n4013), .A3(n4012), .ZN(n5034) );
  XOR2_X1 U4471 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n4029), .Z(n6316) );
  AOI22_X1 U4472 ( .A1(n4427), .A2(EAX_REG_9__SCAN_IN), .B1(n5191), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4027) );
  AOI22_X1 U4473 ( .A1(n4405), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3430), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4019) );
  AOI22_X1 U4474 ( .A1(n4412), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3622), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4018) );
  AOI22_X1 U4475 ( .A1(n3428), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U4476 ( .A1(n4371), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4301), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4016) );
  NAND4_X1 U4477 ( .A1(n4019), .A2(n4018), .A3(n4017), .A4(n4016), .ZN(n4025)
         );
  AOI22_X1 U4478 ( .A1(n3427), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4023) );
  AOI22_X1 U4479 ( .A1(n3429), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4022) );
  AOI22_X1 U4480 ( .A1(n3627), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4021) );
  AOI22_X1 U4481 ( .A1(n4342), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4020) );
  NAND4_X1 U4482 ( .A1(n4023), .A2(n4022), .A3(n4021), .A4(n4020), .ZN(n4024)
         );
  OAI21_X1 U4483 ( .B1(n4025), .B2(n4024), .A(n4274), .ZN(n4026) );
  OAI211_X1 U4484 ( .C1(n6316), .C2(n4425), .A(n4027), .B(n4026), .ZN(n4028)
         );
  INV_X1 U4485 ( .A(n4028), .ZN(n5104) );
  NAND2_X1 U4486 ( .A1(n4029), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4045)
         );
  INV_X1 U4487 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5119) );
  XNOR2_X1 U4488 ( .A(n4045), .B(n5119), .ZN(n5134) );
  NAND2_X1 U4489 ( .A1(n5134), .A2(n4562), .ZN(n4044) );
  AOI22_X1 U4490 ( .A1(n3430), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4342), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4033) );
  AOI22_X1 U4491 ( .A1(n4405), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4032) );
  AOI22_X1 U4492 ( .A1(n3627), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4031) );
  AOI22_X1 U4493 ( .A1(n4371), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4030) );
  NAND4_X1 U4494 ( .A1(n4033), .A2(n4032), .A3(n4031), .A4(n4030), .ZN(n4039)
         );
  AOI22_X1 U4495 ( .A1(n4412), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4037) );
  AOI22_X1 U4496 ( .A1(n3427), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3622), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4036) );
  AOI22_X1 U4497 ( .A1(n3544), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4035) );
  AOI22_X1 U4498 ( .A1(n3429), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4301), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4034) );
  NAND4_X1 U4499 ( .A1(n4037), .A2(n4036), .A3(n4035), .A4(n4034), .ZN(n4038)
         );
  OAI21_X1 U4500 ( .B1(n4039), .B2(n4038), .A(n4274), .ZN(n4042) );
  NAND2_X1 U4501 ( .A1(n4427), .A2(EAX_REG_10__SCAN_IN), .ZN(n4041) );
  NAND2_X1 U4502 ( .A1(n5191), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4040)
         );
  AND3_X1 U4503 ( .A1(n4042), .A2(n4041), .A3(n4040), .ZN(n4043) );
  NAND2_X1 U4504 ( .A1(n4044), .A2(n4043), .ZN(n5114) );
  AND2_X2 U4505 ( .A1(n3445), .A2(n5114), .ZN(n5113) );
  XOR2_X1 U4506 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n4058), .Z(n6103) );
  AOI22_X1 U4507 ( .A1(n4427), .A2(EAX_REG_11__SCAN_IN), .B1(n5191), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4057) );
  AOI22_X1 U4508 ( .A1(n3429), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3627), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4049) );
  AOI22_X1 U4509 ( .A1(n3427), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3622), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4048) );
  AOI22_X1 U4510 ( .A1(n4342), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4047) );
  AOI22_X1 U4511 ( .A1(n4371), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4046) );
  NAND4_X1 U4512 ( .A1(n4049), .A2(n4048), .A3(n4047), .A4(n4046), .ZN(n4055)
         );
  AOI22_X1 U4513 ( .A1(n4412), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4053) );
  AOI22_X1 U4514 ( .A1(n4405), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4052) );
  AOI22_X1 U4515 ( .A1(n3430), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4051) );
  AOI22_X1 U4516 ( .A1(n3428), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4301), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4050) );
  NAND4_X1 U4517 ( .A1(n4053), .A2(n4052), .A3(n4051), .A4(n4050), .ZN(n4054)
         );
  OAI21_X1 U4518 ( .B1(n4055), .B2(n4054), .A(n4274), .ZN(n4056) );
  OAI211_X1 U4519 ( .C1(n6103), .C2(n4425), .A(n4057), .B(n4056), .ZN(n5148)
         );
  NAND2_X1 U4520 ( .A1(n4058), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4093)
         );
  XNOR2_X1 U4521 ( .A(n4093), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5167)
         );
  NAND2_X1 U4522 ( .A1(n5167), .A2(n4562), .ZN(n4063) );
  INV_X1 U4523 ( .A(EAX_REG_12__SCAN_IN), .ZN(n4061) );
  INV_X1 U4524 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5164) );
  AOI21_X1 U4525 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n5164), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4059) );
  INV_X1 U4526 ( .A(n4059), .ZN(n4060) );
  OAI21_X1 U4527 ( .B1(n4399), .B2(n4061), .A(n4060), .ZN(n4062) );
  NAND2_X1 U4528 ( .A1(n4063), .A2(n4062), .ZN(n4075) );
  AOI22_X1 U4529 ( .A1(n4405), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4067) );
  AOI22_X1 U4530 ( .A1(n4412), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4342), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4066) );
  AOI22_X1 U4531 ( .A1(n3627), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4065) );
  AOI22_X1 U4532 ( .A1(n4371), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4064) );
  NAND4_X1 U4533 ( .A1(n4067), .A2(n4066), .A3(n4065), .A4(n4064), .ZN(n4073)
         );
  AOI22_X1 U4534 ( .A1(n3427), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4071) );
  AOI22_X1 U4535 ( .A1(n3430), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3622), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4070) );
  AOI22_X1 U4536 ( .A1(n3429), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4069) );
  AOI22_X1 U4537 ( .A1(n4413), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4301), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4068) );
  NAND4_X1 U4538 ( .A1(n4071), .A2(n4070), .A3(n4069), .A4(n4068), .ZN(n4072)
         );
  OAI21_X1 U4539 ( .B1(n4073), .B2(n4072), .A(n4274), .ZN(n4074) );
  NAND2_X1 U4540 ( .A1(n4075), .A2(n4074), .ZN(n5139) );
  AOI22_X1 U4541 ( .A1(n4412), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3622), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4079) );
  AOI22_X1 U4542 ( .A1(n3429), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3430), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4078) );
  AOI22_X1 U4543 ( .A1(n4405), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4077) );
  AOI22_X1 U4544 ( .A1(n3428), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4301), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4076) );
  NAND4_X1 U4545 ( .A1(n4079), .A2(n4078), .A3(n4077), .A4(n4076), .ZN(n4085)
         );
  AOI22_X1 U4546 ( .A1(n3427), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4083) );
  AOI22_X1 U4547 ( .A1(n4342), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4082) );
  AOI22_X1 U4548 ( .A1(n3627), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4081) );
  AOI22_X1 U4549 ( .A1(n4371), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4080) );
  NAND4_X1 U4550 ( .A1(n4083), .A2(n4082), .A3(n4081), .A4(n4080), .ZN(n4084)
         );
  OR2_X1 U4551 ( .A1(n4085), .A2(n4084), .ZN(n4086) );
  AND2_X1 U4552 ( .A1(n4274), .A2(n4086), .ZN(n4088) );
  AND2_X1 U4553 ( .A1(n5139), .A2(n4088), .ZN(n4087) );
  INV_X1 U4554 ( .A(n5139), .ZN(n4090) );
  INV_X1 U4555 ( .A(n4088), .ZN(n4089) );
  NAND2_X1 U4556 ( .A1(n4100), .A2(n4092), .ZN(n5176) );
  INV_X1 U4557 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4096) );
  OAI21_X1 U4558 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n4094), .A(n4265), 
        .ZN(n6332) );
  NAND2_X1 U4559 ( .A1(n6332), .A2(n4562), .ZN(n4095) );
  OAI21_X1 U4560 ( .B1(n4096), .B2(n4283), .A(n4095), .ZN(n4097) );
  AOI21_X1 U4561 ( .B1(n4427), .B2(EAX_REG_13__SCAN_IN), .A(n4097), .ZN(n5175)
         );
  NOR2_X1 U4562 ( .A1(n4665), .A2(n6864), .ZN(n4776) );
  AOI22_X1 U4563 ( .A1(n4307), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4104) );
  AOI22_X1 U4564 ( .A1(n3427), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4342), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4103) );
  AOI22_X1 U4565 ( .A1(n3430), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4102) );
  AOI22_X1 U4566 ( .A1(n3428), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4301), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4101) );
  NAND4_X1 U4567 ( .A1(n4104), .A2(n4103), .A3(n4102), .A4(n4101), .ZN(n4110)
         );
  AOI22_X1 U4568 ( .A1(n4405), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3429), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4108) );
  AOI22_X1 U4569 ( .A1(n3622), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4107) );
  AOI22_X1 U4570 ( .A1(n3627), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4106) );
  AOI22_X1 U4571 ( .A1(n4371), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4105) );
  NAND4_X1 U4572 ( .A1(n4108), .A2(n4107), .A3(n4106), .A4(n4105), .ZN(n4109)
         );
  NOR2_X1 U4573 ( .A1(n4110), .A2(n4109), .ZN(n4284) );
  AOI22_X1 U4574 ( .A1(n3429), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4114) );
  AOI22_X1 U4575 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n3430), .B1(n4406), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4113) );
  AOI22_X1 U4576 ( .A1(n4342), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4112) );
  AOI22_X1 U4577 ( .A1(n4371), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4301), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4111) );
  NAND4_X1 U4578 ( .A1(n4114), .A2(n4113), .A3(n4112), .A4(n4111), .ZN(n4120)
         );
  AOI22_X1 U4579 ( .A1(n4307), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4118) );
  AOI22_X1 U4580 ( .A1(n3427), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3622), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4117) );
  AOI22_X1 U4581 ( .A1(n3627), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4116) );
  AOI22_X1 U4582 ( .A1(n4405), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4115) );
  NAND4_X1 U4583 ( .A1(n4118), .A2(n4117), .A3(n4116), .A4(n4115), .ZN(n4119)
         );
  NOR2_X1 U4584 ( .A1(n4120), .A2(n4119), .ZN(n4285) );
  XNOR2_X1 U4585 ( .A(n4284), .B(n4285), .ZN(n4124) );
  NAND2_X1 U4586 ( .A1(n6657), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4121)
         );
  NAND2_X1 U4587 ( .A1(n4425), .A2(n4121), .ZN(n4122) );
  AOI21_X1 U4588 ( .B1(n4427), .B2(EAX_REG_23__SCAN_IN), .A(n4122), .ZN(n4123)
         );
  OAI21_X1 U4589 ( .B1(n4380), .B2(n4124), .A(n4123), .ZN(n4127) );
  INV_X1 U4590 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6337) );
  INV_X1 U4591 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5613) );
  INV_X1 U4592 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5605) );
  XNOR2_X1 U4593 ( .A(n4281), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5365)
         );
  NAND2_X1 U4594 ( .A1(n5365), .A2(n4562), .ZN(n4126) );
  AND2_X1 U4595 ( .A1(n4127), .A2(n4126), .ZN(n5360) );
  AOI22_X1 U4596 ( .A1(n3691), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4405), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4131) );
  AOI22_X1 U4597 ( .A1(n4412), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4342), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4130) );
  AOI22_X1 U4598 ( .A1(n3430), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4129) );
  AOI22_X1 U4599 ( .A1(n3428), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4128) );
  NAND4_X1 U4600 ( .A1(n4131), .A2(n4130), .A3(n4129), .A4(n4128), .ZN(n4137)
         );
  AOI22_X1 U4601 ( .A1(n3427), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4135) );
  AOI22_X1 U4602 ( .A1(n3429), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4134) );
  AOI22_X1 U4603 ( .A1(n3622), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4133) );
  AOI22_X1 U4604 ( .A1(n4371), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4132) );
  NAND4_X1 U4605 ( .A1(n4135), .A2(n4134), .A3(n4133), .A4(n4132), .ZN(n4136)
         );
  NOR2_X1 U4606 ( .A1(n4137), .A2(n4136), .ZN(n4138) );
  OR2_X1 U4607 ( .A1(n4380), .A2(n4138), .ZN(n4147) );
  NAND2_X1 U4608 ( .A1(n6657), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4139)
         );
  NAND2_X1 U4609 ( .A1(n4425), .A2(n4139), .ZN(n4140) );
  AOI21_X1 U4610 ( .B1(n4427), .B2(EAX_REG_22__SCAN_IN), .A(n4140), .ZN(n4146)
         );
  INV_X1 U4611 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4143) );
  INV_X1 U4612 ( .A(n4141), .ZN(n4142) );
  NAND2_X1 U4613 ( .A1(n4143), .A2(n4142), .ZN(n4144) );
  NAND2_X1 U4614 ( .A1(n4281), .A2(n4144), .ZN(n6396) );
  NOR2_X1 U4615 ( .A1(n6396), .A2(n4425), .ZN(n4145) );
  AOI21_X1 U4616 ( .B1(n4147), .B2(n4146), .A(n4145), .ZN(n5433) );
  INV_X1 U4617 ( .A(n5433), .ZN(n4264) );
  AOI22_X1 U4618 ( .A1(n4412), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4151) );
  AOI22_X1 U4619 ( .A1(n3691), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4405), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4150) );
  AOI22_X1 U4620 ( .A1(n4371), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4149) );
  AOI22_X1 U4621 ( .A1(n3699), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4342), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4148) );
  NAND4_X1 U4622 ( .A1(n4151), .A2(n4150), .A3(n4149), .A4(n4148), .ZN(n4157)
         );
  AOI22_X1 U4623 ( .A1(n3429), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4155) );
  AOI22_X1 U4624 ( .A1(n3430), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4154) );
  AOI22_X1 U4625 ( .A1(n3427), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4153) );
  AOI22_X1 U4626 ( .A1(n4388), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4152) );
  NAND4_X1 U4627 ( .A1(n4155), .A2(n4154), .A3(n4153), .A4(n4152), .ZN(n4156)
         );
  NOR2_X1 U4628 ( .A1(n4157), .A2(n4156), .ZN(n4160) );
  INV_X1 U4629 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5598) );
  AOI21_X1 U4630 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n5598), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4158) );
  AOI21_X1 U4631 ( .B1(n4427), .B2(EAX_REG_21__SCAN_IN), .A(n4158), .ZN(n4159)
         );
  OAI21_X1 U4632 ( .B1(n4380), .B2(n4160), .A(n4159), .ZN(n4162) );
  XNOR2_X1 U4633 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .B(n4177), .ZN(n5600)
         );
  NAND2_X1 U4634 ( .A1(n4562), .A2(n5600), .ZN(n4161) );
  AND2_X1 U4635 ( .A1(n4162), .A2(n4161), .ZN(n5378) );
  INV_X1 U4636 ( .A(n5378), .ZN(n4263) );
  AOI22_X1 U4637 ( .A1(n3627), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4166) );
  AOI22_X1 U4638 ( .A1(n4412), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4165) );
  AOI22_X1 U4639 ( .A1(n3427), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4164) );
  AOI22_X1 U4640 ( .A1(n4371), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4163) );
  NAND4_X1 U4641 ( .A1(n4166), .A2(n4165), .A3(n4164), .A4(n4163), .ZN(n4172)
         );
  AOI22_X1 U4642 ( .A1(n3622), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4342), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4170) );
  AOI22_X1 U4643 ( .A1(n3429), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4169) );
  AOI22_X1 U4644 ( .A1(n3430), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4168) );
  AOI22_X1 U4645 ( .A1(n4405), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4167) );
  NAND4_X1 U4646 ( .A1(n4170), .A2(n4169), .A3(n4168), .A4(n4167), .ZN(n4171)
         );
  NOR2_X1 U4647 ( .A1(n4172), .A2(n4171), .ZN(n4176) );
  OAI21_X1 U4648 ( .B1(PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6670), .A(n6657), 
        .ZN(n4173) );
  INV_X1 U4649 ( .A(n4173), .ZN(n4174) );
  AOI21_X1 U4650 ( .B1(n4427), .B2(EAX_REG_20__SCAN_IN), .A(n4174), .ZN(n4175)
         );
  OAI21_X1 U4651 ( .B1(n4380), .B2(n4176), .A(n4175), .ZN(n4180) );
  OAI21_X1 U4652 ( .B1(PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n4178), .A(n4177), 
        .ZN(n6373) );
  OR2_X1 U4653 ( .A1(n4425), .A2(n6373), .ZN(n4179) );
  NAND2_X1 U4654 ( .A1(n4180), .A2(n4179), .ZN(n5449) );
  INV_X1 U4655 ( .A(n5449), .ZN(n4246) );
  AOI22_X1 U4656 ( .A1(n3429), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3430), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4184) );
  AOI22_X1 U4657 ( .A1(n4405), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4183) );
  AOI22_X1 U4658 ( .A1(n4342), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4182) );
  AOI22_X1 U4659 ( .A1(n3428), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4181) );
  NAND4_X1 U4660 ( .A1(n4184), .A2(n4183), .A3(n4182), .A4(n4181), .ZN(n4190)
         );
  AOI22_X1 U4661 ( .A1(n4412), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4188) );
  AOI22_X1 U4662 ( .A1(n3427), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3622), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4187) );
  AOI22_X1 U4663 ( .A1(n3627), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4186) );
  AOI22_X1 U4664 ( .A1(n4371), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4185) );
  NAND4_X1 U4665 ( .A1(n4188), .A2(n4187), .A3(n4186), .A4(n4185), .ZN(n4189)
         );
  NOR2_X1 U4666 ( .A1(n4190), .A2(n4189), .ZN(n4193) );
  AOI21_X1 U4667 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n5605), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4191) );
  AOI21_X1 U4668 ( .B1(n4427), .B2(EAX_REG_19__SCAN_IN), .A(n4191), .ZN(n4192)
         );
  OAI21_X1 U4669 ( .B1(n4380), .B2(n4193), .A(n4192), .ZN(n4195) );
  XNOR2_X1 U4670 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .B(n4210), .ZN(n5607)
         );
  NAND2_X1 U4671 ( .A1(n4562), .A2(n5607), .ZN(n4194) );
  NAND2_X1 U4672 ( .A1(n4195), .A2(n4194), .ZN(n5389) );
  INV_X1 U4673 ( .A(n5389), .ZN(n4245) );
  AOI22_X1 U4674 ( .A1(n4412), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3427), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4199) );
  AOI22_X1 U4675 ( .A1(n3622), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4342), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4198) );
  AOI22_X1 U4676 ( .A1(n3627), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4197) );
  AOI22_X1 U4677 ( .A1(n4371), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4301), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4196) );
  NAND4_X1 U4678 ( .A1(n4199), .A2(n4198), .A3(n4197), .A4(n4196), .ZN(n4205)
         );
  AOI22_X1 U4679 ( .A1(n4405), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4203) );
  AOI22_X1 U4680 ( .A1(n3429), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4202) );
  AOI22_X1 U4681 ( .A1(n3430), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4201) );
  AOI22_X1 U4682 ( .A1(n4366), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4200) );
  NAND4_X1 U4683 ( .A1(n4203), .A2(n4202), .A3(n4201), .A4(n4200), .ZN(n4204)
         );
  NOR2_X1 U4684 ( .A1(n4205), .A2(n4204), .ZN(n4209) );
  NAND2_X1 U4685 ( .A1(n6657), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4206)
         );
  NAND2_X1 U4686 ( .A1(n4425), .A2(n4206), .ZN(n4207) );
  AOI21_X1 U4687 ( .B1(n4427), .B2(EAX_REG_18__SCAN_IN), .A(n4207), .ZN(n4208)
         );
  OAI21_X1 U4688 ( .B1(n4380), .B2(n4209), .A(n4208), .ZN(n4213) );
  OAI21_X1 U4689 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n4211), .A(n4210), 
        .ZN(n6363) );
  OR2_X1 U4690 ( .A1(n4425), .A2(n6363), .ZN(n4212) );
  NAND2_X1 U4691 ( .A1(n4213), .A2(n4212), .ZN(n5455) );
  INV_X1 U4692 ( .A(n5455), .ZN(n4244) );
  XNOR2_X1 U4693 ( .A(n4214), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5615)
         );
  AOI22_X1 U4694 ( .A1(n3427), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4218) );
  AOI22_X1 U4695 ( .A1(n3622), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4342), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4217) );
  AOI22_X1 U4696 ( .A1(n4405), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4216) );
  AOI22_X1 U4697 ( .A1(n3430), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4215) );
  NAND4_X1 U4698 ( .A1(n4218), .A2(n4217), .A3(n4216), .A4(n4215), .ZN(n4224)
         );
  AOI22_X1 U4699 ( .A1(n3429), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3627), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4222) );
  AOI22_X1 U4700 ( .A1(n4412), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4221) );
  AOI22_X1 U4701 ( .A1(n3428), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4220) );
  AOI22_X1 U4702 ( .A1(n4371), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4301), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4219) );
  NAND4_X1 U4703 ( .A1(n4222), .A2(n4221), .A3(n4220), .A4(n4219), .ZN(n4223)
         );
  OR2_X1 U4704 ( .A1(n4224), .A2(n4223), .ZN(n4227) );
  NAND2_X1 U4705 ( .A1(n4427), .A2(EAX_REG_17__SCAN_IN), .ZN(n4225) );
  OAI211_X1 U4706 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n5613), .A(n4225), .B(
        n4425), .ZN(n4226) );
  AOI21_X1 U4707 ( .B1(n4422), .B2(n4227), .A(n4226), .ZN(n4228) );
  AOI21_X1 U4708 ( .B1(n5615), .B2(n4562), .A(n4228), .ZN(n5403) );
  XOR2_X1 U4709 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n4229), .Z(n6353) );
  AOI22_X1 U4710 ( .A1(n4412), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3622), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4233) );
  AOI22_X1 U4711 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n3429), .B1(n4342), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4232) );
  AOI22_X1 U4712 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4405), .B1(n4413), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4231) );
  AOI22_X1 U4713 ( .A1(n3428), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4301), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4230) );
  NAND4_X1 U4714 ( .A1(n4233), .A2(n4232), .A3(n4231), .A4(n4230), .ZN(n4239)
         );
  AOI22_X1 U4715 ( .A1(n3427), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4237) );
  AOI22_X1 U4716 ( .A1(n3430), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4236) );
  AOI22_X1 U4717 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n3627), .B1(n4406), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4235) );
  AOI22_X1 U4718 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4371), .B1(n4308), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4234) );
  NAND4_X1 U4719 ( .A1(n4237), .A2(n4236), .A3(n4235), .A4(n4234), .ZN(n4238)
         );
  OR2_X1 U4720 ( .A1(n4239), .A2(n4238), .ZN(n4242) );
  INV_X1 U4721 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4240) );
  INV_X1 U4722 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5626) );
  OAI22_X1 U4723 ( .A1(n4399), .A2(n4240), .B1(n4283), .B2(n5626), .ZN(n4241)
         );
  AOI21_X1 U4724 ( .B1(n4422), .B2(n4242), .A(n4241), .ZN(n4243) );
  OAI21_X1 U4725 ( .B1(n6353), .B2(n4425), .A(n4243), .ZN(n5469) );
  AND2_X1 U4726 ( .A1(n5403), .A2(n5469), .ZN(n5402) );
  AND2_X1 U4727 ( .A1(n4244), .A2(n5402), .ZN(n5388) );
  AND2_X1 U4728 ( .A1(n4245), .A2(n5388), .ZN(n5387) );
  NAND2_X1 U4729 ( .A1(n4246), .A2(n5387), .ZN(n4262) );
  XNOR2_X1 U4730 ( .A(n4247), .B(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5639)
         );
  AOI22_X1 U4731 ( .A1(n3429), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4251) );
  AOI22_X1 U4732 ( .A1(n4366), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4250) );
  AOI22_X1 U4733 ( .A1(n3627), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4249) );
  AOI22_X1 U4734 ( .A1(n3428), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4248) );
  NAND4_X1 U4735 ( .A1(n4251), .A2(n4250), .A3(n4249), .A4(n4248), .ZN(n4257)
         );
  AOI22_X1 U4736 ( .A1(n4412), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3427), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4255) );
  AOI22_X1 U4737 ( .A1(n4405), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3430), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4254) );
  AOI22_X1 U4738 ( .A1(n3622), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4342), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4253) );
  AOI22_X1 U4739 ( .A1(n4371), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4301), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4252) );
  NAND4_X1 U4740 ( .A1(n4255), .A2(n4254), .A3(n4253), .A4(n4252), .ZN(n4256)
         );
  OAI21_X1 U4741 ( .B1(n4257), .B2(n4256), .A(n4274), .ZN(n4260) );
  NAND2_X1 U4742 ( .A1(n4427), .A2(EAX_REG_15__SCAN_IN), .ZN(n4259) );
  NAND2_X1 U4743 ( .A1(n5191), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4258)
         );
  NAND3_X1 U4744 ( .A1(n4260), .A2(n4259), .A3(n4258), .ZN(n4261) );
  AOI21_X1 U4745 ( .B1(n5639), .B2(n4562), .A(n4261), .ZN(n5413) );
  OR2_X1 U4746 ( .A1(n4262), .A2(n5413), .ZN(n5375) );
  NOR2_X1 U4747 ( .A1(n4264), .A2(n5376), .ZN(n5358) );
  AND2_X1 U4748 ( .A1(n5360), .A2(n5358), .ZN(n4279) );
  XOR2_X1 U4749 ( .A(n6337), .B(n4265), .Z(n6341) );
  AOI22_X1 U4750 ( .A1(n4427), .A2(EAX_REG_14__SCAN_IN), .B1(n5191), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4278) );
  AOI22_X1 U4751 ( .A1(n3429), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3691), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4269) );
  AOI22_X1 U4752 ( .A1(n4412), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3427), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4268) );
  AOI22_X1 U4753 ( .A1(n4342), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4267) );
  AOI22_X1 U4754 ( .A1(n4405), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4266) );
  NAND4_X1 U4755 ( .A1(n4269), .A2(n4268), .A3(n4267), .A4(n4266), .ZN(n4276)
         );
  AOI22_X1 U4756 ( .A1(n4366), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3699), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4273) );
  AOI22_X1 U4757 ( .A1(n3428), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4272) );
  AOI22_X1 U4758 ( .A1(n3430), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4271) );
  AOI22_X1 U4759 ( .A1(n4371), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4301), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4270) );
  NAND4_X1 U4760 ( .A1(n4273), .A2(n4272), .A3(n4271), .A4(n4270), .ZN(n4275)
         );
  OAI21_X1 U4761 ( .B1(n4276), .B2(n4275), .A(n4274), .ZN(n4277) );
  OAI211_X1 U4762 ( .C1(n6341), .C2(n4425), .A(n4278), .B(n4277), .ZN(n5482)
         );
  XNOR2_X1 U4763 ( .A(n4299), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5574)
         );
  INV_X1 U4764 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5576) );
  OAI22_X1 U4765 ( .A1(n5574), .A2(n4425), .B1(n5576), .B2(n4283), .ZN(n4298)
         );
  OR2_X1 U4766 ( .A1(n4285), .A2(n4284), .ZN(n4316) );
  AOI22_X1 U4767 ( .A1(n4307), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4342), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4289) );
  AOI22_X1 U4768 ( .A1(n3429), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3430), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4288) );
  AOI22_X1 U4769 ( .A1(n3427), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3699), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4287) );
  AOI22_X1 U4770 ( .A1(n4371), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4301), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4286) );
  NAND4_X1 U4771 ( .A1(n4289), .A2(n4288), .A3(n4287), .A4(n4286), .ZN(n4295)
         );
  AOI22_X1 U4772 ( .A1(n3627), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4405), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4293) );
  AOI22_X1 U4773 ( .A1(n3428), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4292) );
  AOI22_X1 U4774 ( .A1(n4366), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4291) );
  AOI22_X1 U4775 ( .A1(n3544), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4290) );
  NAND4_X1 U4776 ( .A1(n4293), .A2(n4292), .A3(n4291), .A4(n4290), .ZN(n4294)
         );
  NOR2_X1 U4777 ( .A1(n4295), .A2(n4294), .ZN(n4315) );
  XNOR2_X1 U4778 ( .A(n4316), .B(n4315), .ZN(n4296) );
  NOR2_X1 U4779 ( .A1(n4380), .A2(n4296), .ZN(n4297) );
  AOI211_X1 U4780 ( .C1(n4427), .C2(EAX_REG_24__SCAN_IN), .A(n4298), .B(n4297), 
        .ZN(n5345) );
  NOR2_X2 U4781 ( .A1(n5361), .A2(n5345), .ZN(n5330) );
  XNOR2_X1 U4782 ( .A(n4321), .B(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5559)
         );
  AOI22_X1 U4783 ( .A1(n4405), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4305) );
  AOI22_X1 U4784 ( .A1(n3430), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4304) );
  AOI22_X1 U4785 ( .A1(n3699), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4303) );
  AOI22_X1 U4786 ( .A1(n3428), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4301), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4302) );
  NAND4_X1 U4787 ( .A1(n4305), .A2(n4304), .A3(n4303), .A4(n4302), .ZN(n4314)
         );
  AOI22_X1 U4788 ( .A1(n4307), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4312) );
  AOI22_X1 U4789 ( .A1(n3429), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3691), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4311) );
  AOI22_X1 U4790 ( .A1(n3427), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4342), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4310) );
  AOI22_X1 U4791 ( .A1(n4371), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4309) );
  NAND4_X1 U4792 ( .A1(n4312), .A2(n4311), .A3(n4310), .A4(n4309), .ZN(n4313)
         );
  NOR2_X1 U4793 ( .A1(n4314), .A2(n4313), .ZN(n4327) );
  OR2_X1 U4794 ( .A1(n4316), .A2(n4315), .ZN(n4326) );
  XOR2_X1 U4795 ( .A(n4327), .B(n4326), .Z(n4319) );
  INV_X1 U4796 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5337) );
  NAND2_X1 U4797 ( .A1(n4427), .A2(EAX_REG_25__SCAN_IN), .ZN(n4317) );
  OAI211_X1 U4798 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n5337), .A(n4317), .B(
        n4425), .ZN(n4318) );
  AOI21_X1 U4799 ( .B1(n4319), .B2(n4422), .A(n4318), .ZN(n4320) );
  AOI21_X1 U4800 ( .B1(n4562), .B2(n5559), .A(n4320), .ZN(n5331) );
  NAND2_X1 U4801 ( .A1(n5330), .A2(n5331), .ZN(n5315) );
  INV_X1 U4802 ( .A(n4321), .ZN(n4322) );
  INV_X1 U4803 ( .A(n4323), .ZN(n4324) );
  INV_X1 U4804 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5318) );
  NAND2_X1 U4805 ( .A1(n4324), .A2(n5318), .ZN(n4325) );
  NAND2_X1 U4806 ( .A1(n4359), .A2(n4325), .ZN(n5552) );
  NOR2_X1 U4807 ( .A1(n4327), .A2(n4326), .ZN(n4354) );
  AOI22_X1 U4808 ( .A1(n4412), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4331) );
  AOI22_X1 U4809 ( .A1(n3427), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3622), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4330) );
  AOI22_X1 U4810 ( .A1(n3430), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4329) );
  AOI22_X1 U4811 ( .A1(n4342), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4328) );
  NAND4_X1 U4812 ( .A1(n4331), .A2(n4330), .A3(n4329), .A4(n4328), .ZN(n4337)
         );
  AOI22_X1 U4813 ( .A1(n3429), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3691), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4335) );
  AOI22_X1 U4814 ( .A1(n4405), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4334) );
  AOI22_X1 U4815 ( .A1(n3428), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4333) );
  AOI22_X1 U4816 ( .A1(n4371), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4332) );
  NAND4_X1 U4817 ( .A1(n4335), .A2(n4334), .A3(n4333), .A4(n4332), .ZN(n4336)
         );
  OR2_X1 U4818 ( .A1(n4337), .A2(n4336), .ZN(n4353) );
  XNOR2_X1 U4819 ( .A(n4354), .B(n4353), .ZN(n4340) );
  AOI21_X1 U4820 ( .B1(PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6657), .A(n4562), 
        .ZN(n4339) );
  NAND2_X1 U4821 ( .A1(n4427), .A2(EAX_REG_26__SCAN_IN), .ZN(n4338) );
  OAI211_X1 U4822 ( .C1(n4340), .C2(n4380), .A(n4339), .B(n4338), .ZN(n4341)
         );
  OAI21_X1 U4823 ( .B1(n4425), .B2(n5552), .A(n4341), .ZN(n5317) );
  AOI22_X1 U4824 ( .A1(n4366), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4342), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4346) );
  AOI22_X1 U4825 ( .A1(n4405), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4345) );
  AOI22_X1 U4826 ( .A1(n3429), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4344) );
  AOI22_X1 U4827 ( .A1(n3430), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4343) );
  NAND4_X1 U4828 ( .A1(n4346), .A2(n4345), .A3(n4344), .A4(n4343), .ZN(n4352)
         );
  AOI22_X1 U4829 ( .A1(n4412), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3427), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4350) );
  AOI22_X1 U4830 ( .A1(n3691), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3699), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4349) );
  AOI22_X1 U4831 ( .A1(n3428), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4348) );
  AOI22_X1 U4832 ( .A1(n4371), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4347) );
  NAND4_X1 U4833 ( .A1(n4350), .A2(n4349), .A3(n4348), .A4(n4347), .ZN(n4351)
         );
  NOR2_X1 U4834 ( .A1(n4352), .A2(n4351), .ZN(n4365) );
  NAND2_X1 U4835 ( .A1(n4354), .A2(n4353), .ZN(n4364) );
  XOR2_X1 U4836 ( .A(n4365), .B(n4364), .Z(n4355) );
  NAND2_X1 U4837 ( .A1(n4355), .A2(n4422), .ZN(n4358) );
  INV_X1 U4838 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5308) );
  NOR2_X1 U4839 ( .A1(n5308), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4356) );
  AOI211_X1 U4840 ( .C1(n4427), .C2(EAX_REG_27__SCAN_IN), .A(n4562), .B(n4356), 
        .ZN(n4357) );
  XNOR2_X1 U4841 ( .A(n4359), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5307)
         );
  AOI22_X1 U4842 ( .A1(n4358), .A2(n4357), .B1(n4562), .B2(n5307), .ZN(n5301)
         );
  NAND2_X1 U4843 ( .A1(n5300), .A2(n5301), .ZN(n5289) );
  INV_X1 U4844 ( .A(n4359), .ZN(n4360) );
  INV_X1 U4845 ( .A(n4361), .ZN(n4362) );
  INV_X1 U4846 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5292) );
  NAND2_X1 U4847 ( .A1(n4362), .A2(n5292), .ZN(n4363) );
  NAND2_X1 U4848 ( .A1(n4428), .A2(n4363), .ZN(n5535) );
  NOR2_X1 U4849 ( .A1(n4365), .A2(n4364), .ZN(n4396) );
  AOI22_X1 U4850 ( .A1(n4412), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4366), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4370) );
  AOI22_X1 U4851 ( .A1(n3427), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3699), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4369) );
  AOI22_X1 U4852 ( .A1(n3430), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4368) );
  AOI22_X1 U4853 ( .A1(n4342), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4367) );
  NAND4_X1 U4854 ( .A1(n4370), .A2(n4369), .A3(n4368), .A4(n4367), .ZN(n4377)
         );
  AOI22_X1 U4855 ( .A1(n3429), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3627), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4375) );
  AOI22_X1 U4856 ( .A1(n4405), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4374) );
  AOI22_X1 U4857 ( .A1(n3428), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4373) );
  AOI22_X1 U4858 ( .A1(n4371), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4372) );
  NAND4_X1 U4859 ( .A1(n4375), .A2(n4374), .A3(n4373), .A4(n4372), .ZN(n4376)
         );
  OR2_X1 U4860 ( .A1(n4377), .A2(n4376), .ZN(n4395) );
  XNOR2_X1 U4861 ( .A(n4396), .B(n4395), .ZN(n4381) );
  AOI21_X1 U4862 ( .B1(PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6657), .A(n4562), 
        .ZN(n4379) );
  NAND2_X1 U4863 ( .A1(n4427), .A2(EAX_REG_28__SCAN_IN), .ZN(n4378) );
  OAI211_X1 U4864 ( .C1(n4381), .C2(n4380), .A(n4379), .B(n4378), .ZN(n4382)
         );
  OAI21_X1 U4865 ( .B1(n4425), .B2(n5535), .A(n4382), .ZN(n5291) );
  NOR2_X2 U4866 ( .A1(n5289), .A2(n5291), .ZN(n5271) );
  XNOR2_X1 U4867 ( .A(n4428), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5275)
         );
  AOI22_X1 U4868 ( .A1(n3429), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3691), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4387) );
  AOI22_X1 U4869 ( .A1(n4405), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4386) );
  AOI22_X1 U4870 ( .A1(n3430), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4385) );
  AOI22_X1 U4871 ( .A1(n4371), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4384) );
  NAND4_X1 U4872 ( .A1(n4387), .A2(n4386), .A3(n4385), .A4(n4384), .ZN(n4394)
         );
  AOI22_X1 U4873 ( .A1(n4412), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4392) );
  AOI22_X1 U4874 ( .A1(n3427), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3699), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4391) );
  AOI22_X1 U4875 ( .A1(n4342), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4390) );
  AOI22_X1 U4876 ( .A1(n4413), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4389) );
  NAND4_X1 U4877 ( .A1(n4392), .A2(n4391), .A3(n4390), .A4(n4389), .ZN(n4393)
         );
  NOR2_X1 U4878 ( .A1(n4394), .A2(n4393), .ZN(n4404) );
  NAND2_X1 U4879 ( .A1(n4396), .A2(n4395), .ZN(n4403) );
  XOR2_X1 U4880 ( .A(n4404), .B(n4403), .Z(n4401) );
  INV_X1 U4881 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4398) );
  NAND2_X1 U4882 ( .A1(n6657), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4397)
         );
  OAI211_X1 U4883 ( .C1(n4399), .C2(n4398), .A(n4425), .B(n4397), .ZN(n4400)
         );
  AOI21_X1 U4884 ( .B1(n4401), .B2(n4422), .A(n4400), .ZN(n4402) );
  AOI21_X1 U4885 ( .B1(n4562), .B2(n5275), .A(n4402), .ZN(n5270) );
  AND2_X2 U4886 ( .A1(n5271), .A2(n5270), .ZN(n5272) );
  NOR2_X1 U4887 ( .A1(n4404), .A2(n4403), .ZN(n4421) );
  AOI22_X1 U4888 ( .A1(n4405), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4411) );
  AOI22_X1 U4889 ( .A1(n3430), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4410) );
  AOI22_X1 U4890 ( .A1(n4342), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4409) );
  AOI22_X1 U4891 ( .A1(n4371), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4301), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4408) );
  NAND4_X1 U4892 ( .A1(n4411), .A2(n4410), .A3(n4409), .A4(n4408), .ZN(n4419)
         );
  AOI22_X1 U4893 ( .A1(n4412), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4417) );
  AOI22_X1 U4894 ( .A1(n3429), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3691), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4416) );
  AOI22_X1 U4895 ( .A1(n3427), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3699), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4415) );
  AOI22_X1 U4896 ( .A1(n4413), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4414) );
  NAND4_X1 U4897 ( .A1(n4417), .A2(n4416), .A3(n4415), .A4(n4414), .ZN(n4418)
         );
  NOR2_X1 U4898 ( .A1(n4419), .A2(n4418), .ZN(n4420) );
  XNOR2_X1 U4899 ( .A(n4421), .B(n4420), .ZN(n4423) );
  NAND2_X1 U4900 ( .A1(n4423), .A2(n4422), .ZN(n4431) );
  NAND2_X1 U4901 ( .A1(n6657), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4424)
         );
  NAND2_X1 U4902 ( .A1(n4425), .A2(n4424), .ZN(n4426) );
  AOI21_X1 U4903 ( .B1(n4427), .B2(EAX_REG_30__SCAN_IN), .A(n4426), .ZN(n4430)
         );
  INV_X1 U4904 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5276) );
  XNOR2_X1 U4905 ( .A(n4567), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4574)
         );
  AND2_X1 U4906 ( .A1(n4574), .A2(n4562), .ZN(n4429) );
  AOI21_X1 U4907 ( .B1(n4431), .B2(n4430), .A(n4429), .ZN(n5190) );
  NOR2_X1 U4908 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6655) );
  NAND2_X1 U4909 ( .A1(n6491), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4622) );
  INV_X1 U4910 ( .A(n4622), .ZN(n4561) );
  NAND2_X1 U4911 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n4561), .ZN(n6144) );
  INV_X1 U4912 ( .A(n6144), .ZN(n4432) );
  AND2_X2 U4913 ( .A1(n6655), .A2(n4432), .ZN(n6969) );
  INV_X1 U4914 ( .A(n6969), .ZN(n6862) );
  INV_X1 U4915 ( .A(n6655), .ZN(n6622) );
  NAND2_X1 U4916 ( .A1(n6622), .A2(n4433), .ZN(n6151) );
  NAND2_X1 U4917 ( .A1(n6151), .A2(n6491), .ZN(n4434) );
  NAND2_X1 U4918 ( .A1(n6491), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4436) );
  NAND2_X1 U4919 ( .A1(n6670), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4435) );
  NAND2_X1 U4920 ( .A1(n4436), .A2(n4435), .ZN(n4638) );
  INV_X1 U4921 ( .A(n4638), .ZN(n4437) );
  NAND2_X1 U4922 ( .A1(n6655), .A2(n6440), .ZN(n6134) );
  OR2_X2 U4923 ( .A1(n6134), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6247) );
  INV_X1 U4924 ( .A(REIP_REG_30__SCAN_IN), .ZN(n5951) );
  NOR2_X1 U4925 ( .A1(n6247), .A2(n5951), .ZN(n5660) );
  INV_X1 U4926 ( .A(n6119), .ZN(n5627) );
  INV_X1 U4927 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4566) );
  NOR2_X1 U4928 ( .A1(n5627), .A2(n4566), .ZN(n4438) );
  AOI211_X1 U4929 ( .C1(n4574), .C2(n6104), .A(n5660), .B(n4438), .ZN(n4439)
         );
  NAND3_X1 U4930 ( .A1(n4441), .A2(n4440), .A3(n4439), .ZN(U2956) );
  NAND2_X4 U4931 ( .A1(n6780), .A2(n4831), .ZN(n4543) );
  NAND2_X1 U4932 ( .A1(n4448), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4442)
         );
  NAND2_X1 U4933 ( .A1(n4543), .A2(n4442), .ZN(n4447) );
  NAND2_X1 U4934 ( .A1(n4444), .A2(n4443), .ZN(n4455) );
  INV_X1 U4935 ( .A(n4455), .ZN(n4449) );
  NAND2_X1 U4936 ( .A1(n4449), .A2(n4445), .ZN(n4446) );
  INV_X2 U4937 ( .A(n4448), .ZN(n4645) );
  NAND2_X2 U4938 ( .A1(n4645), .A2(n4449), .ZN(n4547) );
  OR2_X1 U4939 ( .A1(n4547), .A2(EBX_REG_1__SCAN_IN), .ZN(n4450) );
  NAND2_X1 U4940 ( .A1(n4543), .A2(EBX_REG_0__SCAN_IN), .ZN(n4454) );
  INV_X1 U4941 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4452) );
  NAND2_X1 U4942 ( .A1(n4448), .A2(n4452), .ZN(n4453) );
  NAND2_X1 U4943 ( .A1(n4454), .A2(n4453), .ZN(n4739) );
  XNOR2_X1 U4944 ( .A(n4456), .B(n4739), .ZN(n4671) );
  NAND2_X1 U4945 ( .A1(n4669), .A2(n4456), .ZN(n6078) );
  MUX2_X1 U4946 ( .A(n4539), .B(n3431), .S(EBX_REG_3__SCAN_IN), .Z(n4458) );
  OR2_X1 U4947 ( .A1(n5184), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4457)
         );
  OR2_X1 U4948 ( .A1(n4547), .A2(EBX_REG_2__SCAN_IN), .ZN(n4462) );
  INV_X1 U4949 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4459) );
  NAND2_X1 U4950 ( .A1(n4543), .A2(n4459), .ZN(n4460) );
  OAI211_X1 U4951 ( .C1(n4518), .C2(EBX_REG_2__SCAN_IN), .A(n4460), .B(n3431), 
        .ZN(n4461) );
  NAND2_X1 U4952 ( .A1(n4462), .A2(n4461), .ZN(n6077) );
  NAND2_X1 U4953 ( .A1(n4823), .A2(n6077), .ZN(n4463) );
  NOR2_X2 U4954 ( .A1(n6078), .A2(n4463), .ZN(n4825) );
  OR2_X1 U4955 ( .A1(n4547), .A2(EBX_REG_4__SCAN_IN), .ZN(n4467) );
  NAND2_X1 U4956 ( .A1(n3431), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4464)
         );
  NAND2_X1 U4957 ( .A1(n4543), .A2(n4464), .ZN(n4465) );
  OAI21_X1 U4958 ( .B1(EBX_REG_4__SCAN_IN), .B2(n4518), .A(n4465), .ZN(n4466)
         );
  NAND2_X1 U4959 ( .A1(n4467), .A2(n4466), .ZN(n4595) );
  NAND2_X1 U4960 ( .A1(n4825), .A2(n4595), .ZN(n4594) );
  INV_X1 U4961 ( .A(n4594), .ZN(n4470) );
  MUX2_X1 U4962 ( .A(n4539), .B(n3431), .S(EBX_REG_5__SCAN_IN), .Z(n4468) );
  OAI21_X1 U4963 ( .B1(n3432), .B2(INSTADDRPOINTER_REG_5__SCAN_IN), .A(n4468), 
        .ZN(n4938) );
  INV_X1 U4964 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6291) );
  NAND2_X1 U4965 ( .A1(n4524), .A2(n6291), .ZN(n4474) );
  NAND2_X1 U4966 ( .A1(n4543), .A2(n4471), .ZN(n4472) );
  OAI211_X1 U4967 ( .C1(n4518), .C2(EBX_REG_6__SCAN_IN), .A(n4472), .B(n3431), 
        .ZN(n4473) );
  MUX2_X1 U4968 ( .A(n4539), .B(n3431), .S(EBX_REG_7__SCAN_IN), .Z(n4477) );
  OAI21_X1 U4969 ( .B1(n3432), .B2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n4477), 
        .ZN(n4980) );
  INV_X1 U4970 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5053) );
  NAND2_X1 U4971 ( .A1(n4524), .A2(n5053), .ZN(n4481) );
  NAND2_X1 U4972 ( .A1(n4543), .A2(n4478), .ZN(n4479) );
  OAI211_X1 U4973 ( .C1(n4518), .C2(EBX_REG_8__SCAN_IN), .A(n4479), .B(n3431), 
        .ZN(n4480) );
  NAND2_X1 U4974 ( .A1(n4481), .A2(n4480), .ZN(n5026) );
  AND2_X2 U4975 ( .A1(n5027), .A2(n5026), .ZN(n5025) );
  OR2_X1 U4976 ( .A1(n3432), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4483)
         );
  MUX2_X1 U4977 ( .A(n4539), .B(n3431), .S(EBX_REG_9__SCAN_IN), .Z(n4482) );
  AND2_X1 U4978 ( .A1(n4483), .A2(n4482), .ZN(n5127) );
  INV_X1 U4979 ( .A(EBX_REG_10__SCAN_IN), .ZN(n4484) );
  NAND2_X1 U4980 ( .A1(n4524), .A2(n4484), .ZN(n4488) );
  NAND2_X1 U4981 ( .A1(n4543), .A2(n4485), .ZN(n4486) );
  OAI211_X1 U4982 ( .C1(n4518), .C2(EBX_REG_10__SCAN_IN), .A(n4486), .B(n3431), 
        .ZN(n4487) );
  MUX2_X1 U4983 ( .A(n4539), .B(n3431), .S(EBX_REG_11__SCAN_IN), .Z(n4492) );
  OR2_X1 U4984 ( .A1(n3432), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4491)
         );
  NAND2_X1 U4985 ( .A1(n4492), .A2(n4491), .ZN(n5152) );
  NOR2_X2 U4986 ( .A1(n5153), .A2(n5152), .ZN(n5154) );
  OR2_X1 U4987 ( .A1(n4547), .A2(EBX_REG_12__SCAN_IN), .ZN(n4496) );
  NAND2_X1 U4988 ( .A1(n3431), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4493) );
  NAND2_X1 U4989 ( .A1(n4543), .A2(n4493), .ZN(n4494) );
  OAI21_X1 U4990 ( .B1(EBX_REG_12__SCAN_IN), .B2(n4518), .A(n4494), .ZN(n4495)
         );
  NAND2_X1 U4991 ( .A1(n4496), .A2(n4495), .ZN(n5095) );
  MUX2_X1 U4992 ( .A(n4539), .B(n3431), .S(EBX_REG_13__SCAN_IN), .Z(n4497) );
  OAI21_X1 U4993 ( .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n3432), .A(n4497), 
        .ZN(n5181) );
  INV_X1 U4994 ( .A(EBX_REG_14__SCAN_IN), .ZN(n6336) );
  NAND2_X1 U4995 ( .A1(n4524), .A2(n6336), .ZN(n4502) );
  NAND2_X1 U4996 ( .A1(n4543), .A2(n5644), .ZN(n4500) );
  OAI211_X1 U4997 ( .C1(n4518), .C2(EBX_REG_14__SCAN_IN), .A(n4500), .B(n3431), 
        .ZN(n4501) );
  AND2_X1 U4998 ( .A1(n4502), .A2(n4501), .ZN(n5483) );
  OR2_X2 U4999 ( .A1(n5484), .A2(n5483), .ZN(n5486) );
  MUX2_X1 U5000 ( .A(n4539), .B(n3431), .S(EBX_REG_15__SCAN_IN), .Z(n4503) );
  OAI21_X1 U5001 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n3432), .A(n4503), 
        .ZN(n5415) );
  INV_X1 U5002 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5475) );
  NAND2_X1 U5003 ( .A1(n4524), .A2(n5475), .ZN(n4506) );
  NAND2_X1 U5004 ( .A1(n4543), .A2(n6230), .ZN(n4504) );
  OAI211_X1 U5005 ( .C1(n4518), .C2(EBX_REG_16__SCAN_IN), .A(n4504), .B(n3431), 
        .ZN(n4505) );
  NAND2_X1 U5006 ( .A1(n4506), .A2(n4505), .ZN(n5471) );
  NAND2_X1 U5007 ( .A1(n5472), .A2(n5471), .ZN(n5474) );
  MUX2_X1 U5008 ( .A(n4539), .B(n3431), .S(EBX_REG_17__SCAN_IN), .Z(n4508) );
  OR2_X1 U5009 ( .A1(n3432), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4507)
         );
  NAND2_X1 U5010 ( .A1(n4508), .A2(n4507), .ZN(n5404) );
  INV_X1 U5011 ( .A(n4509), .ZN(n5460) );
  INV_X1 U5012 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5463) );
  NAND2_X1 U5013 ( .A1(n4524), .A2(n5463), .ZN(n4512) );
  INV_X1 U5014 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5751) );
  NAND2_X1 U5015 ( .A1(n4543), .A2(n5751), .ZN(n4510) );
  OAI211_X1 U5016 ( .C1(n4518), .C2(EBX_REG_18__SCAN_IN), .A(n4510), .B(n3431), 
        .ZN(n4511) );
  AND2_X1 U5017 ( .A1(n4512), .A2(n4511), .ZN(n5459) );
  NOR2_X2 U5018 ( .A1(n5460), .A2(n5459), .ZN(n5461) );
  OR2_X1 U5019 ( .A1(n4539), .A2(EBX_REG_19__SCAN_IN), .ZN(n4515) );
  NAND2_X1 U5020 ( .A1(n3431), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4513) );
  OAI211_X1 U5021 ( .C1(n4518), .C2(EBX_REG_19__SCAN_IN), .A(n4543), .B(n4513), 
        .ZN(n4514) );
  AND2_X1 U5022 ( .A1(n4515), .A2(n4514), .ZN(n5391) );
  AND2_X2 U5023 ( .A1(n5461), .A2(n5391), .ZN(n5447) );
  OR2_X1 U5024 ( .A1(n4547), .A2(EBX_REG_20__SCAN_IN), .ZN(n4520) );
  NAND2_X1 U5025 ( .A1(n3431), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4516) );
  NAND2_X1 U5026 ( .A1(n4543), .A2(n4516), .ZN(n4517) );
  OAI21_X1 U5027 ( .B1(EBX_REG_20__SCAN_IN), .B2(n4518), .A(n4517), .ZN(n4519)
         );
  NAND2_X1 U5028 ( .A1(n4520), .A2(n4519), .ZN(n5446) );
  NAND2_X1 U5029 ( .A1(n5447), .A2(n5446), .ZN(n5382) );
  OR2_X1 U5030 ( .A1(n4539), .A2(EBX_REG_21__SCAN_IN), .ZN(n4523) );
  NAND2_X1 U5031 ( .A1(n3431), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4521) );
  OAI211_X1 U5032 ( .C1(n4518), .C2(EBX_REG_21__SCAN_IN), .A(n4543), .B(n4521), 
        .ZN(n4522) );
  NAND2_X1 U5033 ( .A1(n4523), .A2(n4522), .ZN(n5383) );
  OR2_X2 U5034 ( .A1(n5382), .A2(n5383), .ZN(n5438) );
  INV_X1 U5035 ( .A(EBX_REG_22__SCAN_IN), .ZN(n6383) );
  NAND2_X1 U5036 ( .A1(n4524), .A2(n6383), .ZN(n4527) );
  INV_X1 U5037 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5589) );
  NAND2_X1 U5038 ( .A1(n4543), .A2(n5589), .ZN(n4525) );
  OAI211_X1 U5039 ( .C1(n4518), .C2(EBX_REG_22__SCAN_IN), .A(n4525), .B(n3431), 
        .ZN(n4526) );
  AND2_X1 U5040 ( .A1(n4527), .A2(n4526), .ZN(n5437) );
  OR2_X2 U5041 ( .A1(n5438), .A2(n5437), .ZN(n5440) );
  MUX2_X1 U5042 ( .A(n4539), .B(n3431), .S(EBX_REG_23__SCAN_IN), .Z(n4529) );
  OR2_X1 U5043 ( .A1(n3432), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4528)
         );
  NAND2_X1 U5044 ( .A1(n4529), .A2(n4528), .ZN(n5366) );
  NOR2_X4 U5045 ( .A1(n5440), .A2(n5366), .ZN(n5368) );
  MUX2_X1 U5046 ( .A(n4539), .B(n3431), .S(EBX_REG_25__SCAN_IN), .Z(n4531) );
  OR2_X1 U5047 ( .A1(n3432), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4530)
         );
  NAND2_X1 U5048 ( .A1(n4531), .A2(n4530), .ZN(n5333) );
  OR2_X1 U5049 ( .A1(n4547), .A2(EBX_REG_24__SCAN_IN), .ZN(n4534) );
  INV_X1 U5050 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5713) );
  NAND2_X1 U5051 ( .A1(n4543), .A2(n5713), .ZN(n4532) );
  OAI211_X1 U5052 ( .C1(n4518), .C2(EBX_REG_24__SCAN_IN), .A(n4532), .B(n3431), 
        .ZN(n4533) );
  AND2_X1 U5053 ( .A1(n4534), .A2(n4533), .ZN(n5346) );
  NOR2_X1 U5054 ( .A1(n5333), .A2(n5346), .ZN(n4535) );
  NAND2_X1 U5055 ( .A1(n5368), .A2(n4535), .ZN(n5324) );
  OR2_X1 U5056 ( .A1(n4547), .A2(EBX_REG_26__SCAN_IN), .ZN(n4538) );
  NAND2_X1 U5057 ( .A1(n4543), .A2(n5693), .ZN(n4536) );
  OAI211_X1 U5058 ( .C1(EBX_REG_26__SCAN_IN), .C2(n4518), .A(n4536), .B(n3431), 
        .ZN(n4537) );
  AND2_X1 U5059 ( .A1(n4538), .A2(n4537), .ZN(n5327) );
  OR2_X2 U5060 ( .A1(n5324), .A2(n5327), .ZN(n5325) );
  MUX2_X1 U5061 ( .A(n4539), .B(n3431), .S(EBX_REG_27__SCAN_IN), .Z(n4541) );
  OR2_X1 U5062 ( .A1(n3432), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4540)
         );
  NAND2_X1 U5063 ( .A1(n4541), .A2(n4540), .ZN(n5303) );
  OR2_X1 U5064 ( .A1(n4547), .A2(EBX_REG_28__SCAN_IN), .ZN(n4546) );
  NAND2_X1 U5065 ( .A1(n3431), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4542) );
  NAND2_X1 U5066 ( .A1(n4543), .A2(n4542), .ZN(n4544) );
  OAI21_X1 U5067 ( .B1(EBX_REG_28__SCAN_IN), .B2(n4518), .A(n4544), .ZN(n4545)
         );
  NAND2_X1 U5068 ( .A1(n4546), .A2(n4545), .ZN(n5286) );
  OAI22_X1 U5069 ( .A1(n3432), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        EBX_REG_29__SCAN_IN), .B2(n4518), .ZN(n4548) );
  OAI22_X1 U5070 ( .A1(n4548), .A2(n4645), .B1(EBX_REG_29__SCAN_IN), .B2(n4547), .ZN(n5281) );
  INV_X1 U5071 ( .A(n5288), .ZN(n4549) );
  OAI22_X1 U5072 ( .A1(n3432), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        EBX_REG_30__SCAN_IN), .B2(n4518), .ZN(n5186) );
  INV_X1 U5073 ( .A(n5186), .ZN(n4552) );
  OR3_X1 U5074 ( .A1(n4556), .A2(n4555), .A3(n4554), .ZN(n4557) );
  NAND2_X1 U5075 ( .A1(n4558), .A2(n4557), .ZN(n4560) );
  NAND2_X1 U5076 ( .A1(n4560), .A2(n4559), .ZN(n5259) );
  INV_X1 U5077 ( .A(n5259), .ZN(n5265) );
  OR3_X1 U5078 ( .A1(n5264), .A2(n5265), .A3(n6428), .ZN(n4610) );
  AND2_X1 U5079 ( .A1(n4562), .A2(n4561), .ZN(n6437) );
  INV_X1 U5080 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6678) );
  NOR2_X1 U5081 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n6445) );
  INV_X1 U5082 ( .A(n6445), .ZN(n6148) );
  NOR3_X1 U5083 ( .A1(n6491), .A2(n6678), .A3(n6148), .ZN(n6447) );
  NOR2_X1 U5084 ( .A1(n6437), .A2(n6447), .ZN(n4563) );
  NAND2_X1 U5085 ( .A1(n4563), .A2(n6247), .ZN(n4564) );
  INV_X1 U5086 ( .A(READY_N), .ZN(n6462) );
  NAND2_X1 U5087 ( .A1(n6670), .A2(n6462), .ZN(n4577) );
  NAND2_X1 U5088 ( .A1(EBX_REG_31__SCAN_IN), .A2(n4577), .ZN(n4565) );
  NOR2_X1 U5089 ( .A1(n4576), .A2(n4565), .ZN(n6254) );
  INV_X1 U5090 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5200) );
  XNOR2_X1 U5091 ( .A(n4568), .B(n5200), .ZN(n5239) );
  NOR2_X1 U5092 ( .A1(n5239), .A2(n6440), .ZN(n4569) );
  INV_X1 U5093 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6463) );
  NAND2_X1 U5094 ( .A1(n6458), .A2(n6463), .ZN(n6141) );
  NOR2_X1 U5095 ( .A1(n6141), .A2(n4577), .ZN(n5197) );
  INV_X1 U5096 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5189) );
  NAND3_X1 U5097 ( .A1(n4831), .A2(n4577), .A3(n5189), .ZN(n4570) );
  OAI21_X1 U5098 ( .B1(n3659), .B2(n5197), .A(n4570), .ZN(n4571) );
  INV_X1 U5099 ( .A(n4571), .ZN(n4572) );
  INV_X1 U5100 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5244) );
  AND2_X1 U5101 ( .A1(n5239), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4573) );
  AOI22_X1 U5102 ( .A1(n6354), .A2(n4574), .B1(n6370), .B2(
        PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4575) );
  OAI21_X1 U5103 ( .B1(n6382), .B2(n5244), .A(n4575), .ZN(n4590) );
  INV_X1 U5104 ( .A(n6141), .ZN(n4764) );
  INV_X1 U5105 ( .A(n4577), .ZN(n4578) );
  OAI211_X1 U5106 ( .C1(n4837), .C2(n4764), .A(n4831), .B(n4578), .ZN(n4579)
         );
  INV_X1 U5107 ( .A(n4579), .ZN(n4580) );
  INV_X1 U5108 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6381) );
  INV_X1 U5109 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6380) );
  NOR2_X1 U5110 ( .A1(n6381), .A2(n6380), .ZN(n6379) );
  AND2_X1 U5111 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6379), .ZN(n4586) );
  NAND2_X1 U5112 ( .A1(REIP_REG_11__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .ZN(
        n5142) );
  NAND3_X1 U5113 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .A3(
        REIP_REG_3__SCAN_IN), .ZN(n4601) );
  INV_X1 U5114 ( .A(REIP_REG_4__SCAN_IN), .ZN(n4853) );
  NOR2_X1 U5115 ( .A1(n4601), .A2(n4853), .ZN(n6281) );
  NAND2_X1 U5116 ( .A1(n6281), .A2(REIP_REG_5__SCAN_IN), .ZN(n6290) );
  INV_X1 U5117 ( .A(n6290), .ZN(n6284) );
  NAND2_X1 U5118 ( .A1(n6284), .A2(REIP_REG_6__SCAN_IN), .ZN(n6300) );
  INV_X1 U5119 ( .A(n6300), .ZN(n4581) );
  NAND2_X1 U5120 ( .A1(n4581), .A2(REIP_REG_7__SCAN_IN), .ZN(n5050) );
  INV_X1 U5121 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6019) );
  NOR2_X1 U5122 ( .A1(n5050), .A2(n6019), .ZN(n6315) );
  NAND2_X1 U5123 ( .A1(n6315), .A2(REIP_REG_9__SCAN_IN), .ZN(n5120) );
  NOR2_X1 U5124 ( .A1(n5142), .A2(n5120), .ZN(n5140) );
  NAND2_X1 U5125 ( .A1(REIP_REG_12__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .ZN(
        n6335) );
  INV_X1 U5126 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6177) );
  NOR2_X1 U5127 ( .A1(n6335), .A2(n6177), .ZN(n5418) );
  NAND4_X1 U5128 ( .A1(n5140), .A2(n5418), .A3(REIP_REG_15__SCAN_IN), .A4(
        REIP_REG_16__SCAN_IN), .ZN(n5363) );
  INV_X1 U5129 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6031) );
  NOR2_X1 U5130 ( .A1(n5363), .A2(n6031), .ZN(n5396) );
  NAND4_X1 U5131 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .A3(
        REIP_REG_19__SCAN_IN), .A4(n5396), .ZN(n4585) );
  INV_X1 U5132 ( .A(n4585), .ZN(n4582) );
  NAND2_X1 U5133 ( .A1(n4586), .A2(n4582), .ZN(n4583) );
  NOR2_X1 U5134 ( .A1(n6301), .A2(n4583), .ZN(n5347) );
  NAND2_X1 U5135 ( .A1(n5347), .A2(REIP_REG_24__SCAN_IN), .ZN(n5338) );
  INV_X1 U5136 ( .A(REIP_REG_26__SCAN_IN), .ZN(n5868) );
  INV_X1 U5137 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6043) );
  OR3_X1 U5138 ( .A1(n5338), .A2(n5868), .A3(n6043), .ZN(n5312) );
  INV_X1 U5139 ( .A(n5312), .ZN(n5293) );
  NAND2_X1 U5140 ( .A1(REIP_REG_27__SCAN_IN), .A2(REIP_REG_28__SCAN_IN), .ZN(
        n4587) );
  INV_X1 U5141 ( .A(n4587), .ZN(n4584) );
  NAND2_X1 U5142 ( .A1(n5293), .A2(n4584), .ZN(n5279) );
  INV_X1 U5143 ( .A(REIP_REG_29__SCAN_IN), .ZN(n5955) );
  OAI21_X1 U5144 ( .B1(n5279), .B2(n5955), .A(n5951), .ZN(n4588) );
  NOR2_X1 U5145 ( .A1(n5951), .A2(n5955), .ZN(n5195) );
  INV_X1 U5146 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6041) );
  INV_X1 U5147 ( .A(n6283), .ZN(n5070) );
  NOR2_X1 U5148 ( .A1(n5070), .A2(n4585), .ZN(n5379) );
  NAND2_X1 U5149 ( .A1(n4586), .A2(n5379), .ZN(n5348) );
  NOR2_X1 U5150 ( .A1(n6041), .A2(n5348), .ZN(n5336) );
  AND2_X1 U5151 ( .A1(n5336), .A2(REIP_REG_25__SCAN_IN), .ZN(n5321) );
  NAND2_X1 U5152 ( .A1(n5321), .A2(REIP_REG_26__SCAN_IN), .ZN(n5306) );
  NAND2_X1 U5153 ( .A1(n6301), .A2(n6283), .ZN(n5349) );
  OAI21_X1 U5154 ( .B1(n5306), .B2(n4587), .A(n5349), .ZN(n5295) );
  OAI21_X1 U5155 ( .B1(n5195), .B2(n6301), .A(n5295), .ZN(n5203) );
  NAND2_X1 U5156 ( .A1(n3440), .A2(n4593), .ZN(U2797) );
  OR2_X1 U5157 ( .A1(n4825), .A2(n4595), .ZN(n4596) );
  NAND2_X1 U5158 ( .A1(n4939), .A2(n4596), .ZN(n4920) );
  OAI21_X1 U5159 ( .B1(n5070), .B2(n4601), .A(n5349), .ZN(n5068) );
  OAI22_X1 U5160 ( .A1(n6389), .A2(n4920), .B1(n4853), .B2(n5068), .ZN(n4609)
         );
  INV_X1 U5161 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4921) );
  INV_X1 U5162 ( .A(n6610), .ZN(n4597) );
  NOR2_X1 U5163 ( .A1(n4598), .A2(n4597), .ZN(n4599) );
  XNOR2_X1 U5164 ( .A(n4599), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4903)
         );
  NAND2_X1 U5165 ( .A1(n6492), .A2(n4837), .ZN(n5268) );
  INV_X1 U5166 ( .A(n5268), .ZN(n4600) );
  NAND2_X1 U5167 ( .A1(n5198), .A2(n4600), .ZN(n6264) );
  OAI22_X1 U5168 ( .A1(n4921), .A2(n6382), .B1(n4903), .B2(n6264), .ZN(n4608)
         );
  INV_X1 U5169 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4603) );
  NOR2_X1 U5170 ( .A1(n5070), .A2(n6134), .ZN(n6362) );
  INV_X1 U5171 ( .A(n6362), .ZN(n6343) );
  OR3_X1 U5172 ( .A1(n6301), .A2(n4601), .A3(REIP_REG_4__SCAN_IN), .ZN(n4602)
         );
  OAI211_X1 U5173 ( .C1(n6384), .C2(n4603), .A(n6343), .B(n4602), .ZN(n4607)
         );
  OR2_X1 U5174 ( .A1(n4819), .A2(n4820), .ZN(n4822) );
  AOI21_X1 U5175 ( .B1(n4604), .B2(n4822), .A(n4952), .ZN(n4961) );
  INV_X1 U5176 ( .A(n4961), .ZN(n4922) );
  NAND2_X1 U5177 ( .A1(n5198), .A2(n4673), .ZN(n4605) );
  NAND2_X1 U5178 ( .A1(n4605), .A2(n6390), .ZN(n6271) );
  INV_X1 U5179 ( .A(n6271), .ZN(n6277) );
  OAI22_X1 U5180 ( .A1(n4922), .A2(n6277), .B1(n4959), .B2(n6395), .ZN(n4606)
         );
  OR4_X1 U5181 ( .A1(n4609), .A2(n4608), .A3(n4607), .A4(n4606), .ZN(U2823) );
  INV_X1 U5182 ( .A(n4610), .ZN(n4611) );
  INV_X1 U5183 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n6473) );
  OAI211_X1 U5184 ( .C1(n4611), .C2(n6473), .A(n4612), .B(n6134), .ZN(U2788)
         );
  INV_X1 U5185 ( .A(EAX_REG_11__SCAN_IN), .ZN(n5998) );
  INV_X1 U5186 ( .A(n4612), .ZN(n4615) );
  NOR2_X1 U5187 ( .A1(n4746), .A2(n4518), .ZN(n4847) );
  NAND2_X1 U5188 ( .A1(n4847), .A2(n6449), .ZN(n4614) );
  NAND2_X1 U5189 ( .A1(n4736), .A2(DATAI_11_), .ZN(n4699) );
  OAI21_X1 U5190 ( .B1(n6147), .B2(n6462), .A(n4615), .ZN(n4689) );
  NAND2_X1 U5191 ( .A1(n4689), .A2(LWORD_REG_11__SCAN_IN), .ZN(n4616) );
  OAI211_X1 U5192 ( .C1(n5998), .C2(n4738), .A(n4699), .B(n4616), .ZN(U2950)
         );
  NAND2_X1 U5193 ( .A1(n4736), .A2(DATAI_12_), .ZN(n4685) );
  NAND2_X1 U5194 ( .A1(n4689), .A2(LWORD_REG_12__SCAN_IN), .ZN(n4617) );
  OAI211_X1 U5195 ( .C1(n4061), .C2(n4738), .A(n4685), .B(n4617), .ZN(U2951)
         );
  INV_X1 U5196 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6003) );
  NAND2_X1 U5197 ( .A1(n4736), .A2(DATAI_14_), .ZN(n4695) );
  NAND2_X1 U5198 ( .A1(n4689), .A2(LWORD_REG_14__SCAN_IN), .ZN(n4618) );
  OAI211_X1 U5199 ( .C1(n6003), .C2(n4738), .A(n4695), .B(n4618), .ZN(U2953)
         );
  INV_X1 U5200 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6001) );
  NAND2_X1 U5201 ( .A1(n4736), .A2(DATAI_13_), .ZN(n4688) );
  NAND2_X1 U5202 ( .A1(n4689), .A2(LWORD_REG_13__SCAN_IN), .ZN(n4619) );
  OAI211_X1 U5203 ( .C1(n6001), .C2(n4738), .A(n4688), .B(n4619), .ZN(U2952)
         );
  INV_X1 U5204 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4702) );
  NAND2_X1 U5205 ( .A1(n4613), .A2(n6147), .ZN(n6430) );
  OR2_X1 U5206 ( .A1(n5264), .A2(n6691), .ZN(n4890) );
  AND2_X1 U5207 ( .A1(n6430), .A2(n4890), .ZN(n4621) );
  OR2_X1 U5208 ( .A1(n6428), .A2(n6141), .ZN(n4620) );
  OR2_X1 U5209 ( .A1(n6007), .A2(n6492), .ZN(n4817) );
  OR2_X1 U5210 ( .A1(n6657), .A2(n4622), .ZN(n6427) );
  INV_X1 U5213 ( .A(n6007), .ZN(n4623) );
  AOI22_X1 U5214 ( .A1(n6152), .A2(UWORD_REG_7__SCAN_IN), .B1(n5777), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4624) );
  OAI21_X1 U5215 ( .B1(n4702), .B2(n4817), .A(n4624), .ZN(U2900) );
  INV_X1 U5216 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4719) );
  AOI22_X1 U5217 ( .A1(n6152), .A2(UWORD_REG_5__SCAN_IN), .B1(n5777), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4625) );
  OAI21_X1 U5218 ( .B1(n4719), .B2(n4817), .A(n4625), .ZN(U2902) );
  INV_X1 U5219 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4734) );
  AOI22_X1 U5220 ( .A1(n6152), .A2(UWORD_REG_6__SCAN_IN), .B1(n5777), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4626) );
  OAI21_X1 U5221 ( .B1(n4734), .B2(n4817), .A(n4626), .ZN(U2901) );
  INV_X1 U5222 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4713) );
  AOI22_X1 U5223 ( .A1(n6152), .A2(UWORD_REG_8__SCAN_IN), .B1(n5777), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4627) );
  OAI21_X1 U5224 ( .B1(n4713), .B2(n4817), .A(n4627), .ZN(U2899) );
  AOI22_X1 U5225 ( .A1(n6152), .A2(UWORD_REG_13__SCAN_IN), .B1(n5777), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4628) );
  OAI21_X1 U5226 ( .B1(n4398), .B2(n4817), .A(n4628), .ZN(U2894) );
  INV_X1 U5227 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4686) );
  AOI22_X1 U5228 ( .A1(n6152), .A2(UWORD_REG_12__SCAN_IN), .B1(n5777), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4629) );
  OAI21_X1 U5229 ( .B1(n4686), .B2(n4817), .A(n4629), .ZN(U2895) );
  INV_X1 U5230 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4700) );
  AOI22_X1 U5231 ( .A1(n6152), .A2(UWORD_REG_11__SCAN_IN), .B1(n5777), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4630) );
  OAI21_X1 U5232 ( .B1(n4700), .B2(n4817), .A(n4630), .ZN(U2896) );
  INV_X1 U5233 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4693) );
  AOI22_X1 U5234 ( .A1(n6152), .A2(UWORD_REG_10__SCAN_IN), .B1(n5777), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4631) );
  OAI21_X1 U5235 ( .B1(n4693), .B2(n4817), .A(n4631), .ZN(U2897) );
  INV_X1 U5236 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4729) );
  AOI22_X1 U5237 ( .A1(n6152), .A2(UWORD_REG_4__SCAN_IN), .B1(n5777), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4632) );
  OAI21_X1 U5238 ( .B1(n4729), .B2(n4817), .A(n4632), .ZN(U2903) );
  INV_X1 U5239 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4716) );
  AOI22_X1 U5240 ( .A1(n6152), .A2(UWORD_REG_9__SCAN_IN), .B1(n5777), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4633) );
  OAI21_X1 U5241 ( .B1(n4716), .B2(n4817), .A(n4633), .ZN(U2898) );
  XOR2_X1 U5242 ( .A(n4635), .B(n4634), .Z(n5047) );
  INV_X1 U5243 ( .A(n5047), .ZN(n4740) );
  AOI21_X1 U5244 ( .B1(n4637), .B2(n5763), .A(n4636), .ZN(n5770) );
  INV_X1 U5245 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6075) );
  NOR2_X1 U5246 ( .A1(n6247), .A2(n6075), .ZN(n5769) );
  OAI21_X1 U5247 ( .B1(n4638), .B2(n6119), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4639) );
  INV_X1 U5248 ( .A(n4639), .ZN(n4640) );
  AOI211_X1 U5249 ( .C1(n6121), .C2(n5770), .A(n5769), .B(n4640), .ZN(n4641)
         );
  OAI21_X1 U5250 ( .B1(n4740), .B2(n6862), .A(n4641), .ZN(U2986) );
  OAI21_X1 U5251 ( .B1(n4643), .B2(n4642), .A(n4784), .ZN(n6087) );
  NOR2_X1 U5252 ( .A1(n5268), .A2(n4839), .ZN(n4758) );
  OAI21_X1 U5253 ( .B1(n4758), .B2(n3432), .A(n4644), .ZN(n4648) );
  NAND2_X1 U5254 ( .A1(n4646), .A2(n4645), .ZN(n4647) );
  OAI211_X1 U5255 ( .C1(n6732), .C2(n4649), .A(n4648), .B(n4647), .ZN(n4653)
         );
  NAND3_X1 U5256 ( .A1(n4650), .A2(n4831), .A3(n4681), .ZN(n4652) );
  OR2_X1 U5257 ( .A1(n4681), .A2(n3659), .ZN(n4651) );
  NAND2_X1 U5258 ( .A1(n4652), .A2(n4651), .ZN(n4767) );
  NOR2_X1 U5259 ( .A1(n4653), .A2(n4767), .ZN(n4655) );
  NAND2_X1 U5260 ( .A1(n4655), .A2(n4654), .ZN(n4743) );
  NOR2_X1 U5261 ( .A1(n4656), .A2(n4831), .ZN(n4657) );
  NAND2_X1 U5262 ( .A1(n4776), .A2(n4657), .ZN(n4891) );
  INV_X1 U5263 ( .A(n4658), .ZN(n4659) );
  NAND2_X1 U5264 ( .A1(n4660), .A2(n4659), .ZN(n4661) );
  OAI211_X1 U5265 ( .C1(n4744), .C2(n4662), .A(n4891), .B(n4661), .ZN(n4663)
         );
  NOR2_X1 U5266 ( .A1(n4743), .A2(n4663), .ZN(n4850) );
  NOR2_X1 U5267 ( .A1(n4665), .A2(n4664), .ZN(n4834) );
  AND2_X1 U5268 ( .A1(n4850), .A2(n4834), .ZN(n4852) );
  NAND2_X1 U5269 ( .A1(n5262), .A2(n4852), .ZN(n4760) );
  INV_X1 U5270 ( .A(n5494), .ZN(n6965) );
  NAND3_X1 U5271 ( .A1(n6965), .A2(n6822), .A3(n3941), .ZN(n4677) );
  INV_X1 U5272 ( .A(n4677), .ZN(n4666) );
  NAND4_X1 U5273 ( .A1(n4666), .A2(n3529), .A3(n6780), .A4(n4670), .ZN(n4667)
         );
  NAND2_X1 U5274 ( .A1(n4760), .A2(n4667), .ZN(n4668) );
  OAI21_X1 U5275 ( .B1(n4671), .B2(n4670), .A(n4669), .ZN(n4884) );
  INV_X1 U5276 ( .A(n4884), .ZN(n4672) );
  OAI222_X1 U5277 ( .A1(n6087), .A2(n5489), .B1(n6086), .B2(n4445), .C1(n5479), 
        .C2(n4672), .ZN(U2858) );
  NAND2_X1 U5278 ( .A1(n4769), .A2(n4673), .ZN(n4845) );
  OR2_X1 U5279 ( .A1(n5262), .A2(n4845), .ZN(n4676) );
  INV_X1 U5280 ( .A(n4901), .ZN(n4674) );
  NAND3_X1 U5281 ( .A1(n4674), .A2(n6462), .A3(n5259), .ZN(n4675) );
  NAND2_X1 U5282 ( .A1(n4676), .A2(n4675), .ZN(n4762) );
  NOR2_X1 U5283 ( .A1(n4744), .A2(n4677), .ZN(n4678) );
  OAI21_X1 U5284 ( .B1(n4762), .B2(n4678), .A(n6449), .ZN(n4680) );
  NAND2_X1 U5285 ( .A1(n4681), .A2(n5494), .ZN(n4682) );
  NAND2_X2 U5286 ( .A1(n5520), .A2(n4682), .ZN(n6475) );
  INV_X1 U5287 ( .A(n4682), .ZN(n4683) );
  NAND2_X1 U5288 ( .A1(n5520), .A2(n4683), .ZN(n5521) );
  INV_X1 U5289 ( .A(DATAI_0_), .ZN(n6488) );
  INV_X1 U5290 ( .A(EAX_REG_0__SCAN_IN), .ZN(n5977) );
  OAI222_X1 U5291 ( .A1(n6475), .A2(n4740), .B1(n5521), .B2(n6488), .C1(n5520), 
        .C2(n5977), .ZN(U2891) );
  INV_X1 U5292 ( .A(DATAI_1_), .ZN(n6690) );
  INV_X1 U5293 ( .A(EAX_REG_1__SCAN_IN), .ZN(n5979) );
  OAI222_X1 U5294 ( .A1(n6087), .A2(n6475), .B1(n5521), .B2(n6690), .C1(n5520), 
        .C2(n5979), .ZN(U2890) );
  NAND2_X1 U5295 ( .A1(n4689), .A2(UWORD_REG_12__SCAN_IN), .ZN(n4684) );
  OAI211_X1 U5296 ( .C1(n4686), .C2(n4738), .A(n4685), .B(n4684), .ZN(U2936)
         );
  NAND2_X1 U5297 ( .A1(n4689), .A2(UWORD_REG_13__SCAN_IN), .ZN(n4687) );
  OAI211_X1 U5298 ( .C1(n4398), .C2(n4738), .A(n4688), .B(n4687), .ZN(U2937)
         );
  INV_X1 U5299 ( .A(EAX_REG_4__SCAN_IN), .ZN(n5985) );
  NAND2_X1 U5300 ( .A1(n4736), .A2(DATAI_4_), .ZN(n4728) );
  NAND2_X1 U5301 ( .A1(n4735), .A2(LWORD_REG_4__SCAN_IN), .ZN(n4690) );
  OAI211_X1 U5302 ( .C1(n4738), .C2(n5985), .A(n4728), .B(n4690), .ZN(U2943)
         );
  INV_X1 U5303 ( .A(EAX_REG_3__SCAN_IN), .ZN(n5983) );
  NAND2_X1 U5304 ( .A1(n4736), .A2(DATAI_3_), .ZN(n4726) );
  NAND2_X1 U5305 ( .A1(n4735), .A2(LWORD_REG_3__SCAN_IN), .ZN(n4691) );
  OAI211_X1 U5306 ( .C1(n5983), .C2(n4738), .A(n4726), .B(n4691), .ZN(U2942)
         );
  NAND2_X1 U5307 ( .A1(n4736), .A2(DATAI_10_), .ZN(n4704) );
  NAND2_X1 U5308 ( .A1(n4735), .A2(UWORD_REG_10__SCAN_IN), .ZN(n4692) );
  OAI211_X1 U5309 ( .C1(n4693), .C2(n4738), .A(n4704), .B(n4692), .ZN(U2934)
         );
  INV_X1 U5310 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4810) );
  NAND2_X1 U5311 ( .A1(n4735), .A2(UWORD_REG_14__SCAN_IN), .ZN(n4694) );
  OAI211_X1 U5312 ( .C1(n4810), .C2(n4738), .A(n4695), .B(n4694), .ZN(U2938)
         );
  NAND2_X1 U5313 ( .A1(n4736), .A2(DATAI_1_), .ZN(n4722) );
  NAND2_X1 U5314 ( .A1(n4735), .A2(LWORD_REG_1__SCAN_IN), .ZN(n4696) );
  OAI211_X1 U5315 ( .C1(n5979), .C2(n4738), .A(n4722), .B(n4696), .ZN(U2940)
         );
  INV_X1 U5316 ( .A(EAX_REG_5__SCAN_IN), .ZN(n5987) );
  NAND2_X1 U5317 ( .A1(n4736), .A2(DATAI_5_), .ZN(n4718) );
  NAND2_X1 U5318 ( .A1(n4735), .A2(LWORD_REG_5__SCAN_IN), .ZN(n4697) );
  OAI211_X1 U5319 ( .C1(n5987), .C2(n4738), .A(n4718), .B(n4697), .ZN(U2944)
         );
  NAND2_X1 U5320 ( .A1(n4735), .A2(UWORD_REG_11__SCAN_IN), .ZN(n4698) );
  OAI211_X1 U5321 ( .C1(n4700), .C2(n4738), .A(n4699), .B(n4698), .ZN(U2935)
         );
  NAND2_X1 U5322 ( .A1(n4736), .A2(DATAI_7_), .ZN(n4708) );
  NAND2_X1 U5323 ( .A1(n4735), .A2(UWORD_REG_7__SCAN_IN), .ZN(n4701) );
  OAI211_X1 U5324 ( .C1(n4702), .C2(n4738), .A(n4708), .B(n4701), .ZN(U2931)
         );
  INV_X1 U5325 ( .A(EAX_REG_10__SCAN_IN), .ZN(n5996) );
  NAND2_X1 U5326 ( .A1(n4735), .A2(LWORD_REG_10__SCAN_IN), .ZN(n4703) );
  OAI211_X1 U5327 ( .C1(n5996), .C2(n4738), .A(n4704), .B(n4703), .ZN(U2949)
         );
  INV_X1 U5328 ( .A(EAX_REG_9__SCAN_IN), .ZN(n5994) );
  NAND2_X1 U5329 ( .A1(n4736), .A2(DATAI_9_), .ZN(n4715) );
  NAND2_X1 U5330 ( .A1(n4735), .A2(LWORD_REG_9__SCAN_IN), .ZN(n4705) );
  OAI211_X1 U5331 ( .C1(n5994), .C2(n4738), .A(n4715), .B(n4705), .ZN(U2948)
         );
  INV_X1 U5332 ( .A(EAX_REG_8__SCAN_IN), .ZN(n5992) );
  NAND2_X1 U5333 ( .A1(n4736), .A2(DATAI_8_), .ZN(n4712) );
  NAND2_X1 U5334 ( .A1(n4735), .A2(LWORD_REG_8__SCAN_IN), .ZN(n4706) );
  OAI211_X1 U5335 ( .C1(n5992), .C2(n4738), .A(n4712), .B(n4706), .ZN(U2947)
         );
  NAND2_X1 U5336 ( .A1(n4735), .A2(LWORD_REG_7__SCAN_IN), .ZN(n4707) );
  OAI211_X1 U5337 ( .C1(n3997), .C2(n4738), .A(n4708), .B(n4707), .ZN(U2946)
         );
  INV_X1 U5338 ( .A(EAX_REG_6__SCAN_IN), .ZN(n5989) );
  NAND2_X1 U5339 ( .A1(n4736), .A2(DATAI_6_), .ZN(n4733) );
  NAND2_X1 U5340 ( .A1(n4735), .A2(LWORD_REG_6__SCAN_IN), .ZN(n4709) );
  OAI211_X1 U5341 ( .C1(n4738), .C2(n5989), .A(n4733), .B(n4709), .ZN(U2945)
         );
  NAND2_X1 U5342 ( .A1(n4736), .A2(DATAI_0_), .ZN(n4731) );
  NAND2_X1 U5343 ( .A1(n4735), .A2(LWORD_REG_0__SCAN_IN), .ZN(n4710) );
  OAI211_X1 U5344 ( .C1(n5977), .C2(n4738), .A(n4731), .B(n4710), .ZN(U2939)
         );
  NAND2_X1 U5345 ( .A1(n4735), .A2(UWORD_REG_8__SCAN_IN), .ZN(n4711) );
  OAI211_X1 U5346 ( .C1(n4713), .C2(n4738), .A(n4712), .B(n4711), .ZN(U2932)
         );
  NAND2_X1 U5347 ( .A1(n4735), .A2(UWORD_REG_9__SCAN_IN), .ZN(n4714) );
  OAI211_X1 U5348 ( .C1(n4716), .C2(n4738), .A(n4715), .B(n4714), .ZN(U2933)
         );
  NAND2_X1 U5349 ( .A1(n4735), .A2(UWORD_REG_5__SCAN_IN), .ZN(n4717) );
  OAI211_X1 U5350 ( .C1(n4719), .C2(n4738), .A(n4718), .B(n4717), .ZN(U2929)
         );
  INV_X1 U5351 ( .A(EAX_REG_2__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U5352 ( .A1(n4736), .A2(DATAI_2_), .ZN(n4724) );
  NAND2_X1 U5353 ( .A1(n4735), .A2(LWORD_REG_2__SCAN_IN), .ZN(n4720) );
  OAI211_X1 U5354 ( .C1(n5981), .C2(n4738), .A(n4724), .B(n4720), .ZN(U2941)
         );
  INV_X1 U5355 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4813) );
  NAND2_X1 U5356 ( .A1(n4735), .A2(UWORD_REG_1__SCAN_IN), .ZN(n4721) );
  OAI211_X1 U5357 ( .C1(n4813), .C2(n4738), .A(n4722), .B(n4721), .ZN(U2925)
         );
  INV_X1 U5358 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4815) );
  NAND2_X1 U5359 ( .A1(n4735), .A2(UWORD_REG_2__SCAN_IN), .ZN(n4723) );
  OAI211_X1 U5360 ( .C1(n4815), .C2(n4738), .A(n4724), .B(n4723), .ZN(U2926)
         );
  INV_X1 U5361 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4818) );
  NAND2_X1 U5362 ( .A1(n4735), .A2(UWORD_REG_3__SCAN_IN), .ZN(n4725) );
  OAI211_X1 U5363 ( .C1(n4818), .C2(n4738), .A(n4726), .B(n4725), .ZN(U2927)
         );
  NAND2_X1 U5364 ( .A1(n4735), .A2(UWORD_REG_4__SCAN_IN), .ZN(n4727) );
  OAI211_X1 U5365 ( .C1(n4738), .C2(n4729), .A(n4728), .B(n4727), .ZN(U2928)
         );
  NAND2_X1 U5366 ( .A1(n4735), .A2(UWORD_REG_0__SCAN_IN), .ZN(n4730) );
  OAI211_X1 U5367 ( .C1(n4240), .C2(n4738), .A(n4731), .B(n4730), .ZN(U2924)
         );
  NAND2_X1 U5368 ( .A1(n4735), .A2(UWORD_REG_6__SCAN_IN), .ZN(n4732) );
  OAI211_X1 U5369 ( .C1(n4734), .C2(n4738), .A(n4733), .B(n4732), .ZN(U2930)
         );
  INV_X1 U5370 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6008) );
  AOI22_X1 U5371 ( .A1(n4736), .A2(DATAI_15_), .B1(n4735), .B2(
        LWORD_REG_15__SCAN_IN), .ZN(n4737) );
  OAI21_X1 U5372 ( .B1(n6008), .B2(n4738), .A(n4737), .ZN(U2954) );
  OAI21_X1 U5373 ( .B1(n3432), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4739), 
        .ZN(n5767) );
  OAI222_X1 U5374 ( .A1(n5479), .A2(n5767), .B1(n4452), .B2(n6086), .C1(n5489), 
        .C2(n4740), .ZN(U2859) );
  INV_X1 U5375 ( .A(n4743), .ZN(n4748) );
  AND4_X1 U5376 ( .A1(n4901), .A2(n4746), .A3(n4745), .A4(n4744), .ZN(n4747)
         );
  NAND2_X1 U5377 ( .A1(n4748), .A2(n4747), .ZN(n4888) );
  INV_X1 U5378 ( .A(n4888), .ZN(n4804) );
  INV_X1 U5379 ( .A(n4890), .ZN(n6407) );
  INV_X1 U5380 ( .A(n4749), .ZN(n4752) );
  INV_X1 U5381 ( .A(n4750), .ZN(n4751) );
  NAND2_X1 U5382 ( .A1(n4752), .A2(n4751), .ZN(n4755) );
  AOI22_X1 U5383 ( .A1(n6407), .A2(n4753), .B1(n4776), .B2(n4755), .ZN(n4754)
         );
  OAI21_X1 U5384 ( .B1(n4742), .B2(n4804), .A(n4754), .ZN(n6408) );
  INV_X1 U5385 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5229) );
  AOI22_X1 U5386 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5229), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n3669), .ZN(n5246) );
  NOR2_X1 U5387 ( .A1(n6440), .A2(n5763), .ZN(n4779) );
  INV_X1 U5388 ( .A(n5248), .ZN(n6444) );
  AOI222_X1 U5389 ( .A1(n6408), .A2(n6434), .B1(n5246), .B2(n4779), .C1(n4755), 
        .C2(n6444), .ZN(n4775) );
  NOR2_X1 U5390 ( .A1(n4890), .A2(n6141), .ZN(n4756) );
  NOR2_X1 U5391 ( .A1(n4847), .A2(n4756), .ZN(n4757) );
  NOR2_X1 U5392 ( .A1(n4766), .A2(n4757), .ZN(n4763) );
  INV_X1 U5393 ( .A(n4758), .ZN(n4759) );
  NAND2_X1 U5394 ( .A1(n4760), .A2(n4759), .ZN(n4761) );
  NOR3_X1 U5395 ( .A1(n4763), .A2(n4762), .A3(n4761), .ZN(n4773) );
  NAND2_X1 U5396 ( .A1(n4613), .A2(n4764), .ZN(n4765) );
  INV_X1 U5397 ( .A(n4767), .ZN(n4768) );
  NAND2_X1 U5398 ( .A1(n4769), .A2(n4768), .ZN(n4770) );
  NAND2_X1 U5399 ( .A1(n4770), .A2(n5264), .ZN(n4771) );
  NOR2_X1 U5400 ( .A1(n6657), .A2(n6440), .ZN(n6438) );
  NAND2_X1 U5401 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6438), .ZN(n6441) );
  INV_X1 U5402 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6398) );
  OAI22_X1 U5403 ( .A1(n6410), .A2(n6428), .B1(n6441), .B2(n6398), .ZN(n6402)
         );
  AOI21_X1 U5404 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6491), .A(n6402), .ZN(
        n5253) );
  NAND2_X1 U5405 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n5253), .ZN(n4774) );
  OAI21_X1 U5406 ( .B1(n4775), .B2(n5253), .A(n4774), .ZN(U3460) );
  INV_X1 U5407 ( .A(n6529), .ZN(n6573) );
  INV_X1 U5408 ( .A(n4776), .ZN(n4777) );
  OAI22_X1 U5409 ( .A1(n6573), .A2(n4804), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n4777), .ZN(n6406) );
  INV_X1 U5410 ( .A(n6406), .ZN(n4778) );
  OAI21_X1 U5411 ( .B1(n4778), .B2(STATE2_REG_3__SCAN_IN), .A(n6440), .ZN(
        n4780) );
  INV_X1 U5412 ( .A(n4779), .ZN(n5245) );
  AOI22_X1 U5413 ( .A1(n4780), .A2(n5245), .B1(n6444), .B2(n4781), .ZN(n4783)
         );
  AOI21_X1 U5414 ( .B1(n6407), .B2(n6434), .A(n5253), .ZN(n4782) );
  OAI22_X1 U5415 ( .A1(n4783), .A2(n5253), .B1(n4782), .B2(n4781), .ZN(U3461)
         );
  NAND3_X1 U5416 ( .A1(n4786), .A2(n4785), .A3(n4784), .ZN(n4787) );
  AND2_X1 U5417 ( .A1(n4819), .A2(n4787), .ZN(n6272) );
  INV_X1 U5418 ( .A(n6272), .ZN(n4788) );
  INV_X1 U5419 ( .A(DATAI_2_), .ZN(n6731) );
  OAI222_X1 U5420 ( .A1(n4788), .A2(n6475), .B1(n5521), .B2(n6731), .C1(n5520), 
        .C2(n5981), .ZN(U2889) );
  INV_X1 U5421 ( .A(n6574), .ZN(n6638) );
  INV_X1 U5422 ( .A(n4891), .ZN(n4796) );
  INV_X1 U5423 ( .A(n4791), .ZN(n4792) );
  OAI211_X1 U5424 ( .C1(n4790), .C2(n4807), .A(n4793), .B(n4792), .ZN(n4805)
         );
  NAND2_X1 U5425 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4794) );
  XNOR2_X1 U5426 ( .A(n4794), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4795)
         );
  AOI22_X1 U5427 ( .A1(n4796), .A2(n4805), .B1(n6407), .B2(n4795), .ZN(n4803)
         );
  INV_X1 U5428 ( .A(n4845), .ZN(n4797) );
  OR2_X1 U5429 ( .A1(n4852), .A2(n4797), .ZN(n4894) );
  INV_X1 U5430 ( .A(n4798), .ZN(n4904) );
  INV_X1 U5431 ( .A(n4799), .ZN(n4800) );
  MUX2_X1 U5432 ( .A(n4800), .B(n4807), .S(n4790), .Z(n4801) );
  NAND3_X1 U5433 ( .A1(n4894), .A2(n4904), .A3(n4801), .ZN(n4802) );
  OAI211_X1 U5434 ( .C1(n6638), .C2(n4804), .A(n4803), .B(n4802), .ZN(n4900)
         );
  AOI22_X1 U5435 ( .A1(n4900), .A2(n6434), .B1(n6444), .B2(n4805), .ZN(n4806)
         );
  INV_X1 U5436 ( .A(n5253), .ZN(n6405) );
  MUX2_X1 U5437 ( .A(n4807), .B(n4806), .S(n6405), .Z(n4808) );
  INV_X1 U5438 ( .A(n4808), .ZN(U3456) );
  AOI22_X1 U5439 ( .A1(n6152), .A2(UWORD_REG_14__SCAN_IN), .B1(n6004), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4809) );
  OAI21_X1 U5440 ( .B1(n4810), .B2(n4817), .A(n4809), .ZN(U2893) );
  AOI22_X1 U5441 ( .A1(n6152), .A2(UWORD_REG_0__SCAN_IN), .B1(n6004), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4811) );
  OAI21_X1 U5442 ( .B1(n4240), .B2(n4817), .A(n4811), .ZN(U2907) );
  AOI22_X1 U5443 ( .A1(n6152), .A2(UWORD_REG_1__SCAN_IN), .B1(n6004), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4812) );
  OAI21_X1 U5444 ( .B1(n4813), .B2(n4817), .A(n4812), .ZN(U2906) );
  AOI22_X1 U5445 ( .A1(n6152), .A2(UWORD_REG_2__SCAN_IN), .B1(n6004), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4814) );
  OAI21_X1 U5446 ( .B1(n4815), .B2(n4817), .A(n4814), .ZN(U2905) );
  AOI22_X1 U5447 ( .A1(n6152), .A2(UWORD_REG_3__SCAN_IN), .B1(n6004), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4816) );
  OAI21_X1 U5448 ( .B1(n4818), .B2(n4817), .A(n4816), .ZN(U2904) );
  NAND2_X1 U5449 ( .A1(n4820), .A2(n4819), .ZN(n4821) );
  AND2_X1 U5450 ( .A1(n4822), .A2(n4821), .ZN(n5073) );
  INV_X1 U5451 ( .A(n5073), .ZN(n4828) );
  INV_X1 U5452 ( .A(DATAI_3_), .ZN(n6779) );
  OAI222_X1 U5453 ( .A1(n4828), .A2(n6475), .B1(n5521), .B2(n6779), .C1(n5520), 
        .C2(n5983), .ZN(U2888) );
  INV_X1 U5454 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4827) );
  INV_X1 U5455 ( .A(n6078), .ZN(n4824) );
  AOI21_X1 U5456 ( .B1(n4824), .B2(n6077), .A(n4823), .ZN(n4826) );
  OR2_X1 U5457 ( .A1(n4826), .A2(n4825), .ZN(n5067) );
  OAI222_X1 U5458 ( .A1(n4828), .A2(n5489), .B1(n4827), .B2(n6086), .C1(n5067), 
        .C2(n5479), .ZN(U2856) );
  XNOR2_X1 U5459 ( .A(n4830), .B(n4829), .ZN(n4963) );
  AND2_X1 U5460 ( .A1(n4837), .A2(n6462), .ZN(n4833) );
  AOI21_X1 U5461 ( .B1(n5491), .B2(n4831), .A(n4839), .ZN(n4832) );
  AOI21_X1 U5462 ( .B1(n4613), .B2(n4833), .A(n4832), .ZN(n4836) );
  INV_X1 U5463 ( .A(n4834), .ZN(n4835) );
  MUX2_X1 U5464 ( .A(n4836), .B(n4835), .S(n5262), .Z(n4841) );
  NAND2_X1 U5465 ( .A1(n4837), .A2(n6141), .ZN(n4838) );
  NAND4_X1 U5466 ( .A1(n5259), .A2(n6462), .A3(n4839), .A4(n4838), .ZN(n4840)
         );
  NAND3_X1 U5467 ( .A1(n4842), .A2(n4841), .A3(n4840), .ZN(n4843) );
  NAND2_X1 U5468 ( .A1(n4845), .A2(n4844), .ZN(n5256) );
  OAI21_X1 U5469 ( .B1(n4854), .B2(n6822), .A(n4901), .ZN(n4846) );
  OR2_X1 U5470 ( .A1(n4847), .A2(n4846), .ZN(n4848) );
  NOR2_X1 U5471 ( .A1(n5256), .A2(n4848), .ZN(n4849) );
  OR2_X1 U5472 ( .A1(n4858), .A2(n4850), .ZN(n5090) );
  NAND2_X1 U5473 ( .A1(n5090), .A2(n5765), .ZN(n5086) );
  NAND2_X1 U5474 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4861) );
  NAND2_X1 U5475 ( .A1(n6247), .A2(n4858), .ZN(n5764) );
  INV_X1 U5476 ( .A(n5090), .ZN(n4881) );
  NAND2_X1 U5477 ( .A1(n4881), .A2(n5763), .ZN(n4851) );
  NAND2_X1 U5478 ( .A1(n5764), .A2(n4851), .ZN(n5085) );
  AOI21_X1 U5479 ( .B1(n5086), .B2(n4861), .A(n5085), .ZN(n6178) );
  INV_X1 U5480 ( .A(n4852), .ZN(n5258) );
  AOI21_X1 U5481 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n4944) );
  NAND2_X1 U5482 ( .A1(n5089), .A2(n4944), .ZN(n6185) );
  NAND2_X1 U5483 ( .A1(n6178), .A2(n6185), .ZN(n4983) );
  NOR2_X1 U5484 ( .A1(n6247), .A2(n4853), .ZN(n4957) );
  INV_X1 U5485 ( .A(n4854), .ZN(n4855) );
  NAND2_X1 U5486 ( .A1(n4855), .A2(n6822), .ZN(n4856) );
  AND2_X1 U5487 ( .A1(n6430), .A2(n4856), .ZN(n4857) );
  NOR2_X1 U5488 ( .A1(n6224), .A2(n4920), .ZN(n4859) );
  AOI211_X1 U5489 ( .C1(n4983), .C2(INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4957), 
        .B(n4859), .ZN(n4863) );
  AND2_X1 U5490 ( .A1(n5765), .A2(n5763), .ZN(n4878) );
  INV_X1 U5491 ( .A(n4878), .ZN(n4860) );
  NAND2_X1 U5492 ( .A1(n4860), .A2(n5086), .ZN(n6183) );
  NOR2_X1 U5493 ( .A1(n6183), .A2(n4861), .ZN(n4941) );
  INV_X1 U5494 ( .A(n4944), .ZN(n5088) );
  OAI21_X1 U5495 ( .B1(n5089), .B2(n4941), .A(n5088), .ZN(n4993) );
  INV_X1 U5496 ( .A(n4993), .ZN(n4869) );
  NAND2_X1 U5497 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4943) );
  OAI211_X1 U5498 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A(n4869), .B(n4943), .ZN(n4862) );
  OAI211_X1 U5499 ( .C1(n4963), .C2(n6225), .A(n4863), .B(n4862), .ZN(U3014)
         );
  NAND2_X1 U5500 ( .A1(n4865), .A2(n4864), .ZN(n4867) );
  XNOR2_X1 U5501 ( .A(n4867), .B(n4866), .ZN(n4968) );
  INV_X1 U5502 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4868) );
  AOI22_X1 U5503 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n4983), .B1(n4869), 
        .B2(n4868), .ZN(n4872) );
  INV_X1 U5504 ( .A(REIP_REG_3__SCAN_IN), .ZN(n4870) );
  NOR2_X1 U5505 ( .A1(n6247), .A2(n4870), .ZN(n4964) );
  INV_X1 U5506 ( .A(n4964), .ZN(n4871) );
  OAI211_X1 U5507 ( .C1(n6224), .C2(n5067), .A(n4872), .B(n4871), .ZN(n4873)
         );
  INV_X1 U5508 ( .A(n4873), .ZN(n4874) );
  OAI21_X1 U5509 ( .B1(n4968), .B2(n6225), .A(n4874), .ZN(U3015) );
  XNOR2_X1 U5510 ( .A(n4875), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4876)
         );
  XNOR2_X1 U5511 ( .A(n4877), .B(n4876), .ZN(n6088) );
  INV_X1 U5512 ( .A(n6247), .ZN(n6235) );
  INV_X1 U5513 ( .A(n5086), .ZN(n4947) );
  NAND2_X1 U5514 ( .A1(n4947), .A2(n6179), .ZN(n6214) );
  INV_X1 U5515 ( .A(n6214), .ZN(n6194) );
  NOR3_X1 U5516 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4878), .A3(n6194), 
        .ZN(n4879) );
  AOI21_X1 U5517 ( .B1(n6235), .B2(REIP_REG_1__SCAN_IN), .A(n4879), .ZN(n4880)
         );
  INV_X1 U5518 ( .A(n4880), .ZN(n4883) );
  OAI21_X1 U5519 ( .B1(n5089), .B2(n4881), .A(n5763), .ZN(n5771) );
  AOI21_X1 U5520 ( .B1(n5771), .B2(n5764), .A(n3669), .ZN(n4882) );
  AOI211_X1 U5521 ( .C1(n6243), .C2(n4884), .A(n4883), .B(n4882), .ZN(n4885)
         );
  OAI21_X1 U5522 ( .B1(n6088), .B2(n6225), .A(n4885), .ZN(U3017) );
  NAND2_X1 U5523 ( .A1(n6518), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4923) );
  XNOR2_X1 U5524 ( .A(n6537), .B(n4923), .ZN(n4916) );
  INV_X1 U5525 ( .A(n6410), .ZN(n4897) );
  NAND2_X1 U5526 ( .A1(n4887), .A2(n4888), .ZN(n4896) );
  XNOR2_X1 U5527 ( .A(n4790), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4893)
         );
  XNOR2_X1 U5528 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4889) );
  OAI22_X1 U5529 ( .A1(n4891), .A2(n4893), .B1(n4890), .B2(n4889), .ZN(n4892)
         );
  AOI21_X1 U5530 ( .B1(n4894), .B2(n4893), .A(n4892), .ZN(n4895) );
  NAND2_X1 U5531 ( .A1(n4896), .A2(n4895), .ZN(n5250) );
  NAND2_X1 U5532 ( .A1(n4897), .A2(n5250), .ZN(n4899) );
  NAND2_X1 U5533 ( .A1(n6410), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4898) );
  AND2_X1 U5534 ( .A1(n4899), .A2(n4898), .ZN(n6415) );
  MUX2_X1 U5535 ( .A(n4900), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6410), 
        .Z(n6417) );
  NAND2_X1 U5536 ( .A1(n6440), .A2(n6417), .ZN(n4909) );
  NAND2_X1 U5537 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6398), .ZN(n4905) );
  OR2_X1 U5538 ( .A1(n4901), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4902) );
  OR2_X1 U5539 ( .A1(n4903), .A2(n4902), .ZN(n6400) );
  OAI21_X1 U5540 ( .B1(n4905), .B2(n4904), .A(n6400), .ZN(n4906) );
  INV_X1 U5541 ( .A(n4906), .ZN(n4908) );
  MUX2_X1 U5542 ( .A(n6410), .B(n6398), .S(STATE2_REG_1__SCAN_IN), .Z(n4907)
         );
  NAND2_X1 U5543 ( .A1(n4907), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4910) );
  OAI211_X1 U5544 ( .C1(n6415), .C2(n4909), .A(n4908), .B(n4910), .ZN(n6424)
         );
  NAND2_X1 U5545 ( .A1(n3451), .A2(n4910), .ZN(n4911) );
  NAND2_X1 U5546 ( .A1(n6424), .A2(n4911), .ZN(n4928) );
  NAND2_X1 U5547 ( .A1(n4928), .A2(n6398), .ZN(n4913) );
  INV_X1 U5548 ( .A(n6441), .ZN(n4912) );
  NAND2_X1 U5549 ( .A1(n4913), .A2(n4912), .ZN(n4914) );
  INV_X1 U5550 ( .A(n6963), .ZN(n6541) );
  NAND2_X1 U5551 ( .A1(n4914), .A2(n6963), .ZN(n4924) );
  NAND2_X1 U5552 ( .A1(n4924), .A2(n6655), .ZN(n4932) );
  INV_X1 U5553 ( .A(n4887), .ZN(n4915) );
  OAI21_X1 U5554 ( .B1(n6440), .B2(STATE2_REG_3__SCAN_IN), .A(n4924), .ZN(
        n4929) );
  OAI222_X1 U5555 ( .A1(n4916), .A2(n4932), .B1(n4915), .B2(n4929), .C1(n6619), 
        .C2(n4924), .ZN(U3463) );
  INV_X1 U5556 ( .A(n4923), .ZN(n4917) );
  NAND2_X1 U5557 ( .A1(n4917), .A2(n6585), .ZN(n4918) );
  NOR2_X1 U5558 ( .A1(n4918), .A2(n6560), .ZN(n6576) );
  AOI21_X1 U5559 ( .B1(n6632), .B2(n4918), .A(n6576), .ZN(n4919) );
  OAI222_X1 U5560 ( .A1(n4924), .A2(n6499), .B1(n4932), .B2(n4919), .C1(n4929), 
        .C2(n6638), .ZN(U3462) );
  INV_X1 U5561 ( .A(DATAI_4_), .ZN(n6821) );
  OAI222_X1 U5562 ( .A1(n4922), .A2(n6475), .B1(n5521), .B2(n6821), .C1(n5985), 
        .C2(n5520), .ZN(U2887) );
  OAI222_X1 U5563 ( .A1(n4922), .A2(n5489), .B1(n6086), .B2(n4921), .C1(n4920), 
        .C2(n5479), .ZN(U2855) );
  OAI21_X1 U5564 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n6518), .A(n4923), .ZN(
        n4927) );
  INV_X1 U5565 ( .A(n4924), .ZN(n5776) );
  INV_X1 U5566 ( .A(n4742), .ZN(n6551) );
  INV_X1 U5567 ( .A(n4929), .ZN(n4925) );
  AOI22_X1 U5568 ( .A1(n5776), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n6551), .B2(n4925), .ZN(n4926) );
  OAI21_X1 U5569 ( .B1(n4932), .B2(n4927), .A(n4926), .ZN(U3464) );
  NAND2_X1 U5570 ( .A1(n4928), .A2(n6438), .ZN(n6452) );
  OAI22_X1 U5571 ( .A1(n5776), .A2(n6452), .B1(n4929), .B2(n6573), .ZN(n4930)
         );
  AOI21_X1 U5572 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n5776), .A(n4930), 
        .ZN(n4931) );
  OAI21_X1 U5573 ( .B1(n6645), .B2(n4932), .A(n4931), .ZN(U3465) );
  NAND2_X1 U5574 ( .A1(n4935), .A2(n4934), .ZN(n4936) );
  XNOR2_X1 U5575 ( .A(n4937), .B(n4936), .ZN(n4973) );
  NAND2_X1 U5576 ( .A1(n4939), .A2(n4938), .ZN(n4940) );
  AND2_X1 U5577 ( .A1(n4976), .A2(n4940), .ZN(n6280) );
  INV_X1 U5578 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6013) );
  NOR2_X1 U5579 ( .A1(n6247), .A2(n6013), .ZN(n4942) );
  INV_X1 U5580 ( .A(n4943), .ZN(n4946) );
  AND3_X1 U5581 ( .A1(n4946), .A2(n4941), .A3(n3800), .ZN(n4996) );
  AOI211_X1 U5582 ( .C1(n6243), .C2(n6280), .A(n4942), .B(n4996), .ZN(n4950)
         );
  NOR3_X1 U5583 ( .A1(n4944), .A2(n4943), .A3(n6179), .ZN(n4948) );
  NAND2_X1 U5584 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n4946), .ZN(n4994)
         );
  AOI21_X1 U5585 ( .B1(n5089), .B2(n4994), .A(n4983), .ZN(n4945) );
  OAI21_X1 U5586 ( .B1(n4947), .B2(n4946), .A(n4945), .ZN(n4995) );
  OAI21_X1 U5587 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n4948), .A(n4995), 
        .ZN(n4949) );
  OAI211_X1 U5588 ( .C1(n6225), .C2(n4973), .A(n4950), .B(n4949), .ZN(U3013)
         );
  INV_X1 U5589 ( .A(n4951), .ZN(n4955) );
  INV_X1 U5590 ( .A(n4952), .ZN(n4954) );
  AOI21_X1 U5591 ( .B1(n4955), .B2(n4954), .A(n4953), .ZN(n4971) );
  INV_X1 U5592 ( .A(n4971), .ZN(n6278) );
  INV_X1 U5593 ( .A(n6086), .ZN(n5487) );
  AOI22_X1 U5594 ( .A1(n6082), .A2(n6280), .B1(EBX_REG_5__SCAN_IN), .B2(n5487), 
        .ZN(n4956) );
  OAI21_X1 U5595 ( .B1(n6278), .B2(n5489), .A(n4956), .ZN(U2854) );
  AOI21_X1 U5596 ( .B1(n6119), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n4957), 
        .ZN(n4958) );
  OAI21_X1 U5597 ( .B1(n6125), .B2(n4959), .A(n4958), .ZN(n4960) );
  AOI21_X1 U5598 ( .B1(n4961), .B2(n6969), .A(n4960), .ZN(n4962) );
  OAI21_X1 U5599 ( .B1(n4963), .B2(n6397), .A(n4962), .ZN(U2982) );
  AOI21_X1 U5600 ( .B1(n6119), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n4964), 
        .ZN(n4965) );
  OAI21_X1 U5601 ( .B1(n6125), .B2(n5062), .A(n4965), .ZN(n4966) );
  AOI21_X1 U5602 ( .B1(n5073), .B2(n6969), .A(n4966), .ZN(n4967) );
  OAI21_X1 U5603 ( .B1(n4968), .B2(n6397), .A(n4967), .ZN(U2983) );
  AOI22_X1 U5604 ( .A1(n6119), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .B1(n6235), 
        .B2(REIP_REG_5__SCAN_IN), .ZN(n4969) );
  OAI21_X1 U5605 ( .B1(n6125), .B2(n6276), .A(n4969), .ZN(n4970) );
  AOI21_X1 U5606 ( .B1(n4971), .B2(n6969), .A(n4970), .ZN(n4972) );
  OAI21_X1 U5607 ( .B1(n6397), .B2(n4973), .A(n4972), .ZN(U2981) );
  INV_X1 U5608 ( .A(DATAI_5_), .ZN(n6863) );
  OAI222_X1 U5609 ( .A1(n6278), .A2(n6475), .B1(n5521), .B2(n6863), .C1(n5520), 
        .C2(n5987), .ZN(U2886) );
  OAI21_X1 U5610 ( .B1(n4953), .B2(n4974), .A(n5003), .ZN(n6294) );
  INV_X1 U5611 ( .A(n4979), .ZN(n4975) );
  AOI21_X1 U5612 ( .B1(n4977), .B2(n4976), .A(n4975), .ZN(n6289) );
  AOI22_X1 U5613 ( .A1(n6082), .A2(n6289), .B1(EBX_REG_6__SCAN_IN), .B2(n5487), 
        .ZN(n4978) );
  OAI21_X1 U5614 ( .B1(n6294), .B2(n5489), .A(n4978), .ZN(U2853) );
  INV_X1 U5615 ( .A(DATAI_6_), .ZN(n6907) );
  OAI222_X1 U5616 ( .A1(n6294), .A2(n6475), .B1(n5521), .B2(n6907), .C1(n5989), 
        .C2(n5520), .ZN(U2885) );
  XNOR2_X1 U5617 ( .A(n5020), .B(n5019), .ZN(n5017) );
  AOI21_X1 U5618 ( .B1(n4980), .B2(n4979), .A(n5027), .ZN(n6299) );
  INV_X1 U5619 ( .A(REIP_REG_7__SCAN_IN), .ZN(n4981) );
  NOR2_X1 U5620 ( .A1(n6247), .A2(n4981), .ZN(n5013) );
  INV_X1 U5621 ( .A(n4994), .ZN(n4982) );
  NAND2_X1 U5622 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4982), .ZN(n5084)
         );
  INV_X1 U5623 ( .A(n5084), .ZN(n4985) );
  INV_X1 U5624 ( .A(n4983), .ZN(n4984) );
  OAI21_X1 U5625 ( .B1(n6194), .B2(n4985), .A(n4984), .ZN(n5018) );
  NOR2_X1 U5626 ( .A1(n5084), .A2(n4993), .ZN(n6188) );
  AOI22_X1 U5627 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n5018), .B1(n6188), 
        .B2(n3835), .ZN(n4986) );
  INV_X1 U5628 ( .A(n4986), .ZN(n4987) );
  AOI211_X1 U5629 ( .C1(n6243), .C2(n6299), .A(n5013), .B(n4987), .ZN(n4988)
         );
  OAI21_X1 U5630 ( .B1(n5017), .B2(n6225), .A(n4988), .ZN(U3011) );
  AND2_X1 U5631 ( .A1(n4990), .A2(n4989), .ZN(n4991) );
  XOR2_X1 U5632 ( .A(n4992), .B(n4991), .Z(n5006) );
  NOR3_X1 U5633 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4994), .A3(n4993), 
        .ZN(n5000) );
  INV_X1 U5634 ( .A(n6289), .ZN(n4998) );
  OAI21_X1 U5635 ( .B1(n4996), .B2(n4995), .A(INSTADDRPOINTER_REG_6__SCAN_IN), 
        .ZN(n4997) );
  NAND2_X1 U5636 ( .A1(n6235), .A2(REIP_REG_6__SCAN_IN), .ZN(n5007) );
  OAI211_X1 U5637 ( .C1(n6224), .C2(n4998), .A(n4997), .B(n5007), .ZN(n4999)
         );
  AOI211_X1 U5638 ( .C1(n5006), .C2(n6244), .A(n5000), .B(n4999), .ZN(n5001)
         );
  INV_X1 U5639 ( .A(n5001), .ZN(U3012) );
  NAND2_X1 U5640 ( .A1(n5003), .A2(n5002), .ZN(n5004) );
  AND2_X1 U5641 ( .A1(n5035), .A2(n5004), .ZN(n6305) );
  INV_X1 U5642 ( .A(n6305), .ZN(n5012) );
  AOI22_X1 U5643 ( .A1(n6299), .A2(n6082), .B1(EBX_REG_7__SCAN_IN), .B2(n5487), 
        .ZN(n5005) );
  OAI21_X1 U5644 ( .B1(n5012), .B2(n5489), .A(n5005), .ZN(U2852) );
  NAND2_X1 U5645 ( .A1(n5006), .A2(n6121), .ZN(n5011) );
  INV_X1 U5646 ( .A(n6293), .ZN(n5009) );
  OAI21_X1 U5647 ( .B1(n5627), .B2(n6292), .A(n5007), .ZN(n5008) );
  AOI21_X1 U5648 ( .B1(n5009), .B2(n6104), .A(n5008), .ZN(n5010) );
  OAI211_X1 U5649 ( .C1(n6862), .C2(n6294), .A(n5011), .B(n5010), .ZN(U2980)
         );
  INV_X1 U5650 ( .A(DATAI_7_), .ZN(n6964) );
  OAI222_X1 U5651 ( .A1(n5012), .A2(n6475), .B1(n5521), .B2(n6964), .C1(n5520), 
        .C2(n3997), .ZN(U2884) );
  AOI21_X1 U5652 ( .B1(n6119), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n5013), 
        .ZN(n5014) );
  OAI21_X1 U5653 ( .B1(n6125), .B2(n6303), .A(n5014), .ZN(n5015) );
  AOI21_X1 U5654 ( .B1(n6305), .B2(n6969), .A(n5015), .ZN(n5016) );
  OAI21_X1 U5655 ( .B1(n5017), .B2(n6397), .A(n5016), .ZN(U2979) );
  INV_X1 U5656 ( .A(n5018), .ZN(n6192) );
  NAND2_X1 U5657 ( .A1(n5020), .A2(n5019), .ZN(n5022) );
  NAND2_X1 U5658 ( .A1(n5022), .A2(n5021), .ZN(n5023) );
  XOR2_X1 U5659 ( .A(n5024), .B(n5023), .Z(n5039) );
  NAND2_X1 U5660 ( .A1(n5039), .A2(n6244), .ZN(n5032) );
  NOR2_X1 U5661 ( .A1(n4478), .A2(n3835), .ZN(n6193) );
  AOI21_X1 U5662 ( .B1(n4478), .B2(n3835), .A(n6193), .ZN(n5030) );
  NOR2_X1 U5663 ( .A1(n6247), .A2(n6019), .ZN(n5041) );
  NOR2_X1 U5664 ( .A1(n5027), .A2(n5026), .ZN(n5028) );
  OR2_X1 U5665 ( .A1(n5025), .A2(n5028), .ZN(n5052) );
  NOR2_X1 U5666 ( .A1(n6224), .A2(n5052), .ZN(n5029) );
  AOI211_X1 U5667 ( .C1(n5030), .C2(n6188), .A(n5041), .B(n5029), .ZN(n5031)
         );
  OAI211_X1 U5668 ( .C1(n6192), .C2(n4478), .A(n5032), .B(n5031), .ZN(U3010)
         );
  INV_X1 U5669 ( .A(n5033), .ZN(n5105) );
  NAND2_X1 U5670 ( .A1(n5035), .A2(n5034), .ZN(n5036) );
  NAND2_X1 U5671 ( .A1(n5105), .A2(n5036), .ZN(n5061) );
  INV_X1 U5672 ( .A(n5052), .ZN(n5037) );
  AOI22_X1 U5673 ( .A1(n5037), .A2(n6082), .B1(EBX_REG_8__SCAN_IN), .B2(n5487), 
        .ZN(n5038) );
  OAI21_X1 U5674 ( .B1(n5061), .B2(n5489), .A(n5038), .ZN(U2851) );
  NAND2_X1 U5675 ( .A1(n5039), .A2(n6121), .ZN(n5043) );
  NOR2_X1 U5676 ( .A1(n6125), .A2(n5051), .ZN(n5040) );
  AOI211_X1 U5677 ( .C1(n6119), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n5041), 
        .B(n5040), .ZN(n5042) );
  OAI211_X1 U5678 ( .C1(n6862), .C2(n5061), .A(n5043), .B(n5042), .ZN(U2978)
         );
  INV_X1 U5679 ( .A(DATAI_8_), .ZN(n5876) );
  OAI222_X1 U5680 ( .A1(n5061), .A2(n6475), .B1(n5521), .B2(n5876), .C1(n5520), 
        .C2(n5992), .ZN(U2883) );
  NAND2_X1 U5681 ( .A1(n6369), .A2(EBX_REG_0__SCAN_IN), .ZN(n5045) );
  OAI21_X1 U5682 ( .B1(n6354), .B2(n6370), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5044) );
  OAI211_X1 U5683 ( .C1(n6264), .C2(n6573), .A(n5045), .B(n5044), .ZN(n5046)
         );
  AOI21_X1 U5684 ( .B1(n6271), .B2(n5047), .A(n5046), .ZN(n5049) );
  NAND2_X1 U5685 ( .A1(n5349), .A2(REIP_REG_0__SCAN_IN), .ZN(n5048) );
  OAI211_X1 U5686 ( .C1(n5767), .C2(n6389), .A(n5049), .B(n5048), .ZN(U2827)
         );
  OAI21_X1 U5687 ( .B1(n6301), .B2(n6315), .A(n6283), .ZN(n6312) );
  OAI21_X1 U5688 ( .B1(n6301), .B2(n5050), .A(n6019), .ZN(n5059) );
  INV_X1 U5689 ( .A(n5051), .ZN(n5055) );
  OAI22_X1 U5690 ( .A1(n5053), .A2(n6382), .B1(n6389), .B2(n5052), .ZN(n5054)
         );
  AOI211_X1 U5691 ( .C1(n6354), .C2(n5055), .A(n5054), .B(n6362), .ZN(n5056)
         );
  OAI21_X1 U5692 ( .B1(n5057), .B2(n6384), .A(n5056), .ZN(n5058) );
  AOI21_X1 U5693 ( .B1(n6312), .B2(n5059), .A(n5058), .ZN(n5060) );
  OAI21_X1 U5694 ( .B1(n5061), .B2(n6390), .A(n5060), .ZN(U2819) );
  INV_X1 U5695 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5063) );
  OAI22_X1 U5696 ( .A1(n6384), .A2(n5063), .B1(n5062), .B2(n6395), .ZN(n5065)
         );
  NOR2_X1 U5697 ( .A1(n6264), .A2(n6638), .ZN(n5064) );
  AOI211_X1 U5698 ( .C1(n6369), .C2(EBX_REG_3__SCAN_IN), .A(n5065), .B(n5064), 
        .ZN(n5066) );
  OAI21_X1 U5699 ( .B1(n6389), .B2(n5067), .A(n5066), .ZN(n5072) );
  NAND2_X1 U5700 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .ZN(
        n5069) );
  AOI221_X1 U5701 ( .B1(n5070), .B2(n4870), .C1(n5069), .C2(n4870), .A(n5068), 
        .ZN(n5071) );
  AOI211_X1 U5702 ( .C1(n5073), .C2(n6271), .A(n5072), .B(n5071), .ZN(n5074)
         );
  INV_X1 U5703 ( .A(n5074), .ZN(U2824) );
  NAND2_X1 U5704 ( .A1(n5076), .A2(n5075), .ZN(n5133) );
  NAND2_X1 U5705 ( .A1(n5133), .A2(n5131), .ZN(n6109) );
  NAND2_X1 U5706 ( .A1(n6109), .A2(n5077), .ZN(n5078) );
  AND2_X1 U5707 ( .A1(n5078), .A2(n6098), .ZN(n5082) );
  NAND2_X1 U5708 ( .A1(n5080), .A2(n5079), .ZN(n5081) );
  XNOR2_X1 U5709 ( .A(n5082), .B(n5081), .ZN(n5163) );
  INV_X1 U5710 ( .A(n5163), .ZN(n5101) );
  INV_X1 U5711 ( .A(n6193), .ZN(n5083) );
  NOR4_X1 U5712 ( .A1(n6189), .A2(n4485), .A3(n5084), .A4(n5083), .ZN(n5087)
         );
  NAND3_X1 U5713 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n5087), .ZN(n5093) );
  AOI21_X1 U5714 ( .B1(n5086), .B2(n5093), .A(n5085), .ZN(n5223) );
  NAND2_X1 U5715 ( .A1(n5088), .A2(n5087), .ZN(n5092) );
  NAND2_X1 U5716 ( .A1(n5089), .A2(n5092), .ZN(n5220) );
  NAND2_X1 U5717 ( .A1(n5223), .A2(n5220), .ZN(n6213) );
  INV_X1 U5718 ( .A(n6213), .ZN(n6165) );
  NOR3_X1 U5719 ( .A1(n5763), .A2(n5090), .A3(n5093), .ZN(n5753) );
  INV_X1 U5720 ( .A(n5753), .ZN(n5091) );
  OAI21_X1 U5721 ( .B1(n5092), .B2(n6179), .A(n5091), .ZN(n6164) );
  NAND2_X1 U5722 ( .A1(n3853), .A2(n6233), .ZN(n6211) );
  AOI21_X1 U5723 ( .B1(n6165), .B2(n6211), .A(n6161), .ZN(n5099) );
  NOR3_X1 U5724 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n6215), .A3(n3853), 
        .ZN(n5098) );
  INV_X1 U5725 ( .A(REIP_REG_12__SCAN_IN), .ZN(n5094) );
  NOR2_X1 U5726 ( .A1(n6247), .A2(n5094), .ZN(n5166) );
  OR2_X1 U5727 ( .A1(n5154), .A2(n5095), .ZN(n5096) );
  NAND2_X1 U5728 ( .A1(n5180), .A2(n5096), .ZN(n5174) );
  NOR2_X1 U5729 ( .A1(n5174), .A2(n6224), .ZN(n5097) );
  NOR4_X1 U5730 ( .A1(n5099), .A2(n5098), .A3(n5166), .A4(n5097), .ZN(n5100)
         );
  OAI21_X1 U5731 ( .B1(n5101), .B2(n6225), .A(n5100), .ZN(U3006) );
  XOR2_X1 U5732 ( .A(n5103), .B(n5102), .Z(n6202) );
  INV_X1 U5733 ( .A(n6202), .ZN(n5112) );
  AND2_X1 U5734 ( .A1(n5105), .A2(n5104), .ZN(n5106) );
  NOR2_X1 U5735 ( .A1(n3445), .A2(n5106), .ZN(n6317) );
  INV_X1 U5736 ( .A(n6316), .ZN(n5109) );
  INV_X1 U5737 ( .A(REIP_REG_9__SCAN_IN), .ZN(n5107) );
  NOR2_X1 U5738 ( .A1(n6247), .A2(n5107), .ZN(n6200) );
  AOI21_X1 U5739 ( .B1(n6119), .B2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6200), 
        .ZN(n5108) );
  OAI21_X1 U5740 ( .B1(n6125), .B2(n5109), .A(n5108), .ZN(n5110) );
  AOI21_X1 U5741 ( .B1(n6317), .B2(n6969), .A(n5110), .ZN(n5111) );
  OAI21_X1 U5742 ( .B1(n5112), .B2(n6397), .A(n5111), .ZN(U2977) );
  INV_X1 U5743 ( .A(n5113), .ZN(n5150) );
  OAI21_X1 U5744 ( .B1(n3445), .B2(n5114), .A(n5150), .ZN(n5138) );
  INV_X1 U5745 ( .A(n5153), .ZN(n5115) );
  AOI21_X1 U5746 ( .B1(n5116), .B2(n5126), .A(n5115), .ZN(n6191) );
  AOI22_X1 U5747 ( .A1(n6191), .A2(n6082), .B1(EBX_REG_10__SCAN_IN), .B2(n5487), .ZN(n5117) );
  OAI21_X1 U5748 ( .B1(n5138), .B2(n5489), .A(n5117), .ZN(U2849) );
  AOI22_X1 U5749 ( .A1(EBX_REG_10__SCAN_IN), .A2(n6369), .B1(n6334), .B2(n6191), .ZN(n5118) );
  OAI211_X1 U5750 ( .C1(n6384), .C2(n5119), .A(n5118), .B(n6343), .ZN(n5124)
         );
  NOR2_X1 U5751 ( .A1(n6301), .A2(REIP_REG_9__SCAN_IN), .ZN(n6314) );
  OAI21_X1 U5752 ( .B1(n6312), .B2(n6314), .A(REIP_REG_10__SCAN_IN), .ZN(n5122) );
  NOR2_X1 U5753 ( .A1(n6301), .A2(n5120), .ZN(n5157) );
  INV_X1 U5754 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6021) );
  NAND2_X1 U5755 ( .A1(n5157), .A2(n6021), .ZN(n5121) );
  OAI211_X1 U5756 ( .C1(n5134), .C2(n6395), .A(n5122), .B(n5121), .ZN(n5123)
         );
  NOR2_X1 U5757 ( .A1(n5124), .A2(n5123), .ZN(n5125) );
  OAI21_X1 U5758 ( .B1(n5138), .B2(n6390), .A(n5125), .ZN(U2817) );
  INV_X1 U5759 ( .A(n6317), .ZN(n5130) );
  INV_X1 U5760 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5128) );
  OAI21_X1 U5761 ( .B1(n5025), .B2(n5127), .A(n5126), .ZN(n6199) );
  OAI222_X1 U5762 ( .A1(n5130), .A2(n5489), .B1(n5128), .B2(n6086), .C1(n5479), 
        .C2(n6199), .ZN(U2850) );
  INV_X1 U5763 ( .A(DATAI_9_), .ZN(n5129) );
  OAI222_X1 U5764 ( .A1(n5130), .A2(n6475), .B1(n5521), .B2(n5129), .C1(n5520), 
        .C2(n5994), .ZN(U2882) );
  NAND2_X1 U5765 ( .A1(n6100), .A2(n5131), .ZN(n5132) );
  XNOR2_X1 U5766 ( .A(n5133), .B(n5132), .ZN(n6195) );
  NAND2_X1 U5767 ( .A1(n6195), .A2(n6121), .ZN(n5137) );
  AND2_X1 U5768 ( .A1(n6235), .A2(REIP_REG_10__SCAN_IN), .ZN(n6190) );
  NOR2_X1 U5769 ( .A1(n6125), .A2(n5134), .ZN(n5135) );
  AOI211_X1 U5770 ( .C1(n6119), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6190), 
        .B(n5135), .ZN(n5136) );
  OAI211_X1 U5771 ( .C1(n6862), .C2(n5138), .A(n5137), .B(n5136), .ZN(U2976)
         );
  INV_X1 U5772 ( .A(DATAI_10_), .ZN(n5915) );
  OAI222_X1 U5773 ( .A1(n5138), .A2(n6475), .B1(n5521), .B2(n5915), .C1(n5520), 
        .C2(n5996), .ZN(U2881) );
  XNOR2_X1 U5774 ( .A(n5149), .B(n5139), .ZN(n5172) );
  OR2_X1 U5775 ( .A1(n6301), .A2(n5140), .ZN(n5141) );
  NAND2_X1 U5776 ( .A1(n5141), .A2(n6283), .ZN(n6328) );
  INV_X1 U5777 ( .A(n6328), .ZN(n5416) );
  OAI22_X1 U5778 ( .A1(n5416), .A2(n5094), .B1(n6389), .B2(n5174), .ZN(n5146)
         );
  INV_X1 U5779 ( .A(n5142), .ZN(n5143) );
  AND2_X1 U5780 ( .A1(n5157), .A2(n5143), .ZN(n6339) );
  INV_X1 U5781 ( .A(n6339), .ZN(n6322) );
  NOR2_X1 U5782 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6322), .ZN(n6329) );
  AOI211_X1 U5783 ( .C1(n6369), .C2(EBX_REG_12__SCAN_IN), .A(n6362), .B(n6329), 
        .ZN(n5144) );
  OAI21_X1 U5784 ( .B1(n5164), .B2(n6384), .A(n5144), .ZN(n5145) );
  AOI211_X1 U5785 ( .C1(n6354), .C2(n5167), .A(n5146), .B(n5145), .ZN(n5147)
         );
  OAI21_X1 U5786 ( .B1(n5172), .B2(n6390), .A(n5147), .ZN(U2815) );
  INV_X1 U5787 ( .A(n5148), .ZN(n5151) );
  AOI21_X1 U5788 ( .B1(n5151), .B2(n5150), .A(n5149), .ZN(n6105) );
  INV_X1 U5789 ( .A(n6105), .ZN(n5171) );
  AND2_X1 U5790 ( .A1(n5153), .A2(n5152), .ZN(n5155) );
  OR2_X1 U5791 ( .A1(n5155), .A2(n5154), .ZN(n6207) );
  AOI21_X1 U5792 ( .B1(n6354), .B2(n6103), .A(n6362), .ZN(n5156) );
  OAI21_X1 U5793 ( .B1(n6207), .B2(n6389), .A(n5156), .ZN(n5161) );
  NAND2_X1 U5794 ( .A1(REIP_REG_10__SCAN_IN), .A2(n5157), .ZN(n5159) );
  AOI22_X1 U5795 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n6370), .B1(
        EBX_REG_11__SCAN_IN), .B2(n6369), .ZN(n5158) );
  OAI21_X1 U5796 ( .B1(REIP_REG_11__SCAN_IN), .B2(n5159), .A(n5158), .ZN(n5160) );
  AOI211_X1 U5797 ( .C1(REIP_REG_11__SCAN_IN), .C2(n6328), .A(n5161), .B(n5160), .ZN(n5162) );
  OAI21_X1 U5798 ( .B1(n5171), .B2(n6390), .A(n5162), .ZN(U2816) );
  NAND2_X1 U5799 ( .A1(n5163), .A2(n6121), .ZN(n5169) );
  NOR2_X1 U5800 ( .A1(n5627), .A2(n5164), .ZN(n5165) );
  AOI211_X1 U5801 ( .C1(n6104), .C2(n5167), .A(n5166), .B(n5165), .ZN(n5168)
         );
  OAI211_X1 U5802 ( .C1(n5172), .C2(n6862), .A(n5169), .B(n5168), .ZN(U2974)
         );
  INV_X1 U5803 ( .A(DATAI_11_), .ZN(n5909) );
  OAI222_X1 U5804 ( .A1(n5171), .A2(n6475), .B1(n5521), .B2(n5909), .C1(n5520), 
        .C2(n5998), .ZN(U2880) );
  INV_X1 U5805 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5170) );
  OAI222_X1 U5806 ( .A1(n5171), .A2(n5489), .B1(n5170), .B2(n6086), .C1(n5479), 
        .C2(n6207), .ZN(U2848) );
  INV_X1 U5807 ( .A(DATAI_12_), .ZN(n5910) );
  OAI222_X1 U5808 ( .A1(n6475), .A2(n5172), .B1(n5521), .B2(n5910), .C1(n5520), 
        .C2(n4061), .ZN(U2879) );
  INV_X1 U5809 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5173) );
  OAI222_X1 U5810 ( .A1(n5174), .A2(n5479), .B1(n6086), .B2(n5173), .C1(n5489), 
        .C2(n5172), .ZN(U2847) );
  NAND2_X1 U5811 ( .A1(n5176), .A2(n5175), .ZN(n5177) );
  AND2_X1 U5812 ( .A1(n5178), .A2(n5177), .ZN(n6327) );
  INV_X1 U5813 ( .A(n6327), .ZN(n5183) );
  INV_X1 U5814 ( .A(n5484), .ZN(n5179) );
  AOI21_X1 U5815 ( .B1(n5181), .B2(n5180), .A(n5179), .ZN(n6323) );
  AOI22_X1 U5816 ( .A1(n6323), .A2(n6082), .B1(EBX_REG_13__SCAN_IN), .B2(n5487), .ZN(n5182) );
  OAI21_X1 U5817 ( .B1(n5183), .B2(n5489), .A(n5182), .ZN(U2846) );
  INV_X1 U5818 ( .A(DATAI_13_), .ZN(n5902) );
  OAI222_X1 U5819 ( .A1(n5183), .A2(n6475), .B1(n5521), .B2(n5902), .C1(n5520), 
        .C2(n6001), .ZN(U2878) );
  OAI22_X1 U5820 ( .A1(n3432), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4518), .ZN(n5188) );
  OAI22_X1 U5821 ( .A1(n5234), .A2(n5479), .B1(n6086), .B2(n5189), .ZN(U2828)
         );
  NAND2_X1 U5822 ( .A1(n5272), .A2(n5190), .ZN(n5194) );
  AOI22_X1 U5823 ( .A1(n4427), .A2(EAX_REG_31__SCAN_IN), .B1(n5191), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5192) );
  INV_X1 U5824 ( .A(n5192), .ZN(n5193) );
  NAND2_X1 U5825 ( .A1(n5490), .A2(n6375), .ZN(n5205) );
  INV_X1 U5826 ( .A(n5195), .ZN(n5196) );
  NOR3_X1 U5827 ( .A1(n5279), .A2(REIP_REG_31__SCAN_IN), .A3(n5196), .ZN(n5202) );
  INV_X1 U5828 ( .A(n5197), .ZN(n6429) );
  NAND4_X1 U5829 ( .A1(n5198), .A2(n6147), .A3(EBX_REG_31__SCAN_IN), .A4(n6429), .ZN(n5199) );
  OAI21_X1 U5830 ( .B1(n6384), .B2(n5200), .A(n5199), .ZN(n5201) );
  AOI211_X1 U5831 ( .C1(n5203), .C2(REIP_REG_31__SCAN_IN), .A(n5202), .B(n5201), .ZN(n5204) );
  OAI211_X1 U5832 ( .C1(n5234), .C2(n6389), .A(n5205), .B(n5204), .ZN(U2796)
         );
  INV_X1 U5833 ( .A(n5539), .ZN(n5206) );
  OAI21_X1 U5834 ( .B1(n5748), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5206), 
        .ZN(n5531) );
  XOR2_X1 U5835 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .B(n3851), .Z(n5524) );
  INV_X1 U5836 ( .A(n5524), .ZN(n5207) );
  INV_X1 U5837 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5665) );
  NAND2_X1 U5838 ( .A1(n5209), .A2(n5665), .ZN(n5212) );
  NAND2_X1 U5839 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5210) );
  NAND2_X1 U5840 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n5210), .ZN(n5211) );
  NOR3_X1 U5841 ( .A1(n5215), .A2(n6161), .A3(n3853), .ZN(n6174) );
  NAND2_X1 U5842 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6174), .ZN(n6216) );
  NOR3_X1 U5843 ( .A1(n6230), .A2(n6222), .A3(n6216), .ZN(n5758) );
  NAND3_X1 U5844 ( .A1(n5219), .A2(n5758), .A3(n6233), .ZN(n6160) );
  INV_X1 U5845 ( .A(n5740), .ZN(n5224) );
  NOR2_X1 U5846 ( .A1(n6160), .A2(n5224), .ZN(n6251) );
  NAND2_X1 U5847 ( .A1(n6251), .A2(n5216), .ZN(n5721) );
  AND2_X1 U5848 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5692) );
  INV_X1 U5849 ( .A(n5692), .ZN(n5217) );
  NOR2_X1 U5850 ( .A1(n5703), .A2(n5217), .ZN(n5656) );
  INV_X1 U5851 ( .A(n5656), .ZN(n5687) );
  NOR4_X1 U5852 ( .A1(n5687), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n5654), 
        .A4(n3875), .ZN(n5232) );
  INV_X1 U5853 ( .A(n5675), .ZN(n5666) );
  NAND2_X1 U5854 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5218) );
  NAND2_X1 U5855 ( .A1(n6251), .A2(n5218), .ZN(n5731) );
  NAND3_X1 U5856 ( .A1(n5220), .A2(n5219), .A3(n5758), .ZN(n5221) );
  NAND2_X1 U5857 ( .A1(n6214), .A2(n5221), .ZN(n5222) );
  NAND2_X1 U5858 ( .A1(n5223), .A2(n5222), .ZN(n6155) );
  AND2_X1 U5859 ( .A1(n6214), .A2(n5224), .ZN(n5225) );
  NOR2_X1 U5860 ( .A1(n6155), .A2(n5225), .ZN(n6246) );
  NAND2_X1 U5861 ( .A1(n5731), .A2(n6246), .ZN(n5726) );
  INV_X1 U5862 ( .A(n5226), .ZN(n5227) );
  AOI21_X1 U5863 ( .B1(n6183), .B2(n6179), .A(n5227), .ZN(n5228) );
  NOR2_X1 U5864 ( .A1(n5726), .A2(n5228), .ZN(n5711) );
  OAI21_X1 U5865 ( .B1(n6194), .B2(n5692), .A(n5711), .ZN(n5689) );
  AOI211_X1 U5866 ( .C1(n5666), .C2(n6214), .A(n5665), .B(n5689), .ZN(n5664)
         );
  INV_X1 U5867 ( .A(n5711), .ZN(n5697) );
  NOR2_X1 U5868 ( .A1(n5697), .A2(n6214), .ZN(n5658) );
  AOI211_X1 U5869 ( .C1(n5664), .C2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5658), .B(n5229), .ZN(n5230) );
  INV_X1 U5870 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6054) );
  NOR2_X1 U5871 ( .A1(n6247), .A2(n6054), .ZN(n5237) );
  OAI21_X1 U5872 ( .B1(n5242), .B2(n6225), .A(n5236), .ZN(U2987) );
  AOI21_X1 U5873 ( .B1(n6119), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5237), 
        .ZN(n5238) );
  OAI21_X1 U5874 ( .B1(n6125), .B2(n5239), .A(n5238), .ZN(n5240) );
  OAI21_X1 U5875 ( .B1(n5242), .B2(n6397), .A(n5241), .ZN(U2955) );
  OAI222_X1 U5876 ( .A1(n5243), .A2(n5489), .B1(n5244), .B2(n6086), .C1(n5479), 
        .C2(n5653), .ZN(U2829) );
  NAND2_X1 U5877 ( .A1(n4790), .A2(n3446), .ZN(n5247) );
  OAI22_X1 U5878 ( .A1(n5248), .A2(n5247), .B1(n5246), .B2(n5245), .ZN(n5249)
         );
  AOI21_X1 U5879 ( .B1(n5250), .B2(n6434), .A(n5249), .ZN(n5254) );
  INV_X1 U5880 ( .A(n4790), .ZN(n5251) );
  AOI21_X1 U5881 ( .B1(n6444), .B2(n5251), .A(n5253), .ZN(n5252) );
  OAI22_X1 U5882 ( .A1(n5254), .A2(n5253), .B1(n5252), .B2(n3446), .ZN(U3459)
         );
  INV_X1 U5883 ( .A(n5263), .ZN(n5255) );
  NOR2_X1 U5884 ( .A1(n5256), .A2(n5255), .ZN(n5257) );
  MUX2_X1 U5885 ( .A(n5258), .B(n5257), .S(n5262), .Z(n5261) );
  OR2_X1 U5886 ( .A1(n5264), .A2(n5259), .ZN(n5260) );
  AND2_X1 U5887 ( .A1(n5261), .A2(n5260), .ZN(n6420) );
  INV_X1 U5888 ( .A(n6420), .ZN(n5269) );
  NAND2_X1 U5889 ( .A1(n5262), .A2(n3882), .ZN(n5267) );
  OAI21_X1 U5890 ( .B1(n5265), .B2(n5264), .A(n5263), .ZN(n5266) );
  NAND2_X1 U5891 ( .A1(n5267), .A2(n5266), .ZN(n6126) );
  NAND2_X1 U5892 ( .A1(n3659), .A2(n5268), .ZN(n6131) );
  AOI21_X1 U5893 ( .B1(n6131), .B2(n6141), .A(READY_N), .ZN(n6145) );
  OR2_X1 U5894 ( .A1(n6126), .A2(n6145), .ZN(n6421) );
  AND2_X1 U5895 ( .A1(n6421), .A2(n6449), .ZN(n6399) );
  MUX2_X1 U5896 ( .A(MORE_REG_SCAN_IN), .B(n5269), .S(n6399), .Z(U3471) );
  INV_X1 U5897 ( .A(n5270), .ZN(n5274) );
  INV_X1 U5898 ( .A(n5290), .ZN(n5273) );
  AOI21_X1 U5899 ( .B1(n5274), .B2(n5273), .A(n5272), .ZN(n5528) );
  INV_X1 U5900 ( .A(n5528), .ZN(n5500) );
  INV_X1 U5901 ( .A(n5295), .ZN(n5284) );
  INV_X1 U5902 ( .A(n5275), .ZN(n5526) );
  OAI22_X1 U5903 ( .A1(n6384), .A2(n5276), .B1(n5526), .B2(n6395), .ZN(n5277)
         );
  AOI21_X1 U5904 ( .B1(n6369), .B2(EBX_REG_29__SCAN_IN), .A(n5277), .ZN(n5278)
         );
  OAI21_X1 U5905 ( .B1(n5279), .B2(REIP_REG_29__SCAN_IN), .A(n5278), .ZN(n5283) );
  OAI21_X1 U5906 ( .B1(n5288), .B2(n5281), .A(n5280), .ZN(n5667) );
  NOR2_X1 U5907 ( .A1(n5667), .A2(n6389), .ZN(n5282) );
  AOI211_X1 U5908 ( .C1(n5284), .C2(REIP_REG_29__SCAN_IN), .A(n5283), .B(n5282), .ZN(n5285) );
  OAI21_X1 U5909 ( .B1(n5500), .B2(n6390), .A(n5285), .ZN(U2798) );
  NOR2_X1 U5910 ( .A1(n5302), .A2(n5286), .ZN(n5287) );
  OR2_X1 U5911 ( .A1(n5288), .A2(n5287), .ZN(n5674) );
  AOI21_X1 U5912 ( .B1(n5291), .B2(n5289), .A(n5290), .ZN(n5537) );
  NAND2_X1 U5913 ( .A1(n5537), .A2(n6375), .ZN(n5299) );
  OAI22_X1 U5914 ( .A1(n6384), .A2(n5292), .B1(n5535), .B2(n6395), .ZN(n5297)
         );
  AOI21_X1 U5915 ( .B1(n5293), .B2(REIP_REG_27__SCAN_IN), .A(
        REIP_REG_28__SCAN_IN), .ZN(n5294) );
  NOR2_X1 U5916 ( .A1(n5295), .A2(n5294), .ZN(n5296) );
  AOI211_X1 U5917 ( .C1(EBX_REG_28__SCAN_IN), .C2(n6369), .A(n5297), .B(n5296), 
        .ZN(n5298) );
  OAI211_X1 U5918 ( .C1(n6389), .C2(n5674), .A(n5299), .B(n5298), .ZN(U2799)
         );
  OAI21_X1 U5919 ( .B1(n5316), .B2(n5301), .A(n5289), .ZN(n5543) );
  INV_X1 U5920 ( .A(n5302), .ZN(n5305) );
  NAND2_X1 U5921 ( .A1(n5325), .A2(n5303), .ZN(n5304) );
  NAND2_X1 U5922 ( .A1(n5305), .A2(n5304), .ZN(n5427) );
  INV_X1 U5923 ( .A(n5427), .ZN(n5685) );
  NAND3_X1 U5924 ( .A1(n5306), .A2(REIP_REG_27__SCAN_IN), .A3(n5349), .ZN(
        n5311) );
  INV_X1 U5925 ( .A(n5307), .ZN(n5545) );
  OAI22_X1 U5926 ( .A1(n6384), .A2(n5308), .B1(n5545), .B2(n6395), .ZN(n5309)
         );
  AOI21_X1 U5927 ( .B1(n6369), .B2(EBX_REG_27__SCAN_IN), .A(n5309), .ZN(n5310)
         );
  OAI211_X1 U5928 ( .C1(REIP_REG_27__SCAN_IN), .C2(n5312), .A(n5311), .B(n5310), .ZN(n5313) );
  AOI21_X1 U5929 ( .B1(n5685), .B2(n6334), .A(n5313), .ZN(n5314) );
  OAI21_X1 U5930 ( .B1(n5543), .B2(n6390), .A(n5314), .ZN(U2800) );
  AOI21_X1 U5931 ( .B1(n5317), .B2(n5315), .A(n5316), .ZN(n5554) );
  INV_X1 U5932 ( .A(n5554), .ZN(n5508) );
  OAI22_X1 U5933 ( .A1(n6384), .A2(n5318), .B1(n5552), .B2(n6395), .ZN(n5323)
         );
  INV_X1 U5934 ( .A(n5349), .ZN(n5417) );
  INV_X1 U5935 ( .A(n5338), .ZN(n5319) );
  AOI21_X1 U5936 ( .B1(n5319), .B2(REIP_REG_25__SCAN_IN), .A(
        REIP_REG_26__SCAN_IN), .ZN(n5320) );
  AOI211_X1 U5937 ( .C1(n5321), .C2(REIP_REG_26__SCAN_IN), .A(n5417), .B(n5320), .ZN(n5322) );
  AOI211_X1 U5938 ( .C1(EBX_REG_26__SCAN_IN), .C2(n6369), .A(n5323), .B(n5322), 
        .ZN(n5329) );
  INV_X1 U5939 ( .A(n5325), .ZN(n5326) );
  AOI21_X1 U5940 ( .B1(n5327), .B2(n5324), .A(n5326), .ZN(n5696) );
  NAND2_X1 U5941 ( .A1(n5696), .A2(n6334), .ZN(n5328) );
  OAI211_X1 U5942 ( .C1(n5508), .C2(n6390), .A(n5329), .B(n5328), .ZN(U2801)
         );
  OAI21_X1 U5943 ( .B1(n5344), .B2(n5331), .A(n5315), .ZN(n5562) );
  INV_X1 U5944 ( .A(n5346), .ZN(n5332) );
  NAND2_X1 U5945 ( .A1(n5368), .A2(n5332), .ZN(n5334) );
  NAND2_X1 U5946 ( .A1(n5334), .A2(n5333), .ZN(n5335) );
  NAND2_X1 U5947 ( .A1(n5335), .A2(n5324), .ZN(n5430) );
  INV_X1 U5948 ( .A(n5430), .ZN(n5702) );
  INV_X1 U5949 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5431) );
  NOR3_X1 U5950 ( .A1(n5417), .A2(n5336), .A3(n6043), .ZN(n5340) );
  OAI22_X1 U5951 ( .A1(REIP_REG_25__SCAN_IN), .A2(n5338), .B1(n5337), .B2(
        n6384), .ZN(n5339) );
  AOI211_X1 U5952 ( .C1(n6354), .C2(n5559), .A(n5340), .B(n5339), .ZN(n5341)
         );
  OAI21_X1 U5953 ( .B1(n6382), .B2(n5431), .A(n5341), .ZN(n5342) );
  AOI21_X1 U5954 ( .B1(n5702), .B2(n6334), .A(n5342), .ZN(n5343) );
  OAI21_X1 U5955 ( .B1(n5562), .B2(n6390), .A(n5343), .ZN(U2802) );
  AOI21_X1 U5956 ( .B1(n5345), .B2(n5361), .A(n5344), .ZN(n6685) );
  INV_X1 U5957 ( .A(n6685), .ZN(n5356) );
  XNOR2_X1 U5958 ( .A(n5368), .B(n5346), .ZN(n6081) );
  INV_X1 U5959 ( .A(n5347), .ZN(n5353) );
  AND2_X1 U5960 ( .A1(n5349), .A2(n5348), .ZN(n5373) );
  NAND2_X1 U5961 ( .A1(n5373), .A2(REIP_REG_24__SCAN_IN), .ZN(n5352) );
  INV_X1 U5962 ( .A(EBX_REG_24__SCAN_IN), .ZN(n6085) );
  OAI22_X1 U5963 ( .A1(n5576), .A2(n6384), .B1(n6085), .B2(n6382), .ZN(n5350)
         );
  AOI21_X1 U5964 ( .B1(n6354), .B2(n5574), .A(n5350), .ZN(n5351) );
  OAI211_X1 U5965 ( .C1(n5353), .C2(REIP_REG_24__SCAN_IN), .A(n5352), .B(n5351), .ZN(n5354) );
  AOI21_X1 U5966 ( .B1(n6081), .B2(n6334), .A(n5354), .ZN(n5355) );
  OAI21_X1 U5967 ( .B1(n5356), .B2(n6390), .A(n5355), .ZN(U2803) );
  AND2_X1 U5968 ( .A1(n5357), .A2(n5482), .ZN(n5359) );
  AND2_X1 U5969 ( .A1(n5359), .A2(n5358), .ZN(n5436) );
  OR2_X1 U5970 ( .A1(n5436), .A2(n5360), .ZN(n5362) );
  AND2_X1 U5971 ( .A1(n5362), .A2(n5361), .ZN(n5587) );
  INV_X1 U5972 ( .A(n6379), .ZN(n5364) );
  NAND2_X1 U5973 ( .A1(REIP_REG_18__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .ZN(
        n5395) );
  NOR2_X1 U5974 ( .A1(n6301), .A2(n5363), .ZN(n5408) );
  NAND2_X1 U5975 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5408), .ZN(n6360) );
  NOR2_X1 U5976 ( .A1(n5395), .A2(n6360), .ZN(n6368) );
  NAND2_X1 U5977 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6368), .ZN(n6378) );
  INV_X1 U5978 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6039) );
  OAI21_X1 U5979 ( .B1(n5364), .B2(n6378), .A(n6039), .ZN(n5372) );
  INV_X1 U5980 ( .A(n5365), .ZN(n5585) );
  AND2_X1 U5981 ( .A1(n5440), .A2(n5366), .ZN(n5367) );
  NOR2_X1 U5982 ( .A1(n5368), .A2(n5367), .ZN(n5720) );
  NAND2_X1 U5983 ( .A1(n5720), .A2(n6334), .ZN(n5370) );
  AOI22_X1 U5984 ( .A1(PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n6370), .B1(
        EBX_REG_23__SCAN_IN), .B2(n6369), .ZN(n5369) );
  OAI211_X1 U5985 ( .C1(n6395), .C2(n5585), .A(n5370), .B(n5369), .ZN(n5371)
         );
  AOI21_X1 U5986 ( .B1(n5373), .B2(n5372), .A(n5371), .ZN(n5374) );
  OAI21_X1 U5987 ( .B1(n5513), .B2(n6390), .A(n5374), .ZN(U2804) );
  NOR2_X1 U5988 ( .A1(n5481), .A2(n5375), .ZN(n5451) );
  NOR2_X1 U5989 ( .A1(n5481), .A2(n5376), .ZN(n5434) );
  INV_X1 U5990 ( .A(n5434), .ZN(n5377) );
  OAI21_X1 U5991 ( .B1(n5378), .B2(n5451), .A(n5377), .ZN(n5603) );
  NOR2_X1 U5992 ( .A1(n5417), .A2(n5379), .ZN(n6387) );
  INV_X1 U5993 ( .A(n6378), .ZN(n5381) );
  INV_X1 U5994 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5443) );
  OAI22_X1 U5995 ( .A1(n5598), .A2(n6384), .B1(n5443), .B2(n6382), .ZN(n5380)
         );
  AOI221_X1 U5996 ( .B1(n6387), .B2(REIP_REG_21__SCAN_IN), .C1(n5381), .C2(
        n6380), .A(n5380), .ZN(n5386) );
  NAND2_X1 U5997 ( .A1(n5382), .A2(n5383), .ZN(n5384) );
  AND2_X1 U5998 ( .A1(n5438), .A2(n5384), .ZN(n6242) );
  AOI22_X1 U5999 ( .A1(n6242), .A2(n6334), .B1(n6354), .B2(n5600), .ZN(n5385)
         );
  OAI211_X1 U6000 ( .C1(n5603), .C2(n6390), .A(n5386), .B(n5385), .ZN(U2806)
         );
  NAND2_X1 U6001 ( .A1(n5470), .A2(n5387), .ZN(n5450) );
  NAND2_X1 U6002 ( .A1(n5470), .A2(n5388), .ZN(n5458) );
  NAND2_X1 U6003 ( .A1(n5458), .A2(n5389), .ZN(n5390) );
  NAND2_X1 U6004 ( .A1(n5450), .A2(n5390), .ZN(n5610) );
  INV_X1 U6005 ( .A(n5391), .ZN(n5393) );
  INV_X1 U6006 ( .A(n5461), .ZN(n5392) );
  AOI21_X1 U6007 ( .B1(n5393), .B2(n5392), .A(n5447), .ZN(n6156) );
  NAND2_X1 U6008 ( .A1(n6354), .A2(n5607), .ZN(n5394) );
  OAI211_X1 U6009 ( .C1(n6384), .C2(n5605), .A(n5394), .B(n6343), .ZN(n5400)
         );
  OAI21_X1 U6010 ( .B1(REIP_REG_18__SCAN_IN), .B2(REIP_REG_19__SCAN_IN), .A(
        n5395), .ZN(n5398) );
  OAI21_X1 U6011 ( .B1(n6301), .B2(n5396), .A(n6283), .ZN(n6358) );
  AOI22_X1 U6012 ( .A1(EBX_REG_19__SCAN_IN), .A2(n6369), .B1(
        REIP_REG_19__SCAN_IN), .B2(n6358), .ZN(n5397) );
  OAI21_X1 U6013 ( .B1(n6360), .B2(n5398), .A(n5397), .ZN(n5399) );
  AOI211_X1 U6014 ( .C1(n6156), .C2(n6334), .A(n5400), .B(n5399), .ZN(n5401)
         );
  OAI21_X1 U6015 ( .B1(n5610), .B2(n6390), .A(n5401), .ZN(U2808) );
  NAND2_X1 U6016 ( .A1(n5470), .A2(n5402), .ZN(n5456) );
  NAND2_X1 U6017 ( .A1(n5474), .A2(n5404), .ZN(n5405) );
  AND2_X1 U6018 ( .A1(n5460), .A2(n5405), .ZN(n6236) );
  INV_X1 U6019 ( .A(n5615), .ZN(n5407) );
  NAND2_X1 U6020 ( .A1(n6369), .A2(EBX_REG_17__SCAN_IN), .ZN(n5406) );
  OAI211_X1 U6021 ( .C1(n5407), .C2(n6395), .A(n5406), .B(n6343), .ZN(n5411)
         );
  OAI21_X1 U6022 ( .B1(REIP_REG_17__SCAN_IN), .B2(n5408), .A(n6358), .ZN(n5409) );
  OAI21_X1 U6023 ( .B1(n6384), .B2(n5613), .A(n5409), .ZN(n5410) );
  AOI211_X1 U6024 ( .C1(n6236), .C2(n6334), .A(n5411), .B(n5410), .ZN(n5412)
         );
  OAI21_X1 U6025 ( .B1(n5618), .B2(n6390), .A(n5412), .ZN(U2810) );
  AND2_X1 U6026 ( .A1(n5481), .A2(n5413), .ZN(n5414) );
  INV_X1 U6027 ( .A(n5639), .ZN(n5423) );
  NAND2_X1 U6028 ( .A1(n5418), .A2(n6339), .ZN(n6351) );
  AOI21_X1 U6029 ( .B1(n5415), .B2(n5486), .A(n5472), .ZN(n6217) );
  INV_X1 U6030 ( .A(n6217), .ZN(n5478) );
  OAI22_X1 U6031 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6351), .B1(n6389), .B2(
        n5478), .ZN(n5422) );
  INV_X1 U6032 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5420) );
  OAI21_X1 U6033 ( .B1(n5418), .B2(n5417), .A(n5416), .ZN(n6348) );
  AOI22_X1 U6034 ( .A1(EBX_REG_15__SCAN_IN), .A2(n6369), .B1(
        REIP_REG_15__SCAN_IN), .B2(n6348), .ZN(n5419) );
  OAI211_X1 U6035 ( .C1(n6384), .C2(n5420), .A(n5419), .B(n6343), .ZN(n5421)
         );
  AOI211_X1 U6036 ( .C1(n6354), .C2(n5423), .A(n5422), .B(n5421), .ZN(n5424)
         );
  OAI21_X1 U6037 ( .B1(n5637), .B2(n6390), .A(n5424), .ZN(U2812) );
  INV_X1 U6038 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5425) );
  OAI222_X1 U6039 ( .A1(n5489), .A2(n5500), .B1(n5425), .B2(n6086), .C1(n5667), 
        .C2(n5479), .ZN(U2830) );
  INV_X1 U6040 ( .A(n5537), .ZN(n5503) );
  INV_X1 U6041 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5426) );
  OAI222_X1 U6042 ( .A1(n5489), .A2(n5503), .B1(n5426), .B2(n6086), .C1(n5674), 
        .C2(n5479), .ZN(U2831) );
  INV_X1 U6043 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5428) );
  OAI222_X1 U6044 ( .A1(n5489), .A2(n5543), .B1(n5428), .B2(n6086), .C1(n5427), 
        .C2(n5479), .ZN(U2832) );
  AOI22_X1 U6045 ( .A1(n5696), .A2(n6082), .B1(EBX_REG_26__SCAN_IN), .B2(n5487), .ZN(n5429) );
  OAI21_X1 U6046 ( .B1(n5508), .B2(n5489), .A(n5429), .ZN(U2833) );
  OAI222_X1 U6047 ( .A1(n5562), .A2(n5489), .B1(n5431), .B2(n6086), .C1(n5430), 
        .C2(n5479), .ZN(U2834) );
  AOI22_X1 U6048 ( .A1(n5720), .A2(n6082), .B1(EBX_REG_23__SCAN_IN), .B2(n5487), .ZN(n5432) );
  OAI21_X1 U6049 ( .B1(n5513), .B2(n5489), .A(n5432), .ZN(U2836) );
  NOR2_X1 U6050 ( .A1(n5434), .A2(n5433), .ZN(n5435) );
  INV_X1 U6051 ( .A(n6391), .ZN(n6485) );
  INV_X1 U6052 ( .A(n5489), .ZN(n6083) );
  NAND2_X1 U6053 ( .A1(n5438), .A2(n5437), .ZN(n5439) );
  NAND2_X1 U6054 ( .A1(n5440), .A2(n5439), .ZN(n6388) );
  OAI22_X1 U6055 ( .A1(n6388), .A2(n5479), .B1(n6383), .B2(n6086), .ZN(n5441)
         );
  AOI21_X1 U6056 ( .B1(n6485), .B2(n6083), .A(n5441), .ZN(n5442) );
  INV_X1 U6057 ( .A(n5442), .ZN(U2837) );
  NOR2_X1 U6058 ( .A1(n6086), .A2(n5443), .ZN(n5444) );
  AOI21_X1 U6059 ( .B1(n6242), .B2(n6082), .A(n5444), .ZN(n5445) );
  OAI21_X1 U6060 ( .B1(n5603), .B2(n5489), .A(n5445), .ZN(U2838) );
  OR2_X1 U6061 ( .A1(n5447), .A2(n5446), .ZN(n5448) );
  NAND2_X1 U6062 ( .A1(n5382), .A2(n5448), .ZN(n6377) );
  INV_X1 U6063 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5453) );
  AND2_X1 U6064 ( .A1(n5450), .A2(n5449), .ZN(n5452) );
  OAI222_X1 U6065 ( .A1(n5479), .A2(n6377), .B1(n5453), .B2(n6086), .C1(n6120), 
        .C2(n5489), .ZN(U2839) );
  AOI22_X1 U6066 ( .A1(n6156), .A2(n6082), .B1(EBX_REG_19__SCAN_IN), .B2(n5487), .ZN(n5454) );
  OAI21_X1 U6067 ( .B1(n5610), .B2(n5489), .A(n5454), .ZN(U2840) );
  NAND2_X1 U6068 ( .A1(n5456), .A2(n5455), .ZN(n5457) );
  AND2_X1 U6069 ( .A1(n5460), .A2(n5459), .ZN(n5462) );
  OR2_X1 U6070 ( .A1(n5462), .A2(n5461), .ZN(n6367) );
  OAI22_X1 U6071 ( .A1(n6367), .A2(n5479), .B1(n5463), .B2(n6086), .ZN(n5464)
         );
  AOI21_X1 U6072 ( .B1(n6479), .B2(n6083), .A(n5464), .ZN(n5465) );
  INV_X1 U6073 ( .A(n5465), .ZN(U2841) );
  AOI22_X1 U6074 ( .A1(n6236), .A2(n6082), .B1(EBX_REG_17__SCAN_IN), .B2(n5487), .ZN(n5466) );
  OAI21_X1 U6075 ( .B1(n5618), .B2(n5489), .A(n5466), .ZN(U2842) );
  INV_X1 U6076 ( .A(n5467), .ZN(n5468) );
  OAI21_X1 U6077 ( .B1(n5470), .B2(n5469), .A(n5468), .ZN(n5628) );
  INV_X1 U6078 ( .A(n5628), .ZN(n6476) );
  OR2_X1 U6079 ( .A1(n5472), .A2(n5471), .ZN(n5473) );
  NAND2_X1 U6080 ( .A1(n5474), .A2(n5473), .ZN(n6357) );
  OAI22_X1 U6081 ( .A1(n6357), .A2(n5479), .B1(n5475), .B2(n6086), .ZN(n5476)
         );
  AOI21_X1 U6082 ( .B1(n6476), .B2(n6083), .A(n5476), .ZN(n5477) );
  INV_X1 U6083 ( .A(n5477), .ZN(U2843) );
  INV_X1 U6084 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5480) );
  OAI222_X1 U6085 ( .A1(n5637), .A2(n5489), .B1(n5480), .B2(n6086), .C1(n5479), 
        .C2(n5478), .ZN(U2844) );
  OAI21_X1 U6086 ( .B1(n5357), .B2(n5482), .A(n5481), .ZN(n5647) );
  NAND2_X1 U6087 ( .A1(n5484), .A2(n5483), .ZN(n5485) );
  AND2_X1 U6088 ( .A1(n5486), .A2(n5485), .ZN(n6333) );
  AOI22_X1 U6089 ( .A1(n6333), .A2(n6082), .B1(EBX_REG_14__SCAN_IN), .B2(n5487), .ZN(n5488) );
  OAI21_X1 U6090 ( .B1(n5647), .B2(n5489), .A(n5488), .ZN(U2845) );
  NAND3_X1 U6091 ( .A1(n5490), .A2(n6965), .A3(n5520), .ZN(n5493) );
  NOR2_X2 U6092 ( .A1(n6686), .A2(n5491), .ZN(n6683) );
  AOI22_X1 U6093 ( .A1(n6683), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6686), .ZN(n5492) );
  NAND2_X1 U6094 ( .A1(n5493), .A2(n5492), .ZN(U2860) );
  AOI22_X1 U6095 ( .A1(n6683), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n6686), .ZN(n5497) );
  AND2_X1 U6096 ( .A1(n6864), .A2(n5494), .ZN(n5495) );
  NAND2_X1 U6097 ( .A1(n6687), .A2(DATAI_14_), .ZN(n5496) );
  OAI211_X1 U6098 ( .C1(n5243), .C2(n6475), .A(n5497), .B(n5496), .ZN(U2861)
         );
  AOI22_X1 U6099 ( .A1(n6683), .A2(DATAI_29_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n6686), .ZN(n5499) );
  NAND2_X1 U6100 ( .A1(n6687), .A2(DATAI_13_), .ZN(n5498) );
  OAI211_X1 U6101 ( .C1(n5500), .C2(n6475), .A(n5499), .B(n5498), .ZN(U2862)
         );
  AOI22_X1 U6102 ( .A1(n6683), .A2(DATAI_28_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n6686), .ZN(n5502) );
  NAND2_X1 U6103 ( .A1(n6687), .A2(DATAI_12_), .ZN(n5501) );
  OAI211_X1 U6104 ( .C1(n5503), .C2(n6475), .A(n5502), .B(n5501), .ZN(U2863)
         );
  AOI22_X1 U6105 ( .A1(n6683), .A2(DATAI_27_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n6686), .ZN(n5505) );
  NAND2_X1 U6106 ( .A1(n6687), .A2(DATAI_11_), .ZN(n5504) );
  OAI211_X1 U6107 ( .C1(n5543), .C2(n6475), .A(n5505), .B(n5504), .ZN(U2864)
         );
  AOI22_X1 U6108 ( .A1(n6683), .A2(DATAI_26_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n6686), .ZN(n5507) );
  NAND2_X1 U6109 ( .A1(n6687), .A2(DATAI_10_), .ZN(n5506) );
  OAI211_X1 U6110 ( .C1(n5508), .C2(n6475), .A(n5507), .B(n5506), .ZN(U2865)
         );
  AOI22_X1 U6111 ( .A1(n6683), .A2(DATAI_25_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n6686), .ZN(n5510) );
  NAND2_X1 U6112 ( .A1(n6687), .A2(DATAI_9_), .ZN(n5509) );
  OAI211_X1 U6113 ( .C1(n5562), .C2(n6475), .A(n5510), .B(n5509), .ZN(U2866)
         );
  AOI22_X1 U6114 ( .A1(n6683), .A2(DATAI_23_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n6686), .ZN(n5512) );
  NAND2_X1 U6115 ( .A1(n6687), .A2(DATAI_7_), .ZN(n5511) );
  OAI211_X1 U6116 ( .C1(n5513), .C2(n6475), .A(n5512), .B(n5511), .ZN(U2868)
         );
  AOI22_X1 U6117 ( .A1(n6683), .A2(DATAI_21_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n6686), .ZN(n5515) );
  NAND2_X1 U6118 ( .A1(n6687), .A2(DATAI_5_), .ZN(n5514) );
  OAI211_X1 U6119 ( .C1(n5603), .C2(n6475), .A(n5515), .B(n5514), .ZN(U2870)
         );
  AOI22_X1 U6120 ( .A1(n6683), .A2(DATAI_19_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n6686), .ZN(n5517) );
  NAND2_X1 U6121 ( .A1(n6687), .A2(DATAI_3_), .ZN(n5516) );
  OAI211_X1 U6122 ( .C1(n5610), .C2(n6475), .A(n5517), .B(n5516), .ZN(U2872)
         );
  AOI22_X1 U6123 ( .A1(n6683), .A2(DATAI_17_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n6686), .ZN(n5519) );
  NAND2_X1 U6124 ( .A1(n6687), .A2(DATAI_1_), .ZN(n5518) );
  OAI211_X1 U6125 ( .C1(n5618), .C2(n6475), .A(n5519), .B(n5518), .ZN(U2874)
         );
  INV_X1 U6126 ( .A(DATAI_15_), .ZN(n5903) );
  OAI222_X1 U6127 ( .A1(n5637), .A2(n6475), .B1(n5521), .B2(n5903), .C1(n5520), 
        .C2(n6008), .ZN(U2876) );
  INV_X1 U6128 ( .A(DATAI_14_), .ZN(n5900) );
  OAI222_X1 U6129 ( .A1(n5647), .A2(n6475), .B1(n5521), .B2(n5900), .C1(n5520), 
        .C2(n6003), .ZN(U2877) );
  AOI22_X1 U6130 ( .A1(n5531), .A2(n5522), .B1(n3851), .B2(n5676), .ZN(n5523)
         );
  XOR2_X1 U6131 ( .A(n5524), .B(n5523), .Z(n5673) );
  NOR2_X1 U6132 ( .A1(n6247), .A2(n5955), .ZN(n5668) );
  AOI21_X1 U6133 ( .B1(n6119), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5668), 
        .ZN(n5525) );
  OAI21_X1 U6134 ( .B1(n6125), .B2(n5526), .A(n5525), .ZN(n5527) );
  AOI21_X1 U6135 ( .B1(n5528), .B2(n6969), .A(n5527), .ZN(n5529) );
  OAI21_X1 U6136 ( .B1(n6397), .B2(n5673), .A(n5529), .ZN(U2957) );
  NAND2_X1 U6137 ( .A1(n5531), .A2(n5530), .ZN(n5533) );
  XNOR2_X1 U6138 ( .A(n5737), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5532)
         );
  XNOR2_X1 U6139 ( .A(n5533), .B(n5532), .ZN(n5683) );
  INV_X1 U6140 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6050) );
  NOR2_X1 U6141 ( .A1(n6247), .A2(n6050), .ZN(n5679) );
  AOI21_X1 U6142 ( .B1(n6119), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5679), 
        .ZN(n5534) );
  OAI21_X1 U6143 ( .B1(n6125), .B2(n5535), .A(n5534), .ZN(n5536) );
  AOI21_X1 U6144 ( .B1(n5537), .B2(n6969), .A(n5536), .ZN(n5538) );
  OAI21_X1 U6145 ( .B1(n5683), .B2(n6397), .A(n5538), .ZN(U2958) );
  NAND2_X1 U6146 ( .A1(n5541), .A2(n5693), .ZN(n5540) );
  MUX2_X1 U6147 ( .A(n5541), .B(n5540), .S(n5748), .Z(n5542) );
  INV_X1 U6148 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5677) );
  XNOR2_X1 U6149 ( .A(n5542), .B(n5677), .ZN(n5691) );
  INV_X1 U6150 ( .A(n5543), .ZN(n5547) );
  INV_X1 U6151 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6045) );
  NOR2_X1 U6152 ( .A1(n6247), .A2(n6045), .ZN(n5684) );
  AOI21_X1 U6153 ( .B1(n6119), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5684), 
        .ZN(n5544) );
  OAI21_X1 U6154 ( .B1(n6125), .B2(n5545), .A(n5544), .ZN(n5546) );
  AOI21_X1 U6155 ( .B1(n5547), .B2(n6969), .A(n5546), .ZN(n5548) );
  OAI21_X1 U6156 ( .B1(n6397), .B2(n5691), .A(n5548), .ZN(U2959) );
  XNOR2_X1 U6157 ( .A(n5737), .B(n5693), .ZN(n5549) );
  XNOR2_X1 U6158 ( .A(n5550), .B(n5549), .ZN(n5700) );
  NOR2_X1 U6159 ( .A1(n6247), .A2(n5868), .ZN(n5695) );
  AOI21_X1 U6160 ( .B1(n6119), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5695), 
        .ZN(n5551) );
  OAI21_X1 U6161 ( .B1(n6125), .B2(n5552), .A(n5551), .ZN(n5553) );
  AOI21_X1 U6162 ( .B1(n5554), .B2(n6969), .A(n5553), .ZN(n5555) );
  OAI21_X1 U6163 ( .B1(n6397), .B2(n5700), .A(n5555), .ZN(U2960) );
  OAI21_X1 U6164 ( .B1(n5558), .B2(n5557), .A(n5556), .ZN(n5708) );
  NOR2_X1 U6165 ( .A1(n6247), .A2(n6043), .ZN(n5701) );
  AOI21_X1 U6166 ( .B1(n6119), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n5701), 
        .ZN(n5561) );
  NAND2_X1 U6167 ( .A1(n6104), .A2(n5559), .ZN(n5560) );
  OAI211_X1 U6168 ( .C1(n5562), .C2(n6862), .A(n5561), .B(n5560), .ZN(n5563)
         );
  AOI21_X1 U6169 ( .B1(n6121), .B2(n5708), .A(n5563), .ZN(n5564) );
  INV_X1 U6170 ( .A(n5564), .ZN(U2961) );
  XNOR2_X1 U6171 ( .A(n3851), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5604)
         );
  INV_X1 U6172 ( .A(n5735), .ZN(n5568) );
  INV_X1 U6173 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5569) );
  NAND4_X1 U6174 ( .A1(n5568), .A2(n5748), .A3(n5567), .A4(n5569), .ZN(n5582)
         );
  NOR2_X1 U6175 ( .A1(n5737), .A2(n5569), .ZN(n5595) );
  XNOR2_X1 U6176 ( .A(n5748), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5597)
         );
  NOR3_X1 U6177 ( .A1(n5735), .A2(n5595), .A3(n5597), .ZN(n5571) );
  AOI21_X1 U6178 ( .B1(n5740), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5748), 
        .ZN(n5570) );
  NOR2_X1 U6179 ( .A1(n5571), .A2(n5570), .ZN(n5591) );
  NAND4_X1 U6180 ( .A1(n5591), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .A4(n5737), .ZN(n5572) );
  OAI21_X1 U6181 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5582), .A(n5572), 
        .ZN(n5573) );
  XNOR2_X1 U6182 ( .A(n5573), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5717)
         );
  NAND2_X1 U6183 ( .A1(n6104), .A2(n5574), .ZN(n5575) );
  NAND2_X1 U6184 ( .A1(n6235), .A2(REIP_REG_24__SCAN_IN), .ZN(n5710) );
  OAI211_X1 U6185 ( .C1(n5627), .C2(n5576), .A(n5575), .B(n5710), .ZN(n5577)
         );
  AOI21_X1 U6186 ( .B1(n6685), .B2(n6969), .A(n5577), .ZN(n5578) );
  OAI21_X1 U6187 ( .B1(n5717), .B2(n6397), .A(n5578), .ZN(U2962) );
  OR3_X1 U6188 ( .A1(n5580), .A2(n5748), .A3(n5579), .ZN(n5581) );
  NAND2_X1 U6189 ( .A1(n5582), .A2(n5581), .ZN(n5583) );
  XNOR2_X1 U6190 ( .A(n5583), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5718)
         );
  NOR2_X1 U6191 ( .A1(n6247), .A2(n6039), .ZN(n5719) );
  AOI21_X1 U6192 ( .B1(n6119), .B2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n5719), 
        .ZN(n5584) );
  OAI21_X1 U6193 ( .B1(n6125), .B2(n5585), .A(n5584), .ZN(n5586) );
  AOI21_X1 U6194 ( .B1(n5587), .B2(n6969), .A(n5586), .ZN(n5588) );
  OAI21_X1 U6195 ( .B1(n5718), .B2(n6397), .A(n5588), .ZN(U2963) );
  XNOR2_X1 U6196 ( .A(n5737), .B(n5589), .ZN(n5590) );
  XNOR2_X1 U6197 ( .A(n5591), .B(n5590), .ZN(n5733) );
  NAND2_X1 U6198 ( .A1(n5733), .A2(n6121), .ZN(n5594) );
  NOR2_X1 U6199 ( .A1(n6247), .A2(n6381), .ZN(n5727) );
  NOR2_X1 U6200 ( .A1(n6125), .A2(n6396), .ZN(n5592) );
  AOI211_X1 U6201 ( .C1(n6119), .C2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5727), 
        .B(n5592), .ZN(n5593) );
  OAI211_X1 U6202 ( .C1(n6862), .C2(n6391), .A(n5594), .B(n5593), .ZN(U2964)
         );
  OAI22_X1 U6203 ( .A1(n5735), .A2(n5595), .B1(n5748), .B2(n5740), .ZN(n5596)
         );
  XOR2_X1 U6204 ( .A(n5597), .B(n5596), .Z(n6245) );
  NAND2_X1 U6205 ( .A1(n6245), .A2(n6121), .ZN(n5602) );
  OAI22_X1 U6206 ( .A1(n5627), .A2(n5598), .B1(n6247), .B2(n6380), .ZN(n5599)
         );
  AOI21_X1 U6207 ( .B1(n6104), .B2(n5600), .A(n5599), .ZN(n5601) );
  OAI211_X1 U6208 ( .C1(n6862), .C2(n5603), .A(n5602), .B(n5601), .ZN(U2965)
         );
  OAI21_X1 U6209 ( .B1(n5566), .B2(n5604), .A(n5735), .ZN(n6157) );
  NAND2_X1 U6210 ( .A1(n6157), .A2(n6121), .ZN(n5609) );
  OAI22_X1 U6211 ( .A1(n5627), .A2(n5605), .B1(n6247), .B2(n6034), .ZN(n5606)
         );
  AOI21_X1 U6212 ( .B1(n6104), .B2(n5607), .A(n5606), .ZN(n5608) );
  OAI211_X1 U6213 ( .C1(n6862), .C2(n5610), .A(n5609), .B(n5608), .ZN(U2967)
         );
  INV_X1 U6214 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6240) );
  MUX2_X1 U6215 ( .A(n6240), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .S(n5737), 
        .Z(n5612) );
  NAND2_X1 U6216 ( .A1(n5746), .A2(n5619), .ZN(n5747) );
  XOR2_X1 U6217 ( .A(n5612), .B(n5747), .Z(n6237) );
  NAND2_X1 U6218 ( .A1(n6237), .A2(n6121), .ZN(n5617) );
  OAI22_X1 U6219 ( .A1(n5627), .A2(n5613), .B1(n6247), .B2(n6031), .ZN(n5614)
         );
  AOI21_X1 U6220 ( .B1(n6104), .B2(n5615), .A(n5614), .ZN(n5616) );
  OAI211_X1 U6221 ( .C1(n6862), .C2(n5618), .A(n5617), .B(n5616), .ZN(U2969)
         );
  INV_X1 U6222 ( .A(n5619), .ZN(n5621) );
  NOR2_X1 U6223 ( .A1(n5621), .A2(n5620), .ZN(n5624) );
  XOR2_X1 U6224 ( .A(n5624), .B(n5623), .Z(n6226) );
  INV_X1 U6225 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5625) );
  OAI22_X1 U6226 ( .A1(n5627), .A2(n5626), .B1(n6247), .B2(n5625), .ZN(n5630)
         );
  NOR2_X1 U6227 ( .A1(n5628), .A2(n6862), .ZN(n5629) );
  AOI211_X1 U6228 ( .C1(n6104), .C2(n6353), .A(n5630), .B(n5629), .ZN(n5631)
         );
  OAI21_X1 U6229 ( .B1(n6397), .B2(n6226), .A(n5631), .ZN(U2970) );
  INV_X1 U6230 ( .A(n5632), .ZN(n5634) );
  NAND2_X1 U6231 ( .A1(n5634), .A2(n5633), .ZN(n5635) );
  XNOR2_X1 U6232 ( .A(n5636), .B(n5635), .ZN(n6218) );
  INV_X1 U6233 ( .A(n6218), .ZN(n5643) );
  INV_X1 U6234 ( .A(n5637), .ZN(n5641) );
  AOI22_X1 U6235 ( .A1(n6119), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n6235), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n5638) );
  OAI21_X1 U6236 ( .B1(n6125), .B2(n5639), .A(n5638), .ZN(n5640) );
  AOI21_X1 U6237 ( .B1(n5641), .B2(n6969), .A(n5640), .ZN(n5642) );
  OAI21_X1 U6238 ( .B1(n5643), .B2(n6397), .A(n5642), .ZN(U2971) );
  XNOR2_X1 U6239 ( .A(n5737), .B(n5644), .ZN(n5645) );
  XNOR2_X1 U6240 ( .A(n5646), .B(n5645), .ZN(n6171) );
  INV_X1 U6241 ( .A(n5647), .ZN(n6342) );
  INV_X1 U6242 ( .A(n6341), .ZN(n5649) );
  AOI22_X1 U6243 ( .A1(n6119), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n6235), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n5648) );
  OAI21_X1 U6244 ( .B1(n6125), .B2(n5649), .A(n5648), .ZN(n5650) );
  AOI21_X1 U6245 ( .B1(n6342), .B2(n6969), .A(n5650), .ZN(n5651) );
  OAI21_X1 U6246 ( .B1(n6171), .B2(n6397), .A(n5651), .ZN(U2972) );
  INV_X1 U6247 ( .A(n5652), .ZN(n5663) );
  INV_X1 U6248 ( .A(n5653), .ZN(n5661) );
  INV_X1 U6249 ( .A(n5654), .ZN(n5655) );
  AOI21_X1 U6250 ( .B1(n5656), .B2(n5655), .A(INSTADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n5657) );
  AOI211_X1 U6251 ( .C1(n5664), .C2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5658), .B(n5657), .ZN(n5659) );
  AOI211_X1 U6252 ( .C1(n6243), .C2(n5661), .A(n5660), .B(n5659), .ZN(n5662)
         );
  OAI21_X1 U6253 ( .B1(n5663), .B2(n6225), .A(n5662), .ZN(U2988) );
  INV_X1 U6254 ( .A(n5664), .ZN(n5671) );
  OAI21_X1 U6255 ( .B1(n5687), .B2(n5666), .A(n5665), .ZN(n5670) );
  NOR2_X1 U6256 ( .A1(n5667), .A2(n6224), .ZN(n5669) );
  AOI211_X1 U6257 ( .C1(n5671), .C2(n5670), .A(n5669), .B(n5668), .ZN(n5672)
         );
  OAI21_X1 U6258 ( .B1(n5673), .B2(n6225), .A(n5672), .ZN(U2989) );
  INV_X1 U6259 ( .A(n5674), .ZN(n5680) );
  AOI211_X1 U6260 ( .C1(n5677), .C2(n5676), .A(n5675), .B(n5687), .ZN(n5678)
         );
  AOI211_X1 U6261 ( .C1(n6243), .C2(n5680), .A(n5679), .B(n5678), .ZN(n5682)
         );
  NAND2_X1 U6262 ( .A1(n5689), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5681) );
  OAI211_X1 U6263 ( .C1(n5683), .C2(n6225), .A(n5682), .B(n5681), .ZN(U2990)
         );
  AOI21_X1 U6264 ( .B1(n5685), .B2(n6243), .A(n5684), .ZN(n5686) );
  OAI21_X1 U6265 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5687), .A(n5686), 
        .ZN(n5688) );
  AOI21_X1 U6266 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5689), .A(n5688), 
        .ZN(n5690) );
  OAI21_X1 U6267 ( .B1(n5691), .B2(n6225), .A(n5690), .ZN(U2991) );
  AOI211_X1 U6268 ( .C1(n5693), .C2(n5706), .A(n5692), .B(n5703), .ZN(n5694)
         );
  AOI211_X1 U6269 ( .C1(n6243), .C2(n5696), .A(n5695), .B(n5694), .ZN(n5699)
         );
  NAND2_X1 U6270 ( .A1(n5697), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5698) );
  OAI211_X1 U6271 ( .C1(n5700), .C2(n6225), .A(n5699), .B(n5698), .ZN(U2992)
         );
  AOI21_X1 U6272 ( .B1(n5702), .B2(n6243), .A(n5701), .ZN(n5705) );
  OR2_X1 U6273 ( .A1(n5703), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5704)
         );
  OAI211_X1 U6274 ( .C1(n5711), .C2(n5706), .A(n5705), .B(n5704), .ZN(n5707)
         );
  AOI21_X1 U6275 ( .B1(n5708), .B2(n6244), .A(n5707), .ZN(n5709) );
  INV_X1 U6276 ( .A(n5709), .ZN(U2993) );
  INV_X1 U6277 ( .A(n5710), .ZN(n5715) );
  AOI211_X1 U6278 ( .C1(n5713), .C2(n5721), .A(n5712), .B(n5711), .ZN(n5714)
         );
  AOI211_X1 U6279 ( .C1(n6243), .C2(n6081), .A(n5715), .B(n5714), .ZN(n5716)
         );
  OAI21_X1 U6280 ( .B1(n5717), .B2(n6225), .A(n5716), .ZN(U2994) );
  OR2_X1 U6281 ( .A1(n5718), .A2(n6225), .ZN(n5725) );
  AOI21_X1 U6282 ( .B1(n5720), .B2(n6243), .A(n5719), .ZN(n5724) );
  NAND2_X1 U6283 ( .A1(n5726), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5723) );
  OR2_X1 U6284 ( .A1(n5721), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5722)
         );
  NAND4_X1 U6285 ( .A1(n5725), .A2(n5724), .A3(n5723), .A4(n5722), .ZN(U2995)
         );
  INV_X1 U6286 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6250) );
  NAND2_X1 U6287 ( .A1(n5726), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5730) );
  INV_X1 U6288 ( .A(n6388), .ZN(n5728) );
  AOI21_X1 U6289 ( .B1(n5728), .B2(n6243), .A(n5727), .ZN(n5729) );
  OAI211_X1 U6290 ( .C1(n5731), .C2(n6250), .A(n5730), .B(n5729), .ZN(n5732)
         );
  AOI21_X1 U6291 ( .B1(n5733), .B2(n6244), .A(n5732), .ZN(n5734) );
  INV_X1 U6292 ( .A(n5734), .ZN(U2996) );
  NAND2_X1 U6293 ( .A1(n3851), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5736) );
  MUX2_X1 U6294 ( .A(n5737), .B(n5736), .S(n5735), .Z(n5738) );
  XNOR2_X1 U6295 ( .A(n5738), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6122)
         );
  NAND2_X1 U6296 ( .A1(n6155), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5743) );
  NOR3_X1 U6297 ( .A1(n5740), .A2(n5739), .A3(n6160), .ZN(n5741) );
  AOI21_X1 U6298 ( .B1(n6235), .B2(REIP_REG_20__SCAN_IN), .A(n5741), .ZN(n5742) );
  OAI211_X1 U6299 ( .C1(n6224), .C2(n6377), .A(n5743), .B(n5742), .ZN(n5744)
         );
  AOI21_X1 U6300 ( .B1(n6122), .B2(n6244), .A(n5744), .ZN(n5745) );
  INV_X1 U6301 ( .A(n5745), .ZN(U2998) );
  NOR2_X1 U6302 ( .A1(n5746), .A2(n6240), .ZN(n5750) );
  NOR2_X1 U6303 ( .A1(n5747), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5749)
         );
  MUX2_X1 U6304 ( .A(n5750), .B(n5749), .S(n5748), .Z(n5752) );
  XNOR2_X1 U6305 ( .A(n5752), .B(n5751), .ZN(n6116) );
  INV_X1 U6306 ( .A(n6116), .ZN(n5762) );
  INV_X1 U6307 ( .A(n5758), .ZN(n6232) );
  AOI21_X1 U6308 ( .B1(n6232), .B2(n6214), .A(n6213), .ZN(n6241) );
  OAI21_X1 U6309 ( .B1(n6162), .B2(n5753), .A(n6240), .ZN(n5754) );
  OAI211_X1 U6310 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n6179), .A(n6241), .B(n5754), .ZN(n5757) );
  INV_X1 U6311 ( .A(REIP_REG_18__SCAN_IN), .ZN(n5755) );
  OAI22_X1 U6312 ( .A1(n6367), .A2(n6224), .B1(n6247), .B2(n5755), .ZN(n5756)
         );
  AOI21_X1 U6313 ( .B1(n5757), .B2(INSTADDRPOINTER_REG_18__SCAN_IN), .A(n5756), 
        .ZN(n5761) );
  NOR3_X1 U6314 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n6215), .A3(n6240), 
        .ZN(n5759) );
  NAND2_X1 U6315 ( .A1(n5759), .A2(n5758), .ZN(n5760) );
  OAI211_X1 U6316 ( .C1(n5762), .C2(n6225), .A(n5761), .B(n5760), .ZN(U3000)
         );
  AOI21_X1 U6317 ( .B1(n5765), .B2(n5764), .A(n5763), .ZN(n5766) );
  INV_X1 U6318 ( .A(n5766), .ZN(n5773) );
  NOR2_X1 U6319 ( .A1(n6224), .A2(n5767), .ZN(n5768) );
  AOI211_X1 U6320 ( .C1(n5770), .C2(n6244), .A(n5769), .B(n5768), .ZN(n5772)
         );
  NAND3_X1 U6321 ( .A1(n5773), .A2(n5772), .A3(n5771), .ZN(U3018) );
  INV_X1 U6322 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6066) );
  NOR2_X1 U6323 ( .A1(n6140), .A2(STATE_REG_0__SCAN_IN), .ZN(n6474) );
  INV_X1 U6324 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6138) );
  AOI21_X1 U6325 ( .B1(n6138), .B2(STATE_REG_1__SCAN_IN), .A(n6463), .ZN(n5778) );
  NOR2_X1 U6326 ( .A1(n6474), .A2(n5778), .ZN(n6456) );
  INV_X1 U6327 ( .A(n6456), .ZN(n5775) );
  INV_X1 U6328 ( .A(BS16_N), .ZN(n5774) );
  NAND2_X1 U6329 ( .A1(n6138), .A2(n6463), .ZN(n6130) );
  AOI21_X1 U6330 ( .B1(n5774), .B2(n6130), .A(n5775), .ZN(n6453) );
  AOI21_X1 U6331 ( .B1(n6066), .B2(n5775), .A(n6453), .ZN(U3451) );
  AND2_X1 U6332 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n5775), .ZN(U3180) );
  AND2_X1 U6333 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n5775), .ZN(U3179) );
  AND2_X1 U6334 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n5775), .ZN(U3178) );
  AND2_X1 U6335 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n5775), .ZN(U3177) );
  AND2_X1 U6336 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n5775), .ZN(U3176) );
  AND2_X1 U6337 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n5775), .ZN(U3175) );
  AND2_X1 U6338 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n5775), .ZN(U3174) );
  AND2_X1 U6339 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n5775), .ZN(U3173) );
  AND2_X1 U6340 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n5775), .ZN(U3172) );
  AND2_X1 U6341 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n5775), .ZN(U3171) );
  AND2_X1 U6342 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n5775), .ZN(U3170) );
  AND2_X1 U6343 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n5775), .ZN(U3169) );
  AND2_X1 U6344 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n5775), .ZN(U3168) );
  AND2_X1 U6345 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n5775), .ZN(U3167) );
  AND2_X1 U6346 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n5775), .ZN(U3166) );
  AND2_X1 U6347 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n5775), .ZN(U3165) );
  AND2_X1 U6348 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n5775), .ZN(U3164) );
  AND2_X1 U6349 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n5775), .ZN(U3163) );
  AND2_X1 U6350 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n5775), .ZN(U3162) );
  AND2_X1 U6351 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n5775), .ZN(U3161) );
  AND2_X1 U6352 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n5775), .ZN(U3160) );
  AND2_X1 U6353 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n5775), .ZN(U3159) );
  AND2_X1 U6354 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n5775), .ZN(U3158) );
  AND2_X1 U6355 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n5775), .ZN(U3157) );
  AND2_X1 U6356 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n5775), .ZN(U3156) );
  AND2_X1 U6357 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n5775), .ZN(U3155) );
  AND2_X1 U6358 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n5775), .ZN(U3154) );
  AND2_X1 U6359 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n5775), .ZN(U3153) );
  AND2_X1 U6360 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n5775), .ZN(U3152) );
  AND2_X1 U6361 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n5775), .ZN(U3151) );
  AND2_X1 U6362 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n5776), .ZN(U3019)
         );
  AND2_X1 U6363 ( .A1(n5777), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U6364 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5935) );
  AOI21_X1 U6365 ( .B1(n5778), .B2(n5935), .A(n6474), .ZN(U2789) );
  INV_X1 U6366 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6034) );
  INV_X1 U6367 ( .A(keyinput_62), .ZN(n5865) );
  INV_X1 U6368 ( .A(REIP_REG_20__SCAN_IN), .ZN(n5968) );
  AOI22_X1 U6369 ( .A1(REIP_REG_22__SCAN_IN), .A2(keyinput_60), .B1(
        REIP_REG_23__SCAN_IN), .B2(keyinput_59), .ZN(n5779) );
  OAI221_X1 U6370 ( .B1(REIP_REG_22__SCAN_IN), .B2(keyinput_60), .C1(
        REIP_REG_23__SCAN_IN), .C2(keyinput_59), .A(n5779), .ZN(n5862) );
  INV_X1 U6371 ( .A(keyinput_58), .ZN(n5860) );
  AOI22_X1 U6372 ( .A1(REIP_REG_26__SCAN_IN), .A2(keyinput_56), .B1(n6045), 
        .B2(keyinput_55), .ZN(n5780) );
  OAI221_X1 U6373 ( .B1(REIP_REG_26__SCAN_IN), .B2(keyinput_56), .C1(n6045), 
        .C2(keyinput_55), .A(n5780), .ZN(n5857) );
  INV_X1 U6374 ( .A(keyinput_54), .ZN(n5855) );
  INV_X1 U6375 ( .A(keyinput_53), .ZN(n5853) );
  INV_X1 U6376 ( .A(keyinput_52), .ZN(n5851) );
  INV_X1 U6377 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6136) );
  OAI22_X1 U6378 ( .A1(n6136), .A2(keyinput_46), .B1(BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_49), .ZN(n5781) );
  AOI221_X1 U6379 ( .B1(n6136), .B2(keyinput_46), .C1(keyinput_49), .C2(
        BYTEENABLE_REG_2__SCAN_IN), .A(n5781), .ZN(n5844) );
  INV_X1 U6380 ( .A(keyinput_42), .ZN(n5838) );
  INV_X1 U6381 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6139) );
  INV_X1 U6382 ( .A(keyinput_41), .ZN(n5836) );
  INV_X1 U6383 ( .A(D_C_N_REG_SCAN_IN), .ZN(n6129) );
  INV_X1 U6384 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n6472) );
  INV_X1 U6385 ( .A(keyinput_40), .ZN(n5834) );
  INV_X1 U6386 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6127) );
  INV_X1 U6387 ( .A(keyinput_39), .ZN(n5832) );
  INV_X1 U6388 ( .A(keyinput_38), .ZN(n5830) );
  INV_X1 U6389 ( .A(HOLD), .ZN(n6137) );
  OAI22_X1 U6390 ( .A1(n6137), .A2(keyinput_36), .B1(keyinput_37), .B2(
        READREQUEST_REG_SCAN_IN), .ZN(n5782) );
  AOI221_X1 U6391 ( .B1(n6137), .B2(keyinput_36), .C1(READREQUEST_REG_SCAN_IN), 
        .C2(keyinput_37), .A(n5782), .ZN(n5827) );
  OAI22_X1 U6392 ( .A1(n5876), .A2(keyinput_23), .B1(n6907), .B2(keyinput_25), 
        .ZN(n5783) );
  AOI221_X1 U6393 ( .B1(n5876), .B2(keyinput_23), .C1(keyinput_25), .C2(n6907), 
        .A(n5783), .ZN(n5819) );
  OAI22_X1 U6394 ( .A1(n5910), .A2(keyinput_19), .B1(n5909), .B2(keyinput_20), 
        .ZN(n5784) );
  AOI221_X1 U6395 ( .B1(n5910), .B2(keyinput_19), .C1(keyinput_20), .C2(n5909), 
        .A(n5784), .ZN(n5810) );
  INV_X1 U6396 ( .A(DATAI_21_), .ZN(n6861) );
  AOI22_X1 U6397 ( .A1(DATAI_24_), .A2(keyinput_7), .B1(n6861), .B2(
        keyinput_10), .ZN(n5785) );
  OAI221_X1 U6398 ( .B1(DATAI_24_), .B2(keyinput_7), .C1(n6861), .C2(
        keyinput_10), .A(n5785), .ZN(n5797) );
  INV_X1 U6399 ( .A(DATAI_25_), .ZN(n6692) );
  AOI22_X1 U6400 ( .A1(DATAI_26_), .A2(keyinput_5), .B1(n6692), .B2(keyinput_6), .ZN(n5786) );
  OAI221_X1 U6401 ( .B1(DATAI_26_), .B2(keyinput_5), .C1(n6692), .C2(
        keyinput_6), .A(n5786), .ZN(n5795) );
  INV_X1 U6402 ( .A(DATAI_27_), .ZN(n6781) );
  OAI22_X1 U6403 ( .A1(n6781), .A2(keyinput_4), .B1(keyinput_3), .B2(DATAI_28_), .ZN(n5787) );
  AOI221_X1 U6404 ( .B1(n6781), .B2(keyinput_4), .C1(DATAI_28_), .C2(
        keyinput_3), .A(n5787), .ZN(n5794) );
  INV_X1 U6405 ( .A(keyinput_2), .ZN(n5790) );
  INV_X1 U6406 ( .A(DATAI_29_), .ZN(n5888) );
  AOI22_X1 U6407 ( .A1(DATAI_30_), .A2(keyinput_1), .B1(DATAI_31_), .B2(
        keyinput_0), .ZN(n5788) );
  OAI221_X1 U6408 ( .B1(DATAI_30_), .B2(keyinput_1), .C1(DATAI_31_), .C2(
        keyinput_0), .A(n5788), .ZN(n5789) );
  OAI221_X1 U6409 ( .B1(DATAI_29_), .B2(n5790), .C1(n5888), .C2(keyinput_2), 
        .A(n5789), .ZN(n5793) );
  OAI22_X1 U6410 ( .A1(DATAI_23_), .A2(keyinput_8), .B1(keyinput_9), .B2(
        DATAI_22_), .ZN(n5791) );
  AOI221_X1 U6411 ( .B1(DATAI_23_), .B2(keyinput_8), .C1(DATAI_22_), .C2(
        keyinput_9), .A(n5791), .ZN(n5792) );
  OAI221_X1 U6412 ( .B1(n5795), .B2(n5794), .C1(n5795), .C2(n5793), .A(n5792), 
        .ZN(n5796) );
  OAI22_X1 U6413 ( .A1(n5797), .A2(n5796), .B1(DATAI_20_), .B2(keyinput_11), 
        .ZN(n5798) );
  AOI21_X1 U6414 ( .B1(DATAI_20_), .B2(keyinput_11), .A(n5798), .ZN(n5804) );
  INV_X1 U6415 ( .A(DATAI_19_), .ZN(n5800) );
  OAI22_X1 U6416 ( .A1(n5800), .A2(keyinput_12), .B1(keyinput_13), .B2(
        DATAI_18_), .ZN(n5799) );
  AOI221_X1 U6417 ( .B1(n5800), .B2(keyinput_12), .C1(DATAI_18_), .C2(
        keyinput_13), .A(n5799), .ZN(n5803) );
  INV_X1 U6418 ( .A(DATAI_17_), .ZN(n5878) );
  AOI22_X1 U6419 ( .A1(DATAI_16_), .A2(keyinput_15), .B1(n5878), .B2(
        keyinput_14), .ZN(n5801) );
  OAI221_X1 U6420 ( .B1(DATAI_16_), .B2(keyinput_15), .C1(n5878), .C2(
        keyinput_14), .A(n5801), .ZN(n5802) );
  AOI21_X1 U6421 ( .B1(n5804), .B2(n5803), .A(n5802), .ZN(n5807) );
  AOI22_X1 U6422 ( .A1(DATAI_14_), .A2(keyinput_17), .B1(n5902), .B2(
        keyinput_18), .ZN(n5805) );
  OAI221_X1 U6423 ( .B1(DATAI_14_), .B2(keyinput_17), .C1(n5902), .C2(
        keyinput_18), .A(n5805), .ZN(n5806) );
  AOI211_X1 U6424 ( .C1(DATAI_15_), .C2(keyinput_16), .A(n5807), .B(n5806), 
        .ZN(n5808) );
  OAI21_X1 U6425 ( .B1(DATAI_15_), .B2(keyinput_16), .A(n5808), .ZN(n5809) );
  AOI22_X1 U6426 ( .A1(DATAI_10_), .A2(keyinput_21), .B1(n5810), .B2(n5809), 
        .ZN(n5813) );
  AOI22_X1 U6427 ( .A1(DATAI_7_), .A2(keyinput_24), .B1(DATAI_9_), .B2(
        keyinput_22), .ZN(n5811) );
  OAI221_X1 U6428 ( .B1(DATAI_7_), .B2(keyinput_24), .C1(DATAI_9_), .C2(
        keyinput_22), .A(n5811), .ZN(n5812) );
  AOI221_X1 U6429 ( .B1(DATAI_10_), .B2(n5813), .C1(keyinput_21), .C2(n5813), 
        .A(n5812), .ZN(n5818) );
  AOI22_X1 U6430 ( .A1(n6731), .A2(keyinput_29), .B1(n6779), .B2(keyinput_28), 
        .ZN(n5814) );
  OAI221_X1 U6431 ( .B1(n6731), .B2(keyinput_29), .C1(n6779), .C2(keyinput_28), 
        .A(n5814), .ZN(n5817) );
  AOI22_X1 U6432 ( .A1(DATAI_4_), .A2(keyinput_27), .B1(DATAI_5_), .B2(
        keyinput_26), .ZN(n5815) );
  OAI221_X1 U6433 ( .B1(DATAI_4_), .B2(keyinput_27), .C1(DATAI_5_), .C2(
        keyinput_26), .A(n5815), .ZN(n5816) );
  AOI211_X1 U6434 ( .C1(n5819), .C2(n5818), .A(n5817), .B(n5816), .ZN(n5825)
         );
  XOR2_X1 U6435 ( .A(n6690), .B(keyinput_30), .Z(n5824) );
  INV_X1 U6436 ( .A(NA_N), .ZN(n6465) );
  OAI22_X1 U6437 ( .A1(n6465), .A2(keyinput_33), .B1(keyinput_32), .B2(
        MEMORYFETCH_REG_SCAN_IN), .ZN(n5820) );
  AOI221_X1 U6438 ( .B1(n6465), .B2(keyinput_33), .C1(MEMORYFETCH_REG_SCAN_IN), 
        .C2(keyinput_32), .A(n5820), .ZN(n5823) );
  OAI22_X1 U6439 ( .A1(DATAI_0_), .A2(keyinput_31), .B1(keyinput_34), .B2(
        BS16_N), .ZN(n5821) );
  AOI221_X1 U6440 ( .B1(DATAI_0_), .B2(keyinput_31), .C1(BS16_N), .C2(
        keyinput_34), .A(n5821), .ZN(n5822) );
  OAI211_X1 U6441 ( .C1(n5825), .C2(n5824), .A(n5823), .B(n5822), .ZN(n5826)
         );
  OAI211_X1 U6442 ( .C1(READY_N), .C2(keyinput_35), .A(n5827), .B(n5826), .ZN(
        n5828) );
  AOI21_X1 U6443 ( .B1(READY_N), .B2(keyinput_35), .A(n5828), .ZN(n5829) );
  AOI221_X1 U6444 ( .B1(ADS_N_REG_SCAN_IN), .B2(n5830), .C1(n5935), .C2(
        keyinput_38), .A(n5829), .ZN(n5831) );
  AOI221_X1 U6445 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(keyinput_39), .C1(n6127), 
        .C2(n5832), .A(n5831), .ZN(n5833) );
  AOI221_X1 U6446 ( .B1(M_IO_N_REG_SCAN_IN), .B2(keyinput_40), .C1(n6472), 
        .C2(n5834), .A(n5833), .ZN(n5835) );
  AOI221_X1 U6447 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5836), .C1(n6129), .C2(
        keyinput_41), .A(n5835), .ZN(n5837) );
  AOI221_X1 U6448 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(n5838), .C1(n6139), 
        .C2(keyinput_42), .A(n5837), .ZN(n5841) );
  AOI22_X1 U6449 ( .A1(MORE_REG_SCAN_IN), .A2(keyinput_44), .B1(n6398), .B2(
        keyinput_45), .ZN(n5839) );
  OAI221_X1 U6450 ( .B1(MORE_REG_SCAN_IN), .B2(keyinput_44), .C1(n6398), .C2(
        keyinput_45), .A(n5839), .ZN(n5840) );
  AOI211_X1 U6451 ( .C1(STATEBS16_REG_SCAN_IN), .C2(keyinput_43), .A(n5841), 
        .B(n5840), .ZN(n5842) );
  OAI21_X1 U6452 ( .B1(STATEBS16_REG_SCAN_IN), .B2(keyinput_43), .A(n5842), 
        .ZN(n5843) );
  OAI211_X1 U6453 ( .C1(BYTEENABLE_REG_1__SCAN_IN), .C2(keyinput_48), .A(n5844), .B(n5843), .ZN(n5845) );
  AOI21_X1 U6454 ( .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_48), .A(n5845), 
        .ZN(n5849) );
  INV_X1 U6455 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6074) );
  OAI22_X1 U6456 ( .A1(n6074), .A2(keyinput_47), .B1(keyinput_50), .B2(
        BYTEENABLE_REG_3__SCAN_IN), .ZN(n5846) );
  AOI221_X1 U6457 ( .B1(n6074), .B2(keyinput_47), .C1(
        BYTEENABLE_REG_3__SCAN_IN), .C2(keyinput_50), .A(n5846), .ZN(n5848) );
  NOR2_X1 U6458 ( .A1(REIP_REG_31__SCAN_IN), .A2(keyinput_51), .ZN(n5847) );
  AOI221_X1 U6459 ( .B1(n5849), .B2(n5848), .C1(keyinput_51), .C2(
        REIP_REG_31__SCAN_IN), .A(n5847), .ZN(n5850) );
  AOI221_X1 U6460 ( .B1(REIP_REG_30__SCAN_IN), .B2(keyinput_52), .C1(n5951), 
        .C2(n5851), .A(n5850), .ZN(n5852) );
  AOI221_X1 U6461 ( .B1(REIP_REG_29__SCAN_IN), .B2(keyinput_53), .C1(n5955), 
        .C2(n5853), .A(n5852), .ZN(n5854) );
  AOI221_X1 U6462 ( .B1(REIP_REG_28__SCAN_IN), .B2(n5855), .C1(n6050), .C2(
        keyinput_54), .A(n5854), .ZN(n5856) );
  OAI22_X1 U6463 ( .A1(n5857), .A2(n5856), .B1(keyinput_57), .B2(
        REIP_REG_25__SCAN_IN), .ZN(n5858) );
  AOI21_X1 U6464 ( .B1(keyinput_57), .B2(REIP_REG_25__SCAN_IN), .A(n5858), 
        .ZN(n5859) );
  AOI221_X1 U6465 ( .B1(REIP_REG_24__SCAN_IN), .B2(n5860), .C1(n6041), .C2(
        keyinput_58), .A(n5859), .ZN(n5861) );
  OAI22_X1 U6466 ( .A1(keyinput_61), .A2(n6380), .B1(n5862), .B2(n5861), .ZN(
        n5863) );
  AOI21_X1 U6467 ( .B1(keyinput_61), .B2(n6380), .A(n5863), .ZN(n5864) );
  AOI221_X1 U6468 ( .B1(REIP_REG_20__SCAN_IN), .B2(n5865), .C1(n5968), .C2(
        keyinput_62), .A(n5864), .ZN(n5973) );
  INV_X1 U6469 ( .A(keyinput_127), .ZN(n5970) );
  INV_X1 U6470 ( .A(keyinput_126), .ZN(n5967) );
  OAI22_X1 U6471 ( .A1(n6381), .A2(keyinput_124), .B1(REIP_REG_23__SCAN_IN), 
        .B2(keyinput_123), .ZN(n5866) );
  AOI221_X1 U6472 ( .B1(n6381), .B2(keyinput_124), .C1(keyinput_123), .C2(
        REIP_REG_23__SCAN_IN), .A(n5866), .ZN(n5964) );
  INV_X1 U6473 ( .A(keyinput_122), .ZN(n5962) );
  AOI22_X1 U6474 ( .A1(n5868), .A2(keyinput_120), .B1(n6045), .B2(keyinput_119), .ZN(n5867) );
  OAI221_X1 U6475 ( .B1(n5868), .B2(keyinput_120), .C1(n6045), .C2(
        keyinput_119), .A(n5867), .ZN(n5960) );
  INV_X1 U6476 ( .A(keyinput_118), .ZN(n5957) );
  INV_X1 U6477 ( .A(keyinput_117), .ZN(n5954) );
  INV_X1 U6478 ( .A(keyinput_116), .ZN(n5952) );
  AOI22_X1 U6479 ( .A1(keyinput_113), .A2(BYTEENABLE_REG_2__SCAN_IN), .B1(
        n6074), .B2(keyinput_111), .ZN(n5869) );
  OAI221_X1 U6480 ( .B1(keyinput_113), .B2(BYTEENABLE_REG_2__SCAN_IN), .C1(
        n6074), .C2(keyinput_111), .A(n5869), .ZN(n5872) );
  AOI22_X1 U6481 ( .A1(BYTEENABLE_REG_1__SCAN_IN), .A2(keyinput_112), .B1(
        n6136), .B2(keyinput_110), .ZN(n5870) );
  OAI221_X1 U6482 ( .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_112), .C1(
        n6136), .C2(keyinput_110), .A(n5870), .ZN(n5871) );
  AOI211_X1 U6483 ( .C1(keyinput_114), .C2(BYTEENABLE_REG_3__SCAN_IN), .A(
        n5872), .B(n5871), .ZN(n5873) );
  OAI21_X1 U6484 ( .B1(keyinput_114), .B2(BYTEENABLE_REG_3__SCAN_IN), .A(n5873), .ZN(n5948) );
  OAI22_X1 U6485 ( .A1(n6398), .A2(keyinput_109), .B1(keyinput_108), .B2(
        MORE_REG_SCAN_IN), .ZN(n5874) );
  AOI221_X1 U6486 ( .B1(n6398), .B2(keyinput_109), .C1(MORE_REG_SCAN_IN), .C2(
        keyinput_108), .A(n5874), .ZN(n5945) );
  INV_X1 U6487 ( .A(keyinput_106), .ZN(n5943) );
  INV_X1 U6488 ( .A(keyinput_105), .ZN(n5941) );
  INV_X1 U6489 ( .A(keyinput_104), .ZN(n5939) );
  INV_X1 U6490 ( .A(keyinput_103), .ZN(n5937) );
  INV_X1 U6491 ( .A(keyinput_102), .ZN(n5934) );
  XOR2_X1 U6492 ( .A(n6690), .B(keyinput_94), .Z(n5928) );
  AOI22_X1 U6493 ( .A1(n6907), .A2(keyinput_89), .B1(n5876), .B2(keyinput_87), 
        .ZN(n5875) );
  OAI221_X1 U6494 ( .B1(n6907), .B2(keyinput_89), .C1(n5876), .C2(keyinput_87), 
        .A(n5875), .ZN(n5922) );
  OAI22_X1 U6495 ( .A1(n5878), .A2(keyinput_78), .B1(DATAI_16_), .B2(
        keyinput_79), .ZN(n5877) );
  AOI221_X1 U6496 ( .B1(n5878), .B2(keyinput_78), .C1(keyinput_79), .C2(
        DATAI_16_), .A(n5877), .ZN(n5907) );
  INV_X1 U6497 ( .A(DATAI_22_), .ZN(n5881) );
  INV_X1 U6498 ( .A(DATAI_24_), .ZN(n5880) );
  AOI22_X1 U6499 ( .A1(n5881), .A2(keyinput_73), .B1(n5880), .B2(keyinput_71), 
        .ZN(n5879) );
  OAI221_X1 U6500 ( .B1(n5881), .B2(keyinput_73), .C1(n5880), .C2(keyinput_71), 
        .A(n5879), .ZN(n5899) );
  INV_X1 U6501 ( .A(DATAI_26_), .ZN(n5883) );
  AOI22_X1 U6502 ( .A1(n6692), .A2(keyinput_70), .B1(n5883), .B2(keyinput_69), 
        .ZN(n5882) );
  OAI221_X1 U6503 ( .B1(n6692), .B2(keyinput_70), .C1(n5883), .C2(keyinput_69), 
        .A(n5882), .ZN(n5893) );
  OAI22_X1 U6504 ( .A1(n6781), .A2(keyinput_68), .B1(DATAI_28_), .B2(
        keyinput_67), .ZN(n5884) );
  AOI221_X1 U6505 ( .B1(n6781), .B2(keyinput_68), .C1(keyinput_67), .C2(
        DATAI_28_), .A(n5884), .ZN(n5892) );
  INV_X1 U6506 ( .A(keyinput_66), .ZN(n5887) );
  AOI22_X1 U6507 ( .A1(DATAI_30_), .A2(keyinput_65), .B1(DATAI_31_), .B2(
        keyinput_64), .ZN(n5885) );
  OAI221_X1 U6508 ( .B1(DATAI_30_), .B2(keyinput_65), .C1(DATAI_31_), .C2(
        keyinput_64), .A(n5885), .ZN(n5886) );
  OAI221_X1 U6509 ( .B1(DATAI_29_), .B2(keyinput_66), .C1(n5888), .C2(n5887), 
        .A(n5886), .ZN(n5891) );
  OAI22_X1 U6510 ( .A1(n6861), .A2(keyinput_74), .B1(DATAI_23_), .B2(
        keyinput_72), .ZN(n5889) );
  AOI221_X1 U6511 ( .B1(n6861), .B2(keyinput_74), .C1(keyinput_72), .C2(
        DATAI_23_), .A(n5889), .ZN(n5890) );
  OAI221_X1 U6512 ( .B1(n5893), .B2(n5892), .C1(n5893), .C2(n5891), .A(n5890), 
        .ZN(n5898) );
  INV_X1 U6513 ( .A(DATAI_20_), .ZN(n5895) );
  OAI22_X1 U6514 ( .A1(n5895), .A2(keyinput_75), .B1(DATAI_19_), .B2(
        keyinput_76), .ZN(n5894) );
  AOI221_X1 U6515 ( .B1(n5895), .B2(keyinput_75), .C1(keyinput_76), .C2(
        DATAI_19_), .A(n5894), .ZN(n5897) );
  XNOR2_X1 U6516 ( .A(DATAI_18_), .B(keyinput_77), .ZN(n5896) );
  OAI211_X1 U6517 ( .C1(n5899), .C2(n5898), .A(n5897), .B(n5896), .ZN(n5906)
         );
  XOR2_X1 U6518 ( .A(n5900), .B(keyinput_81), .Z(n5905) );
  AOI22_X1 U6519 ( .A1(n5903), .A2(keyinput_80), .B1(n5902), .B2(keyinput_82), 
        .ZN(n5901) );
  OAI221_X1 U6520 ( .B1(n5903), .B2(keyinput_80), .C1(n5902), .C2(keyinput_82), 
        .A(n5901), .ZN(n5904) );
  AOI211_X1 U6521 ( .C1(n5907), .C2(n5906), .A(n5905), .B(n5904), .ZN(n5912)
         );
  AOI22_X1 U6522 ( .A1(n5910), .A2(keyinput_83), .B1(keyinput_84), .B2(n5909), 
        .ZN(n5908) );
  OAI221_X1 U6523 ( .B1(n5910), .B2(keyinput_83), .C1(n5909), .C2(keyinput_84), 
        .A(n5908), .ZN(n5911) );
  OAI22_X1 U6524 ( .A1(n5912), .A2(n5911), .B1(keyinput_85), .B2(n5915), .ZN(
        n5916) );
  OAI22_X1 U6525 ( .A1(DATAI_9_), .A2(keyinput_86), .B1(keyinput_88), .B2(
        DATAI_7_), .ZN(n5913) );
  AOI221_X1 U6526 ( .B1(DATAI_9_), .B2(keyinput_86), .C1(DATAI_7_), .C2(
        keyinput_88), .A(n5913), .ZN(n5914) );
  OAI221_X1 U6527 ( .B1(n5916), .B2(keyinput_85), .C1(n5916), .C2(n5915), .A(
        n5914), .ZN(n5921) );
  OAI22_X1 U6528 ( .A1(n6821), .A2(keyinput_91), .B1(keyinput_92), .B2(
        DATAI_3_), .ZN(n5917) );
  AOI221_X1 U6529 ( .B1(n6821), .B2(keyinput_91), .C1(DATAI_3_), .C2(
        keyinput_92), .A(n5917), .ZN(n5920) );
  OAI22_X1 U6530 ( .A1(DATAI_5_), .A2(keyinput_90), .B1(DATAI_2_), .B2(
        keyinput_93), .ZN(n5918) );
  AOI221_X1 U6531 ( .B1(DATAI_5_), .B2(keyinput_90), .C1(keyinput_93), .C2(
        DATAI_2_), .A(n5918), .ZN(n5919) );
  OAI211_X1 U6532 ( .C1(n5922), .C2(n5921), .A(n5920), .B(n5919), .ZN(n5927)
         );
  AOI22_X1 U6533 ( .A1(keyinput_96), .A2(MEMORYFETCH_REG_SCAN_IN), .B1(n6465), 
        .B2(keyinput_97), .ZN(n5923) );
  OAI221_X1 U6534 ( .B1(keyinput_96), .B2(MEMORYFETCH_REG_SCAN_IN), .C1(n6465), 
        .C2(keyinput_97), .A(n5923), .ZN(n5926) );
  AOI22_X1 U6535 ( .A1(BS16_N), .A2(keyinput_98), .B1(DATAI_0_), .B2(
        keyinput_95), .ZN(n5924) );
  OAI221_X1 U6536 ( .B1(BS16_N), .B2(keyinput_98), .C1(DATAI_0_), .C2(
        keyinput_95), .A(n5924), .ZN(n5925) );
  AOI211_X1 U6537 ( .C1(n5928), .C2(n5927), .A(n5926), .B(n5925), .ZN(n5931)
         );
  AOI22_X1 U6538 ( .A1(READREQUEST_REG_SCAN_IN), .A2(keyinput_101), .B1(n6462), 
        .B2(keyinput_99), .ZN(n5929) );
  OAI221_X1 U6539 ( .B1(READREQUEST_REG_SCAN_IN), .B2(keyinput_101), .C1(n6462), .C2(keyinput_99), .A(n5929), .ZN(n5930) );
  AOI211_X1 U6540 ( .C1(n6137), .C2(keyinput_100), .A(n5931), .B(n5930), .ZN(
        n5932) );
  OAI21_X1 U6541 ( .B1(n6137), .B2(keyinput_100), .A(n5932), .ZN(n5933) );
  OAI221_X1 U6542 ( .B1(keyinput_102), .B2(n5935), .C1(n5934), .C2(
        ADS_N_REG_SCAN_IN), .A(n5933), .ZN(n5936) );
  OAI221_X1 U6543 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(keyinput_103), .C1(n6127), 
        .C2(n5937), .A(n5936), .ZN(n5938) );
  OAI221_X1 U6544 ( .B1(M_IO_N_REG_SCAN_IN), .B2(n5939), .C1(n6472), .C2(
        keyinput_104), .A(n5938), .ZN(n5940) );
  OAI221_X1 U6545 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5941), .C1(n6129), .C2(
        keyinput_105), .A(n5940), .ZN(n5942) );
  OAI221_X1 U6546 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(n5943), .C1(n6139), 
        .C2(keyinput_106), .A(n5942), .ZN(n5944) );
  OAI211_X1 U6547 ( .C1(STATEBS16_REG_SCAN_IN), .C2(keyinput_107), .A(n5945), 
        .B(n5944), .ZN(n5946) );
  AOI21_X1 U6548 ( .B1(STATEBS16_REG_SCAN_IN), .B2(keyinput_107), .A(n5946), 
        .ZN(n5947) );
  OAI22_X1 U6549 ( .A1(keyinput_115), .A2(n6054), .B1(n5948), .B2(n5947), .ZN(
        n5949) );
  AOI21_X1 U6550 ( .B1(keyinput_115), .B2(n6054), .A(n5949), .ZN(n5950) );
  AOI221_X1 U6551 ( .B1(REIP_REG_30__SCAN_IN), .B2(n5952), .C1(n5951), .C2(
        keyinput_116), .A(n5950), .ZN(n5953) );
  AOI221_X1 U6552 ( .B1(REIP_REG_29__SCAN_IN), .B2(keyinput_117), .C1(n5955), 
        .C2(n5954), .A(n5953), .ZN(n5956) );
  AOI221_X1 U6553 ( .B1(REIP_REG_28__SCAN_IN), .B2(n5957), .C1(n6050), .C2(
        keyinput_118), .A(n5956), .ZN(n5959) );
  NAND2_X1 U6554 ( .A1(n6043), .A2(keyinput_121), .ZN(n5958) );
  OAI221_X1 U6555 ( .B1(n5960), .B2(n5959), .C1(n6043), .C2(keyinput_121), .A(
        n5958), .ZN(n5961) );
  OAI221_X1 U6556 ( .B1(REIP_REG_24__SCAN_IN), .B2(keyinput_122), .C1(n6041), 
        .C2(n5962), .A(n5961), .ZN(n5963) );
  AOI22_X1 U6557 ( .A1(keyinput_125), .A2(n6380), .B1(n5964), .B2(n5963), .ZN(
        n5965) );
  OAI21_X1 U6558 ( .B1(n6380), .B2(keyinput_125), .A(n5965), .ZN(n5966) );
  OAI221_X1 U6559 ( .B1(REIP_REG_20__SCAN_IN), .B2(keyinput_126), .C1(n5968), 
        .C2(n5967), .A(n5966), .ZN(n5969) );
  OAI221_X1 U6560 ( .B1(REIP_REG_19__SCAN_IN), .B2(keyinput_127), .C1(n6034), 
        .C2(n5970), .A(n5969), .ZN(n5971) );
  OAI21_X1 U6561 ( .B1(n6034), .B2(keyinput_63), .A(n5971), .ZN(n5972) );
  AOI211_X1 U6562 ( .C1(n6034), .C2(keyinput_63), .A(n5973), .B(n5972), .ZN(
        n5975) );
  NAND2_X1 U6563 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6474), .ZN(n6049) );
  INV_X1 U6564 ( .A(n6049), .ZN(n6051) );
  NAND2_X1 U6565 ( .A1(n6138), .A2(n6474), .ZN(n6053) );
  INV_X1 U6566 ( .A(n6053), .ZN(n6047) );
  AOI222_X1 U6567 ( .A1(n6471), .A2(ADDRESS_REG_28__SCAN_IN), .B1(
        REIP_REG_29__SCAN_IN), .B2(n6051), .C1(REIP_REG_30__SCAN_IN), .C2(
        n6047), .ZN(n5974) );
  XNOR2_X1 U6568 ( .A(n5975), .B(n5974), .ZN(U3212) );
  AOI22_X1 U6569 ( .A1(n6152), .A2(LWORD_REG_0__SCAN_IN), .B1(n6004), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n5976) );
  OAI21_X1 U6570 ( .B1(n5977), .B2(n6007), .A(n5976), .ZN(U2923) );
  AOI22_X1 U6571 ( .A1(n6152), .A2(LWORD_REG_1__SCAN_IN), .B1(n6004), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n5978) );
  OAI21_X1 U6572 ( .B1(n5979), .B2(n6007), .A(n5978), .ZN(U2922) );
  AOI22_X1 U6573 ( .A1(n6152), .A2(LWORD_REG_2__SCAN_IN), .B1(n6004), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n5980) );
  OAI21_X1 U6574 ( .B1(n5981), .B2(n6007), .A(n5980), .ZN(U2921) );
  AOI22_X1 U6575 ( .A1(n6152), .A2(LWORD_REG_3__SCAN_IN), .B1(n6004), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n5982) );
  OAI21_X1 U6576 ( .B1(n5983), .B2(n6007), .A(n5982), .ZN(U2920) );
  AOI22_X1 U6577 ( .A1(n6152), .A2(LWORD_REG_4__SCAN_IN), .B1(n6004), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n5984) );
  OAI21_X1 U6578 ( .B1(n5985), .B2(n6007), .A(n5984), .ZN(U2919) );
  AOI22_X1 U6579 ( .A1(n6152), .A2(LWORD_REG_5__SCAN_IN), .B1(n6004), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n5986) );
  OAI21_X1 U6580 ( .B1(n5987), .B2(n6007), .A(n5986), .ZN(U2918) );
  AOI22_X1 U6581 ( .A1(n6152), .A2(LWORD_REG_6__SCAN_IN), .B1(n6004), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n5988) );
  OAI21_X1 U6582 ( .B1(n5989), .B2(n6007), .A(n5988), .ZN(U2917) );
  AOI22_X1 U6583 ( .A1(n6152), .A2(LWORD_REG_7__SCAN_IN), .B1(n6004), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n5990) );
  OAI21_X1 U6584 ( .B1(n3997), .B2(n6007), .A(n5990), .ZN(U2916) );
  AOI22_X1 U6585 ( .A1(n6152), .A2(LWORD_REG_8__SCAN_IN), .B1(n6004), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n5991) );
  OAI21_X1 U6586 ( .B1(n5992), .B2(n6007), .A(n5991), .ZN(U2915) );
  AOI22_X1 U6587 ( .A1(n6152), .A2(LWORD_REG_9__SCAN_IN), .B1(n6004), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n5993) );
  OAI21_X1 U6588 ( .B1(n5994), .B2(n6007), .A(n5993), .ZN(U2914) );
  AOI22_X1 U6589 ( .A1(n6152), .A2(LWORD_REG_10__SCAN_IN), .B1(n6004), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n5995) );
  OAI21_X1 U6590 ( .B1(n5996), .B2(n6007), .A(n5995), .ZN(U2913) );
  AOI22_X1 U6591 ( .A1(n6152), .A2(LWORD_REG_11__SCAN_IN), .B1(n6004), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n5997) );
  OAI21_X1 U6592 ( .B1(n5998), .B2(n6007), .A(n5997), .ZN(U2912) );
  AOI22_X1 U6593 ( .A1(n6152), .A2(LWORD_REG_12__SCAN_IN), .B1(n6004), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n5999) );
  OAI21_X1 U6594 ( .B1(n4061), .B2(n6007), .A(n5999), .ZN(U2911) );
  AOI22_X1 U6595 ( .A1(n6152), .A2(LWORD_REG_13__SCAN_IN), .B1(n6004), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6000) );
  OAI21_X1 U6596 ( .B1(n6001), .B2(n6007), .A(n6000), .ZN(U2910) );
  AOI22_X1 U6597 ( .A1(n6152), .A2(LWORD_REG_14__SCAN_IN), .B1(n6004), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6002) );
  OAI21_X1 U6598 ( .B1(n6003), .B2(n6007), .A(n6002), .ZN(U2909) );
  AOI22_X1 U6599 ( .A1(n6152), .A2(LWORD_REG_15__SCAN_IN), .B1(n6004), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6006) );
  OAI21_X1 U6600 ( .B1(n6008), .B2(n6007), .A(n6006), .ZN(U2908) );
  INV_X1 U6601 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6261) );
  AOI22_X1 U6602 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6047), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6471), .ZN(n6009) );
  OAI21_X1 U6603 ( .B1(n6261), .B2(n6049), .A(n6009), .ZN(U3184) );
  AOI22_X1 U6604 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6051), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6471), .ZN(n6010) );
  OAI21_X1 U6605 ( .B1(n4870), .B2(n6053), .A(n6010), .ZN(U3185) );
  AOI22_X1 U6606 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6047), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6471), .ZN(n6011) );
  OAI21_X1 U6607 ( .B1(n4870), .B2(n6049), .A(n6011), .ZN(U3186) );
  AOI22_X1 U6608 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6051), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6471), .ZN(n6012) );
  OAI21_X1 U6609 ( .B1(n6013), .B2(n6053), .A(n6012), .ZN(U3187) );
  INV_X1 U6610 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6016) );
  AOI22_X1 U6611 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6051), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6471), .ZN(n6014) );
  OAI21_X1 U6612 ( .B1(n6016), .B2(n6053), .A(n6014), .ZN(U3188) );
  AOI22_X1 U6613 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6047), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6471), .ZN(n6015) );
  OAI21_X1 U6614 ( .B1(n6016), .B2(n6049), .A(n6015), .ZN(U3189) );
  AOI22_X1 U6615 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6051), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6471), .ZN(n6017) );
  OAI21_X1 U6616 ( .B1(n6019), .B2(n6053), .A(n6017), .ZN(U3190) );
  AOI22_X1 U6617 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6047), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6471), .ZN(n6018) );
  OAI21_X1 U6618 ( .B1(n6019), .B2(n6049), .A(n6018), .ZN(U3191) );
  AOI22_X1 U6619 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6051), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6471), .ZN(n6020) );
  OAI21_X1 U6620 ( .B1(n6021), .B2(n6053), .A(n6020), .ZN(U3192) );
  INV_X1 U6621 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6206) );
  AOI22_X1 U6622 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6051), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6471), .ZN(n6022) );
  OAI21_X1 U6623 ( .B1(n6206), .B2(n6053), .A(n6022), .ZN(U3193) );
  AOI22_X1 U6624 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6051), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6471), .ZN(n6023) );
  OAI21_X1 U6625 ( .B1(n5094), .B2(n6053), .A(n6023), .ZN(U3194) );
  AOI22_X1 U6626 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6047), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6471), .ZN(n6024) );
  OAI21_X1 U6627 ( .B1(n5094), .B2(n6049), .A(n6024), .ZN(U3195) );
  AOI22_X1 U6628 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6051), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6471), .ZN(n6025) );
  OAI21_X1 U6629 ( .B1(n6177), .B2(n6053), .A(n6025), .ZN(U3196) );
  AOI22_X1 U6630 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6047), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6471), .ZN(n6026) );
  OAI21_X1 U6631 ( .B1(n6177), .B2(n6049), .A(n6026), .ZN(U3197) );
  INV_X1 U6632 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6028) );
  AOI22_X1 U6633 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6047), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6471), .ZN(n6027) );
  OAI21_X1 U6634 ( .B1(n6028), .B2(n6049), .A(n6027), .ZN(U3198) );
  AOI22_X1 U6635 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6051), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6471), .ZN(n6029) );
  OAI21_X1 U6636 ( .B1(n6031), .B2(n6053), .A(n6029), .ZN(U3199) );
  AOI22_X1 U6637 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6047), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6471), .ZN(n6030) );
  OAI21_X1 U6638 ( .B1(n6031), .B2(n6049), .A(n6030), .ZN(U3200) );
  AOI22_X1 U6639 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6051), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6471), .ZN(n6032) );
  OAI21_X1 U6640 ( .B1(n6034), .B2(n6053), .A(n6032), .ZN(U3201) );
  AOI22_X1 U6641 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6047), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6471), .ZN(n6033) );
  OAI21_X1 U6642 ( .B1(n6034), .B2(n6049), .A(n6033), .ZN(U3202) );
  AOI22_X1 U6643 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6051), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6471), .ZN(n6035) );
  OAI21_X1 U6644 ( .B1(n6380), .B2(n6053), .A(n6035), .ZN(U3203) );
  AOI22_X1 U6645 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6047), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6471), .ZN(n6036) );
  OAI21_X1 U6646 ( .B1(n6380), .B2(n6049), .A(n6036), .ZN(U3204) );
  AOI22_X1 U6647 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6047), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6471), .ZN(n6037) );
  OAI21_X1 U6648 ( .B1(n6381), .B2(n6049), .A(n6037), .ZN(U3205) );
  AOI22_X1 U6649 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6047), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6471), .ZN(n6038) );
  OAI21_X1 U6650 ( .B1(n6039), .B2(n6049), .A(n6038), .ZN(U3206) );
  AOI22_X1 U6651 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6047), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6471), .ZN(n6040) );
  OAI21_X1 U6652 ( .B1(n6041), .B2(n6049), .A(n6040), .ZN(U3207) );
  AOI22_X1 U6653 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6047), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6471), .ZN(n6042) );
  OAI21_X1 U6654 ( .B1(n6043), .B2(n6049), .A(n6042), .ZN(U3208) );
  AOI22_X1 U6655 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6051), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6471), .ZN(n6044) );
  OAI21_X1 U6656 ( .B1(n6045), .B2(n6053), .A(n6044), .ZN(U3209) );
  AOI22_X1 U6657 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6051), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6471), .ZN(n6046) );
  OAI21_X1 U6658 ( .B1(n6050), .B2(n6053), .A(n6046), .ZN(U3210) );
  AOI22_X1 U6659 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6047), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6471), .ZN(n6048) );
  OAI21_X1 U6660 ( .B1(n6050), .B2(n6049), .A(n6048), .ZN(U3211) );
  AOI22_X1 U6661 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6051), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6471), .ZN(n6052) );
  OAI21_X1 U6662 ( .B1(n6054), .B2(n6053), .A(n6052), .ZN(U3213) );
  MUX2_X1 U6663 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n6471), .Z(U3445) );
  NOR4_X1 U6664 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(
        DATAWIDTH_REG_12__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(
        DATAWIDTH_REG_10__SCAN_IN), .ZN(n6058) );
  NOR4_X1 U6665 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(
        DATAWIDTH_REG_16__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(
        DATAWIDTH_REG_14__SCAN_IN), .ZN(n6057) );
  NOR4_X1 U6666 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_2__SCAN_IN), .ZN(
        n6056) );
  NOR4_X1 U6667 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), 
        .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_6__SCAN_IN), .ZN(
        n6055) );
  NAND4_X1 U6668 ( .A1(n6058), .A2(n6057), .A3(n6056), .A4(n6055), .ZN(n6064)
         );
  NOR4_X1 U6669 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_27__SCAN_IN), .A4(
        DATAWIDTH_REG_26__SCAN_IN), .ZN(n6062) );
  AOI211_X1 U6670 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_31__SCAN_IN), .B(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n6061) );
  NOR4_X1 U6671 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_19__SCAN_IN), .A4(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n6060) );
  NOR4_X1 U6672 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(
        DATAWIDTH_REG_24__SCAN_IN), .A3(DATAWIDTH_REG_23__SCAN_IN), .A4(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n6059) );
  NAND4_X1 U6673 ( .A1(n6062), .A2(n6061), .A3(n6060), .A4(n6059), .ZN(n6063)
         );
  NOR2_X1 U6674 ( .A1(n6064), .A2(n6063), .ZN(n6068) );
  INV_X1 U6675 ( .A(n6068), .ZN(n6073) );
  NOR2_X1 U6676 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6073), .ZN(n6076) );
  INV_X1 U6677 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6455) );
  AOI22_X1 U6678 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(n6073), .B1(n6076), 
        .B2(n6455), .ZN(n6065) );
  NAND4_X1 U6679 ( .A1(n6068), .A2(n6075), .A3(n6455), .A4(n6066), .ZN(n6072)
         );
  NAND2_X1 U6680 ( .A1(n6065), .A2(n6072), .ZN(U2795) );
  MUX2_X1 U6681 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6471), .Z(U3446) );
  OAI211_X1 U6682 ( .C1(n6066), .C2(n6075), .A(n6455), .B(n6076), .ZN(n6070)
         );
  OAI21_X1 U6683 ( .B1(n6261), .B2(n6075), .A(n6068), .ZN(n6067) );
  OAI21_X1 U6684 ( .B1(BYTEENABLE_REG_2__SCAN_IN), .B2(n6068), .A(n6067), .ZN(
        n6069) );
  NAND2_X1 U6685 ( .A1(n6070), .A2(n6069), .ZN(U3468) );
  MUX2_X1 U6686 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6471), .Z(U3447) );
  INV_X1 U6687 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6071) );
  AOI22_X1 U6688 ( .A1(n6076), .A2(n6072), .B1(n6071), .B2(n6073), .ZN(U2794)
         );
  MUX2_X1 U6689 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6471), .Z(U3448) );
  AOI22_X1 U6690 ( .A1(n6076), .A2(n6075), .B1(n6074), .B2(n6073), .ZN(U3469)
         );
  INV_X1 U6691 ( .A(EBX_REG_2__SCAN_IN), .ZN(n6080) );
  XNOR2_X1 U6692 ( .A(n6078), .B(n6077), .ZN(n6263) );
  AOI22_X1 U6693 ( .A1(n6272), .A2(n6083), .B1(n6082), .B2(n6263), .ZN(n6079)
         );
  OAI21_X1 U6694 ( .B1(n6086), .B2(n6080), .A(n6079), .ZN(U2857) );
  AOI22_X1 U6695 ( .A1(n6685), .A2(n6083), .B1(n6082), .B2(n6081), .ZN(n6084)
         );
  OAI21_X1 U6696 ( .B1(n6086), .B2(n6085), .A(n6084), .ZN(U2835) );
  AOI22_X1 U6697 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n6119), .B1(n6235), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n6091) );
  INV_X1 U6698 ( .A(n6087), .ZN(n6258) );
  INV_X1 U6699 ( .A(n6088), .ZN(n6089) );
  AOI22_X1 U6700 ( .A1(n6969), .A2(n6258), .B1(n6089), .B2(n6121), .ZN(n6090)
         );
  OAI211_X1 U6701 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n6125), .A(n6091), 
        .B(n6090), .ZN(U2985) );
  AOI22_X1 U6702 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n6119), .B1(n6235), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U6703 ( .A1(n6093), .A2(n6092), .ZN(n6094) );
  XOR2_X1 U6704 ( .A(n6095), .B(n6094), .Z(n6181) );
  AOI22_X1 U6705 ( .A1(n6181), .A2(n6121), .B1(n6969), .B2(n6272), .ZN(n6096)
         );
  OAI211_X1 U6706 ( .C1(n6125), .C2(n6275), .A(n6097), .B(n6096), .ZN(U2984)
         );
  NAND2_X1 U6707 ( .A1(n6099), .A2(n6098), .ZN(n6102) );
  NAND2_X1 U6708 ( .A1(n6109), .A2(n6100), .ZN(n6101) );
  XOR2_X1 U6709 ( .A(n6102), .B(n6101), .Z(n6208) );
  AOI22_X1 U6710 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n6119), .B1(n6235), 
        .B2(REIP_REG_11__SCAN_IN), .ZN(n6107) );
  AOI22_X1 U6711 ( .A1(n6105), .A2(n6969), .B1(n6104), .B2(n6103), .ZN(n6106)
         );
  OAI211_X1 U6712 ( .C1(n6208), .C2(n6397), .A(n6107), .B(n6106), .ZN(U2975)
         );
  AOI22_X1 U6713 ( .A1(PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n6119), .B1(n6235), 
        .B2(REIP_REG_13__SCAN_IN), .ZN(n6115) );
  NAND2_X1 U6714 ( .A1(n6109), .A2(n6108), .ZN(n6111) );
  NAND2_X1 U6715 ( .A1(n6111), .A2(n6110), .ZN(n6113) );
  XNOR2_X1 U6716 ( .A(n6113), .B(n6112), .ZN(n6166) );
  AOI22_X1 U6717 ( .A1(n6166), .A2(n6121), .B1(n6969), .B2(n6327), .ZN(n6114)
         );
  OAI211_X1 U6718 ( .C1(n6125), .C2(n6332), .A(n6115), .B(n6114), .ZN(U2973)
         );
  AOI22_X1 U6719 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n6119), .B1(n6235), 
        .B2(REIP_REG_18__SCAN_IN), .ZN(n6118) );
  AOI22_X1 U6720 ( .A1(n6116), .A2(n6121), .B1(n6969), .B2(n6479), .ZN(n6117)
         );
  OAI211_X1 U6721 ( .C1(n6125), .C2(n6363), .A(n6118), .B(n6117), .ZN(U2968)
         );
  AOI22_X1 U6722 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n6119), .B1(n6235), 
        .B2(REIP_REG_20__SCAN_IN), .ZN(n6124) );
  AOI22_X1 U6723 ( .A1(n6122), .A2(n6121), .B1(n6969), .B2(n6482), .ZN(n6123)
         );
  OAI211_X1 U6724 ( .C1(n6125), .C2(n6373), .A(n6124), .B(n6123), .ZN(U2966)
         );
  NOR2_X1 U6725 ( .A1(n6126), .A2(n6428), .ZN(n6128) );
  OAI22_X1 U6726 ( .A1(n6128), .A2(n6127), .B1(n6491), .B2(n6134), .ZN(U2790)
         );
  OAI222_X1 U6727 ( .A1(n6474), .A2(n6130), .B1(n6474), .B2(n6129), .C1(
        CODEFETCH_REG_SCAN_IN), .C2(n6471), .ZN(U2791) );
  INV_X1 U6728 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6135) );
  INV_X1 U6729 ( .A(n6131), .ZN(n6132) );
  NAND2_X1 U6730 ( .A1(n6150), .A2(n6132), .ZN(n6133) );
  OAI211_X1 U6731 ( .C1(n6150), .C2(n6135), .A(n6134), .B(n6133), .ZN(U3474)
         );
  AOI22_X1 U6732 ( .A1(n6474), .A2(READREQUEST_REG_SCAN_IN), .B1(n6136), .B2(
        n6471), .ZN(U3470) );
  NOR2_X1 U6733 ( .A1(n6138), .A2(n6137), .ZN(n6457) );
  NOR2_X1 U6734 ( .A1(n6463), .A2(n6139), .ZN(n6466) );
  AOI21_X1 U6735 ( .B1(HOLD), .B2(STATE_REG_1__SCAN_IN), .A(n6466), .ZN(n6142)
         );
  NOR2_X1 U6736 ( .A1(n6140), .A2(n6462), .ZN(n6459) );
  INV_X1 U6737 ( .A(n6459), .ZN(n6467) );
  OAI211_X1 U6738 ( .C1(n6457), .C2(n6142), .A(n6141), .B(n6467), .ZN(U3182)
         );
  NOR2_X1 U6739 ( .A1(READY_N), .A2(n6491), .ZN(n6433) );
  OAI211_X1 U6740 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6433), .A(n6441), .B(
        n6148), .ZN(n6143) );
  NAND2_X1 U6741 ( .A1(n6144), .A2(n6143), .ZN(U3150) );
  INV_X1 U6742 ( .A(n6145), .ZN(n6146) );
  AOI211_X1 U6743 ( .C1(n6147), .C2(n6670), .A(n6657), .B(n6146), .ZN(n6149)
         );
  OAI21_X1 U6744 ( .B1(n6149), .B2(n6491), .A(n6148), .ZN(n6154) );
  AOI211_X1 U6745 ( .C1(n6152), .C2(n6462), .A(n6151), .B(n6150), .ZN(n6153)
         );
  MUX2_X1 U6746 ( .A(n6154), .B(REQUESTPENDING_REG_SCAN_IN), .S(n6153), .Z(
        U3472) );
  AOI22_X1 U6747 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n6155), .B1(n6235), .B2(REIP_REG_19__SCAN_IN), .ZN(n6159) );
  AOI22_X1 U6748 ( .A1(n6157), .A2(n6244), .B1(n6243), .B2(n6156), .ZN(n6158)
         );
  OAI211_X1 U6749 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n6160), .A(n6159), .B(n6158), .ZN(U2999) );
  NOR3_X1 U6750 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n6161), .A3(n3853), 
        .ZN(n6163) );
  AOI22_X1 U6751 ( .A1(n6235), .A2(REIP_REG_13__SCAN_IN), .B1(n6162), .B2(
        n6163), .ZN(n6169) );
  AOI22_X1 U6752 ( .A1(n6164), .A2(n6163), .B1(n6243), .B2(n6323), .ZN(n6168)
         );
  OAI21_X1 U6753 ( .B1(n6194), .B2(n6174), .A(n6165), .ZN(n6173) );
  AOI22_X1 U6754 ( .A1(n6166), .A2(n6244), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n6173), .ZN(n6167) );
  NAND3_X1 U6755 ( .A1(n6169), .A2(n6168), .A3(n6167), .ZN(U3005) );
  INV_X1 U6756 ( .A(n6333), .ZN(n6170) );
  OAI22_X1 U6757 ( .A1(n6171), .A2(n6225), .B1(n6224), .B2(n6170), .ZN(n6172)
         );
  AOI21_X1 U6758 ( .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n6173), .A(n6172), 
        .ZN(n6176) );
  NAND3_X1 U6759 ( .A1(n6174), .A2(n5644), .A3(n6233), .ZN(n6175) );
  OAI211_X1 U6760 ( .C1(n6177), .C2(n6247), .A(n6176), .B(n6175), .ZN(U3004)
         );
  AOI22_X1 U6761 ( .A1(n6243), .A2(n6263), .B1(n6235), .B2(REIP_REG_2__SCAN_IN), .ZN(n6187) );
  NAND2_X1 U6762 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6180) );
  OAI21_X1 U6763 ( .B1(n6180), .B2(n6179), .A(n6178), .ZN(n6182) );
  AOI22_X1 U6764 ( .A1(n6182), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n6244), 
        .B2(n6181), .ZN(n6186) );
  OR3_X1 U6765 ( .A1(n3669), .A2(n6183), .A3(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6184) );
  NAND4_X1 U6766 ( .A1(n6187), .A2(n6186), .A3(n6185), .A4(n6184), .ZN(U3016)
         );
  NAND2_X1 U6767 ( .A1(n6193), .A2(n6188), .ZN(n6205) );
  AOI22_X1 U6768 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n4485), .B1(
        INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6189), .ZN(n6198) );
  AOI21_X1 U6769 ( .B1(n6191), .B2(n6243), .A(n6190), .ZN(n6197) );
  OAI21_X1 U6770 ( .B1(n6194), .B2(n6193), .A(n6192), .ZN(n6201) );
  AOI22_X1 U6771 ( .A1(n6195), .A2(n6244), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6201), .ZN(n6196) );
  OAI211_X1 U6772 ( .C1(n6205), .C2(n6198), .A(n6197), .B(n6196), .ZN(U3008)
         );
  INV_X1 U6773 ( .A(n6199), .ZN(n6313) );
  AOI21_X1 U6774 ( .B1(n6243), .B2(n6313), .A(n6200), .ZN(n6204) );
  AOI22_X1 U6775 ( .A1(n6202), .A2(n6244), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6201), .ZN(n6203) );
  OAI211_X1 U6776 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6205), .A(n6204), 
        .B(n6203), .ZN(U3009) );
  OAI22_X1 U6777 ( .A1(n6207), .A2(n6224), .B1(n6206), .B2(n6247), .ZN(n6210)
         );
  NOR2_X1 U6778 ( .A1(n6208), .A2(n6225), .ZN(n6209) );
  AOI211_X1 U6779 ( .C1(INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n6213), .A(n6210), .B(n6209), .ZN(n6212) );
  NAND2_X1 U6780 ( .A1(n6212), .A2(n6211), .ZN(U3007) );
  AOI21_X1 U6781 ( .B1(n6216), .B2(n6214), .A(n6213), .ZN(n6231) );
  NOR2_X1 U6782 ( .A1(n6216), .A2(n6215), .ZN(n6221) );
  AOI22_X1 U6783 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6235), .B1(n6221), .B2(
        n6222), .ZN(n6220) );
  AOI22_X1 U6784 ( .A1(n6218), .A2(n6244), .B1(n6243), .B2(n6217), .ZN(n6219)
         );
  OAI211_X1 U6785 ( .C1(n6231), .C2(n6222), .A(n6220), .B(n6219), .ZN(U3003)
         );
  OAI221_X1 U6786 ( .B1(n6230), .B2(n6222), .C1(
        INSTADDRPOINTER_REG_16__SCAN_IN), .C2(INSTADDRPOINTER_REG_15__SCAN_IN), 
        .A(n6221), .ZN(n6223) );
  INV_X1 U6787 ( .A(n6223), .ZN(n6228) );
  OAI22_X1 U6788 ( .A1(n6226), .A2(n6225), .B1(n6224), .B2(n6357), .ZN(n6227)
         );
  AOI211_X1 U6789 ( .C1(REIP_REG_16__SCAN_IN), .C2(n6235), .A(n6228), .B(n6227), .ZN(n6229) );
  OAI21_X1 U6790 ( .B1(n6231), .B2(n6230), .A(n6229), .ZN(U3002) );
  NOR2_X1 U6791 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n6232), .ZN(n6234)
         );
  AOI22_X1 U6792 ( .A1(n6235), .A2(REIP_REG_17__SCAN_IN), .B1(n6234), .B2(
        n6233), .ZN(n6239) );
  AOI22_X1 U6793 ( .A1(n6237), .A2(n6244), .B1(n6243), .B2(n6236), .ZN(n6238)
         );
  OAI211_X1 U6794 ( .C1(n6241), .C2(n6240), .A(n6239), .B(n6238), .ZN(U3001)
         );
  AOI22_X1 U6795 ( .A1(n6245), .A2(n6244), .B1(n6243), .B2(n6242), .ZN(n6253)
         );
  INV_X1 U6796 ( .A(n6246), .ZN(n6249) );
  NOR2_X1 U6797 ( .A1(n6247), .A2(n6380), .ZN(n6248) );
  AOI221_X1 U6798 ( .B1(n6251), .B2(n6250), .C1(n6249), .C2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .A(n6248), .ZN(n6252) );
  NAND2_X1 U6799 ( .A1(n6253), .A2(n6252), .ZN(U2997) );
  AOI22_X1 U6800 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n6370), .B1(
        EBX_REG_1__SCAN_IN), .B2(n6369), .ZN(n6260) );
  INV_X1 U6801 ( .A(n6254), .ZN(n6255) );
  OAI22_X1 U6802 ( .A1(n6255), .A2(n4669), .B1(PHYADDRPOINTER_REG_1__SCAN_IN), 
        .B2(n6395), .ZN(n6257) );
  OAI22_X1 U6803 ( .A1(n4742), .A2(n6264), .B1(n6301), .B2(REIP_REG_1__SCAN_IN), .ZN(n6256) );
  AOI211_X1 U6804 ( .C1(n6258), .C2(n6271), .A(n6257), .B(n6256), .ZN(n6259)
         );
  OAI211_X1 U6805 ( .C1(n6283), .C2(n6261), .A(n6260), .B(n6259), .ZN(U2826)
         );
  OAI21_X1 U6806 ( .B1(n6301), .B2(REIP_REG_1__SCAN_IN), .A(n6283), .ZN(n6262)
         );
  AOI22_X1 U6807 ( .A1(n6334), .A2(n6263), .B1(REIP_REG_2__SCAN_IN), .B2(n6262), .ZN(n6274) );
  INV_X1 U6808 ( .A(n6264), .ZN(n6265) );
  AOI22_X1 U6809 ( .A1(n6265), .A2(n4887), .B1(n6369), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n6268) );
  INV_X1 U6810 ( .A(n6301), .ZN(n6282) );
  INV_X1 U6811 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6266) );
  NAND3_X1 U6812 ( .A1(n6282), .A2(n6266), .A3(REIP_REG_1__SCAN_IN), .ZN(n6267) );
  OAI211_X1 U6813 ( .C1(n6384), .C2(n6269), .A(n6268), .B(n6267), .ZN(n6270)
         );
  AOI21_X1 U6814 ( .B1(n6272), .B2(n6271), .A(n6270), .ZN(n6273) );
  OAI211_X1 U6815 ( .C1(n6275), .C2(n6395), .A(n6274), .B(n6273), .ZN(U2825)
         );
  AOI22_X1 U6816 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n6370), .B1(
        EBX_REG_5__SCAN_IN), .B2(n6369), .ZN(n6288) );
  OAI22_X1 U6817 ( .A1(n6278), .A2(n6277), .B1(n6276), .B2(n6395), .ZN(n6279)
         );
  AOI21_X1 U6818 ( .B1(n6334), .B2(n6280), .A(n6279), .ZN(n6287) );
  AND2_X1 U6819 ( .A1(n6282), .A2(n6281), .ZN(n6285) );
  OAI21_X1 U6820 ( .B1(n6301), .B2(n6284), .A(n6283), .ZN(n6306) );
  OAI21_X1 U6821 ( .B1(n6285), .B2(REIP_REG_5__SCAN_IN), .A(n6306), .ZN(n6286)
         );
  NAND4_X1 U6822 ( .A1(n6288), .A2(n6287), .A3(n6343), .A4(n6286), .ZN(U2822)
         );
  AOI22_X1 U6823 ( .A1(n6334), .A2(n6289), .B1(REIP_REG_6__SCAN_IN), .B2(n6306), .ZN(n6298) );
  NOR3_X1 U6824 ( .A1(n6301), .A2(REIP_REG_6__SCAN_IN), .A3(n6290), .ZN(n6307)
         );
  OAI22_X1 U6825 ( .A1(n6292), .A2(n6384), .B1(n6291), .B2(n6382), .ZN(n6296)
         );
  OAI22_X1 U6826 ( .A1(n6294), .A2(n6390), .B1(n6293), .B2(n6395), .ZN(n6295)
         );
  NOR4_X1 U6827 ( .A1(n6362), .A2(n6307), .A3(n6296), .A4(n6295), .ZN(n6297)
         );
  NAND2_X1 U6828 ( .A1(n6298), .A2(n6297), .ZN(U2821) );
  AOI22_X1 U6829 ( .A1(EBX_REG_7__SCAN_IN), .A2(n6369), .B1(n6334), .B2(n6299), 
        .ZN(n6311) );
  NOR3_X1 U6830 ( .A1(n6301), .A2(REIP_REG_7__SCAN_IN), .A3(n6300), .ZN(n6302)
         );
  AOI211_X1 U6831 ( .C1(n6370), .C2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n6362), 
        .B(n6302), .ZN(n6310) );
  NOR2_X1 U6832 ( .A1(n6395), .A2(n6303), .ZN(n6304) );
  AOI21_X1 U6833 ( .B1(n6305), .B2(n6375), .A(n6304), .ZN(n6309) );
  OAI21_X1 U6834 ( .B1(n6307), .B2(n6306), .A(REIP_REG_7__SCAN_IN), .ZN(n6308)
         );
  NAND4_X1 U6835 ( .A1(n6311), .A2(n6310), .A3(n6309), .A4(n6308), .ZN(U2820)
         );
  AOI22_X1 U6836 ( .A1(n6334), .A2(n6313), .B1(REIP_REG_9__SCAN_IN), .B2(n6312), .ZN(n6321) );
  AOI22_X1 U6837 ( .A1(PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n6370), .B1(n6315), 
        .B2(n6314), .ZN(n6320) );
  AOI21_X1 U6838 ( .B1(n6369), .B2(EBX_REG_9__SCAN_IN), .A(n6362), .ZN(n6319)
         );
  AOI22_X1 U6839 ( .A1(n6317), .A2(n6375), .B1(n6354), .B2(n6316), .ZN(n6318)
         );
  NAND4_X1 U6840 ( .A1(n6321), .A2(n6320), .A3(n6319), .A4(n6318), .ZN(U2818)
         );
  NOR3_X1 U6841 ( .A1(n6322), .A2(REIP_REG_13__SCAN_IN), .A3(n5094), .ZN(n6326) );
  AOI22_X1 U6842 ( .A1(EBX_REG_13__SCAN_IN), .A2(n6369), .B1(n6334), .B2(n6323), .ZN(n6324) );
  OAI211_X1 U6843 ( .C1(n6384), .C2(n4096), .A(n6324), .B(n6343), .ZN(n6325)
         );
  AOI211_X1 U6844 ( .C1(n6327), .C2(n6375), .A(n6326), .B(n6325), .ZN(n6331)
         );
  OAI21_X1 U6845 ( .B1(n6329), .B2(n6328), .A(REIP_REG_13__SCAN_IN), .ZN(n6330) );
  OAI211_X1 U6846 ( .C1(n6395), .C2(n6332), .A(n6331), .B(n6330), .ZN(U2814)
         );
  AOI22_X1 U6847 ( .A1(n6334), .A2(n6333), .B1(REIP_REG_14__SCAN_IN), .B2(
        n6348), .ZN(n6346) );
  NOR2_X1 U6848 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6335), .ZN(n6340) );
  OAI22_X1 U6849 ( .A1(n6337), .A2(n6384), .B1(n6336), .B2(n6382), .ZN(n6338)
         );
  AOI21_X1 U6850 ( .B1(n6340), .B2(n6339), .A(n6338), .ZN(n6345) );
  AOI22_X1 U6851 ( .A1(n6342), .A2(n6375), .B1(n6354), .B2(n6341), .ZN(n6344)
         );
  NAND4_X1 U6852 ( .A1(n6346), .A2(n6345), .A3(n6344), .A4(n6343), .ZN(U2813)
         );
  NAND2_X1 U6853 ( .A1(REIP_REG_15__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .ZN(
        n6347) );
  OAI21_X1 U6854 ( .B1(REIP_REG_15__SCAN_IN), .B2(REIP_REG_16__SCAN_IN), .A(
        n6347), .ZN(n6350) );
  AOI22_X1 U6855 ( .A1(EBX_REG_16__SCAN_IN), .A2(n6369), .B1(
        REIP_REG_16__SCAN_IN), .B2(n6348), .ZN(n6349) );
  OAI21_X1 U6856 ( .B1(n6351), .B2(n6350), .A(n6349), .ZN(n6352) );
  AOI211_X1 U6857 ( .C1(n6370), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6362), 
        .B(n6352), .ZN(n6356) );
  AOI22_X1 U6858 ( .A1(n6476), .A2(n6375), .B1(n6354), .B2(n6353), .ZN(n6355)
         );
  OAI211_X1 U6859 ( .C1(n6389), .C2(n6357), .A(n6356), .B(n6355), .ZN(U2811)
         );
  AOI22_X1 U6860 ( .A1(EBX_REG_18__SCAN_IN), .A2(n6369), .B1(
        REIP_REG_18__SCAN_IN), .B2(n6358), .ZN(n6359) );
  OAI21_X1 U6861 ( .B1(REIP_REG_18__SCAN_IN), .B2(n6360), .A(n6359), .ZN(n6361) );
  AOI211_X1 U6862 ( .C1(n6370), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6362), 
        .B(n6361), .ZN(n6366) );
  NOR2_X1 U6863 ( .A1(n6395), .A2(n6363), .ZN(n6364) );
  AOI21_X1 U6864 ( .B1(n6479), .B2(n6375), .A(n6364), .ZN(n6365) );
  OAI211_X1 U6865 ( .C1(n6367), .C2(n6389), .A(n6366), .B(n6365), .ZN(U2809)
         );
  OAI21_X1 U6866 ( .B1(REIP_REG_20__SCAN_IN), .B2(n6368), .A(n6387), .ZN(n6372) );
  AOI22_X1 U6867 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n6370), .B1(
        EBX_REG_20__SCAN_IN), .B2(n6369), .ZN(n6371) );
  OAI211_X1 U6868 ( .C1(n6373), .C2(n6395), .A(n6372), .B(n6371), .ZN(n6374)
         );
  AOI21_X1 U6869 ( .B1(n6482), .B2(n6375), .A(n6374), .ZN(n6376) );
  OAI21_X1 U6870 ( .B1(n6377), .B2(n6389), .A(n6376), .ZN(U2807) );
  AOI211_X1 U6871 ( .C1(n6381), .C2(n6380), .A(n6379), .B(n6378), .ZN(n6386)
         );
  OAI22_X1 U6872 ( .A1(n4143), .A2(n6384), .B1(n6383), .B2(n6382), .ZN(n6385)
         );
  AOI211_X1 U6873 ( .C1(n6387), .C2(REIP_REG_22__SCAN_IN), .A(n6386), .B(n6385), .ZN(n6394) );
  OAI22_X1 U6874 ( .A1(n6391), .A2(n6390), .B1(n6389), .B2(n6388), .ZN(n6392)
         );
  INV_X1 U6875 ( .A(n6392), .ZN(n6393) );
  OAI211_X1 U6876 ( .C1(n6396), .C2(n6395), .A(n6394), .B(n6393), .ZN(U2805)
         );
  OAI21_X1 U6877 ( .B1(n6399), .B2(n6398), .A(n6397), .ZN(U2793) );
  INV_X1 U6878 ( .A(n6400), .ZN(n6401) );
  NAND3_X1 U6879 ( .A1(n6402), .A2(n6401), .A3(n6678), .ZN(n6403) );
  OAI21_X1 U6880 ( .B1(n6405), .B2(n6404), .A(n6403), .ZN(U3455) );
  AOI211_X1 U6881 ( .C1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n6407), .A(n6647), .B(n6406), .ZN(n6411) );
  INV_X1 U6882 ( .A(n6411), .ZN(n6413) );
  INV_X1 U6883 ( .A(n6408), .ZN(n6409) );
  OAI22_X1 U6884 ( .A1(n6411), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n6410), .B2(n6409), .ZN(n6412) );
  OAI21_X1 U6885 ( .B1(n6413), .B2(n6621), .A(n6412), .ZN(n6414) );
  AOI222_X1 U6886 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6415), .B1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6414), .C1(n6415), .C2(n6414), 
        .ZN(n6416) );
  AOI222_X1 U6887 ( .A1(n6499), .A2(n6417), .B1(n6499), .B2(n6416), .C1(n6417), 
        .C2(n6416), .ZN(n6418) );
  OR2_X1 U6888 ( .A1(n6418), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6426)
         );
  NOR2_X1 U6889 ( .A1(FLUSH_REG_SCAN_IN), .A2(MORE_REG_SCAN_IN), .ZN(n6422) );
  OAI211_X1 U6890 ( .C1(n6422), .C2(n6421), .A(n6420), .B(n6419), .ZN(n6423)
         );
  NOR2_X1 U6891 ( .A1(n6424), .A2(n6423), .ZN(n6425) );
  NAND2_X1 U6892 ( .A1(n6426), .A2(n6425), .ZN(n6448) );
  OAI22_X1 U6893 ( .A1(n6448), .A2(n6428), .B1(n6462), .B2(n6427), .ZN(n6432)
         );
  OR2_X1 U6894 ( .A1(n6430), .A2(n6429), .ZN(n6431) );
  OAI221_X1 U6895 ( .B1(n6443), .B2(READY_N), .C1(n6443), .C2(n6657), .A(
        STATE2_REG_0__SCAN_IN), .ZN(n6450) );
  AOI21_X1 U6896 ( .B1(n6434), .B2(n6433), .A(n6449), .ZN(n6435) );
  NOR2_X1 U6897 ( .A1(n6435), .A2(n6443), .ZN(n6436) );
  AOI211_X1 U6898 ( .C1(n6443), .C2(n6438), .A(n6437), .B(n6436), .ZN(n6439)
         );
  OAI21_X1 U6899 ( .B1(n6440), .B2(n6450), .A(n6439), .ZN(U3149) );
  INV_X1 U6900 ( .A(n6443), .ZN(n6442) );
  OAI221_X1 U6901 ( .B1(n6678), .B2(STATE2_REG_0__SCAN_IN), .C1(n6678), .C2(
        n6442), .A(n6441), .ZN(U3453) );
  AOI211_X1 U6902 ( .C1(n6445), .C2(n6444), .A(STATE2_REG_0__SCAN_IN), .B(
        n6443), .ZN(n6446) );
  AOI211_X1 U6903 ( .C1(n6449), .C2(n6448), .A(n6447), .B(n6446), .ZN(n6451)
         );
  OAI211_X1 U6904 ( .C1(n6491), .C2(n6452), .A(n6451), .B(n6450), .ZN(U3148)
         );
  INV_X1 U6905 ( .A(n6453), .ZN(n6454) );
  OAI21_X1 U6906 ( .B1(n6456), .B2(n6670), .A(n6454), .ZN(U2792) );
  OAI21_X1 U6907 ( .B1(n6456), .B2(n6455), .A(n6454), .ZN(U3452) );
  NAND2_X1 U6908 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6461) );
  AOI221_X1 U6909 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6465), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6469) );
  AOI221_X1 U6910 ( .B1(n6459), .B2(n6458), .C1(n6457), .C2(n6458), .A(n6469), 
        .ZN(n6460) );
  OAI221_X1 U6911 ( .B1(n6474), .B2(REQUESTPENDING_REG_SCAN_IN), .C1(n6474), 
        .C2(n6461), .A(n6460), .ZN(U3181) );
  AOI221_X1 U6912 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6462), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6464) );
  AOI221_X1 U6913 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6464), .C2(HOLD), .A(n6463), .ZN(n6470) );
  AOI21_X1 U6914 ( .B1(n6466), .B2(n6465), .A(STATE_REG_2__SCAN_IN), .ZN(n6468) );
  OAI22_X1 U6915 ( .A1(n6470), .A2(n6469), .B1(n6468), .B2(n6467), .ZN(U3183)
         );
  AOI22_X1 U6916 ( .A1(n6474), .A2(n6473), .B1(n6472), .B2(n6471), .ZN(U3473)
         );
  INV_X1 U6917 ( .A(n6475), .ZN(n6684) );
  AOI22_X1 U6918 ( .A1(n6476), .A2(n6684), .B1(n6683), .B2(DATAI_16_), .ZN(
        n6478) );
  AOI22_X1 U6919 ( .A1(n6687), .A2(DATAI_0_), .B1(n6686), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6477) );
  NAND2_X1 U6920 ( .A1(n6478), .A2(n6477), .ZN(U2875) );
  AOI22_X1 U6921 ( .A1(n6479), .A2(n6684), .B1(n6683), .B2(DATAI_18_), .ZN(
        n6481) );
  AOI22_X1 U6922 ( .A1(n6687), .A2(DATAI_2_), .B1(n6686), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6480) );
  NAND2_X1 U6923 ( .A1(n6481), .A2(n6480), .ZN(U2873) );
  AOI22_X1 U6924 ( .A1(n6482), .A2(n6684), .B1(n6683), .B2(DATAI_20_), .ZN(
        n6484) );
  AOI22_X1 U6925 ( .A1(n6687), .A2(DATAI_4_), .B1(n6686), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n6483) );
  NAND2_X1 U6926 ( .A1(n6484), .A2(n6483), .ZN(U2871) );
  AOI22_X1 U6927 ( .A1(n6485), .A2(n6684), .B1(n6683), .B2(DATAI_22_), .ZN(
        n6487) );
  AOI22_X1 U6928 ( .A1(n6687), .A2(DATAI_6_), .B1(n6686), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n6486) );
  NAND2_X1 U6929 ( .A1(n6487), .A2(n6486), .ZN(U2869) );
  AND2_X1 U6930 ( .A1(n6969), .A2(DATAI_16_), .ZN(n6679) );
  INV_X1 U6931 ( .A(n6679), .ZN(n6662) );
  NAND2_X1 U6932 ( .A1(n6585), .A2(n6518), .ZN(n6561) );
  INV_X1 U6933 ( .A(n6560), .ZN(n6584) );
  NOR2_X2 U6934 ( .A1(n6488), .A2(n6963), .ZN(n6669) );
  AND2_X1 U6935 ( .A1(n6574), .A2(n6529), .ZN(n6552) );
  NOR2_X1 U6936 ( .A1(n6489), .A2(n6499), .ZN(n6967) );
  AOI21_X1 U6937 ( .B1(n6552), .B2(n6575), .A(n6967), .ZN(n6494) );
  NAND3_X1 U6938 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n6500) );
  OAI22_X1 U6939 ( .A1(n6494), .A2(n6622), .B1(n6500), .B2(n6657), .ZN(n6968)
         );
  NOR2_X2 U6940 ( .A1(n6966), .A2(n6492), .ZN(n6668) );
  AOI22_X1 U6941 ( .A1(n6669), .A2(n6968), .B1(n6668), .B2(n6967), .ZN(n6498)
         );
  AOI21_X1 U6942 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6647), .A(n6963), .ZN(
        n6653) );
  NOR2_X1 U6943 ( .A1(n6622), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6635) );
  INV_X1 U6944 ( .A(n6635), .ZN(n6527) );
  OAI21_X1 U6945 ( .B1(n6496), .B2(n6862), .A(n6527), .ZN(n6493) );
  AOI22_X1 U6946 ( .A1(n6494), .A2(n6493), .B1(n6622), .B2(n6500), .ZN(n6495)
         );
  NAND2_X1 U6947 ( .A1(n6653), .A2(n6495), .ZN(n6970) );
  AND2_X1 U6948 ( .A1(n6969), .A2(DATAI_24_), .ZN(n6648) );
  NAND2_X1 U6949 ( .A1(n6496), .A2(n6645), .ZN(n6869) );
  AOI22_X1 U6950 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n6970), .B1(n6648), 
        .B2(n6975), .ZN(n6497) );
  OAI211_X1 U6951 ( .C1(n6662), .C2(n7072), .A(n6498), .B(n6497), .ZN(U3140)
         );
  NAND2_X1 U6952 ( .A1(n6574), .A2(n6655), .ZN(n6672) );
  INV_X1 U6953 ( .A(n6575), .ZN(n6587) );
  NOR2_X1 U6954 ( .A1(n6606), .A2(n6499), .ZN(n6501) );
  INV_X1 U6955 ( .A(n6501), .ZN(n6545) );
  NAND2_X1 U6956 ( .A1(n6502), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6608) );
  OAI22_X1 U6957 ( .A1(n6672), .A2(n6587), .B1(n6545), .B2(n6608), .ZN(n6974)
         );
  NOR2_X1 U6958 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6500), .ZN(n6973)
         );
  AOI22_X1 U6959 ( .A1(n6669), .A2(n6974), .B1(n6668), .B2(n6973), .ZN(n6509)
         );
  INV_X1 U6960 ( .A(n6973), .ZN(n6504) );
  NOR2_X1 U6961 ( .A1(n6501), .A2(n6657), .ZN(n6542) );
  INV_X1 U6962 ( .A(n6502), .ZN(n6503) );
  NAND2_X1 U6963 ( .A1(n6503), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6664) );
  NAND2_X1 U6964 ( .A1(n6541), .A2(n6664), .ZN(n6612) );
  AOI211_X1 U6965 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6504), .A(n6542), .B(
        n6612), .ZN(n6507) );
  NOR2_X1 U6966 ( .A1(n6574), .A2(n6622), .ZN(n6564) );
  NOR2_X1 U6967 ( .A1(n6575), .A2(n6622), .ZN(n6589) );
  AND3_X1 U6968 ( .A1(n6585), .A2(n6583), .A3(n6560), .ZN(n6510) );
  NAND2_X1 U6969 ( .A1(n6510), .A2(n6634), .ZN(n6984) );
  OAI21_X1 U6970 ( .B1(n6975), .B2(n6913), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6505) );
  OAI21_X1 U6971 ( .B1(n6564), .B2(n6589), .A(n6505), .ZN(n6506) );
  NAND2_X1 U6972 ( .A1(n6507), .A2(n6506), .ZN(n6976) );
  AOI22_X1 U6973 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n6976), .B1(n6648), 
        .B2(n6913), .ZN(n6508) );
  OAI211_X1 U6974 ( .C1(n6662), .C2(n6869), .A(n6509), .B(n6508), .ZN(U3132)
         );
  INV_X1 U6975 ( .A(n6648), .ZN(n6682) );
  NAND3_X1 U6976 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6621), .ZN(n6517) );
  NOR2_X1 U6977 ( .A1(n6647), .A2(n6517), .ZN(n6979) );
  AOI22_X1 U6978 ( .A1(n6913), .A2(n6679), .B1(n6668), .B2(n6979), .ZN(n6516)
         );
  NAND2_X1 U6979 ( .A1(n4887), .A2(n4742), .ZN(n6611) );
  INV_X1 U6980 ( .A(n6611), .ZN(n6596) );
  AOI21_X1 U6981 ( .B1(n6552), .B2(n6596), .A(n6979), .ZN(n6513) );
  AOI21_X1 U6982 ( .B1(n6510), .B2(STATEBS16_REG_SCAN_IN), .A(n6622), .ZN(
        n6512) );
  AOI22_X1 U6983 ( .A1(n6513), .A2(n6512), .B1(n6622), .B2(n6517), .ZN(n6511)
         );
  NAND2_X1 U6984 ( .A1(n6653), .A2(n6511), .ZN(n6981) );
  INV_X1 U6985 ( .A(n6512), .ZN(n6514) );
  OAI22_X1 U6986 ( .A1(n6514), .A2(n6513), .B1(n6657), .B2(n6517), .ZN(n6980)
         );
  AOI22_X1 U6987 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n6981), .B1(n6669), 
        .B2(n6980), .ZN(n6515) );
  OAI211_X1 U6988 ( .C1(n6682), .C2(n6916), .A(n6516), .B(n6515), .ZN(U3124)
         );
  NAND2_X1 U6989 ( .A1(n6605), .A2(n6606), .ZN(n6562) );
  OAI22_X1 U6990 ( .A1(n6672), .A2(n6611), .B1(n6608), .B2(n6562), .ZN(n6986)
         );
  NOR2_X1 U6991 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6517), .ZN(n6985)
         );
  AOI22_X1 U6992 ( .A1(n6669), .A2(n6986), .B1(n6668), .B2(n6985), .ZN(n6525)
         );
  INV_X1 U6993 ( .A(n6985), .ZN(n6522) );
  NAND2_X1 U6994 ( .A1(n6537), .A2(n6518), .ZN(n6604) );
  INV_X1 U6995 ( .A(n6604), .ZN(n6519) );
  NAND2_X1 U6996 ( .A1(n6519), .A2(n6632), .ZN(n6526) );
  AOI21_X1 U6997 ( .B1(n6996), .B2(n6916), .A(n6670), .ZN(n6520) );
  AOI211_X1 U6998 ( .C1(n6596), .C2(n6610), .A(n6622), .B(n6520), .ZN(n6521)
         );
  AOI211_X1 U6999 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6522), .A(n6612), .B(
        n6521), .ZN(n6523) );
  NAND2_X1 U7000 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6562), .ZN(n6567) );
  NAND2_X1 U7001 ( .A1(n6523), .A2(n6567), .ZN(n6988) );
  INV_X1 U7002 ( .A(n6996), .ZN(n6872) );
  AOI22_X1 U7003 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n6988), .B1(n6648), 
        .B2(n6872), .ZN(n6524) );
  OAI211_X1 U7004 ( .C1(n6662), .C2(n6916), .A(n6525), .B(n6524), .ZN(U3116)
         );
  INV_X1 U7005 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6619) );
  NAND3_X1 U7006 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6619), .ZN(n6539) );
  NOR2_X1 U7007 ( .A1(n6647), .A2(n6539), .ZN(n6991) );
  AOI22_X1 U7008 ( .A1(n6998), .A2(n6648), .B1(n6668), .B2(n6991), .ZN(n6536)
         );
  INV_X1 U7009 ( .A(n6526), .ZN(n6528) );
  OAI21_X1 U7010 ( .B1(n6528), .B2(n6622), .A(n6527), .ZN(n6532) );
  OR2_X1 U7011 ( .A1(n4887), .A2(n4742), .ZN(n6630) );
  INV_X1 U7012 ( .A(n6630), .ZN(n6637) );
  NAND2_X1 U7013 ( .A1(n6637), .A2(n6574), .ZN(n6546) );
  INV_X1 U7014 ( .A(n6546), .ZN(n6530) );
  AOI21_X1 U7015 ( .B1(n6530), .B2(n6529), .A(n6991), .ZN(n6533) );
  AOI22_X1 U7016 ( .A1(n6532), .A2(n6533), .B1(n6539), .B2(n6622), .ZN(n6531)
         );
  NAND2_X1 U7017 ( .A1(n6653), .A2(n6531), .ZN(n6993) );
  INV_X1 U7018 ( .A(n6532), .ZN(n6534) );
  OAI22_X1 U7019 ( .A1(n6534), .A2(n6533), .B1(n6539), .B2(n6657), .ZN(n6992)
         );
  AOI22_X1 U7020 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6993), .B1(n6669), 
        .B2(n6992), .ZN(n6535) );
  OAI211_X1 U7021 ( .C1(n6662), .C2(n6996), .A(n6536), .B(n6535), .ZN(U3108)
         );
  NAND2_X1 U7022 ( .A1(n6537), .A2(n6583), .ZN(n6633) );
  INV_X1 U7023 ( .A(n6633), .ZN(n6538) );
  NAND2_X1 U7024 ( .A1(n6538), .A2(n6632), .ZN(n6550) );
  INV_X1 U7025 ( .A(n7009), .ZN(n6879) );
  NOR2_X1 U7026 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6539), .ZN(n6997)
         );
  AOI22_X1 U7027 ( .A1(n6879), .A2(n6648), .B1(n6668), .B2(n6997), .ZN(n6549)
         );
  AOI21_X1 U7028 ( .B1(n6924), .B2(n7009), .A(n6670), .ZN(n6540) );
  NOR2_X1 U7029 ( .A1(n6540), .A2(n6622), .ZN(n6544) );
  NAND2_X1 U7030 ( .A1(n6541), .A2(n6608), .ZN(n6640) );
  AOI211_X1 U7031 ( .C1(n6544), .C2(n6546), .A(n6640), .B(n6542), .ZN(n6543)
         );
  OAI21_X1 U7032 ( .B1(n6997), .B2(n6678), .A(n6543), .ZN(n7000) );
  INV_X1 U7033 ( .A(n6544), .ZN(n6547) );
  OAI22_X1 U7034 ( .A1(n6547), .A2(n6546), .B1(n6664), .B2(n6545), .ZN(n6999)
         );
  AOI22_X1 U7035 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n7000), .B1(n6669), 
        .B2(n6999), .ZN(n6548) );
  OAI211_X1 U7036 ( .C1(n6924), .C2(n6662), .A(n6549), .B(n6548), .ZN(U3100)
         );
  NOR3_X1 U7037 ( .A1(n6499), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6555) );
  INV_X1 U7038 ( .A(n6555), .ZN(n6563) );
  NOR2_X1 U7039 ( .A1(n6647), .A2(n6563), .ZN(n7003) );
  AOI22_X1 U7040 ( .A1(n7004), .A2(n6648), .B1(n6668), .B2(n7003), .ZN(n6559)
         );
  OAI21_X1 U7041 ( .B1(n6550), .B2(n6670), .A(n6655), .ZN(n6557) );
  INV_X1 U7042 ( .A(n6557), .ZN(n6553) );
  INV_X1 U7043 ( .A(n6665), .ZN(n6650) );
  AOI21_X1 U7044 ( .B1(n6552), .B2(n6650), .A(n7003), .ZN(n6556) );
  NAND2_X1 U7045 ( .A1(n6553), .A2(n6556), .ZN(n6554) );
  OAI211_X1 U7046 ( .C1(n6655), .C2(n6555), .A(n6653), .B(n6554), .ZN(n7006)
         );
  OAI22_X1 U7047 ( .A1(n6557), .A2(n6556), .B1(n6657), .B2(n6563), .ZN(n7005)
         );
  AOI22_X1 U7048 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n7006), .B1(n6669), 
        .B2(n7005), .ZN(n6558) );
  OAI211_X1 U7049 ( .C1(n6662), .C2(n7009), .A(n6559), .B(n6558), .ZN(U3092)
         );
  NOR2_X1 U7050 ( .A1(n6561), .A2(n6560), .ZN(n6571) );
  NAND2_X1 U7051 ( .A1(n6571), .A2(n6634), .ZN(n7023) );
  OAI22_X1 U7052 ( .A1(n6672), .A2(n6665), .B1(n6664), .B2(n6562), .ZN(n7011)
         );
  NOR2_X1 U7053 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6563), .ZN(n7010)
         );
  AOI22_X1 U7054 ( .A1(n6669), .A2(n7011), .B1(n6668), .B2(n7010), .ZN(n6570)
         );
  INV_X1 U7055 ( .A(n6564), .ZN(n6666) );
  NAND2_X1 U7056 ( .A1(n6665), .A2(n6655), .ZN(n6673) );
  AOI21_X1 U7057 ( .B1(n7016), .B2(n7023), .A(n6670), .ZN(n6565) );
  AOI21_X1 U7058 ( .B1(n6666), .B2(n6673), .A(n6565), .ZN(n6566) );
  NOR2_X1 U7059 ( .A1(n6566), .A2(n6640), .ZN(n6568) );
  OAI211_X1 U7060 ( .C1(n7010), .C2(n6678), .A(n6568), .B(n6567), .ZN(n7013)
         );
  AOI22_X1 U7061 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n7013), .B1(n6679), 
        .B2(n7004), .ZN(n6569) );
  OAI211_X1 U7062 ( .C1(n6682), .C2(n7023), .A(n6570), .B(n6569), .ZN(U3084)
         );
  INV_X1 U7063 ( .A(n6572), .ZN(n7017) );
  AOI22_X1 U7064 ( .A1(n7018), .A2(n6648), .B1(n7017), .B2(n6668), .ZN(n6582)
         );
  AOI21_X1 U7065 ( .B1(n3435), .B2(n6575), .A(n7017), .ZN(n6580) );
  NOR2_X1 U7066 ( .A1(n6576), .A2(n6622), .ZN(n6578) );
  NAND3_X1 U7067 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6499), .ZN(n6588) );
  AOI22_X1 U7068 ( .A1(n6580), .A2(n6578), .B1(n6622), .B2(n6588), .ZN(n6577)
         );
  NAND2_X1 U7069 ( .A1(n6653), .A2(n6577), .ZN(n7020) );
  INV_X1 U7070 ( .A(n6578), .ZN(n6579) );
  OAI22_X1 U7071 ( .A1(n6580), .A2(n6579), .B1(n6657), .B2(n6588), .ZN(n7019)
         );
  AOI22_X1 U7072 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n7020), .B1(n6669), 
        .B2(n7019), .ZN(n6581) );
  OAI211_X1 U7073 ( .C1(n6662), .C2(n7023), .A(n6582), .B(n6581), .ZN(U3076)
         );
  INV_X1 U7074 ( .A(n7031), .ZN(n6759) );
  INV_X1 U7075 ( .A(n6606), .ZN(n6586) );
  NAND2_X1 U7076 ( .A1(n6586), .A2(n6499), .ZN(n6629) );
  OAI22_X1 U7077 ( .A1(n6666), .A2(n6587), .B1(n6608), .B2(n6629), .ZN(n7025)
         );
  NOR2_X1 U7078 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6588), .ZN(n7024)
         );
  AOI22_X1 U7079 ( .A1(n6669), .A2(n7025), .B1(n6668), .B2(n7024), .ZN(n6595)
         );
  OAI21_X1 U7080 ( .B1(n7018), .B2(n7031), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6592) );
  INV_X1 U7081 ( .A(n6589), .ZN(n6590) );
  NAND2_X1 U7082 ( .A1(n6590), .A2(n6672), .ZN(n6591) );
  AOI21_X1 U7083 ( .B1(n6592), .B2(n6591), .A(n6612), .ZN(n6593) );
  NAND2_X1 U7084 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6629), .ZN(n6641) );
  OAI211_X1 U7085 ( .C1(n7024), .C2(n6678), .A(n6593), .B(n6641), .ZN(n7026)
         );
  AOI22_X1 U7086 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n7026), .B1(n6679), 
        .B2(n7018), .ZN(n6594) );
  OAI211_X1 U7087 ( .C1(n6682), .C2(n6759), .A(n6595), .B(n6594), .ZN(U3068)
         );
  NAND2_X1 U7088 ( .A1(n6597), .A2(n6645), .ZN(n7036) );
  NAND3_X1 U7089 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6499), .A3(n6621), .ZN(n6609) );
  NOR2_X1 U7090 ( .A1(n6647), .A2(n6609), .ZN(n7030) );
  AOI22_X1 U7091 ( .A1(n7031), .A2(n6679), .B1(n6668), .B2(n7030), .ZN(n6603)
         );
  AOI21_X1 U7092 ( .B1(n3435), .B2(n6596), .A(n7030), .ZN(n6601) );
  AOI21_X1 U7093 ( .B1(n6597), .B2(STATEBS16_REG_SCAN_IN), .A(n6622), .ZN(
        n6599) );
  AOI22_X1 U7094 ( .A1(n6601), .A2(n6599), .B1(n6622), .B2(n6609), .ZN(n6598)
         );
  NAND2_X1 U7095 ( .A1(n6653), .A2(n6598), .ZN(n7033) );
  INV_X1 U7096 ( .A(n6599), .ZN(n6600) );
  OAI22_X1 U7097 ( .A1(n6601), .A2(n6600), .B1(n6657), .B2(n6609), .ZN(n7032)
         );
  AOI22_X1 U7098 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n7033), .B1(n6669), 
        .B2(n7032), .ZN(n6602) );
  OAI211_X1 U7099 ( .C1(n6682), .C2(n7036), .A(n6603), .B(n6602), .ZN(U3060)
         );
  INV_X1 U7100 ( .A(n6605), .ZN(n6607) );
  NAND2_X1 U7101 ( .A1(n6607), .A2(n6606), .ZN(n6663) );
  OAI22_X1 U7102 ( .A1(n6666), .A2(n6611), .B1(n6608), .B2(n6663), .ZN(n7038)
         );
  NOR2_X1 U7103 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6609), .ZN(n7037)
         );
  AOI22_X1 U7104 ( .A1(n6669), .A2(n7038), .B1(n6668), .B2(n7037), .ZN(n6618)
         );
  AOI21_X1 U7105 ( .B1(n7048), .B2(n7036), .A(n6670), .ZN(n6616) );
  OAI21_X1 U7106 ( .B1(n6611), .B2(n6610), .A(n6655), .ZN(n6615) );
  INV_X1 U7107 ( .A(n7037), .ZN(n6613) );
  AND2_X1 U7108 ( .A1(n6663), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6674) );
  AOI211_X1 U7109 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6613), .A(n6674), .B(
        n6612), .ZN(n6614) );
  OAI21_X1 U7110 ( .B1(n6616), .B2(n6615), .A(n6614), .ZN(n7040) );
  AOI22_X1 U7111 ( .A1(n7040), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n7039), 
        .B2(n6679), .ZN(n6617) );
  OAI211_X1 U7112 ( .C1(n6682), .C2(n7048), .A(n6618), .B(n6617), .ZN(U3052)
         );
  NAND2_X1 U7113 ( .A1(n6499), .A2(n6619), .ZN(n6667) );
  NOR2_X1 U7114 ( .A1(n6620), .A2(n6667), .ZN(n7043) );
  AOI22_X1 U7115 ( .A1(n7051), .A2(n6648), .B1(n6668), .B2(n7043), .ZN(n6628)
         );
  AOI21_X1 U7116 ( .B1(n3435), .B2(n6637), .A(n7043), .ZN(n6625) );
  AOI21_X1 U7117 ( .B1(n3437), .B2(STATEBS16_REG_SCAN_IN), .A(n6622), .ZN(
        n6624) );
  OR2_X1 U7118 ( .A1(n6621), .A2(n6667), .ZN(n6631) );
  AOI22_X1 U7119 ( .A1(n6625), .A2(n6624), .B1(n6622), .B2(n6631), .ZN(n6623)
         );
  NAND2_X1 U7120 ( .A1(n6653), .A2(n6623), .ZN(n7045) );
  INV_X1 U7121 ( .A(n6624), .ZN(n6626) );
  OAI22_X1 U7122 ( .A1(n6626), .A2(n6625), .B1(n6657), .B2(n6631), .ZN(n7044)
         );
  AOI22_X1 U7123 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n7045), .B1(n6669), 
        .B2(n7044), .ZN(n6627) );
  OAI211_X1 U7124 ( .C1(n6662), .C2(n7048), .A(n6628), .B(n6627), .ZN(U3044)
         );
  OAI22_X1 U7125 ( .A1(n6666), .A2(n6630), .B1(n6664), .B2(n6629), .ZN(n7050)
         );
  NOR2_X1 U7126 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6631), .ZN(n7049)
         );
  AOI22_X1 U7127 ( .A1(n6669), .A2(n7050), .B1(n6668), .B2(n7049), .ZN(n6644)
         );
  AOI21_X1 U7128 ( .B1(n6947), .B2(n7062), .A(n6635), .ZN(n6636) );
  AOI21_X1 U7129 ( .B1(n6638), .B2(n6637), .A(n6636), .ZN(n6639) );
  NOR2_X1 U7130 ( .A1(n6639), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6642) );
  INV_X1 U7131 ( .A(n6640), .ZN(n6677) );
  OAI211_X1 U7132 ( .C1(n6642), .C2(n7049), .A(n6641), .B(n6677), .ZN(n7052)
         );
  INV_X1 U7133 ( .A(n7062), .ZN(n6898) );
  AOI22_X1 U7134 ( .A1(INSTQUEUE_REG_2__0__SCAN_IN), .A2(n7052), .B1(n6648), 
        .B2(n6898), .ZN(n6643) );
  OAI211_X1 U7135 ( .C1(n6662), .C2(n6947), .A(n6644), .B(n6643), .ZN(U3036)
         );
  NAND2_X1 U7136 ( .A1(n6646), .A2(n6645), .ZN(n6956) );
  NOR2_X1 U7137 ( .A1(n6667), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6654)
         );
  INV_X1 U7138 ( .A(n6654), .ZN(n6656) );
  NOR2_X1 U7139 ( .A1(n6647), .A2(n6656), .ZN(n7055) );
  AOI22_X1 U7140 ( .A1(n7067), .A2(n6648), .B1(n6668), .B2(n7055), .ZN(n6661)
         );
  OAI21_X1 U7141 ( .B1(n6649), .B2(n6670), .A(n6655), .ZN(n6658) );
  INV_X1 U7142 ( .A(n6658), .ZN(n6651) );
  AOI21_X1 U7143 ( .B1(n3435), .B2(n6650), .A(n7055), .ZN(n6659) );
  NAND2_X1 U7144 ( .A1(n6651), .A2(n6659), .ZN(n6652) );
  OAI211_X1 U7145 ( .C1(n6655), .C2(n6654), .A(n6653), .B(n6652), .ZN(n7058)
         );
  OAI22_X1 U7146 ( .A1(n6659), .A2(n6658), .B1(n6657), .B2(n6656), .ZN(n7057)
         );
  AOI22_X1 U7147 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n7058), .B1(n6669), 
        .B2(n7057), .ZN(n6660) );
  OAI211_X1 U7148 ( .C1(n6662), .C2(n7062), .A(n6661), .B(n6660), .ZN(U3028)
         );
  OAI22_X1 U7149 ( .A1(n6666), .A2(n6665), .B1(n6664), .B2(n6663), .ZN(n7065)
         );
  AOI22_X1 U7150 ( .A1(n6669), .A2(n7065), .B1(n6668), .B2(n7063), .ZN(n6681)
         );
  AOI21_X1 U7151 ( .B1(n6956), .B2(n7072), .A(n6670), .ZN(n6671) );
  AOI21_X1 U7152 ( .B1(n6673), .B2(n6672), .A(n6671), .ZN(n6675) );
  NOR2_X1 U7153 ( .A1(n6675), .A2(n6674), .ZN(n6676) );
  OAI211_X1 U7154 ( .C1(n7063), .C2(n6678), .A(n6677), .B(n6676), .ZN(n7069)
         );
  AOI22_X1 U7155 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n7069), .B1(n6679), 
        .B2(n7067), .ZN(n6680) );
  OAI211_X1 U7156 ( .C1(n6682), .C2(n7072), .A(n6681), .B(n6680), .ZN(U3020)
         );
  AOI22_X1 U7157 ( .A1(n6685), .A2(n6684), .B1(n6683), .B2(DATAI_24_), .ZN(
        n6689) );
  AOI22_X1 U7158 ( .A1(n6687), .A2(DATAI_8_), .B1(n6686), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n6688) );
  NAND2_X1 U7159 ( .A1(n6689), .A2(n6688), .ZN(U2867) );
  AND2_X1 U7160 ( .A1(n6969), .A2(DATAI_17_), .ZN(n6727) );
  INV_X1 U7161 ( .A(n6727), .ZN(n6720) );
  NOR2_X2 U7162 ( .A1(n6690), .A2(n6963), .ZN(n6726) );
  NOR2_X2 U7163 ( .A1(n6966), .A2(n6691), .ZN(n6725) );
  AOI22_X1 U7164 ( .A1(n6726), .A2(n6968), .B1(n6725), .B2(n6967), .ZN(n6694)
         );
  NOR2_X1 U7165 ( .A1(n6862), .A2(n6692), .ZN(n6717) );
  AOI22_X1 U7166 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n6970), .B1(n6717), 
        .B2(n6975), .ZN(n6693) );
  OAI211_X1 U7167 ( .C1(n6720), .C2(n7072), .A(n6694), .B(n6693), .ZN(U3141)
         );
  INV_X1 U7168 ( .A(n6717), .ZN(n6730) );
  AOI22_X1 U7169 ( .A1(n6726), .A2(n6974), .B1(n6725), .B2(n6973), .ZN(n6696)
         );
  AOI22_X1 U7170 ( .A1(INSTQUEUE_REG_14__1__SCAN_IN), .A2(n6976), .B1(n6727), 
        .B2(n6975), .ZN(n6695) );
  OAI211_X1 U7171 ( .C1(n6730), .C2(n6984), .A(n6696), .B(n6695), .ZN(U3133)
         );
  AOI22_X1 U7172 ( .A1(n6987), .A2(n6717), .B1(n6725), .B2(n6979), .ZN(n6698)
         );
  AOI22_X1 U7173 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n6981), .B1(n6726), 
        .B2(n6980), .ZN(n6697) );
  OAI211_X1 U7174 ( .C1(n6720), .C2(n6984), .A(n6698), .B(n6697), .ZN(U3125)
         );
  AOI22_X1 U7175 ( .A1(n6726), .A2(n6986), .B1(n6725), .B2(n6985), .ZN(n6700)
         );
  AOI22_X1 U7176 ( .A1(INSTQUEUE_REG_12__1__SCAN_IN), .A2(n6988), .B1(n6727), 
        .B2(n6987), .ZN(n6699) );
  OAI211_X1 U7177 ( .C1(n6730), .C2(n6996), .A(n6700), .B(n6699), .ZN(U3117)
         );
  AOI22_X1 U7178 ( .A1(n6872), .A2(n6727), .B1(n6725), .B2(n6991), .ZN(n6702)
         );
  AOI22_X1 U7179 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6993), .B1(n6726), 
        .B2(n6992), .ZN(n6701) );
  OAI211_X1 U7180 ( .C1(n6924), .C2(n6730), .A(n6702), .B(n6701), .ZN(U3109)
         );
  AOI22_X1 U7181 ( .A1(n6998), .A2(n6727), .B1(n6725), .B2(n6997), .ZN(n6704)
         );
  AOI22_X1 U7182 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(n7000), .B1(n6726), 
        .B2(n6999), .ZN(n6703) );
  OAI211_X1 U7183 ( .C1(n7009), .C2(n6730), .A(n6704), .B(n6703), .ZN(U3101)
         );
  AOI22_X1 U7184 ( .A1(n7004), .A2(n6717), .B1(n6725), .B2(n7003), .ZN(n6706)
         );
  AOI22_X1 U7185 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n7006), .B1(n6726), 
        .B2(n7005), .ZN(n6705) );
  OAI211_X1 U7186 ( .C1(n7009), .C2(n6720), .A(n6706), .B(n6705), .ZN(U3093)
         );
  AOI22_X1 U7187 ( .A1(n6726), .A2(n7011), .B1(n6725), .B2(n7010), .ZN(n6708)
         );
  AOI22_X1 U7188 ( .A1(INSTQUEUE_REG_8__1__SCAN_IN), .A2(n7013), .B1(n6727), 
        .B2(n7004), .ZN(n6707) );
  OAI211_X1 U7189 ( .C1(n6730), .C2(n7023), .A(n6708), .B(n6707), .ZN(U3085)
         );
  AOI22_X1 U7190 ( .A1(n7018), .A2(n6717), .B1(n7017), .B2(n6725), .ZN(n6710)
         );
  AOI22_X1 U7191 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n7020), .B1(n6726), 
        .B2(n7019), .ZN(n6709) );
  OAI211_X1 U7192 ( .C1(n6720), .C2(n7023), .A(n6710), .B(n6709), .ZN(U3077)
         );
  AOI22_X1 U7193 ( .A1(n6726), .A2(n7025), .B1(n6725), .B2(n7024), .ZN(n6712)
         );
  AOI22_X1 U7194 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(n7026), .B1(n6727), 
        .B2(n7018), .ZN(n6711) );
  OAI211_X1 U7195 ( .C1(n6730), .C2(n6759), .A(n6712), .B(n6711), .ZN(U3069)
         );
  AOI22_X1 U7196 ( .A1(n7031), .A2(n6727), .B1(n6725), .B2(n7030), .ZN(n6714)
         );
  AOI22_X1 U7197 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n7033), .B1(n6726), 
        .B2(n7032), .ZN(n6713) );
  OAI211_X1 U7198 ( .C1(n6730), .C2(n7036), .A(n6714), .B(n6713), .ZN(U3061)
         );
  AOI22_X1 U7199 ( .A1(n6726), .A2(n7038), .B1(n6725), .B2(n7037), .ZN(n6716)
         );
  AOI22_X1 U7200 ( .A1(n7040), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n7039), 
        .B2(n6727), .ZN(n6715) );
  OAI211_X1 U7201 ( .C1(n6730), .C2(n7048), .A(n6716), .B(n6715), .ZN(U3053)
         );
  AOI22_X1 U7202 ( .A1(n7051), .A2(n6717), .B1(n6725), .B2(n7043), .ZN(n6719)
         );
  AOI22_X1 U7203 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n7045), .B1(n6726), 
        .B2(n7044), .ZN(n6718) );
  OAI211_X1 U7204 ( .C1(n6720), .C2(n7048), .A(n6719), .B(n6718), .ZN(U3045)
         );
  AOI22_X1 U7205 ( .A1(n6726), .A2(n7050), .B1(n6725), .B2(n7049), .ZN(n6722)
         );
  AOI22_X1 U7206 ( .A1(INSTQUEUE_REG_2__1__SCAN_IN), .A2(n7052), .B1(n7051), 
        .B2(n6727), .ZN(n6721) );
  OAI211_X1 U7207 ( .C1(n7062), .C2(n6730), .A(n6722), .B(n6721), .ZN(U3037)
         );
  AOI22_X1 U7208 ( .A1(n6898), .A2(n6727), .B1(n6725), .B2(n7055), .ZN(n6724)
         );
  AOI22_X1 U7209 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n7058), .B1(n6726), 
        .B2(n7057), .ZN(n6723) );
  OAI211_X1 U7210 ( .C1(n6730), .C2(n6956), .A(n6724), .B(n6723), .ZN(U3029)
         );
  AOI22_X1 U7211 ( .A1(n6726), .A2(n7065), .B1(n6725), .B2(n7063), .ZN(n6729)
         );
  AOI22_X1 U7212 ( .A1(INSTQUEUE_REG_0__1__SCAN_IN), .A2(n7069), .B1(n6727), 
        .B2(n7067), .ZN(n6728) );
  OAI211_X1 U7213 ( .C1(n6730), .C2(n7072), .A(n6729), .B(n6728), .ZN(U3021)
         );
  AND2_X1 U7214 ( .A1(n6969), .A2(DATAI_26_), .ZN(n6765) );
  INV_X1 U7215 ( .A(n6765), .ZN(n6778) );
  NOR2_X2 U7216 ( .A1(n6731), .A2(n6963), .ZN(n6774) );
  NOR2_X1 U7217 ( .A1(n6966), .A2(n6732), .ZN(n6773) );
  AOI22_X1 U7218 ( .A1(n6774), .A2(n6968), .B1(n6773), .B2(n6967), .ZN(n6735)
         );
  AND2_X1 U7219 ( .A1(n6969), .A2(DATAI_18_), .ZN(n6775) );
  INV_X1 U7220 ( .A(n7072), .ZN(n6733) );
  AOI22_X1 U7221 ( .A1(INSTQUEUE_REG_15__2__SCAN_IN), .A2(n6970), .B1(n6775), 
        .B2(n6733), .ZN(n6734) );
  OAI211_X1 U7222 ( .C1(n6778), .C2(n6869), .A(n6735), .B(n6734), .ZN(U3142)
         );
  INV_X1 U7223 ( .A(n6775), .ZN(n6769) );
  AOI22_X1 U7224 ( .A1(n6774), .A2(n6974), .B1(n6773), .B2(n6973), .ZN(n6737)
         );
  AOI22_X1 U7225 ( .A1(INSTQUEUE_REG_14__2__SCAN_IN), .A2(n6976), .B1(n6765), 
        .B2(n6913), .ZN(n6736) );
  OAI211_X1 U7226 ( .C1(n6769), .C2(n6869), .A(n6737), .B(n6736), .ZN(U3134)
         );
  AOI22_X1 U7227 ( .A1(n6913), .A2(n6775), .B1(n6773), .B2(n6979), .ZN(n6739)
         );
  AOI22_X1 U7228 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n6981), .B1(n6774), 
        .B2(n6980), .ZN(n6738) );
  OAI211_X1 U7229 ( .C1(n6778), .C2(n6916), .A(n6739), .B(n6738), .ZN(U3126)
         );
  AOI22_X1 U7230 ( .A1(n6774), .A2(n6986), .B1(n6773), .B2(n6985), .ZN(n6741)
         );
  AOI22_X1 U7231 ( .A1(INSTQUEUE_REG_12__2__SCAN_IN), .A2(n6988), .B1(n6765), 
        .B2(n6872), .ZN(n6740) );
  OAI211_X1 U7232 ( .C1(n6769), .C2(n6916), .A(n6741), .B(n6740), .ZN(U3118)
         );
  INV_X1 U7233 ( .A(n6773), .ZN(n6768) );
  INV_X1 U7234 ( .A(n6991), .ZN(n6919) );
  OAI22_X1 U7235 ( .A1(n6996), .A2(n6769), .B1(n6768), .B2(n6919), .ZN(n6742)
         );
  INV_X1 U7236 ( .A(n6742), .ZN(n6744) );
  AOI22_X1 U7237 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6993), .B1(n6774), 
        .B2(n6992), .ZN(n6743) );
  OAI211_X1 U7238 ( .C1(n6924), .C2(n6778), .A(n6744), .B(n6743), .ZN(U3110)
         );
  INV_X1 U7239 ( .A(n6997), .ZN(n6923) );
  OAI22_X1 U7240 ( .A1(n7009), .A2(n6778), .B1(n6768), .B2(n6923), .ZN(n6745)
         );
  INV_X1 U7241 ( .A(n6745), .ZN(n6747) );
  AOI22_X1 U7242 ( .A1(INSTQUEUE_REG_10__2__SCAN_IN), .A2(n7000), .B1(n6774), 
        .B2(n6999), .ZN(n6746) );
  OAI211_X1 U7243 ( .C1(n6924), .C2(n6769), .A(n6747), .B(n6746), .ZN(U3102)
         );
  INV_X1 U7244 ( .A(n7003), .ZN(n6928) );
  OAI22_X1 U7245 ( .A1(n7016), .A2(n6778), .B1(n6768), .B2(n6928), .ZN(n6748)
         );
  INV_X1 U7246 ( .A(n6748), .ZN(n6750) );
  AOI22_X1 U7247 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n7006), .B1(n6774), 
        .B2(n7005), .ZN(n6749) );
  OAI211_X1 U7248 ( .C1(n7009), .C2(n6769), .A(n6750), .B(n6749), .ZN(U3094)
         );
  AOI22_X1 U7249 ( .A1(n6774), .A2(n7011), .B1(n6773), .B2(n7010), .ZN(n6752)
         );
  AOI22_X1 U7250 ( .A1(INSTQUEUE_REG_8__2__SCAN_IN), .A2(n7013), .B1(n6775), 
        .B2(n7004), .ZN(n6751) );
  OAI211_X1 U7251 ( .C1(n6778), .C2(n7023), .A(n6752), .B(n6751), .ZN(U3086)
         );
  AOI22_X1 U7252 ( .A1(n7012), .A2(n6775), .B1(n7017), .B2(n6773), .ZN(n6754)
         );
  AOI22_X1 U7253 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n7020), .B1(n6774), 
        .B2(n7019), .ZN(n6753) );
  OAI211_X1 U7254 ( .C1(n6778), .C2(n7029), .A(n6754), .B(n6753), .ZN(U3078)
         );
  AOI22_X1 U7255 ( .A1(n6774), .A2(n7025), .B1(n6773), .B2(n7024), .ZN(n6756)
         );
  AOI22_X1 U7256 ( .A1(INSTQUEUE_REG_6__2__SCAN_IN), .A2(n7026), .B1(n6765), 
        .B2(n7031), .ZN(n6755) );
  OAI211_X1 U7257 ( .C1(n6769), .C2(n7029), .A(n6756), .B(n6755), .ZN(U3070)
         );
  AOI22_X1 U7258 ( .A1(n7039), .A2(n6765), .B1(n6773), .B2(n7030), .ZN(n6758)
         );
  AOI22_X1 U7259 ( .A1(INSTQUEUE_REG_5__2__SCAN_IN), .A2(n7033), .B1(n6774), 
        .B2(n7032), .ZN(n6757) );
  OAI211_X1 U7260 ( .C1(n6769), .C2(n6759), .A(n6758), .B(n6757), .ZN(U3062)
         );
  AOI22_X1 U7261 ( .A1(n6774), .A2(n7038), .B1(n6773), .B2(n7037), .ZN(n6761)
         );
  AOI22_X1 U7262 ( .A1(n7040), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n7039), 
        .B2(n6775), .ZN(n6760) );
  OAI211_X1 U7263 ( .C1(n6778), .C2(n7048), .A(n6761), .B(n6760), .ZN(U3054)
         );
  INV_X1 U7264 ( .A(n7043), .ZN(n6943) );
  OAI22_X1 U7265 ( .A1(n6947), .A2(n6778), .B1(n6768), .B2(n6943), .ZN(n6762)
         );
  INV_X1 U7266 ( .A(n6762), .ZN(n6764) );
  AOI22_X1 U7267 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n7045), .B1(n6774), 
        .B2(n7044), .ZN(n6763) );
  OAI211_X1 U7268 ( .C1(n6769), .C2(n7048), .A(n6764), .B(n6763), .ZN(U3046)
         );
  AOI22_X1 U7269 ( .A1(n6774), .A2(n7050), .B1(n6773), .B2(n7049), .ZN(n6767)
         );
  AOI22_X1 U7270 ( .A1(INSTQUEUE_REG_2__2__SCAN_IN), .A2(n7052), .B1(n6898), 
        .B2(n6765), .ZN(n6766) );
  OAI211_X1 U7271 ( .C1(n6947), .C2(n6769), .A(n6767), .B(n6766), .ZN(U3038)
         );
  INV_X1 U7272 ( .A(n7055), .ZN(n6950) );
  OAI22_X1 U7273 ( .A1(n7062), .A2(n6769), .B1(n6768), .B2(n6950), .ZN(n6770)
         );
  INV_X1 U7274 ( .A(n6770), .ZN(n6772) );
  AOI22_X1 U7275 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n7058), .B1(n6774), 
        .B2(n7057), .ZN(n6771) );
  OAI211_X1 U7276 ( .C1(n6778), .C2(n6956), .A(n6772), .B(n6771), .ZN(U3030)
         );
  AOI22_X1 U7277 ( .A1(n6774), .A2(n7065), .B1(n6773), .B2(n7063), .ZN(n6777)
         );
  AOI22_X1 U7278 ( .A1(INSTQUEUE_REG_0__2__SCAN_IN), .A2(n7069), .B1(n6775), 
        .B2(n7067), .ZN(n6776) );
  OAI211_X1 U7279 ( .C1(n6778), .C2(n7072), .A(n6777), .B(n6776), .ZN(U3022)
         );
  AND2_X1 U7280 ( .A1(n6969), .A2(DATAI_19_), .ZN(n6817) );
  INV_X1 U7281 ( .A(n6817), .ZN(n6814) );
  NOR2_X2 U7282 ( .A1(n6779), .A2(n6963), .ZN(n6816) );
  NOR2_X2 U7283 ( .A1(n6966), .A2(n6780), .ZN(n6815) );
  AOI22_X1 U7284 ( .A1(n6816), .A2(n6968), .B1(n6815), .B2(n6967), .ZN(n6783)
         );
  NOR2_X1 U7285 ( .A1(n6862), .A2(n6781), .ZN(n6811) );
  AOI22_X1 U7286 ( .A1(INSTQUEUE_REG_15__3__SCAN_IN), .A2(n6970), .B1(n6811), 
        .B2(n6975), .ZN(n6782) );
  OAI211_X1 U7287 ( .C1(n6814), .C2(n7072), .A(n6783), .B(n6782), .ZN(U3143)
         );
  INV_X1 U7288 ( .A(n6811), .ZN(n6820) );
  AOI22_X1 U7289 ( .A1(n6816), .A2(n6974), .B1(n6815), .B2(n6973), .ZN(n6785)
         );
  AOI22_X1 U7290 ( .A1(INSTQUEUE_REG_14__3__SCAN_IN), .A2(n6976), .B1(n6817), 
        .B2(n6975), .ZN(n6784) );
  OAI211_X1 U7291 ( .C1(n6820), .C2(n6984), .A(n6785), .B(n6784), .ZN(U3135)
         );
  AOI22_X1 U7292 ( .A1(n6987), .A2(n6811), .B1(n6815), .B2(n6979), .ZN(n6787)
         );
  AOI22_X1 U7293 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n6981), .B1(n6816), 
        .B2(n6980), .ZN(n6786) );
  OAI211_X1 U7294 ( .C1(n6814), .C2(n6984), .A(n6787), .B(n6786), .ZN(U3127)
         );
  AOI22_X1 U7295 ( .A1(n6816), .A2(n6986), .B1(n6815), .B2(n6985), .ZN(n6789)
         );
  AOI22_X1 U7296 ( .A1(INSTQUEUE_REG_12__3__SCAN_IN), .A2(n6988), .B1(n6817), 
        .B2(n6987), .ZN(n6788) );
  OAI211_X1 U7297 ( .C1(n6820), .C2(n6996), .A(n6789), .B(n6788), .ZN(U3119)
         );
  AOI22_X1 U7298 ( .A1(n6872), .A2(n6817), .B1(n6815), .B2(n6991), .ZN(n6791)
         );
  AOI22_X1 U7299 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6993), .B1(n6816), 
        .B2(n6992), .ZN(n6790) );
  OAI211_X1 U7300 ( .C1(n6924), .C2(n6820), .A(n6791), .B(n6790), .ZN(U3111)
         );
  AOI22_X1 U7301 ( .A1(n6998), .A2(n6817), .B1(n6815), .B2(n6997), .ZN(n6793)
         );
  AOI22_X1 U7302 ( .A1(INSTQUEUE_REG_10__3__SCAN_IN), .A2(n7000), .B1(n6816), 
        .B2(n6999), .ZN(n6792) );
  OAI211_X1 U7303 ( .C1(n7009), .C2(n6820), .A(n6793), .B(n6792), .ZN(U3103)
         );
  AOI22_X1 U7304 ( .A1(n6879), .A2(n6817), .B1(n6815), .B2(n7003), .ZN(n6795)
         );
  AOI22_X1 U7305 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n7006), .B1(n6816), 
        .B2(n7005), .ZN(n6794) );
  OAI211_X1 U7306 ( .C1(n6820), .C2(n7016), .A(n6795), .B(n6794), .ZN(U3095)
         );
  AOI22_X1 U7307 ( .A1(n6816), .A2(n7011), .B1(n6815), .B2(n7010), .ZN(n6797)
         );
  AOI22_X1 U7308 ( .A1(INSTQUEUE_REG_8__3__SCAN_IN), .A2(n7013), .B1(n6811), 
        .B2(n7012), .ZN(n6796) );
  OAI211_X1 U7309 ( .C1(n6814), .C2(n7016), .A(n6797), .B(n6796), .ZN(U3087)
         );
  AOI22_X1 U7310 ( .A1(n7018), .A2(n6811), .B1(n7017), .B2(n6815), .ZN(n6799)
         );
  AOI22_X1 U7311 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n7020), .B1(n6816), 
        .B2(n7019), .ZN(n6798) );
  OAI211_X1 U7312 ( .C1(n6814), .C2(n7023), .A(n6799), .B(n6798), .ZN(U3079)
         );
  AOI22_X1 U7313 ( .A1(n6816), .A2(n7025), .B1(n6815), .B2(n7024), .ZN(n6801)
         );
  AOI22_X1 U7314 ( .A1(INSTQUEUE_REG_6__3__SCAN_IN), .A2(n7026), .B1(n6811), 
        .B2(n7031), .ZN(n6800) );
  OAI211_X1 U7315 ( .C1(n6814), .C2(n7029), .A(n6801), .B(n6800), .ZN(U3071)
         );
  AOI22_X1 U7316 ( .A1(n7031), .A2(n6817), .B1(n6815), .B2(n7030), .ZN(n6803)
         );
  AOI22_X1 U7317 ( .A1(INSTQUEUE_REG_5__3__SCAN_IN), .A2(n7033), .B1(n6816), 
        .B2(n7032), .ZN(n6802) );
  OAI211_X1 U7318 ( .C1(n6820), .C2(n7036), .A(n6803), .B(n6802), .ZN(U3063)
         );
  AOI22_X1 U7319 ( .A1(n6816), .A2(n7038), .B1(n6815), .B2(n7037), .ZN(n6805)
         );
  AOI22_X1 U7320 ( .A1(n7040), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n7039), 
        .B2(n6817), .ZN(n6804) );
  OAI211_X1 U7321 ( .C1(n6820), .C2(n7048), .A(n6805), .B(n6804), .ZN(U3055)
         );
  INV_X1 U7322 ( .A(n7048), .ZN(n6806) );
  AOI22_X1 U7323 ( .A1(n6806), .A2(n6817), .B1(n6815), .B2(n7043), .ZN(n6808)
         );
  AOI22_X1 U7324 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n7045), .B1(n6816), 
        .B2(n7044), .ZN(n6807) );
  OAI211_X1 U7325 ( .C1(n6947), .C2(n6820), .A(n6808), .B(n6807), .ZN(U3047)
         );
  AOI22_X1 U7326 ( .A1(n6816), .A2(n7050), .B1(n6815), .B2(n7049), .ZN(n6810)
         );
  AOI22_X1 U7327 ( .A1(INSTQUEUE_REG_2__3__SCAN_IN), .A2(n7052), .B1(n7051), 
        .B2(n6817), .ZN(n6809) );
  OAI211_X1 U7328 ( .C1(n7062), .C2(n6820), .A(n6810), .B(n6809), .ZN(U3039)
         );
  AOI22_X1 U7329 ( .A1(n7067), .A2(n6811), .B1(n6815), .B2(n7055), .ZN(n6813)
         );
  AOI22_X1 U7330 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n7058), .B1(n6816), 
        .B2(n7057), .ZN(n6812) );
  OAI211_X1 U7331 ( .C1(n7062), .C2(n6814), .A(n6813), .B(n6812), .ZN(U3031)
         );
  AOI22_X1 U7332 ( .A1(n6816), .A2(n7065), .B1(n6815), .B2(n7063), .ZN(n6819)
         );
  AOI22_X1 U7333 ( .A1(INSTQUEUE_REG_0__3__SCAN_IN), .A2(n7069), .B1(n6817), 
        .B2(n7067), .ZN(n6818) );
  OAI211_X1 U7334 ( .C1(n6820), .C2(n7072), .A(n6819), .B(n6818), .ZN(U3023)
         );
  AND2_X1 U7335 ( .A1(n6969), .A2(DATAI_20_), .ZN(n6857) );
  INV_X1 U7336 ( .A(n6857), .ZN(n6854) );
  NOR2_X2 U7337 ( .A1(n6821), .A2(n6963), .ZN(n6856) );
  NOR2_X2 U7338 ( .A1(n6966), .A2(n6822), .ZN(n6855) );
  AOI22_X1 U7339 ( .A1(n6856), .A2(n6968), .B1(n6855), .B2(n6967), .ZN(n6824)
         );
  AND2_X1 U7340 ( .A1(n6969), .A2(DATAI_28_), .ZN(n6851) );
  AOI22_X1 U7341 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n6970), .B1(n6851), 
        .B2(n6975), .ZN(n6823) );
  OAI211_X1 U7342 ( .C1(n6854), .C2(n7072), .A(n6824), .B(n6823), .ZN(U3144)
         );
  INV_X1 U7343 ( .A(n6851), .ZN(n6860) );
  AOI22_X1 U7344 ( .A1(n6856), .A2(n6974), .B1(n6855), .B2(n6973), .ZN(n6826)
         );
  AOI22_X1 U7345 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n6976), .B1(n6857), 
        .B2(n6975), .ZN(n6825) );
  OAI211_X1 U7346 ( .C1(n6860), .C2(n6984), .A(n6826), .B(n6825), .ZN(U3136)
         );
  AOI22_X1 U7347 ( .A1(n6913), .A2(n6857), .B1(n6855), .B2(n6979), .ZN(n6828)
         );
  AOI22_X1 U7348 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n6981), .B1(n6856), 
        .B2(n6980), .ZN(n6827) );
  OAI211_X1 U7349 ( .C1(n6860), .C2(n6916), .A(n6828), .B(n6827), .ZN(U3128)
         );
  AOI22_X1 U7350 ( .A1(n6856), .A2(n6986), .B1(n6855), .B2(n6985), .ZN(n6830)
         );
  AOI22_X1 U7351 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n6988), .B1(n6857), 
        .B2(n6987), .ZN(n6829) );
  OAI211_X1 U7352 ( .C1(n6860), .C2(n6996), .A(n6830), .B(n6829), .ZN(U3120)
         );
  AOI22_X1 U7353 ( .A1(n6998), .A2(n6851), .B1(n6855), .B2(n6991), .ZN(n6832)
         );
  AOI22_X1 U7354 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6993), .B1(n6856), 
        .B2(n6992), .ZN(n6831) );
  OAI211_X1 U7355 ( .C1(n6854), .C2(n6996), .A(n6832), .B(n6831), .ZN(U3112)
         );
  AOI22_X1 U7356 ( .A1(n6998), .A2(n6857), .B1(n6855), .B2(n6997), .ZN(n6834)
         );
  AOI22_X1 U7357 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n7000), .B1(n6856), 
        .B2(n6999), .ZN(n6833) );
  OAI211_X1 U7358 ( .C1(n7009), .C2(n6860), .A(n6834), .B(n6833), .ZN(U3104)
         );
  AOI22_X1 U7359 ( .A1(n6879), .A2(n6857), .B1(n6855), .B2(n7003), .ZN(n6836)
         );
  AOI22_X1 U7360 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n7006), .B1(n6856), 
        .B2(n7005), .ZN(n6835) );
  OAI211_X1 U7361 ( .C1(n6860), .C2(n7016), .A(n6836), .B(n6835), .ZN(U3096)
         );
  AOI22_X1 U7362 ( .A1(n6856), .A2(n7011), .B1(n6855), .B2(n7010), .ZN(n6838)
         );
  AOI22_X1 U7363 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n7013), .B1(n6851), 
        .B2(n7012), .ZN(n6837) );
  OAI211_X1 U7364 ( .C1(n6854), .C2(n7016), .A(n6838), .B(n6837), .ZN(U3088)
         );
  AOI22_X1 U7365 ( .A1(n7018), .A2(n6851), .B1(n7017), .B2(n6855), .ZN(n6840)
         );
  AOI22_X1 U7366 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n7020), .B1(n6856), 
        .B2(n7019), .ZN(n6839) );
  OAI211_X1 U7367 ( .C1(n6854), .C2(n7023), .A(n6840), .B(n6839), .ZN(U3080)
         );
  AOI22_X1 U7368 ( .A1(n6856), .A2(n7025), .B1(n6855), .B2(n7024), .ZN(n6842)
         );
  AOI22_X1 U7369 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n7026), .B1(n6851), 
        .B2(n7031), .ZN(n6841) );
  OAI211_X1 U7370 ( .C1(n6854), .C2(n7029), .A(n6842), .B(n6841), .ZN(U3072)
         );
  AOI22_X1 U7371 ( .A1(n7031), .A2(n6857), .B1(n6855), .B2(n7030), .ZN(n6844)
         );
  AOI22_X1 U7372 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n7033), .B1(n6856), 
        .B2(n7032), .ZN(n6843) );
  OAI211_X1 U7373 ( .C1(n6860), .C2(n7036), .A(n6844), .B(n6843), .ZN(U3064)
         );
  AOI22_X1 U7374 ( .A1(n6856), .A2(n7038), .B1(n6855), .B2(n7037), .ZN(n6846)
         );
  AOI22_X1 U7375 ( .A1(n7040), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n7039), 
        .B2(n6857), .ZN(n6845) );
  OAI211_X1 U7376 ( .C1(n6860), .C2(n7048), .A(n6846), .B(n6845), .ZN(U3056)
         );
  AOI22_X1 U7377 ( .A1(n7051), .A2(n6851), .B1(n6855), .B2(n7043), .ZN(n6848)
         );
  AOI22_X1 U7378 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n7045), .B1(n6856), 
        .B2(n7044), .ZN(n6847) );
  OAI211_X1 U7379 ( .C1(n6854), .C2(n7048), .A(n6848), .B(n6847), .ZN(U3048)
         );
  AOI22_X1 U7380 ( .A1(n6856), .A2(n7050), .B1(n6855), .B2(n7049), .ZN(n6850)
         );
  AOI22_X1 U7381 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n7052), .B1(n7051), 
        .B2(n6857), .ZN(n6849) );
  OAI211_X1 U7382 ( .C1(n7062), .C2(n6860), .A(n6850), .B(n6849), .ZN(U3040)
         );
  AOI22_X1 U7383 ( .A1(n7067), .A2(n6851), .B1(n6855), .B2(n7055), .ZN(n6853)
         );
  AOI22_X1 U7384 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n7058), .B1(n6856), 
        .B2(n7057), .ZN(n6852) );
  OAI211_X1 U7385 ( .C1(n7062), .C2(n6854), .A(n6853), .B(n6852), .ZN(U3032)
         );
  AOI22_X1 U7386 ( .A1(n6856), .A2(n7065), .B1(n6855), .B2(n7063), .ZN(n6859)
         );
  AOI22_X1 U7387 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n7069), .B1(n6857), 
        .B2(n7067), .ZN(n6858) );
  OAI211_X1 U7388 ( .C1(n6860), .C2(n7072), .A(n6859), .B(n6858), .ZN(U3024)
         );
  NOR2_X1 U7389 ( .A1(n6862), .A2(n6861), .ZN(n6903) );
  INV_X1 U7390 ( .A(n6903), .ZN(n6897) );
  NOR2_X2 U7391 ( .A1(n6863), .A2(n6963), .ZN(n6902) );
  NOR2_X2 U7392 ( .A1(n6966), .A2(n6864), .ZN(n6901) );
  AOI22_X1 U7393 ( .A1(n6902), .A2(n6968), .B1(n6901), .B2(n6967), .ZN(n6866)
         );
  AND2_X1 U7394 ( .A1(n6969), .A2(DATAI_29_), .ZN(n6894) );
  AOI22_X1 U7395 ( .A1(INSTQUEUE_REG_15__5__SCAN_IN), .A2(n6970), .B1(n6894), 
        .B2(n6975), .ZN(n6865) );
  OAI211_X1 U7396 ( .C1(n6897), .C2(n7072), .A(n6866), .B(n6865), .ZN(U3145)
         );
  AOI22_X1 U7397 ( .A1(n6902), .A2(n6974), .B1(n6901), .B2(n6973), .ZN(n6868)
         );
  AOI22_X1 U7398 ( .A1(INSTQUEUE_REG_14__5__SCAN_IN), .A2(n6976), .B1(n6894), 
        .B2(n6913), .ZN(n6867) );
  OAI211_X1 U7399 ( .C1(n6897), .C2(n6869), .A(n6868), .B(n6867), .ZN(U3137)
         );
  INV_X1 U7400 ( .A(n6894), .ZN(n6906) );
  AOI22_X1 U7401 ( .A1(n6913), .A2(n6903), .B1(n6901), .B2(n6979), .ZN(n6871)
         );
  AOI22_X1 U7402 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n6981), .B1(n6902), 
        .B2(n6980), .ZN(n6870) );
  OAI211_X1 U7403 ( .C1(n6906), .C2(n6916), .A(n6871), .B(n6870), .ZN(U3129)
         );
  AOI22_X1 U7404 ( .A1(n6902), .A2(n6986), .B1(n6901), .B2(n6985), .ZN(n6874)
         );
  AOI22_X1 U7405 ( .A1(INSTQUEUE_REG_12__5__SCAN_IN), .A2(n6988), .B1(n6894), 
        .B2(n6872), .ZN(n6873) );
  OAI211_X1 U7406 ( .C1(n6897), .C2(n6916), .A(n6874), .B(n6873), .ZN(U3121)
         );
  AOI22_X1 U7407 ( .A1(n6998), .A2(n6894), .B1(n6901), .B2(n6991), .ZN(n6876)
         );
  AOI22_X1 U7408 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6993), .B1(n6902), 
        .B2(n6992), .ZN(n6875) );
  OAI211_X1 U7409 ( .C1(n6897), .C2(n6996), .A(n6876), .B(n6875), .ZN(U3113)
         );
  AOI22_X1 U7410 ( .A1(n6879), .A2(n6894), .B1(n6901), .B2(n6997), .ZN(n6878)
         );
  AOI22_X1 U7411 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(n7000), .B1(n6902), 
        .B2(n6999), .ZN(n6877) );
  OAI211_X1 U7412 ( .C1(n6924), .C2(n6897), .A(n6878), .B(n6877), .ZN(U3105)
         );
  AOI22_X1 U7413 ( .A1(n6879), .A2(n6903), .B1(n6901), .B2(n7003), .ZN(n6881)
         );
  AOI22_X1 U7414 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n7006), .B1(n6902), 
        .B2(n7005), .ZN(n6880) );
  OAI211_X1 U7415 ( .C1(n6906), .C2(n7016), .A(n6881), .B(n6880), .ZN(U3097)
         );
  AOI22_X1 U7416 ( .A1(n6902), .A2(n7011), .B1(n6901), .B2(n7010), .ZN(n6883)
         );
  AOI22_X1 U7417 ( .A1(INSTQUEUE_REG_8__5__SCAN_IN), .A2(n7013), .B1(n6894), 
        .B2(n7012), .ZN(n6882) );
  OAI211_X1 U7418 ( .C1(n6897), .C2(n7016), .A(n6883), .B(n6882), .ZN(U3089)
         );
  AOI22_X1 U7419 ( .A1(n7018), .A2(n6894), .B1(n7017), .B2(n6901), .ZN(n6885)
         );
  AOI22_X1 U7420 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n7020), .B1(n6902), 
        .B2(n7019), .ZN(n6884) );
  OAI211_X1 U7421 ( .C1(n6897), .C2(n7023), .A(n6885), .B(n6884), .ZN(U3081)
         );
  AOI22_X1 U7422 ( .A1(n6902), .A2(n7025), .B1(n6901), .B2(n7024), .ZN(n6887)
         );
  AOI22_X1 U7423 ( .A1(INSTQUEUE_REG_6__5__SCAN_IN), .A2(n7026), .B1(n6894), 
        .B2(n7031), .ZN(n6886) );
  OAI211_X1 U7424 ( .C1(n6897), .C2(n7029), .A(n6887), .B(n6886), .ZN(U3073)
         );
  AOI22_X1 U7425 ( .A1(n7031), .A2(n6903), .B1(n6901), .B2(n7030), .ZN(n6889)
         );
  AOI22_X1 U7426 ( .A1(INSTQUEUE_REG_5__5__SCAN_IN), .A2(n7033), .B1(n6902), 
        .B2(n7032), .ZN(n6888) );
  OAI211_X1 U7427 ( .C1(n6906), .C2(n7036), .A(n6889), .B(n6888), .ZN(U3065)
         );
  AOI22_X1 U7428 ( .A1(n6902), .A2(n7038), .B1(n6901), .B2(n7037), .ZN(n6891)
         );
  AOI22_X1 U7429 ( .A1(n7040), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n7039), 
        .B2(n6903), .ZN(n6890) );
  OAI211_X1 U7430 ( .C1(n6906), .C2(n7048), .A(n6891), .B(n6890), .ZN(U3057)
         );
  AOI22_X1 U7431 ( .A1(n7051), .A2(n6894), .B1(n6901), .B2(n7043), .ZN(n6893)
         );
  AOI22_X1 U7432 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n7045), .B1(n6902), 
        .B2(n7044), .ZN(n6892) );
  OAI211_X1 U7433 ( .C1(n6897), .C2(n7048), .A(n6893), .B(n6892), .ZN(U3049)
         );
  AOI22_X1 U7434 ( .A1(n6902), .A2(n7050), .B1(n6901), .B2(n7049), .ZN(n6896)
         );
  AOI22_X1 U7435 ( .A1(INSTQUEUE_REG_2__5__SCAN_IN), .A2(n7052), .B1(n6898), 
        .B2(n6894), .ZN(n6895) );
  OAI211_X1 U7436 ( .C1(n6947), .C2(n6897), .A(n6896), .B(n6895), .ZN(U3041)
         );
  AOI22_X1 U7437 ( .A1(n6898), .A2(n6903), .B1(n6901), .B2(n7055), .ZN(n6900)
         );
  AOI22_X1 U7438 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n7058), .B1(n6902), 
        .B2(n7057), .ZN(n6899) );
  OAI211_X1 U7439 ( .C1(n6906), .C2(n6956), .A(n6900), .B(n6899), .ZN(U3033)
         );
  AOI22_X1 U7440 ( .A1(n6902), .A2(n7065), .B1(n6901), .B2(n7063), .ZN(n6905)
         );
  AOI22_X1 U7441 ( .A1(INSTQUEUE_REG_0__5__SCAN_IN), .A2(n7069), .B1(n6903), 
        .B2(n7067), .ZN(n6904) );
  OAI211_X1 U7442 ( .C1(n6906), .C2(n7072), .A(n6905), .B(n6904), .ZN(U3025)
         );
  AND2_X1 U7443 ( .A1(n6969), .A2(DATAI_22_), .ZN(n6959) );
  INV_X1 U7444 ( .A(n6959), .ZN(n6952) );
  NOR2_X2 U7445 ( .A1(n6907), .A2(n6963), .ZN(n6958) );
  NOR2_X1 U7446 ( .A1(n6966), .A2(n6908), .ZN(n6957) );
  AOI22_X1 U7447 ( .A1(n6958), .A2(n6968), .B1(n6957), .B2(n6967), .ZN(n6910)
         );
  AND2_X1 U7448 ( .A1(n6969), .A2(DATAI_30_), .ZN(n6936) );
  AOI22_X1 U7449 ( .A1(INSTQUEUE_REG_15__6__SCAN_IN), .A2(n6970), .B1(n6936), 
        .B2(n6975), .ZN(n6909) );
  OAI211_X1 U7450 ( .C1(n6952), .C2(n7072), .A(n6910), .B(n6909), .ZN(U3146)
         );
  INV_X1 U7451 ( .A(n6936), .ZN(n6962) );
  AOI22_X1 U7452 ( .A1(n6958), .A2(n6974), .B1(n6957), .B2(n6973), .ZN(n6912)
         );
  AOI22_X1 U7453 ( .A1(INSTQUEUE_REG_14__6__SCAN_IN), .A2(n6976), .B1(n6959), 
        .B2(n6975), .ZN(n6911) );
  OAI211_X1 U7454 ( .C1(n6962), .C2(n6984), .A(n6912), .B(n6911), .ZN(U3138)
         );
  AOI22_X1 U7455 ( .A1(n6913), .A2(n6959), .B1(n6957), .B2(n6979), .ZN(n6915)
         );
  AOI22_X1 U7456 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n6981), .B1(n6958), 
        .B2(n6980), .ZN(n6914) );
  OAI211_X1 U7457 ( .C1(n6962), .C2(n6916), .A(n6915), .B(n6914), .ZN(U3130)
         );
  AOI22_X1 U7458 ( .A1(n6958), .A2(n6986), .B1(n6957), .B2(n6985), .ZN(n6918)
         );
  AOI22_X1 U7459 ( .A1(INSTQUEUE_REG_12__6__SCAN_IN), .A2(n6988), .B1(n6959), 
        .B2(n6987), .ZN(n6917) );
  OAI211_X1 U7460 ( .C1(n6962), .C2(n6996), .A(n6918), .B(n6917), .ZN(U3122)
         );
  INV_X1 U7461 ( .A(n6957), .ZN(n6951) );
  OAI22_X1 U7462 ( .A1(n6924), .A2(n6962), .B1(n6951), .B2(n6919), .ZN(n6920)
         );
  INV_X1 U7463 ( .A(n6920), .ZN(n6922) );
  AOI22_X1 U7464 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6993), .B1(n6958), 
        .B2(n6992), .ZN(n6921) );
  OAI211_X1 U7465 ( .C1(n6952), .C2(n6996), .A(n6922), .B(n6921), .ZN(U3114)
         );
  OAI22_X1 U7466 ( .A1(n6924), .A2(n6952), .B1(n6951), .B2(n6923), .ZN(n6925)
         );
  INV_X1 U7467 ( .A(n6925), .ZN(n6927) );
  AOI22_X1 U7468 ( .A1(INSTQUEUE_REG_10__6__SCAN_IN), .A2(n7000), .B1(n6958), 
        .B2(n6999), .ZN(n6926) );
  OAI211_X1 U7469 ( .C1(n7009), .C2(n6962), .A(n6927), .B(n6926), .ZN(U3106)
         );
  OAI22_X1 U7470 ( .A1(n7016), .A2(n6962), .B1(n6951), .B2(n6928), .ZN(n6929)
         );
  INV_X1 U7471 ( .A(n6929), .ZN(n6931) );
  AOI22_X1 U7472 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n7006), .B1(n6958), 
        .B2(n7005), .ZN(n6930) );
  OAI211_X1 U7473 ( .C1(n7009), .C2(n6952), .A(n6931), .B(n6930), .ZN(U3098)
         );
  AOI22_X1 U7474 ( .A1(n6958), .A2(n7011), .B1(n6957), .B2(n7010), .ZN(n6933)
         );
  AOI22_X1 U7475 ( .A1(INSTQUEUE_REG_8__6__SCAN_IN), .A2(n7013), .B1(n6936), 
        .B2(n7012), .ZN(n6932) );
  OAI211_X1 U7476 ( .C1(n6952), .C2(n7016), .A(n6933), .B(n6932), .ZN(U3090)
         );
  AOI22_X1 U7477 ( .A1(n7012), .A2(n6959), .B1(n7017), .B2(n6957), .ZN(n6935)
         );
  AOI22_X1 U7478 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n7020), .B1(n6958), 
        .B2(n7019), .ZN(n6934) );
  OAI211_X1 U7479 ( .C1(n6962), .C2(n7029), .A(n6935), .B(n6934), .ZN(U3082)
         );
  AOI22_X1 U7480 ( .A1(n6958), .A2(n7025), .B1(n6957), .B2(n7024), .ZN(n6938)
         );
  AOI22_X1 U7481 ( .A1(INSTQUEUE_REG_6__6__SCAN_IN), .A2(n7026), .B1(n6936), 
        .B2(n7031), .ZN(n6937) );
  OAI211_X1 U7482 ( .C1(n6952), .C2(n7029), .A(n6938), .B(n6937), .ZN(U3074)
         );
  AOI22_X1 U7483 ( .A1(n7031), .A2(n6959), .B1(n6957), .B2(n7030), .ZN(n6940)
         );
  AOI22_X1 U7484 ( .A1(INSTQUEUE_REG_5__6__SCAN_IN), .A2(n7033), .B1(n6958), 
        .B2(n7032), .ZN(n6939) );
  OAI211_X1 U7485 ( .C1(n6962), .C2(n7036), .A(n6940), .B(n6939), .ZN(U3066)
         );
  AOI22_X1 U7486 ( .A1(n6958), .A2(n7038), .B1(n6957), .B2(n7037), .ZN(n6942)
         );
  AOI22_X1 U7487 ( .A1(n7040), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n7039), 
        .B2(n6959), .ZN(n6941) );
  OAI211_X1 U7488 ( .C1(n6962), .C2(n7048), .A(n6942), .B(n6941), .ZN(U3058)
         );
  OAI22_X1 U7489 ( .A1(n7048), .A2(n6952), .B1(n6951), .B2(n6943), .ZN(n6944)
         );
  INV_X1 U7490 ( .A(n6944), .ZN(n6946) );
  AOI22_X1 U7491 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n7045), .B1(n6958), 
        .B2(n7044), .ZN(n6945) );
  OAI211_X1 U7492 ( .C1(n6947), .C2(n6962), .A(n6946), .B(n6945), .ZN(U3050)
         );
  AOI22_X1 U7493 ( .A1(n6958), .A2(n7050), .B1(n6957), .B2(n7049), .ZN(n6949)
         );
  AOI22_X1 U7494 ( .A1(INSTQUEUE_REG_2__6__SCAN_IN), .A2(n7052), .B1(n7051), 
        .B2(n6959), .ZN(n6948) );
  OAI211_X1 U7495 ( .C1(n7062), .C2(n6962), .A(n6949), .B(n6948), .ZN(U3042)
         );
  OAI22_X1 U7496 ( .A1(n7062), .A2(n6952), .B1(n6951), .B2(n6950), .ZN(n6953)
         );
  INV_X1 U7497 ( .A(n6953), .ZN(n6955) );
  AOI22_X1 U7498 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n7058), .B1(n6958), 
        .B2(n7057), .ZN(n6954) );
  OAI211_X1 U7499 ( .C1(n6962), .C2(n6956), .A(n6955), .B(n6954), .ZN(U3034)
         );
  AOI22_X1 U7500 ( .A1(n6958), .A2(n7065), .B1(n6957), .B2(n7063), .ZN(n6961)
         );
  AOI22_X1 U7501 ( .A1(INSTQUEUE_REG_0__6__SCAN_IN), .A2(n7069), .B1(n6959), 
        .B2(n7067), .ZN(n6960) );
  OAI211_X1 U7502 ( .C1(n6962), .C2(n7072), .A(n6961), .B(n6960), .ZN(U3026)
         );
  AND2_X1 U7503 ( .A1(n6969), .A2(DATAI_23_), .ZN(n7068) );
  INV_X1 U7504 ( .A(n7068), .ZN(n7061) );
  NOR2_X2 U7505 ( .A1(n6964), .A2(n6963), .ZN(n7066) );
  NOR2_X2 U7506 ( .A1(n6966), .A2(n6965), .ZN(n7064) );
  AOI22_X1 U7507 ( .A1(n7066), .A2(n6968), .B1(n7064), .B2(n6967), .ZN(n6972)
         );
  AND2_X1 U7508 ( .A1(n6969), .A2(DATAI_31_), .ZN(n7056) );
  AOI22_X1 U7509 ( .A1(INSTQUEUE_REG_15__7__SCAN_IN), .A2(n6970), .B1(n7056), 
        .B2(n6975), .ZN(n6971) );
  OAI211_X1 U7510 ( .C1(n7061), .C2(n7072), .A(n6972), .B(n6971), .ZN(U3147)
         );
  INV_X1 U7511 ( .A(n7056), .ZN(n7073) );
  AOI22_X1 U7512 ( .A1(n7066), .A2(n6974), .B1(n7064), .B2(n6973), .ZN(n6978)
         );
  AOI22_X1 U7513 ( .A1(INSTQUEUE_REG_14__7__SCAN_IN), .A2(n6976), .B1(n7068), 
        .B2(n6975), .ZN(n6977) );
  OAI211_X1 U7514 ( .C1(n7073), .C2(n6984), .A(n6978), .B(n6977), .ZN(U3139)
         );
  AOI22_X1 U7515 ( .A1(n6987), .A2(n7056), .B1(n7064), .B2(n6979), .ZN(n6983)
         );
  AOI22_X1 U7516 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n6981), .B1(n7066), 
        .B2(n6980), .ZN(n6982) );
  OAI211_X1 U7517 ( .C1(n7061), .C2(n6984), .A(n6983), .B(n6982), .ZN(U3131)
         );
  AOI22_X1 U7518 ( .A1(n7066), .A2(n6986), .B1(n7064), .B2(n6985), .ZN(n6990)
         );
  AOI22_X1 U7519 ( .A1(INSTQUEUE_REG_12__7__SCAN_IN), .A2(n6988), .B1(n7068), 
        .B2(n6987), .ZN(n6989) );
  OAI211_X1 U7520 ( .C1(n7073), .C2(n6996), .A(n6990), .B(n6989), .ZN(U3123)
         );
  AOI22_X1 U7521 ( .A1(n6998), .A2(n7056), .B1(n7064), .B2(n6991), .ZN(n6995)
         );
  AOI22_X1 U7522 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6993), .B1(n7066), 
        .B2(n6992), .ZN(n6994) );
  OAI211_X1 U7523 ( .C1(n7061), .C2(n6996), .A(n6995), .B(n6994), .ZN(U3115)
         );
  AOI22_X1 U7524 ( .A1(n6998), .A2(n7068), .B1(n7064), .B2(n6997), .ZN(n7002)
         );
  AOI22_X1 U7525 ( .A1(INSTQUEUE_REG_10__7__SCAN_IN), .A2(n7000), .B1(n7066), 
        .B2(n6999), .ZN(n7001) );
  OAI211_X1 U7526 ( .C1(n7009), .C2(n7073), .A(n7002), .B(n7001), .ZN(U3107)
         );
  AOI22_X1 U7527 ( .A1(n7004), .A2(n7056), .B1(n7064), .B2(n7003), .ZN(n7008)
         );
  AOI22_X1 U7528 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n7006), .B1(n7066), 
        .B2(n7005), .ZN(n7007) );
  OAI211_X1 U7529 ( .C1(n7009), .C2(n7061), .A(n7008), .B(n7007), .ZN(U3099)
         );
  AOI22_X1 U7530 ( .A1(n7066), .A2(n7011), .B1(n7064), .B2(n7010), .ZN(n7015)
         );
  AOI22_X1 U7531 ( .A1(INSTQUEUE_REG_8__7__SCAN_IN), .A2(n7013), .B1(n7056), 
        .B2(n7012), .ZN(n7014) );
  OAI211_X1 U7532 ( .C1(n7061), .C2(n7016), .A(n7015), .B(n7014), .ZN(U3091)
         );
  AOI22_X1 U7533 ( .A1(n7018), .A2(n7056), .B1(n7017), .B2(n7064), .ZN(n7022)
         );
  AOI22_X1 U7534 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n7020), .B1(n7066), 
        .B2(n7019), .ZN(n7021) );
  OAI211_X1 U7535 ( .C1(n7061), .C2(n7023), .A(n7022), .B(n7021), .ZN(U3083)
         );
  AOI22_X1 U7536 ( .A1(n7066), .A2(n7025), .B1(n7064), .B2(n7024), .ZN(n7028)
         );
  AOI22_X1 U7537 ( .A1(INSTQUEUE_REG_6__7__SCAN_IN), .A2(n7026), .B1(n7056), 
        .B2(n7031), .ZN(n7027) );
  OAI211_X1 U7538 ( .C1(n7061), .C2(n7029), .A(n7028), .B(n7027), .ZN(U3075)
         );
  AOI22_X1 U7539 ( .A1(n7031), .A2(n7068), .B1(n7064), .B2(n7030), .ZN(n7035)
         );
  AOI22_X1 U7540 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n7033), .B1(n7066), 
        .B2(n7032), .ZN(n7034) );
  OAI211_X1 U7541 ( .C1(n7073), .C2(n7036), .A(n7035), .B(n7034), .ZN(U3067)
         );
  AOI22_X1 U7542 ( .A1(n7066), .A2(n7038), .B1(n7064), .B2(n7037), .ZN(n7042)
         );
  AOI22_X1 U7543 ( .A1(n7040), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n7039), 
        .B2(n7068), .ZN(n7041) );
  OAI211_X1 U7544 ( .C1(n7073), .C2(n7048), .A(n7042), .B(n7041), .ZN(U3059)
         );
  AOI22_X1 U7545 ( .A1(n7051), .A2(n7056), .B1(n7064), .B2(n7043), .ZN(n7047)
         );
  AOI22_X1 U7546 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n7045), .B1(n7066), 
        .B2(n7044), .ZN(n7046) );
  OAI211_X1 U7547 ( .C1(n7061), .C2(n7048), .A(n7047), .B(n7046), .ZN(U3051)
         );
  AOI22_X1 U7548 ( .A1(n7066), .A2(n7050), .B1(n7064), .B2(n7049), .ZN(n7054)
         );
  AOI22_X1 U7549 ( .A1(INSTQUEUE_REG_2__7__SCAN_IN), .A2(n7052), .B1(n7051), 
        .B2(n7068), .ZN(n7053) );
  OAI211_X1 U7550 ( .C1(n7062), .C2(n7073), .A(n7054), .B(n7053), .ZN(U3043)
         );
  AOI22_X1 U7551 ( .A1(n7067), .A2(n7056), .B1(n7064), .B2(n7055), .ZN(n7060)
         );
  AOI22_X1 U7552 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n7058), .B1(n7066), 
        .B2(n7057), .ZN(n7059) );
  OAI211_X1 U7553 ( .C1(n7062), .C2(n7061), .A(n7060), .B(n7059), .ZN(U3035)
         );
  AOI22_X1 U7554 ( .A1(n7066), .A2(n7065), .B1(n7064), .B2(n7063), .ZN(n7071)
         );
  AOI22_X1 U7555 ( .A1(INSTQUEUE_REG_0__7__SCAN_IN), .A2(n7069), .B1(n7068), 
        .B2(n7067), .ZN(n7070) );
  OAI211_X1 U7556 ( .C1(n7073), .C2(n7072), .A(n7071), .B(n7070), .ZN(U3027)
         );
  BUF_X1 U3530 ( .A(n3699), .Z(n3622) );
  CLKBUF_X1 U34710 ( .A(n3544), .Z(n4406) );
  CLKBUF_X1 U34720 ( .A(n3586), .Z(n4656) );
  CLKBUF_X1 U34730 ( .A(n4444), .Z(n4837) );
  CLKBUF_X1 U3478 ( .A(n3564), .Z(n3608) );
  CLKBUF_X1 U3501 ( .A(n5611), .Z(n5746) );
  CLKBUF_X1 U3646 ( .A(n5184), .Z(n3432) );
  CLKBUF_X1 U3739 ( .A(n5777), .Z(n6004) );
  INV_X2 U5211 ( .A(n6427), .ZN(n6152) );
endmodule

