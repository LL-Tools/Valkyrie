

module b20_C_gen_AntiSAT_k_256_9 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, 
        keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, 
        keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, 
        keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, 
        keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, 
        keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, 
        keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, 
        keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, 
        keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104, 
        keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108, 
        keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112, 
        keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116, 
        keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120, 
        keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124, 
        keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, 
        keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, 
        keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, 
        keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, 
        keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, 
        keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, 
        keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, 
        keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, 
        ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, 
        ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, 
        ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, 
        ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, 
        P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, 
        P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, 
        P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, 
        P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, 
        P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, 
        P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, 
        P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, 
        P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, 
        P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, 
        P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, 
        P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, 
        P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, 
        P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, 
        P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, 
        P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, 
        P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, 
        P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, 
        P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, 
        P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, 
        P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, 
        P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, 
        P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, 
        P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, 
        P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, 
        P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, 
        P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, 
        P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, 
        P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, 
        P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, 
        P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, 
        P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703;

  INV_X1 U5011 ( .A(n10067), .ZN(n9139) );
  NAND4_X1 U5012 ( .A1(n6043), .A2(n6042), .A3(n6041), .A4(n6040), .ZN(n6381)
         );
  INV_X1 U5013 ( .A(n10005), .ZN(n10050) );
  CLKBUF_X3 U5014 ( .A(n5355), .Z(n8158) );
  INV_X4 U5015 ( .A(n7471), .ZN(n6070) );
  INV_X2 U5016 ( .A(n6783), .ZN(n5727) );
  XNOR2_X1 U5017 ( .A(n5273), .B(n5272), .ZN(n9909) );
  INV_X1 U5018 ( .A(n8141), .ZN(n7014) );
  INV_X1 U5019 ( .A(n8133), .ZN(n8124) );
  INV_X1 U5020 ( .A(n7936), .ZN(n6270) );
  NAND2_X2 U5021 ( .A1(n5294), .A2(n5322), .ZN(n5346) );
  INV_X1 U5022 ( .A(n5322), .ZN(n5898) );
  AND2_X1 U5023 ( .A1(n6783), .A2(n4506), .ZN(n5355) );
  INV_X1 U5024 ( .A(n8419), .ZN(n4796) );
  NAND2_X1 U5025 ( .A1(n6783), .A2(n6714), .ZN(n6562) );
  INV_X1 U5026 ( .A(n9222), .ZN(n9347) );
  NAND2_X1 U5028 ( .A1(n5155), .A2(n5154), .ZN(n5422) );
  OAI211_X1 U5029 ( .C1(n6562), .C2(n6730), .A(n5313), .B(n5129), .ZN(n10021)
         );
  NAND2_X1 U5030 ( .A1(n5076), .A2(n5075), .ZN(n9023) );
  NAND2_X1 U5031 ( .A1(n5407), .A2(n5406), .ZN(n10067) );
  XNOR2_X1 U5032 ( .A(n5256), .B(P1_IR_REG_21__SCAN_IN), .ZN(n5964) );
  OR4_X1 U5033 ( .A1(n8992), .A2(n5966), .A3(n9919), .A4(n5965), .ZN(n5988) );
  INV_X2 U5034 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X2 U5035 ( .A(n5389), .ZN(n5754) );
  NAND4_X4 U5036 ( .A1(n6051), .A2(n6050), .A3(n6049), .A4(n6048), .ZN(n8420)
         );
  NAND2_X2 U5038 ( .A1(n6572), .A2(n9299), .ZN(n10001) );
  NAND2_X2 U5039 ( .A1(n9900), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5270) );
  BUF_X4 U5040 ( .A(n6071), .Z(n7469) );
  AOI21_X2 U5041 ( .B1(n7127), .B2(n6674), .A(n7106), .ZN(n7258) );
  OAI22_X2 U5042 ( .A1(n7521), .A2(n6531), .B1(n7611), .B2(n9240), .ZN(n7650)
         );
  NAND2_X2 U5043 ( .A1(n6529), .A2(n6528), .ZN(n7521) );
  AND2_X1 U5045 ( .A1(n4989), .A2(n4985), .ZN(n4506) );
  AND2_X1 U5046 ( .A1(n4989), .A2(n4985), .ZN(n4507) );
  INV_X4 U5047 ( .A(n7931), .ZN(n6714) );
  AND2_X1 U5048 ( .A1(n4514), .A2(n4515), .ZN(n6566) );
  CLKBUF_X1 U5049 ( .A(n8248), .Z(n8249) );
  OAI21_X1 U5050 ( .B1(n9058), .B2(n5063), .A(n5060), .ZN(n8989) );
  OAI21_X1 U5051 ( .B1(n9058), .B2(n5059), .A(n5057), .ZN(n8992) );
  AOI21_X1 U5052 ( .B1(n4685), .B2(n10161), .A(n4682), .ZN(n8575) );
  AND2_X1 U5053 ( .A1(n8328), .A2(n8219), .ZN(n5097) );
  OR4_X1 U5054 ( .A1(n8121), .A2(n7971), .A3(n8629), .A4(n7970), .ZN(n7974) );
  AOI21_X1 U5055 ( .B1(n8554), .B2(n8567), .A(n8553), .ZN(n8556) );
  INV_X1 U5056 ( .A(n4975), .ZN(n4974) );
  AOI21_X1 U5057 ( .B1(n4975), .B2(n4973), .A(n4570), .ZN(n4972) );
  NAND2_X1 U5058 ( .A1(n5601), .A2(n9915), .ZN(n9921) );
  INV_X1 U5059 ( .A(n4786), .ZN(n4780) );
  AND2_X1 U5060 ( .A1(n6316), .A2(n8085), .ZN(n4786) );
  NAND2_X1 U5061 ( .A1(n6328), .A2(n6327), .ZN(n8909) );
  NAND2_X1 U5062 ( .A1(n6306), .A2(n6305), .ZN(n8921) );
  AND2_X1 U5063 ( .A1(n5089), .A2(n7870), .ZN(n5087) );
  AND2_X1 U5064 ( .A1(n5116), .A2(n6545), .ZN(n4983) );
  AND2_X1 U5065 ( .A1(n7192), .A2(n5457), .ZN(n7193) );
  AND2_X1 U5066 ( .A1(n7191), .A2(n7248), .ZN(n5458) );
  NAND2_X1 U5067 ( .A1(n4622), .A2(n5440), .ZN(n7192) );
  NAND2_X1 U5068 ( .A1(n5710), .A2(n5709), .ZN(n9743) );
  NAND2_X1 U5069 ( .A1(n6149), .A2(n6148), .ZN(n7718) );
  INV_X1 U5070 ( .A(n9382), .ZN(n9132) );
  INV_X2 U5071 ( .A(n7169), .ZN(n8235) );
  NAND4_X2 U5072 ( .A1(n6062), .A2(n6061), .A3(n6060), .A4(n6059), .ZN(n8418)
         );
  NAND4_X2 U5073 ( .A1(n5365), .A2(n5364), .A3(n5363), .A4(n5362), .ZN(n9384)
         );
  INV_X2 U5074 ( .A(n6744), .ZN(n6834) );
  OAI211_X1 U5075 ( .C1(n6562), .C2(n6717), .A(n5359), .B(n5358), .ZN(n7290)
         );
  NOR2_X2 U5076 ( .A1(n6686), .A2(P2_U3151), .ZN(P2_U3893) );
  OAI211_X1 U5077 ( .C1(n6562), .C2(n6732), .A(n5344), .B(n5343), .ZN(n10005)
         );
  INV_X2 U5078 ( .A(n5360), .ZN(n5928) );
  XNOR2_X1 U5079 ( .A(n6437), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7015) );
  NAND2_X2 U5080 ( .A1(n6025), .A2(n6024), .ZN(n6375) );
  CLKBUF_X1 U5081 ( .A(n6066), .Z(n7936) );
  XNOR2_X1 U5082 ( .A(n5255), .B(n5254), .ZN(n5284) );
  NAND2_X1 U5083 ( .A1(n6436), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6437) );
  INV_X1 U5084 ( .A(n9909), .ZN(n5276) );
  INV_X1 U5085 ( .A(n5963), .ZN(n9351) );
  NAND2_X1 U5086 ( .A1(n6462), .A2(n6463), .ZN(n7767) );
  XNOR2_X1 U5087 ( .A(n6017), .B(n6016), .ZN(n6022) );
  XNOR2_X1 U5088 ( .A(n6465), .B(n6464), .ZN(n8150) );
  XNOR2_X1 U5089 ( .A(n6468), .B(P2_IR_REG_26__SCAN_IN), .ZN(n6727) );
  NAND2_X1 U5090 ( .A1(n5993), .A2(n5992), .ZN(n6208) );
  NAND2_X1 U5091 ( .A1(n4890), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6033) );
  NAND2_X1 U5092 ( .A1(n5257), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5943) );
  NOR2_X1 U5093 ( .A1(n5240), .A2(n5023), .ZN(n5271) );
  NAND2_X1 U5094 ( .A1(n4933), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5230) );
  NAND2_X1 U5095 ( .A1(n5248), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5646) );
  OR2_X1 U5096 ( .A1(n5246), .A2(n9899), .ZN(n5256) );
  XNOR2_X1 U5097 ( .A(n6082), .B(n6081), .ZN(n6974) );
  AND2_X1 U5098 ( .A1(n4541), .A2(n4835), .ZN(n5226) );
  AND3_X1 U5099 ( .A1(n4573), .A2(n5424), .A3(n4648), .ZN(n5246) );
  AND2_X2 U5100 ( .A1(n4989), .A2(n4985), .ZN(n7931) );
  AND2_X1 U5101 ( .A1(n5224), .A2(n5945), .ZN(n4839) );
  AND4_X1 U5102 ( .A1(n5219), .A2(n5218), .A3(n5217), .A4(n5216), .ZN(n5220)
         );
  NAND2_X1 U5103 ( .A1(n5339), .A2(n5213), .ZN(n5375) );
  INV_X4 U5104 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U5105 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5213) );
  INV_X1 U5106 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6004) );
  INV_X1 U5107 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6232) );
  INV_X1 U5108 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6218) );
  INV_X1 U5109 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6005) );
  NOR2_X1 U5110 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n4732) );
  NOR2_X1 U5111 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n4731) );
  NOR2_X1 U5112 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n4730) );
  INV_X1 U5113 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4670) );
  INV_X1 U5114 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6111) );
  INV_X1 U5115 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5214) );
  NOR2_X1 U5116 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5234) );
  INV_X1 U5117 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5685) );
  INV_X1 U5118 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U5119 ( .A1(n6522), .A2(n4511), .ZN(n4508) );
  AND2_X1 U5120 ( .A1(n4508), .A2(n4509), .ZN(n9967) );
  OR2_X1 U5121 ( .A1(n4510), .A2(n9145), .ZN(n4509) );
  INV_X1 U5122 ( .A(n6523), .ZN(n4510) );
  AND2_X1 U5123 ( .A1(n6521), .A2(n6523), .ZN(n4511) );
  INV_X1 U5124 ( .A(n7009), .ZN(n4512) );
  NAND3_X1 U5125 ( .A1(n5335), .A2(n5334), .A3(n5333), .ZN(n6512) );
  INV_X1 U5126 ( .A(n6984), .ZN(n4513) );
  CLKBUF_X2 U5127 ( .A(n6509), .Z(n6984) );
  NAND2_X1 U5128 ( .A1(n5274), .A2(n9909), .ZN(n5361) );
  NAND2_X1 U5129 ( .A1(n5274), .A2(n5276), .ZN(n5969) );
  OR2_X1 U5130 ( .A1(n5361), .A2(n5314), .ZN(n5316) );
  OR2_X1 U5131 ( .A1(n7289), .A2(n7290), .ZN(n9984) );
  INV_X1 U5132 ( .A(n5275), .ZN(n5274) );
  NAND2_X1 U5133 ( .A1(n9590), .A2(n4517), .ZN(n4514) );
  OR2_X1 U5134 ( .A1(n4516), .A2(n6560), .ZN(n4515) );
  INV_X1 U5135 ( .A(n6561), .ZN(n4516) );
  AND2_X1 U5136 ( .A1(n6559), .A2(n6561), .ZN(n4517) );
  CLKBUF_X1 U5137 ( .A(n7178), .Z(n4518) );
  NAND2_X1 U5138 ( .A1(n5624), .A2(n5226), .ZN(n5240) );
  CLKBUF_X1 U5139 ( .A(n9930), .Z(n4519) );
  XNOR2_X1 U5140 ( .A(n5230), .B(n5227), .ZN(n9930) );
  INV_X1 U5141 ( .A(n9983), .ZN(n10063) );
  NAND2_X1 U5142 ( .A1(n5241), .A2(n5240), .ZN(n7770) );
  OR2_X1 U5143 ( .A1(n5271), .A2(n9899), .ZN(n5273) );
  OR2_X1 U5144 ( .A1(n4521), .A2(n9405), .ZN(n5334) );
  BUF_X4 U5145 ( .A(n5969), .Z(n4520) );
  BUF_X2 U5146 ( .A(n5969), .Z(n4521) );
  INV_X1 U5147 ( .A(n4505), .ZN(n6025) );
  AND3_X1 U5148 ( .A1(n4936), .A2(n4934), .A3(n4602), .ZN(n8566) );
  AND2_X1 U5149 ( .A1(n5829), .A2(n5808), .ZN(n5827) );
  OAI21_X1 U5150 ( .B1(n5707), .B2(n5706), .A(n5195), .ZN(n5725) );
  OAI21_X1 U5151 ( .B1(n9291), .B2(n5054), .A(n9348), .ZN(n5053) );
  XNOR2_X1 U5152 ( .A(n5247), .B(n5237), .ZN(n9292) );
  INV_X1 U5153 ( .A(n4964), .ZN(n4963) );
  NAND2_X1 U5154 ( .A1(n5298), .A2(n6046), .ZN(n4954) );
  XNOR2_X1 U5155 ( .A(n5135), .B(n5132), .ZN(n5309) );
  AOI21_X1 U5156 ( .B1(n4525), .B2(n4550), .A(n4771), .ZN(n4770) );
  OAI21_X1 U5157 ( .B1(n4772), .B2(n8038), .A(n4774), .ZN(n4771) );
  INV_X1 U5158 ( .A(n8046), .ZN(n4769) );
  MUX2_X1 U5159 ( .A(n9170), .B(n9169), .S(n9222), .Z(n9176) );
  AOI21_X1 U5160 ( .B1(n4569), .B2(n9181), .A(n9222), .ZN(n4827) );
  BUF_X1 U5161 ( .A(n7169), .Z(n8228) );
  NOR2_X1 U5162 ( .A1(n8121), .A2(n8120), .ZN(n4759) );
  OR2_X1 U5163 ( .A1(n8615), .A2(n6380), .ZN(n8123) );
  OR2_X1 U5164 ( .A1(n7339), .A2(n6646), .ZN(n6648) );
  OR2_X1 U5165 ( .A1(n8955), .A2(n8753), .ZN(n8080) );
  NOR2_X1 U5166 ( .A1(n4794), .A2(n8027), .ZN(n4793) );
  OR2_X1 U5167 ( .A1(n8927), .A2(n8294), .ZN(n7979) );
  NOR2_X1 U5168 ( .A1(n8921), .A2(n8219), .ZN(n8102) );
  NAND2_X1 U5169 ( .A1(n8933), .A2(n8733), .ZN(n8093) );
  OR2_X1 U5170 ( .A1(n8944), .A2(n8754), .ZN(n8085) );
  AOI21_X1 U5171 ( .B1(n4856), .B2(n4858), .A(n4557), .ZN(n4854) );
  OR2_X1 U5172 ( .A1(n7873), .A2(n8409), .ZN(n4864) );
  CLKBUF_X1 U5173 ( .A(n7015), .Z(n4610) );
  NAND2_X1 U5174 ( .A1(n6011), .A2(n4843), .ZN(n4842) );
  NOR2_X1 U5175 ( .A1(n9577), .A2(n9560), .ZN(n8162) );
  OR2_X1 U5176 ( .A1(n9760), .A2(n6592), .ZN(n9282) );
  AND2_X1 U5177 ( .A1(n9259), .A2(n9215), .ZN(n9252) );
  NOR2_X1 U5178 ( .A1(n9607), .A2(n9849), .ZN(n4928) );
  OR2_X1 U5179 ( .A1(n9782), .A2(n6589), .ZN(n9262) );
  NOR2_X1 U5180 ( .A1(n9698), .A2(n4925), .ZN(n4924) );
  INV_X1 U5181 ( .A(n9879), .ZN(n4925) );
  INV_X1 U5182 ( .A(n9171), .ZN(n9316) );
  AND2_X1 U5183 ( .A1(n5220), .A2(n4649), .ZN(n4648) );
  NOR2_X1 U5184 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n4649) );
  NAND2_X1 U5185 ( .A1(n5189), .A2(n5188), .ZN(n5707) );
  OR2_X1 U5186 ( .A1(n5683), .A2(n5186), .ZN(n5189) );
  NAND2_X1 U5187 ( .A1(n4695), .A2(n4694), .ZN(n5623) );
  AOI21_X1 U5188 ( .B1(n4697), .B2(n4699), .A(n4562), .ZN(n4694) );
  NOR2_X1 U5189 ( .A1(n5177), .A2(n4702), .ZN(n4701) );
  INV_X1 U5190 ( .A(n5174), .ZN(n4702) );
  INV_X1 U5191 ( .A(n5577), .ZN(n5177) );
  NAND2_X1 U5192 ( .A1(n8171), .A2(n8170), .ZN(n8258) );
  INV_X1 U5193 ( .A(n8261), .ZN(n8170) );
  AND2_X1 U5194 ( .A1(n8823), .A2(n7976), .ZN(n8135) );
  INV_X1 U5195 ( .A(n6375), .ZN(n6360) );
  AND4_X1 U5196 ( .A1(n6183), .A2(n6182), .A3(n6181), .A4(n6180), .ZN(n7879)
         );
  AND2_X1 U5197 ( .A1(n4505), .A2(n8245), .ZN(n6071) );
  AND3_X1 U5198 ( .A1(n4679), .A2(n4596), .A3(n4678), .ZN(n6703) );
  NAND2_X1 U5199 ( .A1(n4677), .A2(n4676), .ZN(n4675) );
  INV_X1 U5200 ( .A(n7698), .ZN(n4676) );
  NAND2_X1 U5201 ( .A1(n4687), .A2(n4948), .ZN(n8583) );
  NAND2_X1 U5202 ( .A1(n8568), .A2(n4949), .ZN(n4948) );
  NAND2_X1 U5203 ( .A1(n4688), .A2(n4531), .ZN(n4687) );
  NAND2_X1 U5204 ( .A1(n7783), .A2(n6184), .ZN(n4798) );
  NOR2_X1 U5205 ( .A1(n10208), .A2(n4610), .ZN(n6924) );
  NOR2_X1 U5206 ( .A1(n8631), .A2(n4889), .ZN(n8621) );
  AND2_X1 U5207 ( .A1(n8897), .A2(n8645), .ZN(n4889) );
  AOI21_X1 U5208 ( .B1(n8644), .B2(n6433), .A(n6432), .ZN(n8630) );
  XNOR2_X1 U5209 ( .A(n8897), .B(n8386), .ZN(n8629) );
  NAND2_X1 U5210 ( .A1(n8921), .A2(n8219), .ZN(n8674) );
  NOR2_X1 U5211 ( .A1(n8688), .A2(n8102), .ZN(n4785) );
  INV_X1 U5212 ( .A(n8597), .ZN(n6438) );
  AOI21_X1 U5213 ( .B1(n6410), .B2(n6409), .A(n4522), .ZN(n8783) );
  INV_X1 U5214 ( .A(n7963), .ZN(n6409) );
  AOI21_X1 U5215 ( .B1(n4859), .B2(n6406), .A(n4857), .ZN(n4856) );
  INV_X1 U5216 ( .A(n8051), .ZN(n4857) );
  NAND2_X1 U5217 ( .A1(n4863), .A2(n4862), .ZN(n4861) );
  INV_X1 U5218 ( .A(n7836), .ZN(n4863) );
  INV_X1 U5219 ( .A(n6627), .ZN(n6269) );
  AND2_X1 U5220 ( .A1(n5292), .A2(n5976), .ZN(n5293) );
  NAND2_X1 U5221 ( .A1(n5759), .A2(n5760), .ZN(n5079) );
  NAND2_X1 U5222 ( .A1(n9023), .A2(n4667), .ZN(n4659) );
  AND2_X1 U5223 ( .A1(n5875), .A2(n5061), .ZN(n5060) );
  NAND2_X1 U5224 ( .A1(n9031), .A2(n5062), .ZN(n5061) );
  AND2_X1 U5225 ( .A1(n9098), .A2(n9099), .ZN(n5875) );
  INV_X1 U5226 ( .A(n5826), .ZN(n5062) );
  MUX2_X1 U5227 ( .A(n9222), .B(n9221), .S(n9554), .Z(n9228) );
  INV_X1 U5228 ( .A(n5361), .ZN(n5691) );
  NAND2_X1 U5229 ( .A1(n4928), .A2(n4927), .ZN(n9577) );
  INV_X1 U5230 ( .A(n9760), .ZN(n4927) );
  INV_X1 U5231 ( .A(n5860), .ZN(n5858) );
  NOR2_X1 U5232 ( .A1(n6556), .A2(n4979), .ZN(n4978) );
  INV_X1 U5233 ( .A(n6554), .ZN(n4979) );
  INV_X1 U5234 ( .A(n4971), .ZN(n4968) );
  NAND2_X1 U5235 ( .A1(n6595), .A2(n6594), .ZN(n9996) );
  XNOR2_X1 U5236 ( .A(n7935), .B(n7934), .ZN(n8980) );
  NAND2_X1 U5237 ( .A1(n6371), .A2(SI_29_), .ZN(n7925) );
  NAND2_X1 U5238 ( .A1(n5028), .A2(n5805), .ZN(n5828) );
  NAND2_X1 U5239 ( .A1(n5804), .A2(n5803), .ZN(n5028) );
  NAND2_X1 U5240 ( .A1(n4719), .A2(n4721), .ZN(n5743) );
  NAND2_X1 U5241 ( .A1(n5725), .A2(n4723), .ZN(n4719) );
  INV_X1 U5242 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5130) );
  OR2_X1 U5243 ( .A1(n7618), .A2(n7668), .ZN(n4947) );
  XNOR2_X1 U5244 ( .A(n6703), .B(n7630), .ZN(n7618) );
  AOI21_X1 U5245 ( .B1(n9291), .B2(n5051), .A(n9292), .ZN(n5050) );
  OR2_X1 U5246 ( .A1(n9545), .A2(n9225), .ZN(n9355) );
  OR2_X1 U5247 ( .A1(n9383), .A2(n9347), .ZN(n9140) );
  NAND2_X1 U5248 ( .A1(n4802), .A2(n9222), .ZN(n4801) );
  INV_X1 U5249 ( .A(n4775), .ZN(n4772) );
  AND2_X1 U5250 ( .A1(n9305), .A2(n9164), .ZN(n4820) );
  AOI21_X1 U5251 ( .B1(n9154), .B2(n4528), .A(n4819), .ZN(n4818) );
  AOI21_X1 U5252 ( .B1(n4770), .B2(n4773), .A(n4769), .ZN(n4768) );
  NOR2_X1 U5253 ( .A1(n4525), .A2(n4775), .ZN(n4773) );
  OR2_X1 U5254 ( .A1(n4770), .A2(n4769), .ZN(n4766) );
  OR2_X1 U5255 ( .A1(n9943), .A2(n9315), .ZN(n4608) );
  NOR2_X1 U5256 ( .A1(n4834), .A2(n4830), .ZN(n4829) );
  NAND2_X1 U5257 ( .A1(n9181), .A2(n9222), .ZN(n4834) );
  NOR2_X1 U5258 ( .A1(n9179), .A2(n4831), .ZN(n4830) );
  AOI21_X1 U5259 ( .B1(n4827), .B2(n4828), .A(n9182), .ZN(n4826) );
  NAND2_X1 U5260 ( .A1(n4568), .A2(n9181), .ZN(n4828) );
  NAND2_X1 U5261 ( .A1(n4829), .A2(n4832), .ZN(n4823) );
  NAND2_X1 U5262 ( .A1(n4833), .A2(n9296), .ZN(n4832) );
  INV_X1 U5263 ( .A(n9318), .ZN(n4833) );
  NAND2_X1 U5264 ( .A1(n4534), .A2(n4606), .ZN(n4814) );
  INV_X1 U5265 ( .A(n9271), .ZN(n4606) );
  NOR2_X1 U5266 ( .A1(n4744), .A2(n4743), .ZN(n4742) );
  NOR2_X1 U5267 ( .A1(n4746), .A2(n4747), .ZN(n4743) );
  INV_X1 U5268 ( .A(n8096), .ZN(n4747) );
  NAND2_X1 U5269 ( .A1(n4737), .A2(n4741), .ZN(n4740) );
  AND2_X1 U5270 ( .A1(n4745), .A2(n4748), .ZN(n4741) );
  INV_X1 U5271 ( .A(n8089), .ZN(n4748) );
  NAND2_X1 U5272 ( .A1(n9281), .A2(n9222), .ZN(n4803) );
  NOR2_X1 U5273 ( .A1(n9281), .A2(n9213), .ZN(n4805) );
  NAND2_X1 U5274 ( .A1(n9161), .A2(n9148), .ZN(n9152) );
  INV_X1 U5275 ( .A(n5047), .ZN(n5046) );
  OR2_X1 U5276 ( .A1(n8200), .A2(n8356), .ZN(n8201) );
  NAND2_X1 U5277 ( .A1(n4758), .A2(n4757), .ZN(n4756) );
  NOR2_X1 U5278 ( .A1(n5038), .A2(n4589), .ZN(n5037) );
  INV_X1 U5279 ( .A(n5681), .ZN(n5187) );
  AOI21_X1 U5280 ( .B1(n4700), .B2(n4698), .A(n5602), .ZN(n4697) );
  INV_X1 U5281 ( .A(n4701), .ZN(n4698) );
  INV_X1 U5282 ( .A(n4700), .ZN(n4699) );
  AND2_X1 U5283 ( .A1(n5528), .A2(n5532), .ZN(n5166) );
  INV_X1 U5284 ( .A(n5990), .ZN(n4847) );
  NOR2_X1 U5285 ( .A1(n6006), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n4846) );
  NOR2_X1 U5286 ( .A1(n7414), .A2(n5108), .ZN(n5107) );
  INV_X1 U5287 ( .A(n7412), .ZN(n5108) );
  INV_X1 U5288 ( .A(n4756), .ZN(n4752) );
  NOR2_X1 U5289 ( .A1(n8131), .A2(n4610), .ZN(n7972) );
  AOI211_X1 U5290 ( .C1(n7943), .C2(n8123), .A(n8128), .B(n7942), .ZN(n7944)
         );
  NAND2_X1 U5291 ( .A1(n4693), .A2(n4610), .ZN(n4692) );
  NAND2_X1 U5292 ( .A1(n8126), .A2(n8823), .ZN(n4693) );
  OAI21_X1 U5293 ( .B1(n4760), .B2(n4752), .A(n4750), .ZN(n4755) );
  AOI21_X1 U5294 ( .B1(n4751), .B2(n4756), .A(n8633), .ZN(n4750) );
  INV_X1 U5295 ( .A(n4759), .ZN(n4751) );
  INV_X1 U5296 ( .A(n8128), .ZN(n4754) );
  NAND2_X1 U5297 ( .A1(n4760), .A2(n4544), .ZN(n4753) );
  NAND2_X1 U5298 ( .A1(n6964), .A2(n6696), .ZN(n6697) );
  NAND2_X1 U5299 ( .A1(n4953), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4952) );
  NAND2_X1 U5300 ( .A1(n4545), .A2(n6402), .ZN(n4874) );
  INV_X1 U5301 ( .A(n4874), .ZN(n4870) );
  AOI21_X1 U5302 ( .B1(n4879), .B2(n4878), .A(n6398), .ZN(n4877) );
  INV_X1 U5303 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U5304 ( .A1(n4868), .A2(n6386), .ZN(n4866) );
  INV_X1 U5305 ( .A(n6385), .ZN(n4868) );
  OR2_X1 U5306 ( .A1(n8418), .A2(n10186), .ZN(n8003) );
  INV_X1 U5307 ( .A(n7988), .ZN(n6382) );
  NAND2_X1 U5308 ( .A1(n6055), .A2(n7020), .ZN(n7987) );
  NAND2_X1 U5309 ( .A1(n8108), .A2(n8104), .ZN(n4711) );
  NOR2_X1 U5310 ( .A1(n4711), .A2(n4780), .ZN(n4710) );
  NOR2_X1 U5311 ( .A1(n4712), .A2(n8109), .ZN(n4709) );
  INV_X1 U5312 ( .A(n8731), .ZN(n4852) );
  OR2_X1 U5313 ( .A1(n8365), .A2(n8771), .ZN(n8081) );
  OR2_X1 U5314 ( .A1(n7873), .A2(n7907), .ZN(n8045) );
  NOR2_X1 U5315 ( .A1(n5996), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n4765) );
  INV_X1 U5316 ( .A(n7572), .ZN(n5073) );
  NAND2_X1 U5317 ( .A1(n5777), .A2(n4668), .ZN(n4667) );
  INV_X1 U5318 ( .A(n5778), .ZN(n4668) );
  AND2_X1 U5319 ( .A1(n5084), .A2(n5723), .ZN(n5083) );
  NAND2_X1 U5320 ( .A1(n9050), .A2(n5085), .ZN(n5084) );
  AND2_X1 U5321 ( .A1(n9879), .A2(n9369), .ZN(n9327) );
  NOR2_X1 U5322 ( .A1(n6557), .A2(n4976), .ZN(n4975) );
  INV_X1 U5323 ( .A(n4981), .ZN(n4976) );
  NOR2_X1 U5324 ( .A1(n5005), .A2(n5002), .ZN(n5001) );
  INV_X1 U5325 ( .A(n9202), .ZN(n5002) );
  INV_X1 U5326 ( .A(n6590), .ZN(n5005) );
  NOR2_X1 U5327 ( .A1(n9667), .A2(n9862), .ZN(n9636) );
  NOR2_X1 U5328 ( .A1(n9683), .A2(n4923), .ZN(n4922) );
  INV_X1 U5329 ( .A(n4924), .ZN(n4923) );
  INV_X1 U5330 ( .A(n9691), .ZN(n5015) );
  NAND2_X1 U5331 ( .A1(n5020), .A2(n6584), .ZN(n5016) );
  NAND2_X1 U5332 ( .A1(n5018), .A2(n6584), .ZN(n5017) );
  INV_X1 U5333 ( .A(n9723), .ZN(n5018) );
  INV_X1 U5334 ( .A(n9327), .ZN(n6584) );
  AND2_X1 U5335 ( .A1(n9179), .A2(n9178), .ZN(n9244) );
  INV_X1 U5336 ( .A(n6525), .ZN(n4956) );
  AOI21_X1 U5337 ( .B1(n5029), .B2(n5031), .A(n5027), .ZN(n5026) );
  INV_X1 U5338 ( .A(n5829), .ZN(n5027) );
  AND2_X1 U5339 ( .A1(n5119), .A2(n5181), .ZN(n5055) );
  XNOR2_X1 U5340 ( .A(n5167), .B(n10619), .ZN(n5532) );
  NAND2_X1 U5341 ( .A1(n5399), .A2(n5152), .ZN(n4960) );
  OAI21_X1 U5342 ( .B1(n6714), .B2(n5143), .A(n5142), .ZN(n5145) );
  NAND2_X1 U5343 ( .A1(n5911), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5142) );
  INV_X1 U5344 ( .A(n8246), .ZN(n8232) );
  NAND2_X1 U5345 ( .A1(n7013), .A2(n8141), .ZN(n7017) );
  OAI21_X1 U5346 ( .B1(n7015), .B2(n7040), .A(n7014), .ZN(n7016) );
  NAND2_X1 U5347 ( .A1(n8313), .A2(n8312), .ZN(n8180) );
  NAND2_X1 U5348 ( .A1(n5090), .A2(n7820), .ZN(n5089) );
  CLKBUF_X1 U5349 ( .A(n8258), .Z(n8259) );
  NAND2_X1 U5350 ( .A1(n6013), .A2(n5111), .ZN(n4890) );
  OR2_X1 U5351 ( .A1(n7474), .A2(n6661), .ZN(n6050) );
  NAND2_X1 U5352 ( .A1(n4896), .A2(n4895), .ZN(n4894) );
  INV_X1 U5353 ( .A(n6636), .ZN(n4896) );
  NAND2_X1 U5354 ( .A1(n4944), .A2(n4895), .ZN(n4943) );
  INV_X1 U5355 ( .A(n6694), .ZN(n4944) );
  NAND2_X1 U5356 ( .A1(n6694), .A2(n6716), .ZN(n6961) );
  NAND2_X1 U5357 ( .A1(n4894), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4893) );
  OR2_X1 U5358 ( .A1(n6639), .A2(n7101), .ZN(n4909) );
  OR2_X1 U5359 ( .A1(n6697), .A2(n7101), .ZN(n4953) );
  NAND2_X1 U5360 ( .A1(n6697), .A2(n7101), .ZN(n7110) );
  NAND2_X1 U5361 ( .A1(n7798), .A2(n4535), .ZN(n4671) );
  OR2_X1 U5362 ( .A1(n8495), .A2(n4601), .ZN(n4936) );
  NAND2_X1 U5363 ( .A1(n8521), .A2(n4935), .ZN(n4934) );
  INV_X1 U5364 ( .A(n8523), .ZN(n4935) );
  OR2_X1 U5365 ( .A1(n8495), .A2(n8797), .ZN(n4938) );
  OR2_X1 U5366 ( .A1(n8587), .A2(n8560), .ZN(n8562) );
  NOR2_X1 U5367 ( .A1(n8539), .A2(n8775), .ZN(n8569) );
  OR2_X1 U5368 ( .A1(n8531), .A2(n4603), .ZN(n4903) );
  NAND2_X1 U5369 ( .A1(n8550), .A2(n4905), .ZN(n4904) );
  INV_X1 U5370 ( .A(n8551), .ZN(n4905) );
  OR2_X1 U5371 ( .A1(n6347), .A2(n6346), .ZN(n6358) );
  INV_X1 U5372 ( .A(n4620), .ZN(n6273) );
  NAND2_X1 U5373 ( .A1(n6242), .A2(n4779), .ZN(n4778) );
  NOR2_X1 U5374 ( .A1(n6254), .A2(n4736), .ZN(n4779) );
  AND2_X1 U5375 ( .A1(n4774), .A2(n8041), .ZN(n4797) );
  OAI21_X1 U5376 ( .B1(n6126), .B2(n4791), .A(n4787), .ZN(n6172) );
  AOI21_X1 U5377 ( .B1(n4790), .B2(n4789), .A(n4788), .ZN(n4787) );
  INV_X1 U5378 ( .A(n8028), .ZN(n4788) );
  NAND2_X1 U5379 ( .A1(n8040), .A2(n8041), .ZN(n7959) );
  OR2_X1 U5380 ( .A1(n7718), .A2(n7775), .ZN(n8014) );
  NAND2_X1 U5381 ( .A1(n6126), .A2(n4793), .ZN(n4792) );
  NAND2_X1 U5382 ( .A1(n4792), .A2(n4790), .ZN(n7733) );
  NAND2_X1 U5383 ( .A1(n6390), .A2(n6389), .ZN(n7434) );
  NAND2_X1 U5384 ( .A1(n8420), .A2(n7318), .ZN(n7982) );
  NAND2_X1 U5385 ( .A1(n6443), .A2(n7048), .ZN(n7739) );
  AND2_X1 U5386 ( .A1(n8133), .A2(n6499), .ZN(n7044) );
  AND2_X1 U5387 ( .A1(n6907), .A2(n6498), .ZN(n7047) );
  AND2_X1 U5388 ( .A1(n8630), .A2(n8629), .ZN(n8631) );
  OAI21_X1 U5389 ( .B1(n8642), .B2(n8112), .A(n7968), .ZN(n8628) );
  OR2_X1 U5390 ( .A1(n6429), .A2(n6428), .ZN(n6430) );
  OR2_X1 U5391 ( .A1(n6427), .A2(n6426), .ZN(n6428) );
  AND2_X1 U5392 ( .A1(n8108), .A2(n8109), .ZN(n8669) );
  NOR2_X1 U5393 ( .A1(n4785), .A2(n4783), .ZN(n4782) );
  INV_X1 U5394 ( .A(n8101), .ZN(n4783) );
  NAND2_X1 U5395 ( .A1(n8740), .A2(n4786), .ZN(n4784) );
  OR2_X1 U5396 ( .A1(n6315), .A2(n6314), .ZN(n8688) );
  OR2_X1 U5397 ( .A1(n8102), .A2(n7945), .ZN(n8691) );
  OR2_X1 U5398 ( .A1(n8737), .A2(n8745), .ZN(n8719) );
  OR2_X1 U5399 ( .A1(n8737), .A2(n8282), .ZN(n8713) );
  AOI21_X1 U5400 ( .B1(n8726), .B2(n6360), .A(n6297), .ZN(n8733) );
  AND2_X1 U5401 ( .A1(n8713), .A2(n8714), .ZN(n8731) );
  INV_X1 U5402 ( .A(n8813), .ZN(n8765) );
  INV_X1 U5403 ( .A(n8808), .ZN(n8768) );
  OR2_X1 U5404 ( .A1(n7023), .A2(n8133), .ZN(n8770) );
  INV_X1 U5405 ( .A(n4856), .ZN(n4855) );
  INV_X1 U5406 ( .A(n4864), .ZN(n4860) );
  NAND2_X1 U5407 ( .A1(n4861), .A2(n4864), .ZN(n7862) );
  AND2_X1 U5408 ( .A1(n8124), .A2(n7023), .ZN(n8808) );
  INV_X1 U5409 ( .A(n8770), .ZN(n8810) );
  AND2_X1 U5410 ( .A1(n6911), .A2(n6923), .ZN(n7025) );
  OR2_X1 U5411 ( .A1(n6009), .A2(n8145), .ZN(n10208) );
  NAND2_X1 U5412 ( .A1(n6439), .A2(n6487), .ZN(n8813) );
  NAND2_X1 U5413 ( .A1(n4610), .A2(n7014), .ZN(n6439) );
  INV_X1 U5414 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U5415 ( .A1(n4762), .A2(n4761), .ZN(n6436) );
  AOI21_X1 U5416 ( .B1(n4526), .B2(P2_IR_REG_31__SCAN_IN), .A(
        P2_IR_REG_20__SCAN_IN), .ZN(n4761) );
  NAND2_X1 U5417 ( .A1(n6208), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4762) );
  NOR2_X1 U5418 ( .A1(n6105), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n6112) );
  OR2_X1 U5419 ( .A1(n6080), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n6105) );
  INV_X1 U5420 ( .A(n9006), .ZN(n4652) );
  NAND2_X1 U5421 ( .A1(n4658), .A2(n4665), .ZN(n4657) );
  INV_X1 U5422 ( .A(n4660), .ZN(n4658) );
  NAND2_X1 U5423 ( .A1(n4656), .A2(n4655), .ZN(n4654) );
  NAND2_X1 U5424 ( .A1(n4664), .A2(n9022), .ZN(n4655) );
  NAND2_X1 U5425 ( .A1(n4660), .A2(n4663), .ZN(n4656) );
  INV_X1 U5426 ( .A(n4666), .ZN(n4663) );
  NAND2_X1 U5427 ( .A1(n5554), .A2(n5555), .ZN(n7536) );
  NAND2_X1 U5428 ( .A1(n9386), .A2(n5319), .ZN(n5304) );
  NOR2_X1 U5429 ( .A1(n5073), .A2(n5071), .ZN(n5070) );
  INV_X1 U5430 ( .A(n7538), .ZN(n5071) );
  NOR2_X1 U5431 ( .A1(n5073), .A2(n5551), .ZN(n5072) );
  NAND2_X1 U5432 ( .A1(n5262), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5711) );
  INV_X1 U5433 ( .A(n5689), .ZN(n5262) );
  OR2_X1 U5434 ( .A1(n5496), .A2(n10055), .ZN(n5367) );
  OR2_X1 U5435 ( .A1(n5733), .A2(n9018), .ZN(n5747) );
  INV_X1 U5436 ( .A(n5767), .ZN(n5265) );
  AOI21_X1 U5437 ( .B1(n9022), .B2(n4667), .A(n4538), .ZN(n4666) );
  OR2_X1 U5438 ( .A1(n5711), .A2(n7590), .ZN(n5731) );
  NAND2_X1 U5439 ( .A1(n5083), .A2(n4583), .ZN(n4644) );
  NOR2_X1 U5440 ( .A1(n4646), .A2(n9087), .ZN(n4641) );
  NAND2_X1 U5441 ( .A1(n4643), .A2(n5082), .ZN(n4642) );
  NAND2_X1 U5442 ( .A1(n7034), .A2(n5397), .ZN(n4622) );
  NOR4_X1 U5443 ( .A1(n9256), .A2(n9255), .A3(n9254), .A4(n9253), .ZN(n9291)
         );
  OR2_X1 U5444 ( .A1(n5361), .A2(n7330), .ZN(n5300) );
  OAI21_X1 U5445 ( .B1(n6593), .B2(n4546), .A(n4992), .ZN(n4991) );
  NAND2_X1 U5446 ( .A1(n6593), .A2(n4996), .ZN(n4992) );
  NOR2_X1 U5447 ( .A1(n6593), .A2(n4994), .ZN(n4993) );
  INV_X1 U5448 ( .A(n4996), .ZN(n4994) );
  NAND2_X1 U5449 ( .A1(n6593), .A2(n9572), .ZN(n4995) );
  AND2_X1 U5450 ( .A1(n6782), .A2(n9397), .ZN(n9101) );
  NAND2_X1 U5451 ( .A1(n9586), .A2(n9215), .ZN(n9568) );
  AND2_X1 U5452 ( .A1(n9264), .A2(n9207), .ZN(n9620) );
  NAND2_X1 U5453 ( .A1(n6586), .A2(n9199), .ZN(n9663) );
  NAND2_X1 U5454 ( .A1(n9728), .A2(n9879), .ZN(n9712) );
  NAND2_X1 U5455 ( .A1(n5022), .A2(n9192), .ZN(n9707) );
  OR2_X1 U5456 ( .A1(n9722), .A2(n9723), .ZN(n5022) );
  NAND2_X1 U5457 ( .A1(n9747), .A2(n9183), .ZN(n9722) );
  NOR2_X1 U5458 ( .A1(n9045), .A2(n4533), .ZN(n9740) );
  AOI21_X1 U5459 ( .B1(n4967), .B2(n4965), .A(n4554), .ZN(n4964) );
  INV_X1 U5460 ( .A(n4536), .ZN(n4965) );
  OR2_X1 U5461 ( .A1(n9951), .A2(n9374), .ZN(n4971) );
  NOR2_X1 U5462 ( .A1(n7846), .A2(n9172), .ZN(n5011) );
  INV_X1 U5463 ( .A(n9244), .ZN(n7846) );
  OAI21_X1 U5464 ( .B1(n7522), .B2(n5008), .A(n5006), .ZN(n6581) );
  INV_X1 U5465 ( .A(n5007), .ZN(n5006) );
  OAI21_X1 U5466 ( .B1(n4524), .B2(n5008), .A(n9175), .ZN(n5007) );
  NAND2_X1 U5467 ( .A1(n9941), .A2(n9942), .ZN(n9940) );
  NAND2_X1 U5468 ( .A1(n7522), .A2(n4524), .ZN(n7658) );
  OR2_X1 U5469 ( .A1(n7524), .A2(n9240), .ZN(n7522) );
  OR2_X1 U5470 ( .A1(n9962), .A2(n7226), .ZN(n9148) );
  AND2_X1 U5471 ( .A1(n9578), .A2(n9577), .ZN(n9759) );
  NAND2_X1 U5472 ( .A1(n5810), .A2(n5809), .ZN(n9782) );
  AND2_X1 U5473 ( .A1(n9222), .A2(n9292), .ZN(n10122) );
  XNOR2_X1 U5474 ( .A(n7930), .B(n7929), .ZN(n8157) );
  AND3_X1 U5475 ( .A1(n5225), .A2(n4839), .A3(n4837), .ZN(n4836) );
  INV_X1 U5476 ( .A(n5215), .ZN(n4837) );
  INV_X1 U5477 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5227) );
  NAND2_X1 U5478 ( .A1(n5246), .A2(n5238), .ZN(n5242) );
  AND2_X1 U5479 ( .A1(n5805), .A2(n5785), .ZN(n5803) );
  NAND2_X1 U5480 ( .A1(n4584), .A2(n4718), .ZN(n4717) );
  OAI21_X1 U5481 ( .B1(n5725), .B2(n5196), .A(n5198), .ZN(n5283) );
  NAND2_X1 U5482 ( .A1(n5708), .A2(n5252), .ZN(n5066) );
  NAND2_X1 U5483 ( .A1(n5624), .A2(n5233), .ZN(n5248) );
  NAND2_X1 U5484 ( .A1(n5056), .A2(n5181), .ZN(n5645) );
  NAND2_X1 U5485 ( .A1(n4696), .A2(n4700), .ZN(n5603) );
  NAND2_X1 U5486 ( .A1(n5557), .A2(n4701), .ZN(n4696) );
  OAI21_X1 U5487 ( .B1(n5557), .B2(n5556), .A(n5174), .ZN(n5578) );
  NAND2_X1 U5488 ( .A1(n5377), .A2(n5376), .ZN(n5399) );
  NAND2_X1 U5489 ( .A1(n8380), .A2(n8231), .ZN(n8247) );
  AOI21_X1 U5490 ( .B1(n5094), .B2(n5096), .A(n4586), .ZN(n5092) );
  AND2_X1 U5491 ( .A1(n6326), .A2(n6325), .ZN(n8305) );
  XNOR2_X1 U5492 ( .A(n5091), .B(n7820), .ZN(n7822) );
  INV_X2 U5493 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10634) );
  INV_X1 U5494 ( .A(n8645), .ZN(n8386) );
  AND3_X1 U5495 ( .A1(n6278), .A2(n6277), .A3(n6276), .ZN(n8754) );
  AND4_X1 U5496 ( .A1(n6253), .A2(n6252), .A3(n6251), .A4(n6250), .ZN(n8753)
         );
  NAND2_X1 U5497 ( .A1(n7275), .A2(n7274), .ZN(n7411) );
  OAI21_X1 U5498 ( .B1(n4690), .B2(n8135), .A(n7014), .ZN(n4689) );
  OR2_X1 U5499 ( .A1(n7474), .A2(n7055), .ZN(n6040) );
  NAND2_X1 U5500 ( .A1(n4900), .A2(n6647), .ZN(n7626) );
  NAND2_X1 U5501 ( .A1(n4947), .A2(n4946), .ZN(n4677) );
  NAND2_X1 U5502 ( .A1(n6704), .A2(n6765), .ZN(n4946) );
  INV_X1 U5503 ( .A(n7625), .ZN(n4898) );
  INV_X1 U5504 ( .A(n4675), .ZN(n7697) );
  OR2_X1 U5505 ( .A1(P2_U3150), .A2(n6687), .ZN(n8565) );
  AND3_X1 U5506 ( .A1(n4904), .A2(n8577), .A3(n4903), .ZN(n8580) );
  NOR2_X1 U5507 ( .A1(n8583), .A2(n8582), .ZN(n8584) );
  OR2_X1 U5508 ( .A1(n6932), .A2(n8588), .ZN(n10152) );
  XNOR2_X1 U5509 ( .A(n7939), .B(n4758), .ZN(n8619) );
  NAND2_X1 U5510 ( .A1(n6374), .A2(n6373), .ZN(n8615) );
  NAND2_X1 U5511 ( .A1(n6117), .A2(n6116), .ZN(n10201) );
  AND2_X1 U5512 ( .A1(n8141), .A2(n6438), .ZN(n7307) );
  NAND2_X1 U5513 ( .A1(n6924), .A2(n6923), .ZN(n10169) );
  NAND2_X1 U5514 ( .A1(n6345), .A2(n6344), .ZN(n8897) );
  AND2_X1 U5515 ( .A1(n5112), .A2(n6015), .ZN(n4800) );
  NAND2_X1 U5516 ( .A1(n4630), .A2(n9097), .ZN(n4629) );
  INV_X1 U5517 ( .A(n8990), .ZN(n4630) );
  OAI21_X1 U5518 ( .B1(n8990), .B2(n4625), .A(n8995), .ZN(n4624) );
  NAND2_X1 U5519 ( .A1(n4626), .A2(n9097), .ZN(n4625) );
  NAND2_X1 U5520 ( .A1(n4527), .A2(n5058), .ZN(n5057) );
  NAND2_X1 U5521 ( .A1(n4527), .A2(n9031), .ZN(n5059) );
  INV_X1 U5522 ( .A(n5060), .ZN(n5058) );
  OR2_X1 U5523 ( .A1(n6783), .A2(n6795), .ZN(n5129) );
  NAND2_X1 U5524 ( .A1(n4529), .A2(n5079), .ZN(n5075) );
  NAND2_X1 U5525 ( .A1(n4632), .A2(n4556), .ZN(n5076) );
  NAND2_X1 U5526 ( .A1(n5745), .A2(n5744), .ZN(n9698) );
  NAND2_X1 U5527 ( .A1(n5895), .A2(n5894), .ZN(n9104) );
  NAND2_X1 U5528 ( .A1(n8156), .A2(n8155), .ZN(n9545) );
  NAND2_X1 U5529 ( .A1(n4977), .A2(n4981), .ZN(n9606) );
  NAND2_X1 U5530 ( .A1(n6555), .A2(n4978), .ZN(n4977) );
  AND2_X1 U5531 ( .A1(n9752), .A2(n9751), .ZN(n9825) );
  INV_X1 U5532 ( .A(n10019), .ZN(n9699) );
  OR2_X1 U5533 ( .A1(n9907), .A2(n6562), .ZN(n6564) );
  INV_X1 U5534 ( .A(n9743), .ZN(n9887) );
  INV_X1 U5535 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5254) );
  NAND2_X1 U5536 ( .A1(n5065), .A2(n5064), .ZN(n5255) );
  AOI21_X1 U5537 ( .B1(n5067), .B2(n9899), .A(n9899), .ZN(n5064) );
  INV_X1 U5538 ( .A(n9163), .ZN(n4817) );
  INV_X1 U5539 ( .A(n9161), .ZN(n4819) );
  NOR2_X1 U5540 ( .A1(n9126), .A2(n4801), .ZN(n9146) );
  NOR2_X1 U5541 ( .A1(n8037), .A2(n8124), .ZN(n4775) );
  OAI21_X1 U5542 ( .B1(n8043), .B2(n4767), .A(n4566), .ZN(n8054) );
  INV_X1 U5543 ( .A(n4768), .ZN(n4767) );
  NAND2_X1 U5544 ( .A1(n4826), .A2(n4823), .ZN(n4822) );
  AOI21_X1 U5545 ( .B1(n8064), .B2(n8072), .A(n4736), .ZN(n4735) );
  AND2_X1 U5546 ( .A1(n9250), .A2(n9201), .ZN(n4809) );
  NAND2_X1 U5547 ( .A1(n9261), .A2(n9222), .ZN(n4810) );
  NOR2_X1 U5548 ( .A1(n8102), .A2(n4739), .ZN(n4738) );
  NAND2_X1 U5549 ( .A1(n4740), .A2(n4742), .ZN(n8103) );
  INV_X1 U5550 ( .A(SI_8_), .ZN(n10617) );
  INV_X1 U5551 ( .A(n4882), .ZN(n4878) );
  INV_X1 U5552 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n4843) );
  INV_X1 U5553 ( .A(n9040), .ZN(n5085) );
  AND2_X1 U5554 ( .A1(n6577), .A2(n9162), .ZN(n9238) );
  NOR2_X1 U5555 ( .A1(n9152), .A2(n6579), .ZN(n9236) );
  NAND2_X1 U5556 ( .A1(n4930), .A2(n10117), .ZN(n4929) );
  INV_X1 U5557 ( .A(n4931), .ZN(n4930) );
  NAND2_X1 U5558 ( .A1(n7730), .A2(n4932), .ZN(n4931) );
  INV_X1 U5559 ( .A(n5030), .ZN(n5029) );
  OAI21_X1 U5560 ( .B1(n5803), .B2(n5031), .A(n5827), .ZN(n5030) );
  INV_X1 U5561 ( .A(n5805), .ZN(n5031) );
  NAND2_X1 U5562 ( .A1(n5045), .A2(n4555), .ZN(n5044) );
  NAND2_X1 U5563 ( .A1(n5046), .A2(n5166), .ZN(n5045) );
  INV_X1 U5564 ( .A(SI_10_), .ZN(n10619) );
  NOR2_X1 U5565 ( .A1(n5468), .A2(n5048), .ZN(n5047) );
  INV_X1 U5566 ( .A(n5158), .ZN(n5048) );
  INV_X1 U5567 ( .A(SI_15_), .ZN(n10564) );
  INV_X1 U5568 ( .A(SI_18_), .ZN(n10423) );
  INV_X1 U5569 ( .A(SI_24_), .ZN(n10577) );
  INV_X1 U5570 ( .A(SI_11_), .ZN(n10461) );
  AND2_X1 U5571 ( .A1(n8341), .A2(n8201), .ZN(n8211) );
  OR2_X1 U5572 ( .A1(n8205), .A2(n8204), .ZN(n8213) );
  INV_X1 U5573 ( .A(n8213), .ZN(n8214) );
  INV_X1 U5574 ( .A(n5113), .ZN(n5111) );
  NAND2_X1 U5575 ( .A1(n6695), .A2(n6962), .ZN(n6964) );
  NAND2_X1 U5576 ( .A1(n4942), .A2(n6961), .ZN(n6695) );
  NAND2_X1 U5577 ( .A1(n4943), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4942) );
  NAND2_X1 U5578 ( .A1(n4951), .A2(n7110), .ZN(n7112) );
  INV_X1 U5579 ( .A(n4952), .ZN(n4951) );
  INV_X1 U5580 ( .A(n7708), .ZN(n4901) );
  OR2_X1 U5581 ( .A1(n7707), .A2(n6651), .ZN(n6652) );
  NAND2_X1 U5582 ( .A1(n4675), .A2(n6705), .ZN(n7795) );
  AND2_X1 U5583 ( .A1(n4673), .A2(n4672), .ZN(n8472) );
  NAND2_X1 U5584 ( .A1(n8447), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4672) );
  NOR2_X1 U5585 ( .A1(n8494), .A2(n8493), .ZN(n8518) );
  NOR2_X1 U5586 ( .A1(n6307), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n4614) );
  INV_X1 U5587 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10565) );
  NOR2_X1 U5588 ( .A1(n6262), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n4620) );
  INV_X1 U5589 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10660) );
  NOR2_X1 U5590 ( .A1(n6211), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n4619) );
  INV_X1 U5591 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10459) );
  NOR2_X1 U5592 ( .A1(n6177), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n4618) );
  INV_X1 U5593 ( .A(n4793), .ZN(n4789) );
  OR2_X1 U5594 ( .A1(n7819), .A2(n7879), .ZN(n8040) );
  NOR2_X1 U5595 ( .A1(n6396), .A2(n4884), .ZN(n4882) );
  NAND2_X1 U5596 ( .A1(n4883), .A2(n6394), .ZN(n4881) );
  INV_X1 U5597 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10440) );
  NAND2_X1 U5598 ( .A1(n4796), .A2(n7306), .ZN(n6056) );
  NAND2_X1 U5599 ( .A1(n6012), .A2(n5114), .ZN(n5113) );
  INV_X1 U5600 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5114) );
  AOI21_X1 U5601 ( .B1(n4666), .B2(n4662), .A(n4661), .ZN(n4660) );
  INV_X1 U5602 ( .A(n9080), .ZN(n4661) );
  INV_X1 U5603 ( .A(n4667), .ZN(n4662) );
  INV_X1 U5604 ( .A(n9087), .ZN(n4638) );
  AND2_X1 U5605 ( .A1(n5220), .A2(n5233), .ZN(n4647) );
  OR2_X1 U5606 ( .A1(n5470), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5537) );
  AOI21_X1 U5607 ( .B1(n9572), .B2(n4998), .A(n4997), .ZN(n4996) );
  INV_X1 U5608 ( .A(n9215), .ZN(n4998) );
  INV_X1 U5609 ( .A(n9216), .ZN(n4997) );
  OR2_X1 U5610 ( .A1(n9560), .A2(n6565), .ZN(n9283) );
  INV_X1 U5611 ( .A(n4978), .ZN(n4973) );
  NAND2_X1 U5612 ( .A1(n4964), .A2(n4966), .ZN(n4962) );
  INV_X1 U5613 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5610) );
  INV_X1 U5614 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5541) );
  NAND2_X1 U5615 ( .A1(n9302), .A2(n7156), .ZN(n9126) );
  AND2_X1 U5616 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5382) );
  INV_X1 U5617 ( .A(n9289), .ZN(n6782) );
  NAND2_X1 U5618 ( .A1(n6588), .A2(n9202), .ZN(n9646) );
  NOR2_X1 U5619 ( .A1(n7651), .A2(n4931), .ZN(n9954) );
  AND2_X1 U5620 ( .A1(n5963), .A2(n9350), .ZN(n6605) );
  INV_X1 U5621 ( .A(n7929), .ZN(n5033) );
  AND2_X1 U5622 ( .A1(n6369), .A2(n5915), .ZN(n5916) );
  AND2_X1 U5623 ( .A1(n5909), .A2(n5883), .ZN(n5884) );
  AND2_X1 U5624 ( .A1(n5878), .A2(n5855), .ZN(n5876) );
  AOI21_X1 U5625 ( .B1(n5037), .B2(n5040), .A(n4594), .ZN(n5035) );
  INV_X1 U5626 ( .A(n5037), .ZN(n5036) );
  INV_X1 U5627 ( .A(n5706), .ZN(n4718) );
  NOR2_X1 U5628 ( .A1(n4720), .A2(n4592), .ZN(n4715) );
  OAI21_X1 U5629 ( .B1(n4721), .B2(n5040), .A(n5039), .ZN(n4720) );
  INV_X1 U5630 ( .A(n5195), .ZN(n4716) );
  INV_X1 U5631 ( .A(n7931), .ZN(n5911) );
  NOR2_X1 U5632 ( .A1(n5282), .A2(n4724), .ZN(n4723) );
  INV_X1 U5633 ( .A(n5198), .ZN(n4724) );
  AOI21_X1 U5634 ( .B1(n4723), .B2(n5196), .A(n4722), .ZN(n4721) );
  INV_X1 U5635 ( .A(n5203), .ZN(n4722) );
  INV_X1 U5636 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5185) );
  AOI21_X1 U5637 ( .B1(n4701), .B2(n5556), .A(n4563), .ZN(n4700) );
  NAND2_X1 U5638 ( .A1(n5049), .A2(n5047), .ZN(n5529) );
  NAND2_X1 U5639 ( .A1(n5422), .A2(n5156), .ZN(n5049) );
  NAND2_X1 U5640 ( .A1(n4506), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5042) );
  AND2_X1 U5641 ( .A1(n4847), .A2(n4846), .ZN(n4844) );
  INV_X1 U5642 ( .A(n5095), .ZN(n5094) );
  OAI21_X1 U5643 ( .B1(n7875), .B2(n5096), .A(n8167), .ZN(n5095) );
  INV_X1 U5644 ( .A(n7903), .ZN(n5096) );
  NAND2_X1 U5645 ( .A1(n4609), .A2(n4552), .ZN(n5091) );
  AND2_X1 U5646 ( .A1(n8340), .A2(n8188), .ZN(n8277) );
  NAND2_X1 U5647 ( .A1(n7411), .A2(n5107), .ZN(n5110) );
  AND2_X1 U5648 ( .A1(n8376), .A2(n8226), .ZN(n8301) );
  INV_X1 U5649 ( .A(n8664), .ZN(n8306) );
  NOR2_X1 U5650 ( .A1(n8321), .A2(n5100), .ZN(n5099) );
  INV_X1 U5651 ( .A(n8179), .ZN(n5100) );
  AND2_X1 U5652 ( .A1(n8300), .A2(n8222), .ZN(n8329) );
  NAND2_X1 U5653 ( .A1(n7550), .A2(n8020), .ZN(n5109) );
  INV_X1 U5654 ( .A(n7681), .ZN(n5106) );
  OR2_X1 U5655 ( .A1(n7683), .A2(n7684), .ZN(n4609) );
  OR2_X1 U5656 ( .A1(n8199), .A2(n8198), .ZN(n8356) );
  AND2_X1 U5657 ( .A1(n8276), .A2(n8184), .ZN(n8367) );
  INV_X1 U5658 ( .A(n4749), .ZN(n8129) );
  AOI21_X1 U5659 ( .B1(n4760), .B2(n4759), .A(n4752), .ZN(n4749) );
  NOR3_X1 U5660 ( .A1(n7974), .A2(n8126), .A3(n7973), .ZN(n7975) );
  NOR2_X1 U5661 ( .A1(n7944), .A2(n4692), .ZN(n4691) );
  NAND2_X1 U5662 ( .A1(n8136), .A2(n7972), .ZN(n7973) );
  AND3_X1 U5663 ( .A1(n4755), .A2(n4754), .A3(n4753), .ZN(n8137) );
  AND2_X1 U5664 ( .A1(n7478), .A2(n7477), .ZN(n7976) );
  AND2_X1 U5665 ( .A1(n6335), .A2(n6334), .ZN(n8385) );
  CLKBUF_X1 U5666 ( .A(n7474), .Z(n6363) );
  NAND2_X1 U5667 ( .A1(n6930), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n10148) );
  OAI21_X1 U5668 ( .B1(n6036), .B2(n6692), .A(n6691), .ZN(n8428) );
  NAND2_X1 U5669 ( .A1(n6036), .A2(n6692), .ZN(n6691) );
  OR2_X1 U5670 ( .A1(n4893), .A2(n4892), .ZN(n6958) );
  INV_X1 U5671 ( .A(n6956), .ZN(n4892) );
  OAI21_X1 U5672 ( .B1(n6974), .B2(n6074), .A(n4674), .ZN(n6962) );
  NAND2_X1 U5673 ( .A1(n6974), .A2(n6074), .ZN(n4674) );
  NAND2_X1 U5674 ( .A1(n4941), .A2(n6961), .ZN(n6966) );
  INV_X1 U5675 ( .A(n4942), .ZN(n4941) );
  NAND2_X1 U5676 ( .A1(n4952), .A2(n7110), .ZN(n6698) );
  NAND2_X1 U5677 ( .A1(n6701), .A2(n4945), .ZN(n7262) );
  OR2_X1 U5678 ( .A1(n6700), .A2(n6741), .ZN(n4945) );
  NAND2_X1 U5679 ( .A1(n7120), .A2(n4915), .ZN(n4918) );
  AND2_X1 U5680 ( .A1(n7266), .A2(n6642), .ZN(n4915) );
  NAND2_X1 U5681 ( .A1(n4918), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4916) );
  AND2_X1 U5682 ( .A1(n4917), .A2(n4916), .ZN(n7341) );
  OR2_X1 U5683 ( .A1(n7262), .A2(n4680), .ZN(n4679) );
  OR2_X1 U5684 ( .A1(n7332), .A2(n6676), .ZN(n4680) );
  OR2_X1 U5685 ( .A1(n6701), .A2(n7332), .ZN(n4678) );
  OR2_X1 U5686 ( .A1(n7262), .A2(n6676), .ZN(n4681) );
  NAND2_X1 U5687 ( .A1(n4902), .A2(n7630), .ZN(n4900) );
  INV_X1 U5688 ( .A(n6648), .ZN(n4902) );
  AND3_X1 U5689 ( .A1(n4900), .A2(n6647), .A3(P2_REG1_REG_9__SCAN_IN), .ZN(
        n7625) );
  XNOR2_X1 U5690 ( .A(n7795), .B(n7796), .ZN(n6706) );
  AND2_X1 U5691 ( .A1(n6160), .A2(n6005), .ZN(n6185) );
  AOI21_X1 U5692 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n8447), .A(n8438), .ZN(
        n8459) );
  NOR2_X1 U5693 ( .A1(n8478), .A2(n8477), .ZN(n8494) );
  AOI21_X1 U5694 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n8492), .A(n8485), .ZN(
        n8504) );
  AOI21_X1 U5695 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n8537), .A(n8530), .ZN(
        n8548) );
  OR2_X1 U5696 ( .A1(n6329), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6347) );
  NAND2_X1 U5697 ( .A1(n6292), .A2(n6291), .ZN(n6300) );
  INV_X1 U5698 ( .A(n6293), .ZN(n6292) );
  OR2_X1 U5699 ( .A1(n6282), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6293) );
  NAND2_X1 U5700 ( .A1(n4620), .A2(n10565), .ZN(n6282) );
  NAND2_X1 U5701 ( .A1(n6247), .A2(n10660), .ZN(n6262) );
  INV_X1 U5702 ( .A(n6248), .ZN(n6247) );
  OR2_X1 U5703 ( .A1(n6235), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6248) );
  NAND2_X1 U5704 ( .A1(n4619), .A2(n10388), .ZN(n6235) );
  INV_X1 U5705 ( .A(n4619), .ZN(n6223) );
  NAND2_X1 U5706 ( .A1(n6200), .A2(n6199), .ZN(n6211) );
  INV_X1 U5707 ( .A(n6201), .ZN(n6200) );
  NAND2_X1 U5708 ( .A1(n4618), .A2(n10459), .ZN(n6201) );
  INV_X1 U5709 ( .A(n4618), .ZN(n6189) );
  NAND2_X1 U5710 ( .A1(n4869), .A2(n4872), .ZN(n7784) );
  INV_X1 U5711 ( .A(n4873), .ZN(n4872) );
  OAI21_X1 U5712 ( .B1(n7955), .B2(n4874), .A(n6403), .ZN(n4873) );
  OR2_X1 U5713 ( .A1(n6165), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6177) );
  NAND2_X1 U5714 ( .A1(n4615), .A2(n6150), .ZN(n6165) );
  INV_X1 U5715 ( .A(n6151), .ZN(n4615) );
  NAND2_X1 U5716 ( .A1(n4871), .A2(n6402), .ZN(n7735) );
  NAND2_X1 U5717 ( .A1(n7666), .A2(n7955), .ZN(n4871) );
  NAND2_X1 U5718 ( .A1(n6401), .A2(n6400), .ZN(n7666) );
  NAND2_X1 U5719 ( .A1(n4617), .A2(n4616), .ZN(n6151) );
  INV_X1 U5720 ( .A(n6132), .ZN(n4617) );
  INV_X1 U5721 ( .A(n8412), .ZN(n7775) );
  NAND2_X1 U5722 ( .A1(n4876), .A2(n4879), .ZN(n7563) );
  NAND2_X1 U5723 ( .A1(n7462), .A2(n4882), .ZN(n4876) );
  OR2_X1 U5724 ( .A1(n6099), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6120) );
  NAND2_X1 U5725 ( .A1(n6119), .A2(n6118), .ZN(n6132) );
  INV_X1 U5726 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6118) );
  INV_X1 U5727 ( .A(n6120), .ZN(n6119) );
  OAI21_X1 U5728 ( .B1(n7462), .B2(n6394), .A(n4883), .ZN(n7512) );
  NAND2_X1 U5729 ( .A1(n6087), .A2(n6086), .ZN(n6099) );
  INV_X1 U5730 ( .A(n6088), .ZN(n6087) );
  AND2_X1 U5731 ( .A1(n4866), .A2(n6387), .ZN(n4865) );
  NAND2_X1 U5732 ( .A1(n10440), .A2(n10634), .ZN(n6088) );
  NAND2_X1 U5733 ( .A1(n7987), .A2(n7982), .ZN(n7313) );
  NAND2_X1 U5734 ( .A1(n7313), .A2(n7314), .ZN(n7312) );
  INV_X1 U5735 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6929) );
  NAND2_X1 U5736 ( .A1(n8623), .A2(n8810), .ZN(n4887) );
  OR2_X1 U5737 ( .A1(n8112), .A2(n8113), .ZN(n8643) );
  NOR2_X1 U5738 ( .A1(n4782), .A2(n4711), .ZN(n4705) );
  INV_X1 U5739 ( .A(n4708), .ZN(n4704) );
  AOI21_X1 U5740 ( .B1(n8740), .B2(n4710), .A(n4709), .ZN(n4708) );
  INV_X1 U5741 ( .A(n8643), .ZN(n8641) );
  INV_X1 U5742 ( .A(n8669), .ZN(n8662) );
  AND2_X1 U5743 ( .A1(n8662), .A2(n8658), .ZN(n8659) );
  OR2_X1 U5744 ( .A1(n8678), .A2(n8657), .ZN(n8660) );
  NAND2_X1 U5745 ( .A1(n8094), .A2(n4703), .ZN(n8700) );
  INV_X1 U5746 ( .A(n4850), .ZN(n4849) );
  OAI21_X1 U5747 ( .B1(n4537), .B2(n4851), .A(n8718), .ZN(n4850) );
  INV_X1 U5748 ( .A(n8719), .ZN(n4851) );
  INV_X1 U5749 ( .A(n6416), .ZN(n8743) );
  NOR2_X1 U5750 ( .A1(n8755), .A2(n4777), .ZN(n4776) );
  INV_X1 U5751 ( .A(n8066), .ZN(n4777) );
  NAND2_X1 U5752 ( .A1(n6261), .A2(n6260), .ZN(n8365) );
  INV_X1 U5753 ( .A(n8795), .ZN(n8769) );
  AND3_X1 U5754 ( .A1(n6268), .A2(n6267), .A3(n6266), .ZN(n8771) );
  OAI21_X1 U5755 ( .B1(n8791), .B2(n8068), .A(n8063), .ZN(n8780) );
  NAND2_X1 U5756 ( .A1(n4799), .A2(n8056), .ZN(n8791) );
  NAND2_X1 U5757 ( .A1(n8805), .A2(n8057), .ZN(n4799) );
  AND2_X1 U5758 ( .A1(n6486), .A2(n6923), .ZN(n6922) );
  NAND2_X1 U5759 ( .A1(n7739), .A2(n10208), .ZN(n10196) );
  NOR2_X1 U5760 ( .A1(n5113), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n5112) );
  NAND2_X1 U5761 ( .A1(n4764), .A2(n4765), .ZN(n6257) );
  INV_X1 U5762 ( .A(n6208), .ZN(n4764) );
  AND2_X1 U5763 ( .A1(n6142), .A2(n6141), .ZN(n6146) );
  CLKBUF_X1 U5764 ( .A(n6079), .Z(n6080) );
  INV_X1 U5765 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4669) );
  INV_X1 U5766 ( .A(n8991), .ZN(n4626) );
  AOI21_X1 U5767 ( .B1(n5900), .B2(n6984), .A(n5324), .ZN(n5326) );
  INV_X1 U5768 ( .A(n5080), .ZN(n5078) );
  AND2_X1 U5769 ( .A1(n5079), .A2(n9015), .ZN(n5077) );
  NAND2_X1 U5770 ( .A1(n5584), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5611) );
  INV_X1 U5771 ( .A(n9101), .ZN(n9089) );
  INV_X1 U5772 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5497) );
  NAND2_X1 U5773 ( .A1(n4523), .A2(n9015), .ZN(n9014) );
  OR2_X1 U5774 ( .A1(n5765), .A2(n9025), .ZN(n5767) );
  NOR2_X1 U5775 ( .A1(n5542), .A2(n5541), .ZN(n5562) );
  NAND2_X1 U5776 ( .A1(n7537), .A2(n7538), .ZN(n5074) );
  XNOR2_X1 U5777 ( .A(n5349), .B(n5898), .ZN(n5351) );
  NAND2_X1 U5778 ( .A1(n5263), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5733) );
  INV_X1 U5779 ( .A(n4635), .ZN(n4631) );
  OAI21_X1 U5780 ( .B1(n4646), .B2(n4637), .A(n4636), .ZN(n4635) );
  NAND2_X1 U5781 ( .A1(n5081), .A2(n4638), .ZN(n4637) );
  OR2_X1 U5782 ( .A1(n4644), .A2(n9050), .ZN(n4636) );
  NAND2_X1 U5783 ( .A1(n9037), .A2(n4639), .ZN(n4632) );
  NAND2_X1 U5784 ( .A1(n4640), .A2(n4644), .ZN(n4639) );
  INV_X1 U5785 ( .A(n4641), .ZN(n4640) );
  NAND2_X1 U5786 ( .A1(n5261), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5689) );
  INV_X1 U5787 ( .A(n5649), .ZN(n5261) );
  OAI21_X1 U5788 ( .B1(n8161), .B2(n9360), .A(n9257), .ZN(n9338) );
  OR2_X1 U5789 ( .A1(n5361), .A2(n5330), .ZN(n5331) );
  NAND3_X1 U5790 ( .A1(n5318), .A2(n4539), .A3(n5317), .ZN(n6509) );
  OR2_X1 U5791 ( .A1(n5360), .A2(n6794), .ZN(n5317) );
  OR2_X1 U5792 ( .A1(n5969), .A2(n6997), .ZN(n5318) );
  OR2_X1 U5793 ( .A1(n7588), .A2(n7589), .ZN(n7748) );
  OR2_X1 U5794 ( .A1(n7750), .A2(n7751), .ZN(n9521) );
  INV_X1 U5795 ( .A(n8162), .ZN(n9550) );
  INV_X1 U5796 ( .A(n4928), .ZN(n9593) );
  NAND2_X1 U5797 ( .A1(n5788), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5837) );
  NAND2_X1 U5798 ( .A1(n5000), .A2(n5003), .ZN(n9616) );
  AOI21_X1 U5799 ( .B1(n6590), .B2(n9250), .A(n5004), .ZN(n5003) );
  INV_X1 U5800 ( .A(n9262), .ZN(n5004) );
  NAND2_X1 U5801 ( .A1(n9646), .A2(n9653), .ZN(n9648) );
  AND2_X1 U5802 ( .A1(n9262), .A2(n9269), .ZN(n9631) );
  NAND2_X1 U5803 ( .A1(n6551), .A2(n6550), .ZN(n9654) );
  AND2_X1 U5804 ( .A1(n9200), .A2(n9202), .ZN(n9662) );
  NAND2_X1 U5805 ( .A1(n9728), .A2(n4921), .ZN(n9667) );
  AND2_X1 U5806 ( .A1(n4922), .A2(n9867), .ZN(n4921) );
  AOI21_X1 U5807 ( .B1(n5016), .B2(n5017), .A(n5015), .ZN(n5014) );
  NAND2_X1 U5808 ( .A1(n5013), .A2(n5016), .ZN(n9692) );
  OR2_X1 U5809 ( .A1(n9722), .A2(n5017), .ZN(n5013) );
  NAND2_X1 U5810 ( .A1(n9728), .A2(n4924), .ZN(n9696) );
  AND2_X1 U5811 ( .A1(n7888), .A2(n9296), .ZN(n9749) );
  NAND2_X1 U5812 ( .A1(n9749), .A2(n9748), .ZN(n9747) );
  AOI21_X1 U5813 ( .B1(n5011), .B2(n9943), .A(n9321), .ZN(n5009) );
  INV_X1 U5814 ( .A(n5011), .ZN(n5010) );
  OR2_X1 U5815 ( .A1(n5611), .A2(n5610), .ZN(n5629) );
  OR2_X1 U5816 ( .A1(n5629), .A2(n5628), .ZN(n5649) );
  NOR2_X1 U5817 ( .A1(n7651), .A2(n10108), .ZN(n7653) );
  NOR2_X1 U5818 ( .A1(n9969), .A2(n10096), .ZN(n7355) );
  NAND2_X1 U5819 ( .A1(n7355), .A2(n10103), .ZN(n7529) );
  AND2_X1 U5820 ( .A1(n9305), .A2(n9163), .ZN(n9237) );
  INV_X1 U5821 ( .A(n7397), .ZN(n4957) );
  AOI21_X1 U5822 ( .B1(n7397), .B2(n4956), .A(n4558), .ZN(n4955) );
  INV_X1 U5823 ( .A(n9237), .ZN(n7350) );
  NAND2_X1 U5824 ( .A1(n4920), .A2(n4919), .ZN(n9969) );
  NAND2_X1 U5825 ( .A1(n6757), .A2(n5441), .ZN(n4982) );
  NOR2_X1 U5826 ( .A1(n5446), .A2(n6818), .ZN(n5472) );
  NAND2_X1 U5827 ( .A1(n5447), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5446) );
  NOR2_X1 U5828 ( .A1(n9984), .A2(n9983), .ZN(n9987) );
  AND2_X1 U5829 ( .A1(n5382), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U5830 ( .A1(n9131), .A2(n9127), .ZN(n7156) );
  NAND2_X1 U5831 ( .A1(n9991), .A2(n6572), .ZN(n7284) );
  NOR2_X1 U5832 ( .A1(n10021), .A2(n10020), .ZN(n10024) );
  INV_X1 U5833 ( .A(n10116), .ZN(n10095) );
  NAND2_X1 U5834 ( .A1(n5962), .A2(n6605), .ZN(n10116) );
  AND4_X1 U5835 ( .A1(n6613), .A2(n6612), .A3(n6611), .A4(n7147), .ZN(n6620)
         );
  INV_X1 U5836 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5269) );
  INV_X1 U5837 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5272) );
  XNOR2_X1 U5838 ( .A(n5244), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5959) );
  XNOR2_X1 U5839 ( .A(n5946), .B(n5945), .ZN(n9352) );
  INV_X1 U5840 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5942) );
  INV_X1 U5841 ( .A(SI_20_), .ZN(n10419) );
  AOI21_X1 U5842 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_18__SCAN_IN), .ZN(n5067) );
  XNOR2_X1 U5843 ( .A(n5469), .B(n5468), .ZN(n6757) );
  NAND2_X1 U5844 ( .A1(n5049), .A2(n5158), .ZN(n5469) );
  NAND2_X1 U5845 ( .A1(n4960), .A2(n4532), .ZN(n4959) );
  NAND2_X1 U5846 ( .A1(n5147), .A2(n5146), .ZN(n5377) );
  AND2_X1 U5847 ( .A1(n5110), .A2(n5109), .ZN(n7682) );
  OR2_X1 U5848 ( .A1(n6066), .A2(n5131), .ZN(n6054) );
  OR2_X1 U5849 ( .A1(n6065), .A2(n6730), .ZN(n6053) );
  AND2_X1 U5850 ( .A1(n8291), .A2(n8290), .ZN(n8353) );
  NAND2_X1 U5851 ( .A1(n7874), .A2(n7875), .ZN(n7904) );
  AND2_X1 U5852 ( .A1(n6926), .A2(n7025), .ZN(n8337) );
  NAND2_X1 U5853 ( .A1(n5105), .A2(n5103), .ZN(n7683) );
  INV_X1 U5854 ( .A(n5104), .ZN(n5103) );
  NAND2_X1 U5855 ( .A1(n7411), .A2(n4547), .ZN(n5105) );
  OAI22_X1 U5856 ( .A1(n7681), .A2(n5109), .B1(n8413), .B2(n7680), .ZN(n5104)
         );
  INV_X1 U5857 ( .A(n4609), .ZN(n7773) );
  NAND2_X1 U5858 ( .A1(n6198), .A2(n6197), .ZN(n8048) );
  NAND2_X1 U5859 ( .A1(n5088), .A2(n5087), .ZN(n7872) );
  AND2_X1 U5860 ( .A1(n5088), .A2(n5089), .ZN(n7823) );
  INV_X1 U5861 ( .A(n8393), .ZN(n8381) );
  OR2_X1 U5862 ( .A1(n7133), .A2(n7637), .ZN(n8389) );
  NOR2_X1 U5863 ( .A1(n8394), .A2(n5102), .ZN(n5101) );
  INV_X1 U5864 ( .A(n8175), .ZN(n5102) );
  NAND2_X1 U5865 ( .A1(n8259), .A2(n8175), .ZN(n8395) );
  INV_X1 U5866 ( .A(n8384), .ZN(n8402) );
  INV_X1 U5867 ( .A(n7976), .ZN(n8607) );
  NAND2_X1 U5868 ( .A1(n6353), .A2(n6352), .ZN(n8645) );
  INV_X1 U5869 ( .A(n8385), .ZN(n8679) );
  INV_X1 U5870 ( .A(n8305), .ZN(n8693) );
  INV_X1 U5871 ( .A(n8282), .ZN(n8745) );
  INV_X1 U5872 ( .A(n8771), .ZN(n8744) );
  OR2_X1 U5873 ( .A1(n7474), .A2(n6058), .ZN(n6059) );
  OR2_X1 U5874 ( .A1(n6375), .A2(n7319), .ZN(n6049) );
  OR2_X1 U5875 ( .A1(n7471), .A2(n6660), .ZN(n6048) );
  NAND2_X1 U5876 ( .A1(n4894), .A2(n6956), .ZN(n6941) );
  NAND2_X1 U5877 ( .A1(n4943), .A2(n6961), .ZN(n6945) );
  AOI21_X1 U5878 ( .B1(n4895), .B2(n6667), .A(n6937), .ZN(n6954) );
  NAND2_X1 U5879 ( .A1(n4891), .A2(n6955), .ZN(n6960) );
  NAND2_X1 U5880 ( .A1(n4909), .A2(n7116), .ZN(n4908) );
  NAND2_X1 U5881 ( .A1(n4953), .A2(n7110), .ZN(n7094) );
  NAND2_X1 U5882 ( .A1(n4917), .A2(n4918), .ZN(n7256) );
  NOR2_X1 U5883 ( .A1(n4916), .A2(n6644), .ZN(n7255) );
  NAND2_X1 U5884 ( .A1(n4679), .A2(n4678), .ZN(n7331) );
  INV_X1 U5885 ( .A(n4671), .ZN(n7801) );
  INV_X1 U5886 ( .A(n4913), .ZN(n8460) );
  OR2_X1 U5887 ( .A1(n8439), .A2(n8440), .ZN(n4913) );
  INV_X1 U5888 ( .A(n8461), .ZN(n4912) );
  OAI21_X1 U5889 ( .B1(n8439), .B2(n4911), .A(n4910), .ZN(n8485) );
  NAND2_X1 U5890 ( .A1(n4914), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4911) );
  NAND2_X1 U5891 ( .A1(n8461), .A2(n4914), .ZN(n4910) );
  INV_X1 U5892 ( .A(n8462), .ZN(n4914) );
  NAND2_X1 U5893 ( .A1(n4934), .A2(n4936), .ZN(n8538) );
  OR2_X1 U5894 ( .A1(n8531), .A2(n8865), .ZN(n4907) );
  NAND2_X1 U5895 ( .A1(n8573), .A2(n8574), .ZN(n4684) );
  INV_X1 U5896 ( .A(n8572), .ZN(n4683) );
  OR2_X1 U5897 ( .A1(n8569), .A2(n8568), .ZN(n4950) );
  INV_X1 U5898 ( .A(n8583), .ZN(n4686) );
  NAND2_X1 U5899 ( .A1(n4904), .A2(n4903), .ZN(n8578) );
  OAI21_X1 U5900 ( .B1(n8619), .B2(n7739), .A(n6453), .ZN(n6454) );
  XNOR2_X1 U5901 ( .A(n6347), .B(P2_REG3_REG_26__SCAN_IN), .ZN(n8648) );
  NAND2_X1 U5902 ( .A1(n6281), .A2(n6280), .ZN(n8737) );
  NAND2_X1 U5903 ( .A1(n4778), .A2(n8066), .ZN(n8756) );
  OR2_X1 U5904 ( .A1(n10215), .A2(n7307), .ZN(n8815) );
  NAND2_X1 U5905 ( .A1(n4798), .A2(n8041), .ZN(n7833) );
  NAND2_X1 U5906 ( .A1(n6188), .A2(n6187), .ZN(n7873) );
  NAND2_X1 U5907 ( .A1(n6164), .A2(n6163), .ZN(n10212) );
  NAND2_X1 U5908 ( .A1(n4792), .A2(n8022), .ZN(n7670) );
  NAND2_X1 U5909 ( .A1(n6126), .A2(n8026), .ZN(n7562) );
  INV_X1 U5910 ( .A(n10171), .ZN(n8801) );
  INV_X1 U5911 ( .A(n7137), .ZN(n10186) );
  NAND2_X1 U5912 ( .A1(n7300), .A2(n6385), .ZN(n7425) );
  NAND2_X1 U5913 ( .A1(n8817), .A2(n10166), .ZN(n8822) );
  OR2_X1 U5914 ( .A1(n8133), .A2(n7018), .ZN(n7048) );
  NAND2_X1 U5915 ( .A1(n7013), .A2(n7581), .ZN(n10215) );
  NAND2_X1 U5916 ( .A1(n7938), .A2(n7937), .ZN(n8823) );
  AND2_X2 U5917 ( .A1(n7047), .A2(n6503), .ZN(n10233) );
  AOI21_X1 U5918 ( .B1(n8157), .B2(n6139), .A(n7926), .ZN(n8888) );
  NAND2_X1 U5919 ( .A1(n6356), .A2(n6355), .ZN(n8891) );
  AOI21_X1 U5920 ( .B1(n4888), .B2(n8813), .A(n4885), .ZN(n8889) );
  NAND2_X1 U5921 ( .A1(n4887), .A2(n4886), .ZN(n4885) );
  XNOR2_X1 U5922 ( .A(n8621), .B(n7970), .ZN(n4888) );
  NAND2_X1 U5923 ( .A1(n8645), .A2(n8808), .ZN(n4886) );
  AND2_X1 U5924 ( .A1(n8635), .A2(n8634), .ZN(n8896) );
  OR2_X1 U5925 ( .A1(n8632), .A2(n8631), .ZN(n8635) );
  NAND2_X1 U5926 ( .A1(n6337), .A2(n6336), .ZN(n8903) );
  OAI21_X1 U5927 ( .B1(n4707), .B2(n4706), .A(n8104), .ZN(n8670) );
  INV_X1 U5928 ( .A(n4782), .ZN(n4707) );
  NOR2_X1 U5929 ( .A1(n4713), .A2(n4780), .ZN(n4706) );
  NAND2_X1 U5930 ( .A1(n6318), .A2(n6317), .ZN(n8915) );
  AND2_X1 U5931 ( .A1(n4784), .A2(n4781), .ZN(n8675) );
  INV_X1 U5932 ( .A(n4785), .ZN(n4781) );
  AND2_X1 U5933 ( .A1(n8689), .A2(n8688), .ZN(n8690) );
  NAND2_X1 U5934 ( .A1(n6299), .A2(n6298), .ZN(n8927) );
  NAND2_X1 U5935 ( .A1(n6290), .A2(n6289), .ZN(n8933) );
  NAND2_X1 U5936 ( .A1(n6418), .A2(n6417), .ZN(n8730) );
  NAND2_X1 U5937 ( .A1(n6272), .A2(n6271), .ZN(n8944) );
  NAND2_X1 U5938 ( .A1(n6246), .A2(n6245), .ZN(n8955) );
  NAND2_X1 U5939 ( .A1(n6234), .A2(n6233), .ZN(n8961) );
  AND2_X1 U5940 ( .A1(n8786), .A2(n8785), .ZN(n8960) );
  NAND2_X1 U5941 ( .A1(n6222), .A2(n6221), .ZN(n8967) );
  NAND2_X1 U5942 ( .A1(n6210), .A2(n6209), .ZN(n8974) );
  NAND2_X1 U5943 ( .A1(n4853), .A2(n4856), .ZN(n8807) );
  NAND2_X1 U5944 ( .A1(n7836), .A2(n4859), .ZN(n4853) );
  NAND2_X1 U5945 ( .A1(n4861), .A2(n4859), .ZN(n7864) );
  INV_X1 U5946 ( .A(n8951), .ZN(n8973) );
  INV_X1 U5947 ( .A(n7210), .ZN(n10170) );
  INV_X2 U5948 ( .A(n10223), .ZN(n10221) );
  AND2_X1 U5949 ( .A1(n6630), .A2(n6725), .ZN(n6923) );
  NAND2_X1 U5950 ( .A1(n8982), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6017) );
  INV_X1 U5951 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7639) );
  INV_X1 U5952 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7583) );
  OAI21_X1 U5953 ( .B1(n6208), .B2(n4526), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5997) );
  INV_X1 U5954 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7283) );
  INV_X1 U5955 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7105) );
  INV_X1 U5956 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6766) );
  INV_X1 U5957 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6759) );
  XNOR2_X1 U5958 ( .A(n6129), .B(n6128), .ZN(n6758) );
  XNOR2_X1 U5959 ( .A(n6107), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7127) );
  XNOR2_X1 U5960 ( .A(n4670), .B(n6052), .ZN(n6718) );
  NAND2_X1 U5961 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n6052) );
  NAND2_X1 U5962 ( .A1(n4651), .A2(n4650), .ZN(n9061) );
  NAND2_X1 U5963 ( .A1(n4654), .A2(n4652), .ZN(n4650) );
  AOI21_X1 U5964 ( .B1(n9023), .B2(n4657), .A(n4654), .ZN(n9007) );
  AND2_X1 U5965 ( .A1(n5903), .A2(n5902), .ZN(n5965) );
  NAND2_X1 U5966 ( .A1(n5764), .A2(n5763), .ZN(n9683) );
  NAND2_X1 U5967 ( .A1(n5554), .A2(n5072), .ZN(n5068) );
  NAND2_X1 U5968 ( .A1(n9058), .A2(n5826), .ZN(n9030) );
  NAND2_X1 U5969 ( .A1(n5687), .A2(n5686), .ZN(n9045) );
  NAND2_X1 U5970 ( .A1(n9049), .A2(n9050), .ZN(n9048) );
  NAND2_X1 U5971 ( .A1(n9037), .A2(n9040), .ZN(n9049) );
  NAND2_X1 U5972 ( .A1(n5394), .A2(n5393), .ZN(n7034) );
  NAND2_X1 U5973 ( .A1(n9014), .A2(n5080), .ZN(n9074) );
  NAND2_X1 U5974 ( .A1(n4659), .A2(n4666), .ZN(n9079) );
  OR2_X1 U5975 ( .A1(n9023), .A2(n9022), .ZN(n4653) );
  INV_X1 U5976 ( .A(n9914), .ZN(n9117) );
  INV_X1 U5977 ( .A(n4644), .ZN(n4634) );
  NAND2_X1 U5978 ( .A1(n5729), .A2(n5728), .ZN(n9816) );
  NAND2_X1 U5979 ( .A1(n9030), .A2(n9031), .ZN(n9100) );
  NAND2_X1 U5980 ( .A1(n6890), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9926) );
  NAND2_X1 U5981 ( .A1(n5648), .A2(n5647), .ZN(n9121) );
  NAND2_X1 U5982 ( .A1(n5866), .A2(n5865), .ZN(n9363) );
  OR2_X1 U5983 ( .A1(n5360), .A2(n6797), .ZN(n5365) );
  OR2_X1 U5984 ( .A1(n4520), .A2(n6985), .ZN(n5303) );
  NAND2_X1 U5985 ( .A1(n4551), .A2(n10073), .ZN(n9547) );
  NAND2_X1 U5986 ( .A1(n8160), .A2(n8159), .ZN(n9554) );
  AOI21_X1 U5987 ( .B1(n6603), .B2(n9996), .A(n6602), .ZN(n9566) );
  NAND2_X1 U5988 ( .A1(n5920), .A2(n5919), .ZN(n9760) );
  NAND2_X1 U5989 ( .A1(n9568), .A2(n9572), .ZN(n9567) );
  NAND2_X1 U5990 ( .A1(n6555), .A2(n6554), .ZN(n9621) );
  NAND2_X1 U5991 ( .A1(n4984), .A2(n6545), .ZN(n9690) );
  AND2_X1 U5992 ( .A1(n9711), .A2(n9710), .ZN(n9813) );
  NAND2_X1 U5993 ( .A1(n5022), .A2(n5019), .ZN(n9709) );
  NAND2_X1 U5994 ( .A1(n4961), .A2(n4964), .ZN(n7887) );
  NAND2_X1 U5995 ( .A1(n9944), .A2(n4967), .ZN(n4961) );
  NAND2_X1 U5996 ( .A1(n4969), .A2(n4971), .ZN(n7844) );
  NAND2_X1 U5997 ( .A1(n4970), .A2(n4536), .ZN(n4969) );
  INV_X1 U5998 ( .A(n9944), .ZN(n4970) );
  NAND2_X1 U5999 ( .A1(n9940), .A2(n9177), .ZN(n7845) );
  NAND2_X1 U6000 ( .A1(n5627), .A2(n5626), .ZN(n9951) );
  NAND2_X1 U6001 ( .A1(n7658), .A2(n9312), .ZN(n7641) );
  AND2_X1 U6002 ( .A1(n7522), .A2(n9164), .ZN(n7659) );
  OR2_X1 U6003 ( .A1(n10033), .A2(n5285), .ZN(n9746) );
  INV_X1 U6004 ( .A(n9746), .ZN(n10025) );
  OR2_X1 U6005 ( .A1(n10033), .A2(n7161), .ZN(n10029) );
  AND2_X1 U6006 ( .A1(n5967), .A2(n10122), .ZN(n10019) );
  NAND2_X1 U6007 ( .A1(n5609), .A2(n5608), .ZN(n7694) );
  NAND2_X1 U6008 ( .A1(n5561), .A2(n5560), .ZN(n7614) );
  AND2_X2 U6009 ( .A1(n6614), .A2(n6620), .ZN(n10141) );
  AND2_X1 U6010 ( .A1(n9547), .A2(n9542), .ZN(n9840) );
  NAND2_X1 U6011 ( .A1(n5888), .A2(n5887), .ZN(n9849) );
  NAND2_X1 U6012 ( .A1(n5857), .A2(n5856), .ZN(n9853) );
  NAND2_X1 U6013 ( .A1(n5835), .A2(n5834), .ZN(n9857) );
  NAND2_X1 U6014 ( .A1(n5787), .A2(n5786), .ZN(n9862) );
  AND2_X1 U6015 ( .A1(n5287), .A2(n5286), .ZN(n9879) );
  AND3_X1 U6016 ( .A1(n9826), .A2(n9825), .A3(n9824), .ZN(n9885) );
  AND2_X1 U6017 ( .A1(n6619), .A2(n9897), .ZN(n10036) );
  OR2_X1 U6018 ( .A1(n6371), .A2(SI_29_), .ZN(n6372) );
  NAND2_X1 U6019 ( .A1(n5268), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5229) );
  NOR2_X1 U6020 ( .A1(n5375), .A2(n4560), .ZN(n4838) );
  NAND2_X1 U6021 ( .A1(n5242), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5243) );
  INV_X1 U6022 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n10567) );
  INV_X1 U6023 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7580) );
  INV_X1 U6024 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7559) );
  INV_X1 U6025 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10561) );
  INV_X1 U6026 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10655) );
  CLKBUF_X1 U6027 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n10534) );
  NAND2_X1 U6028 ( .A1(n7411), .A2(n7412), .ZN(n7413) );
  XNOR2_X1 U6029 ( .A(n4726), .B(n8597), .ZN(n8148) );
  NAND2_X1 U6030 ( .A1(n10155), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6934) );
  INV_X1 U6031 ( .A(n4947), .ZN(n7617) );
  INV_X1 U6032 ( .A(n4677), .ZN(n7699) );
  AOI211_X1 U6033 ( .C1(n8601), .C2(n10161), .A(n8600), .B(n8599), .ZN(n8602)
         );
  NAND2_X1 U6034 ( .A1(n4940), .A2(n4939), .ZN(P2_U3295) );
  NAND2_X1 U6035 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_STATE_REG_SCAN_IN), .ZN(
        n4939) );
  NAND2_X1 U6036 ( .A1(n8988), .A2(P2_U3151), .ZN(n4940) );
  NOR2_X1 U6037 ( .A1(n6781), .A2(P1_U3086), .ZN(P1_U3973) );
  INV_X1 U6038 ( .A(n4624), .ZN(n4623) );
  OR2_X1 U6039 ( .A1(n8989), .A2(n4629), .ZN(n4628) );
  AOI21_X1 U6040 ( .B1(n4621), .B2(n4549), .A(n9343), .ZN(n9359) );
  NOR2_X1 U6041 ( .A1(n8967), .A2(n8811), .ZN(n4522) );
  NAND2_X1 U6042 ( .A1(n6342), .A2(n6341), .ZN(n8664) );
  NAND2_X1 U6043 ( .A1(n6418), .A2(n4537), .ZN(n8717) );
  OR2_X1 U6044 ( .A1(n8915), .A2(n8305), .ZN(n8104) );
  NAND2_X1 U6045 ( .A1(n8095), .A2(n8703), .ZN(n4746) );
  AND2_X1 U6046 ( .A1(n4632), .A2(n4631), .ZN(n4523) );
  AND2_X1 U6047 ( .A1(n7660), .A2(n9164), .ZN(n4524) );
  NOR2_X1 U6048 ( .A1(n8042), .A2(n8133), .ZN(n4525) );
  NAND2_X1 U6049 ( .A1(n4765), .A2(n4763), .ZN(n4526) );
  AND2_X1 U6050 ( .A1(n8990), .A2(n8991), .ZN(n4527) );
  XNOR2_X1 U6051 ( .A(n5943), .B(n5942), .ZN(n5963) );
  NAND2_X1 U6052 ( .A1(n5098), .A2(n8328), .ZN(n8268) );
  AND2_X1 U6053 ( .A1(n9155), .A2(n9162), .ZN(n4528) );
  OAI21_X1 U6054 ( .B1(n9037), .B2(n5086), .A(n4634), .ZN(n4633) );
  INV_X1 U6055 ( .A(n9037), .ZN(n4643) );
  INV_X1 U6056 ( .A(n9162), .ZN(n4821) );
  INV_X1 U6057 ( .A(n5040), .ZN(n5034) );
  NOR2_X1 U6058 ( .A1(n5204), .A2(n10419), .ZN(n5040) );
  OR2_X1 U6059 ( .A1(n4585), .A2(n5078), .ZN(n4529) );
  AND2_X1 U6060 ( .A1(n4901), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4530) );
  INV_X1 U6061 ( .A(n9145), .ZN(n4612) );
  INV_X1 U6062 ( .A(n8420), .ZN(n6055) );
  INV_X1 U6063 ( .A(n8570), .ZN(n4949) );
  AND2_X1 U6064 ( .A1(n4949), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4531) );
  XNOR2_X2 U6065 ( .A(n6035), .B(n6034), .ZN(n6036) );
  NAND2_X2 U6066 ( .A1(n5275), .A2(n5276), .ZN(n5360) );
  OR2_X1 U6067 ( .A1(n5151), .A2(n5400), .ZN(n4532) );
  OR3_X1 U6068 ( .A1(n7651), .A2(n9121), .A3(n4929), .ZN(n4533) );
  OR4_X1 U6069 ( .A1(n9195), .A2(n9222), .A3(n9327), .A4(n9328), .ZN(n4534) );
  OR2_X1 U6070 ( .A1(n7797), .A2(n7796), .ZN(n4535) );
  NAND2_X1 U6071 ( .A1(n6627), .A2(n6714), .ZN(n6066) );
  NAND2_X1 U6072 ( .A1(n6564), .A2(n6563), .ZN(n9560) );
  NAND2_X1 U6073 ( .A1(n9951), .A2(n9374), .ZN(n4536) );
  AND2_X1 U6074 ( .A1(n4852), .A2(n6417), .ZN(n4537) );
  INV_X1 U6075 ( .A(n4646), .ZN(n4645) );
  XNOR2_X1 U6076 ( .A(n5322), .B(n5779), .ZN(n4538) );
  AND2_X1 U6077 ( .A1(n5315), .A2(n5316), .ZN(n4539) );
  NAND2_X1 U6078 ( .A1(n6627), .A2(n7931), .ZN(n6065) );
  XNOR2_X1 U6079 ( .A(n8891), .B(n8633), .ZN(n8622) );
  NAND2_X1 U6080 ( .A1(n8123), .A2(n7940), .ZN(n8121) );
  NOR2_X1 U6081 ( .A1(n8823), .A2(n7976), .ZN(n8130) );
  AND2_X1 U6082 ( .A1(n8740), .A2(n8085), .ZN(n8686) );
  INV_X1 U6083 ( .A(n9125), .ZN(n4802) );
  XOR2_X1 U6084 ( .A(n5153), .B(SI_6_), .Z(n4540) );
  INV_X1 U6085 ( .A(n9031), .ZN(n5063) );
  AND4_X1 U6086 ( .A1(n5234), .A2(n5223), .A3(n5222), .A4(n5221), .ZN(n4541)
         );
  INV_X1 U6087 ( .A(n8026), .ZN(n4794) );
  AND2_X1 U6088 ( .A1(n9648), .A2(n6590), .ZN(n4542) );
  OAI211_X1 U6089 ( .C1(n6627), .C2(n6036), .A(n6039), .B(n6038), .ZN(n7306)
         );
  OR2_X1 U6090 ( .A1(n9260), .A2(n9222), .ZN(n4543) );
  AND2_X1 U6091 ( .A1(n4759), .A2(n4757), .ZN(n4544) );
  OR2_X1 U6092 ( .A1(n10212), .A2(n8411), .ZN(n4545) );
  AND2_X1 U6093 ( .A1(n4996), .A2(n4999), .ZN(n4546) );
  AND2_X1 U6094 ( .A1(n5107), .A2(n5106), .ZN(n4547) );
  AND2_X1 U6095 ( .A1(n5397), .A2(n5439), .ZN(n4548) );
  AND2_X1 U6096 ( .A1(n5052), .A2(n5050), .ZN(n4549) );
  NAND2_X1 U6097 ( .A1(n8040), .A2(n8039), .ZN(n4550) );
  INV_X1 U6098 ( .A(n9572), .ZN(n4999) );
  AND2_X1 U6099 ( .A1(n9282), .A2(n9216), .ZN(n9572) );
  INV_X1 U6100 ( .A(n8047), .ZN(n4774) );
  XOR2_X1 U6101 ( .A(n9545), .B(n9548), .Z(n4551) );
  INV_X1 U6102 ( .A(n4884), .ZN(n4883) );
  NAND2_X1 U6103 ( .A1(n7774), .A2(n8412), .ZN(n4552) );
  INV_X1 U6104 ( .A(n6406), .ZN(n4862) );
  OR2_X1 U6105 ( .A1(n8052), .A2(n8050), .ZN(n4553) );
  AND2_X1 U6106 ( .A1(n9121), .A2(n9373), .ZN(n4554) );
  INV_X1 U6107 ( .A(n9245), .ZN(n7891) );
  AND2_X1 U6108 ( .A1(n9181), .A2(n9296), .ZN(n9245) );
  OR2_X1 U6109 ( .A1(n5165), .A2(n5530), .ZN(n4555) );
  AND2_X1 U6110 ( .A1(n4631), .A2(n5077), .ZN(n4556) );
  INV_X1 U6111 ( .A(n4665), .ZN(n4664) );
  NAND2_X1 U6112 ( .A1(n4538), .A2(n4667), .ZN(n4665) );
  NOR2_X1 U6113 ( .A1(n8974), .A2(n8794), .ZN(n4557) );
  NOR2_X1 U6114 ( .A1(n10096), .A2(n9379), .ZN(n4558) );
  INV_X1 U6115 ( .A(n8740), .ZN(n4713) );
  OR2_X1 U6116 ( .A1(n9199), .A2(n9222), .ZN(n4559) );
  OAI21_X1 U6117 ( .B1(n5743), .B2(n5036), .A(n5035), .ZN(n5041) );
  INV_X1 U6118 ( .A(n9172), .ZN(n9177) );
  AND2_X1 U6119 ( .A1(n9951), .A2(n7847), .ZN(n9172) );
  NAND2_X1 U6120 ( .A1(n5227), .A2(n5024), .ZN(n4560) );
  NAND3_X1 U6121 ( .A1(n4573), .A2(n4647), .A3(n5424), .ZN(n4561) );
  AND2_X1 U6122 ( .A1(n5178), .A2(SI_13_), .ZN(n4562) );
  AND2_X1 U6123 ( .A1(n5176), .A2(SI_12_), .ZN(n4563) );
  AND2_X1 U6124 ( .A1(n7891), .A2(n4962), .ZN(n4564) );
  INV_X1 U6125 ( .A(n4791), .ZN(n4790) );
  NAND2_X1 U6126 ( .A1(n4795), .A2(n8022), .ZN(n4791) );
  NAND2_X1 U6127 ( .A1(n4653), .A2(n4664), .ZN(n4565) );
  AND2_X1 U6128 ( .A1(n4766), .A2(n4553), .ZN(n4566) );
  AND2_X1 U6129 ( .A1(n9862), .A2(n9366), .ZN(n4567) );
  NOR2_X1 U6130 ( .A1(n9321), .A2(n9173), .ZN(n4568) );
  NAND2_X1 U6131 ( .A1(n9296), .A2(n9178), .ZN(n4569) );
  NOR2_X1 U6132 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6632) );
  AND2_X1 U6133 ( .A1(n9853), .A2(n9363), .ZN(n4570) );
  OR2_X1 U6134 ( .A1(n8909), .A2(n8385), .ZN(n8108) );
  INV_X1 U6135 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5253) );
  INV_X1 U6136 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6003) );
  OR2_X1 U6137 ( .A1(n8933), .A2(n8733), .ZN(n8094) );
  INV_X1 U6138 ( .A(n5020), .ZN(n5019) );
  NAND2_X1 U6139 ( .A1(n5021), .A2(n9192), .ZN(n5020) );
  INV_X1 U6140 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6011) );
  OR2_X1 U6141 ( .A1(n9275), .A2(n9347), .ZN(n4571) );
  AND3_X1 U6142 ( .A1(n9208), .A2(n9583), .A3(n9620), .ZN(n4572) );
  OR2_X1 U6143 ( .A1(n8961), .A2(n8769), .ZN(n8069) );
  INV_X1 U6144 ( .A(n8069), .ZN(n4736) );
  NOR2_X1 U6145 ( .A1(n5236), .A2(n5235), .ZN(n4573) );
  NAND2_X1 U6146 ( .A1(n8686), .A2(n8699), .ZN(n4574) );
  NAND2_X1 U6147 ( .A1(n5232), .A2(n5231), .ZN(n9669) );
  AND2_X1 U6148 ( .A1(n4532), .A2(n4540), .ZN(n4575) );
  INV_X1 U6149 ( .A(n7266), .ZN(n6741) );
  AND2_X1 U6150 ( .A1(n6127), .A2(n6115), .ZN(n7266) );
  NAND2_X1 U6151 ( .A1(n8714), .A2(n8093), .ZN(n4703) );
  AND2_X1 U6152 ( .A1(n4642), .A2(n4641), .ZN(n4576) );
  AND2_X1 U6153 ( .A1(n7924), .A2(n5033), .ZN(n4577) );
  AND2_X1 U6154 ( .A1(n5166), .A2(n5156), .ZN(n4578) );
  AND2_X1 U6155 ( .A1(n4657), .A2(n4652), .ZN(n4579) );
  AND2_X1 U6156 ( .A1(n4907), .A2(n4906), .ZN(n4580) );
  AND2_X1 U6157 ( .A1(n4938), .A2(n4937), .ZN(n4581) );
  AND2_X1 U6158 ( .A1(n5250), .A2(n5249), .ZN(n4582) );
  INV_X1 U6159 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5233) );
  INV_X1 U6160 ( .A(n4880), .ZN(n4879) );
  OAI21_X1 U6161 ( .B1(n6396), .B2(n4881), .A(n6395), .ZN(n4880) );
  INV_X1 U6162 ( .A(n4746), .ZN(n4745) );
  INV_X1 U6163 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5989) );
  INV_X1 U6164 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5024) );
  INV_X1 U6165 ( .A(n5496), .ZN(n5921) );
  INV_X1 U6166 ( .A(n6716), .ZN(n4895) );
  NAND2_X1 U6167 ( .A1(n5251), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5708) );
  INV_X1 U6168 ( .A(n8411), .ZN(n7820) );
  INV_X1 U6169 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n4763) );
  XOR2_X1 U6170 ( .A(n5738), .B(n5898), .Z(n4583) );
  AND2_X1 U6171 ( .A1(n4723), .A2(n5034), .ZN(n4584) );
  NAND2_X1 U6172 ( .A1(n4610), .A2(n8145), .ZN(n8133) );
  INV_X1 U6173 ( .A(n9312), .ZN(n5008) );
  INV_X1 U6174 ( .A(n9296), .ZN(n4831) );
  INV_X1 U6175 ( .A(n9717), .ZN(n5021) );
  NAND2_X1 U6176 ( .A1(n7904), .A2(n7903), .ZN(n8168) );
  NAND2_X1 U6177 ( .A1(n5066), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5726) );
  AND2_X1 U6178 ( .A1(n9072), .A2(n9071), .ZN(n4585) );
  AND2_X1 U6179 ( .A1(n8169), .A2(n8809), .ZN(n4586) );
  NAND2_X1 U6180 ( .A1(n5093), .A2(n5092), .ZN(n8257) );
  NAND2_X1 U6181 ( .A1(n8180), .A2(n8179), .ZN(n8319) );
  AND2_X1 U6182 ( .A1(n9940), .A2(n5011), .ZN(n4587) );
  AND2_X1 U6183 ( .A1(n4642), .A2(n4645), .ZN(n4588) );
  NAND2_X1 U6184 ( .A1(n9728), .A2(n4922), .ZN(n4926) );
  AND2_X1 U6185 ( .A1(n5761), .A2(n10602), .ZN(n4589) );
  INV_X1 U6186 ( .A(n5082), .ZN(n5081) );
  NOR2_X1 U6187 ( .A1(n5086), .A2(n4583), .ZN(n5082) );
  AND2_X1 U6188 ( .A1(n4913), .A2(n4912), .ZN(n4590) );
  NAND2_X1 U6189 ( .A1(n6366), .A2(n6365), .ZN(n8633) );
  OR2_X1 U6190 ( .A1(n6208), .A2(n5996), .ZN(n4591) );
  AND2_X1 U6191 ( .A1(n4584), .A2(n4716), .ZN(n4592) );
  INV_X1 U6192 ( .A(n9050), .ZN(n5086) );
  INV_X1 U6193 ( .A(n5039), .ZN(n5038) );
  NAND2_X1 U6194 ( .A1(n5204), .A2(n10419), .ZN(n5039) );
  AND2_X1 U6195 ( .A1(n9683), .A2(n9368), .ZN(n4593) );
  NOR2_X1 U6196 ( .A1(n5761), .A2(n10602), .ZN(n4594) );
  NAND2_X1 U6197 ( .A1(n6313), .A2(n6312), .ZN(n8706) );
  AND2_X1 U6198 ( .A1(n8232), .A2(n8231), .ZN(n4595) );
  NAND2_X1 U6199 ( .A1(n6758), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4596) );
  NAND2_X1 U6200 ( .A1(n5260), .A2(n5292), .ZN(n5294) );
  NOR2_X1 U6201 ( .A1(n7229), .A2(n10081), .ZN(n4920) );
  INV_X1 U6202 ( .A(n7015), .ZN(n7013) );
  NAND2_X1 U6203 ( .A1(n4958), .A2(n6525), .ZN(n7393) );
  XNOR2_X1 U6204 ( .A(n5243), .B(P1_IR_REG_24__SCAN_IN), .ZN(n5939) );
  OR2_X1 U6205 ( .A1(n7651), .A2(n4929), .ZN(n4597) );
  INV_X1 U6206 ( .A(n4859), .ZN(n4858) );
  NOR2_X1 U6207 ( .A1(n7961), .A2(n4860), .ZN(n4859) );
  NAND2_X1 U6208 ( .A1(n7034), .A2(n4548), .ZN(n7214) );
  INV_X1 U6209 ( .A(n4967), .ZN(n4966) );
  NOR2_X1 U6210 ( .A1(n6537), .A2(n4968), .ZN(n4967) );
  AND2_X1 U6211 ( .A1(n4898), .A2(n6647), .ZN(n4598) );
  NAND2_X1 U6212 ( .A1(n5702), .A2(n5703), .ZN(n4599) );
  NAND2_X1 U6213 ( .A1(n4844), .A2(n4848), .ZN(n4600) );
  OR2_X1 U6214 ( .A1(n8523), .A2(n8797), .ZN(n4601) );
  NAND2_X1 U6215 ( .A1(n5968), .A2(n9699), .ZN(n9924) );
  INV_X1 U6216 ( .A(n9919), .ZN(n9097) );
  NAND2_X1 U6217 ( .A1(n4982), .A2(n5471), .ZN(n9962) );
  INV_X1 U6218 ( .A(n9962), .ZN(n4919) );
  INV_X1 U6219 ( .A(n7020), .ZN(n7318) );
  OAI211_X1 U6220 ( .C1(n6627), .C2(n6718), .A(n6054), .B(n6053), .ZN(n7020)
         );
  NAND2_X1 U6221 ( .A1(n5583), .A2(n5582), .ZN(n10108) );
  INV_X1 U6222 ( .A(n10108), .ZN(n4932) );
  OR2_X1 U6223 ( .A1(n8527), .A2(n8787), .ZN(n4602) );
  INV_X1 U6224 ( .A(n4725), .ZN(n7423) );
  NAND2_X1 U6225 ( .A1(n7307), .A2(n4610), .ZN(n4725) );
  AND2_X1 U6226 ( .A1(n6643), .A2(n6741), .ZN(n6644) );
  INV_X1 U6227 ( .A(n6644), .ZN(n4917) );
  OR2_X1 U6228 ( .A1(n8551), .A2(n8865), .ZN(n4603) );
  OR2_X1 U6229 ( .A1(n7928), .A2(SI_30_), .ZN(n4604) );
  AND2_X1 U6230 ( .A1(n4681), .A2(n6701), .ZN(n4605) );
  NAND2_X1 U6231 ( .A1(n6436), .A2(n5998), .ZN(n8141) );
  INV_X1 U6232 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n4616) );
  INV_X1 U6233 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5043) );
  XNOR2_X1 U6234 ( .A(n8459), .B(n8473), .ZN(n8439) );
  NAND2_X1 U6235 ( .A1(n4607), .A2(n4572), .ZN(n9209) );
  OAI21_X1 U6236 ( .B1(n9206), .B2(n9205), .A(n9631), .ZN(n4607) );
  AOI21_X1 U6237 ( .B1(n9176), .B2(n9316), .A(n4608), .ZN(n9180) );
  NOR2_X1 U6238 ( .A1(n9146), .A2(n4611), .ZN(n9156) );
  NAND2_X1 U6239 ( .A1(n9974), .A2(n9300), .ZN(n9131) );
  NAND2_X1 U6240 ( .A1(n6571), .A2(n9298), .ZN(n6569) );
  NAND2_X1 U6241 ( .A1(n4808), .A2(n9258), .ZN(n4807) );
  NAND2_X1 U6242 ( .A1(n4813), .A2(n4559), .ZN(n4812) );
  NAND2_X1 U6243 ( .A1(n8269), .A2(n8328), .ZN(n8223) );
  NAND2_X1 U6244 ( .A1(n5097), .A2(n5098), .ZN(n8269) );
  NAND2_X1 U6245 ( .A1(n7822), .A2(n7821), .ZN(n5088) );
  NAND2_X1 U6246 ( .A1(n7017), .A2(n7016), .ZN(n7019) );
  NAND2_X1 U6247 ( .A1(n8218), .A2(n8217), .ZN(n8328) );
  NOR2_X1 U6248 ( .A1(n6079), .A2(n5990), .ZN(n6160) );
  INV_X1 U6249 ( .A(n6195), .ZN(n5993) );
  NAND2_X1 U6250 ( .A1(n6544), .A2(n5115), .ZN(n4984) );
  OAI21_X2 U6251 ( .B1(n9944), .B2(n4963), .A(n4564), .ZN(n6539) );
  OAI21_X2 U6252 ( .B1(n4958), .B2(n4957), .A(n4955), .ZN(n7349) );
  OAI22_X2 U6253 ( .A1(n9738), .A2(n6540), .B1(n9371), .B2(n9743), .ZN(n9721)
         );
  NAND2_X2 U6254 ( .A1(n6553), .A2(n5117), .ZN(n6555) );
  AND2_X1 U6255 ( .A1(n9180), .A2(n4829), .ZN(n4824) );
  NAND2_X1 U6256 ( .A1(n4807), .A2(n9214), .ZN(n4806) );
  NAND2_X1 U6257 ( .A1(n4812), .A2(n9662), .ZN(n4811) );
  NAND2_X1 U6258 ( .A1(n6549), .A2(n5127), .ZN(n6551) );
  NAND4_X1 U6259 ( .A1(n9143), .A2(n9144), .A3(n9142), .A4(n4612), .ZN(n4611)
         );
  NAND2_X2 U6260 ( .A1(n6536), .A2(n6535), .ZN(n9944) );
  OAI21_X1 U6261 ( .B1(n9197), .B2(n4814), .A(n4543), .ZN(n4813) );
  NAND2_X1 U6262 ( .A1(n4613), .A2(n8101), .ZN(n8105) );
  NAND2_X1 U6263 ( .A1(n4738), .A2(n4740), .ZN(n4613) );
  INV_X1 U6264 ( .A(n4614), .ZN(n6319) );
  NAND2_X1 U6265 ( .A1(n4614), .A2(n10413), .ZN(n6329) );
  NOR2_X1 U6266 ( .A1(n4691), .A2(n7975), .ZN(n4690) );
  NAND2_X1 U6267 ( .A1(n4727), .A2(n4689), .ZN(n4726) );
  INV_X1 U6268 ( .A(n4742), .ZN(n4739) );
  NAND2_X1 U6269 ( .A1(n4684), .A2(n4683), .ZN(n4682) );
  INV_X1 U6270 ( .A(n8097), .ZN(n4744) );
  NAND2_X1 U6271 ( .A1(n9209), .A2(n4571), .ZN(n4808) );
  AOI21_X1 U6272 ( .B1(n4811), .B2(n4810), .A(n4809), .ZN(n9206) );
  NAND2_X1 U6273 ( .A1(n4806), .A2(n4805), .ZN(n4804) );
  NAND2_X1 U6274 ( .A1(n4804), .A2(n4803), .ZN(n9218) );
  NAND2_X1 U6275 ( .A1(n9293), .A2(n5964), .ZN(n4621) );
  OAI211_X1 U6276 ( .C1(n4817), .C2(n4818), .A(n4815), .B(n4820), .ZN(n9166)
         );
  NAND2_X1 U6277 ( .A1(n9967), .A2(n9968), .ZN(n4958) );
  INV_X1 U6278 ( .A(n9661), .ZN(n6549) );
  OAI21_X1 U6279 ( .B1(n6555), .B2(n4974), .A(n4972), .ZN(n4980) );
  NAND3_X1 U6280 ( .A1(n5304), .A2(n5305), .A3(n5898), .ZN(n5308) );
  NAND3_X1 U6281 ( .A1(n5304), .A2(n5305), .A3(n5118), .ZN(n6983) );
  NAND3_X1 U6282 ( .A1(n4628), .A2(n4627), .A3(n4623), .ZN(P1_U3214) );
  NAND2_X1 U6283 ( .A1(n8992), .A2(n9097), .ZN(n4627) );
  NOR2_X1 U6284 ( .A1(n5083), .A2(n4583), .ZN(n4646) );
  AND2_X2 U6285 ( .A1(n5423), .A2(n5220), .ZN(n5624) );
  NAND2_X1 U6286 ( .A1(n9023), .A2(n4579), .ZN(n4651) );
  OR2_X2 U6287 ( .A1(n6063), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n6079) );
  NAND3_X1 U6288 ( .A1(n6034), .A2(n4670), .A3(n4669), .ZN(n6063) );
  INV_X2 U6289 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U6290 ( .A1(n6706), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7798) );
  NAND2_X1 U6291 ( .A1(n4671), .A2(n7799), .ZN(n4673) );
  INV_X1 U6292 ( .A(n4673), .ZN(n8446) );
  INV_X1 U6293 ( .A(n4681), .ZN(n7261) );
  OAI21_X1 U6294 ( .B1(n4950), .B2(n4949), .A(n4686), .ZN(n4685) );
  INV_X1 U6295 ( .A(n8539), .ZN(n4688) );
  NAND2_X1 U6296 ( .A1(n5557), .A2(n4697), .ZN(n4695) );
  NOR2_X1 U6297 ( .A1(n4705), .A2(n4704), .ZN(n8642) );
  INV_X1 U6298 ( .A(n8108), .ZN(n4712) );
  OAI21_X1 U6299 ( .B1(n5707), .B2(n4717), .A(n4715), .ZN(n4714) );
  NAND3_X1 U6300 ( .A1(n7985), .A2(n7988), .A3(n4610), .ZN(n7983) );
  NAND2_X1 U6301 ( .A1(n4729), .A2(n4728), .ZN(n4727) );
  NOR2_X1 U6302 ( .A1(n8138), .A2(n7014), .ZN(n4728) );
  NAND2_X1 U6303 ( .A1(n8140), .A2(n8139), .ZN(n4729) );
  NAND4_X1 U6304 ( .A1(n4732), .A2(n4731), .A3(n4730), .A4(n6111), .ZN(n5990)
         );
  NAND2_X1 U6305 ( .A1(n4734), .A2(n4733), .ZN(n8076) );
  INV_X1 U6306 ( .A(n8067), .ZN(n4733) );
  OAI21_X1 U6307 ( .B1(n4735), .B2(n8133), .A(n8766), .ZN(n4734) );
  NAND2_X1 U6308 ( .A1(n8091), .A2(n8090), .ZN(n4737) );
  NAND2_X1 U6309 ( .A1(n8116), .A2(n8115), .ZN(n4760) );
  INV_X1 U6310 ( .A(n8122), .ZN(n4757) );
  INV_X1 U6311 ( .A(n8121), .ZN(n4758) );
  NAND2_X1 U6312 ( .A1(n4778), .A2(n4776), .ZN(n8860) );
  NAND2_X1 U6313 ( .A1(n6242), .A2(n8069), .ZN(n8763) );
  INV_X1 U6314 ( .A(n7955), .ZN(n4795) );
  NAND3_X1 U6315 ( .A1(n7296), .A2(n7988), .A3(n7982), .ZN(n7297) );
  AND2_X2 U6316 ( .A1(n7989), .A2(n6056), .ZN(n7988) );
  NAND2_X1 U6317 ( .A1(n4798), .A2(n4797), .ZN(n7835) );
  NAND2_X1 U6318 ( .A1(n6013), .A2(n5112), .ZN(n6018) );
  INV_X2 U6319 ( .A(n6458), .ZN(n6013) );
  NAND2_X1 U6320 ( .A1(n6013), .A2(n4800), .ZN(n8982) );
  OAI21_X1 U6321 ( .B1(n9156), .B2(n9155), .A(n9154), .ZN(n9160) );
  NAND3_X1 U6322 ( .A1(n9156), .A2(n9154), .A3(n4816), .ZN(n4815) );
  NOR2_X1 U6323 ( .A1(n4817), .A2(n4821), .ZN(n4816) );
  NOR3_X2 U6324 ( .A1(n4825), .A2(n4824), .A3(n4822), .ZN(n9193) );
  AND2_X1 U6325 ( .A1(n9174), .A2(n4827), .ZN(n4825) );
  AND2_X1 U6326 ( .A1(n5225), .A2(n4839), .ZN(n4835) );
  NOR2_X2 U6327 ( .A1(n5375), .A2(n5215), .ZN(n5423) );
  NAND4_X1 U6328 ( .A1(n4838), .A2(n5220), .A3(n4836), .A4(n4541), .ZN(n5268)
         );
  NAND3_X1 U6329 ( .A1(n4841), .A2(n4840), .A3(n4847), .ZN(n6458) );
  NOR2_X1 U6330 ( .A1(n4842), .A2(n6006), .ZN(n4840) );
  NOR2_X1 U6331 ( .A1(n6079), .A2(n6007), .ZN(n4841) );
  NOR2_X1 U6332 ( .A1(n6080), .A2(n6007), .ZN(n4848) );
  NAND2_X1 U6333 ( .A1(n4848), .A2(n4845), .ZN(n6010) );
  NOR2_X1 U6334 ( .A1(n5990), .A2(n6006), .ZN(n4845) );
  OAI21_X2 U6335 ( .B1(n6418), .B2(n4851), .A(n4849), .ZN(n8722) );
  OAI21_X1 U6336 ( .B1(n7836), .B2(n4855), .A(n4854), .ZN(n6408) );
  NAND2_X1 U6337 ( .A1(n4867), .A2(n4865), .ZN(n7205) );
  NAND3_X1 U6338 ( .A1(n6383), .A2(n6386), .A3(n6382), .ZN(n4867) );
  NAND2_X1 U6339 ( .A1(n6383), .A2(n6382), .ZN(n7300) );
  NAND3_X1 U6340 ( .A1(n6401), .A2(n6400), .A3(n4870), .ZN(n4869) );
  NAND2_X1 U6341 ( .A1(n6392), .A2(n6393), .ZN(n7462) );
  NAND2_X1 U6342 ( .A1(n4875), .A2(n4877), .ZN(n6397) );
  NAND3_X1 U6343 ( .A1(n6392), .A2(n6393), .A3(n4879), .ZN(n4875) );
  NOR2_X1 U6344 ( .A1(n7466), .A2(n8415), .ZN(n4884) );
  NAND2_X1 U6345 ( .A1(n8773), .A2(n6412), .ZN(n8751) );
  NAND2_X1 U6346 ( .A1(n6405), .A2(n6404), .ZN(n7836) );
  AOI21_X1 U6347 ( .B1(n10184), .B2(n6457), .A(n8611), .ZN(n6504) );
  OAI21_X1 U6348 ( .B1(n9220), .B2(n9254), .A(n9219), .ZN(n9223) );
  NAND2_X1 U6349 ( .A1(n8764), .A2(n8065), .ZN(n8773) );
  NAND2_X1 U6350 ( .A1(n8722), .A2(n8702), .ZN(n8652) );
  INV_X1 U6351 ( .A(n8792), .ZN(n6410) );
  NAND2_X1 U6352 ( .A1(n6570), .A2(n7002), .ZN(n10011) );
  MUX2_X2 U6353 ( .A(n9223), .B(n9222), .S(n9554), .Z(n9224) );
  NAND2_X1 U6354 ( .A1(n4893), .A2(n6956), .ZN(n4891) );
  NAND2_X1 U6355 ( .A1(n6649), .A2(n4901), .ZN(n4897) );
  NAND2_X1 U6356 ( .A1(n4899), .A2(n4897), .ZN(n7707) );
  NAND3_X1 U6357 ( .A1(n4900), .A2(n6647), .A3(n4530), .ZN(n4899) );
  INV_X1 U6358 ( .A(n4907), .ZN(n8549) );
  INV_X1 U6359 ( .A(n8550), .ZN(n4906) );
  NAND3_X1 U6360 ( .A1(n4909), .A2(P2_REG1_REG_5__SCAN_IN), .A3(n7116), .ZN(
        n7118) );
  NAND2_X1 U6361 ( .A1(n4908), .A2(n6659), .ZN(n7092) );
  NAND2_X1 U6362 ( .A1(n7120), .A2(n6642), .ZN(n6643) );
  INV_X1 U6363 ( .A(n4926), .ZN(n9682) );
  MUX2_X1 U6364 ( .A(n10534), .B(n9910), .S(n6783), .Z(n10020) );
  NAND2_X2 U6365 ( .A1(n9399), .A2(n9930), .ZN(n6783) );
  NAND3_X1 U6366 ( .A1(n5624), .A2(n5024), .A3(n5226), .ZN(n4933) );
  INV_X1 U6367 ( .A(n4938), .ZN(n8520) );
  INV_X1 U6368 ( .A(n8521), .ZN(n4937) );
  NAND2_X1 U6369 ( .A1(n6700), .A2(n6741), .ZN(n6701) );
  NAND2_X1 U6370 ( .A1(n4954), .A2(n5309), .ZN(n5137) );
  XNOR2_X1 U6371 ( .A(n5309), .B(n4954), .ZN(n6730) );
  NAND2_X1 U6372 ( .A1(n4960), .A2(n4575), .ZN(n5155) );
  XNOR2_X1 U6373 ( .A(n4959), .B(n4540), .ZN(n6736) );
  INV_X1 U6374 ( .A(n4980), .ZN(n9592) );
  OR2_X1 U6375 ( .A1(n9857), .A2(n9364), .ZN(n4981) );
  OAI21_X2 U6376 ( .B1(n9681), .B2(n4593), .A(n6548), .ZN(n9661) );
  NAND2_X1 U6377 ( .A1(n4984), .A2(n4983), .ZN(n6547) );
  OAI21_X2 U6378 ( .B1(n9654), .B2(n4567), .A(n6552), .ZN(n9630) );
  INV_X1 U6379 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4988) );
  INV_X1 U6380 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4987) );
  INV_X1 U6381 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4986) );
  NAND3_X1 U6382 ( .A1(n4988), .A2(n4987), .A3(n4986), .ZN(n4985) );
  NAND3_X1 U6383 ( .A1(n5130), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4989) );
  NAND2_X1 U6384 ( .A1(n9386), .A2(n5900), .ZN(n5307) );
  NAND3_X1 U6385 ( .A1(n5124), .A2(n5303), .A3(n5302), .ZN(n9386) );
  NAND2_X1 U6386 ( .A1(n9586), .A2(n4993), .ZN(n4990) );
  OAI211_X1 U6387 ( .C1(n9586), .C2(n4995), .A(n4991), .B(n4990), .ZN(n6603)
         );
  NAND2_X1 U6388 ( .A1(n6588), .A2(n5001), .ZN(n5000) );
  OAI21_X1 U6389 ( .B1(n9941), .B2(n5010), .A(n5009), .ZN(n7890) );
  NAND2_X1 U6390 ( .A1(n9722), .A2(n5016), .ZN(n5012) );
  NAND2_X1 U6391 ( .A1(n5012), .A2(n5014), .ZN(n6585) );
  NAND3_X1 U6392 ( .A1(n5227), .A2(n5024), .A3(n5228), .ZN(n5023) );
  NAND2_X1 U6393 ( .A1(n5804), .A2(n5029), .ZN(n5025) );
  NAND2_X1 U6394 ( .A1(n5025), .A2(n5026), .ZN(n5850) );
  XNOR2_X1 U6395 ( .A(n7923), .B(n7921), .ZN(n6371) );
  NAND2_X1 U6396 ( .A1(n7925), .A2(n4577), .ZN(n5032) );
  NAND2_X1 U6397 ( .A1(n5032), .A2(n4604), .ZN(n7935) );
  NAND2_X1 U6398 ( .A1(n7925), .A2(n7924), .ZN(n7930) );
  INV_X1 U6399 ( .A(n5041), .ZN(n5210) );
  OAI21_X1 U6400 ( .B1(n4507), .B2(n5043), .A(n5042), .ZN(n5135) );
  MUX2_X1 U6401 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n7931), .Z(n5139) );
  AOI21_X1 U6402 ( .B1(n5422), .B2(n4578), .A(n5044), .ZN(n5169) );
  NOR2_X1 U6403 ( .A1(n9339), .A2(n5284), .ZN(n5051) );
  NAND2_X1 U6404 ( .A1(n5053), .A2(n5284), .ZN(n5052) );
  AOI21_X1 U6405 ( .B1(n9290), .B2(n9355), .A(n9289), .ZN(n5054) );
  NAND2_X1 U6406 ( .A1(n5623), .A2(n5179), .ZN(n5056) );
  NAND2_X1 U6407 ( .A1(n5056), .A2(n5055), .ZN(n5184) );
  NAND2_X1 U6408 ( .A1(n5708), .A2(n5067), .ZN(n5065) );
  NAND2_X1 U6409 ( .A1(n7537), .A2(n5070), .ZN(n5069) );
  NAND3_X1 U6410 ( .A1(n5069), .A2(n5068), .A3(n9917), .ZN(n5601) );
  NAND2_X1 U6411 ( .A1(n7571), .A2(n7572), .ZN(n9918) );
  NAND2_X1 U6412 ( .A1(n5074), .A2(n7536), .ZN(n7571) );
  OR2_X1 U6413 ( .A1(n5739), .A2(n5740), .ZN(n5080) );
  NAND2_X1 U6414 ( .A1(n7214), .A2(n7216), .ZN(n7191) );
  NAND2_X1 U6415 ( .A1(n5646), .A2(n4582), .ZN(n5251) );
  NAND2_X1 U6416 ( .A1(n5646), .A2(n5249), .ZN(n5684) );
  INV_X1 U6417 ( .A(n5091), .ZN(n5090) );
  NAND2_X1 U6418 ( .A1(n7874), .A2(n5094), .ZN(n5093) );
  NAND2_X1 U6419 ( .A1(n8208), .A2(n8207), .ZN(n5098) );
  NAND2_X1 U6420 ( .A1(n8320), .A2(n8366), .ZN(n8185) );
  NAND2_X1 U6421 ( .A1(n8180), .A2(n5099), .ZN(n8320) );
  NAND2_X1 U6422 ( .A1(n8258), .A2(n5101), .ZN(n8396) );
  NAND2_X1 U6423 ( .A1(n8380), .A2(n4595), .ZN(n8248) );
  NAND2_X2 U6424 ( .A1(n8229), .A2(n8377), .ZN(n8380) );
  INV_X1 U6425 ( .A(n5110), .ZN(n7549) );
  NAND2_X1 U6426 ( .A1(n6013), .A2(n6012), .ZN(n6467) );
  NAND2_X1 U6427 ( .A1(n6582), .A2(n9245), .ZN(n7888) );
  INV_X1 U6428 ( .A(n7890), .ZN(n6582) );
  CLKBUF_X1 U6429 ( .A(n6569), .Z(n10014) );
  XNOR2_X1 U6430 ( .A(n6566), .B(n9254), .ZN(n9564) );
  NAND2_X2 U6431 ( .A1(n6567), .A2(n5293), .ZN(n5322) );
  INV_X1 U6432 ( .A(n5346), .ZN(n5496) );
  OAI22_X1 U6433 ( .A1(n7861), .A2(n6207), .B1(n7917), .B2(n8809), .ZN(n8805)
         );
  NAND2_X1 U6434 ( .A1(n6431), .A2(n6430), .ZN(n8644) );
  NAND2_X1 U6435 ( .A1(n6032), .A2(n6019), .ZN(n6020) );
  NAND2_X1 U6436 ( .A1(n5512), .A2(n5467), .ZN(n7444) );
  NAND2_X1 U6437 ( .A1(n8210), .A2(n8209), .ZN(n8216) );
  OR2_X1 U6438 ( .A1(n9721), .A2(n6541), .ZN(n6543) );
  NAND2_X1 U6439 ( .A1(n8396), .A2(n8177), .ZN(n8313) );
  XNOR2_X1 U6440 ( .A(n7020), .B(n7169), .ZN(n7058) );
  NAND2_X2 U6441 ( .A1(n7019), .A2(n7018), .ZN(n7169) );
  OAI21_X2 U6442 ( .B1(n9061), .B2(n9060), .A(n9059), .ZN(n9058) );
  NAND2_X1 U6443 ( .A1(n8783), .A2(n8782), .ZN(n8781) );
  NAND2_X4 U6444 ( .A1(n4505), .A2(n6024), .ZN(n7471) );
  INV_X1 U6445 ( .A(n10174), .ZN(n8636) );
  OR2_X1 U6446 ( .A1(n9879), .A2(n9092), .ZN(n5115) );
  OR2_X1 U6447 ( .A1(n9698), .A2(n9024), .ZN(n5116) );
  AND2_X2 U6448 ( .A1(n7151), .A2(n9699), .ZN(n10033) );
  INV_X1 U6449 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6199) );
  OR2_X1 U6450 ( .A1(n9782), .A2(n9365), .ZN(n5117) );
  INV_X1 U6451 ( .A(n9782), .ZN(n6604) );
  OR2_X1 U6452 ( .A1(n5292), .A2(n9929), .ZN(n5118) );
  OR2_X1 U6453 ( .A1(n5182), .A2(n10564), .ZN(n5119) );
  NOR2_X1 U6454 ( .A1(n8212), .A2(n8340), .ZN(n5120) );
  OR2_X1 U6455 ( .A1(n8234), .A2(n8386), .ZN(n5121) );
  OR2_X1 U6456 ( .A1(n6506), .A2(n8864), .ZN(n5122) );
  OR2_X1 U6457 ( .A1(n6506), .A2(n8951), .ZN(n5123) );
  INV_X1 U6458 ( .A(SI_12_), .ZN(n5175) );
  INV_X1 U6459 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5143) );
  AND2_X1 U6460 ( .A1(n5301), .A2(n5300), .ZN(n5124) );
  INV_X1 U6461 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6150) );
  NOR2_X1 U6462 ( .A1(n8909), .A2(n8679), .ZN(n5125) );
  INV_X1 U6463 ( .A(n8706), .ZN(n8219) );
  INV_X1 U6464 ( .A(n9837), .ZN(n6616) );
  NAND2_X1 U6465 ( .A1(n10125), .A2(n10095), .ZN(n9894) );
  INV_X1 U6466 ( .A(n9894), .ZN(n6623) );
  AND3_X1 U6467 ( .A1(n5966), .A2(n9097), .A3(n5965), .ZN(n5126) );
  OR2_X1 U6468 ( .A1(n9669), .A2(n9367), .ZN(n5127) );
  AND2_X1 U6469 ( .A1(n5939), .A2(n5959), .ZN(n5128) );
  INV_X1 U6470 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5224) );
  OR2_X1 U6471 ( .A1(n8169), .A2(n8809), .ZN(n8167) );
  NOR2_X1 U6472 ( .A1(n5120), .A2(n8214), .ZN(n8215) );
  NOR2_X1 U6473 ( .A1(n8482), .A2(n6213), .ZN(n8493) );
  INV_X1 U6474 ( .A(SI_21_), .ZN(n10602) );
  INV_X1 U6475 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5170) );
  NAND2_X1 U6476 ( .A1(n8216), .A2(n8215), .ZN(n8218) );
  INV_X1 U6477 ( .A(n8135), .ZN(n8139) );
  INV_X1 U6478 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10388) );
  OR2_X1 U6479 ( .A1(n8933), .A2(n8707), .ZN(n8702) );
  INV_X1 U6480 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5992) );
  INV_X1 U6481 ( .A(n5731), .ZN(n5263) );
  INV_X1 U6482 ( .A(n9554), .ZN(n8161) );
  INV_X1 U6483 ( .A(n5790), .ZN(n5788) );
  INV_X1 U6484 ( .A(n5747), .ZN(n5264) );
  INV_X1 U6485 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n10335) );
  INV_X1 U6486 ( .A(n5643), .ZN(n5182) );
  INV_X1 U6487 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6692) );
  AND3_X1 U6488 ( .A1(n7041), .A2(n7040), .A3(n6495), .ZN(n6911) );
  NAND2_X1 U6489 ( .A1(n5858), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5924) );
  OR3_X1 U6490 ( .A1(n5837), .A2(n9065), .A3(n5836), .ZN(n5860) );
  NAND2_X1 U6491 ( .A1(n8162), .A2(n8161), .ZN(n9548) );
  INV_X1 U6492 ( .A(n9636), .ZN(n9655) );
  NAND2_X1 U6493 ( .A1(n5265), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5790) );
  NAND2_X1 U6494 ( .A1(n5264), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5765) );
  OR2_X1 U6495 ( .A1(n5498), .A2(n5497), .ZN(n5542) );
  NAND2_X1 U6496 ( .A1(n9636), .A2(n6604), .ZN(n9638) );
  OAI21_X1 U6497 ( .B1(n7351), .B2(n7350), .A(n9163), .ZN(n7524) );
  OR2_X1 U6498 ( .A1(n7923), .A2(n7922), .ZN(n7924) );
  NAND2_X1 U6499 ( .A1(n5171), .A2(n10461), .ZN(n5174) );
  INV_X1 U6500 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5131) );
  AND2_X1 U6501 ( .A1(n8350), .A2(n8197), .ZN(n8290) );
  AND2_X1 U6502 ( .A1(n8289), .A2(n8191), .ZN(n8341) );
  XNOR2_X1 U6503 ( .A(n7058), .B(n8420), .ZN(n7062) );
  INV_X1 U6504 ( .A(n8337), .ZN(n8398) );
  AND2_X1 U6505 ( .A1(n6288), .A2(n6287), .ZN(n8282) );
  NAND2_X1 U6506 ( .A1(n8427), .A2(n8428), .ZN(n8426) );
  INV_X1 U6507 ( .A(n6454), .ZN(n6455) );
  AND2_X1 U6508 ( .A1(n8057), .A2(n8056), .ZN(n8806) );
  INV_X1 U6509 ( .A(n6388), .ZN(n7993) );
  INV_X1 U6510 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n6016) );
  AND2_X1 U6511 ( .A1(n5562), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5584) );
  INV_X1 U6512 ( .A(n7033), .ZN(n5393) );
  OR2_X1 U6513 ( .A1(n5975), .A2(n5962), .ZN(n9914) );
  INV_X1 U6514 ( .A(n4520), .ZN(n5889) );
  INV_X1 U6515 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6818) );
  OR3_X1 U6516 ( .A1(n7496), .A2(n7494), .A3(n7493), .ZN(n7601) );
  OR3_X1 U6517 ( .A1(n7758), .A2(n7756), .A3(n7755), .ZN(n9526) );
  INV_X1 U6518 ( .A(n9252), .ZN(n9591) );
  OAI21_X1 U6519 ( .B1(n9616), .B2(n9211), .A(n9207), .ZN(n9600) );
  INV_X1 U6520 ( .A(n9250), .ZN(n9653) );
  INV_X1 U6521 ( .A(n9182), .ZN(n9748) );
  INV_X1 U6522 ( .A(n9103), .ZN(n9091) );
  AND2_X1 U6523 ( .A1(n6782), .A2(n9399), .ZN(n9103) );
  INV_X1 U6524 ( .A(n10003), .ZN(n10073) );
  INV_X1 U6525 ( .A(n9996), .ZN(n10016) );
  OR2_X1 U6526 ( .A1(n6524), .A2(n9151), .ZN(n9968) );
  AND2_X1 U6527 ( .A1(n5851), .A2(n5833), .ZN(n5849) );
  XNOR2_X1 U6528 ( .A(n5176), .B(n5175), .ZN(n5577) );
  NAND2_X1 U6529 ( .A1(n5488), .A2(n5487), .ZN(n5489) );
  AOI22_X1 U6530 ( .A1(n7273), .A2(n7272), .B1(n7271), .B2(n7270), .ZN(n7275)
         );
  NAND2_X1 U6531 ( .A1(n6925), .A2(n10169), .ZN(n8324) );
  AOI21_X1 U6532 ( .B1(n8710), .B2(n6360), .A(n6304), .ZN(n8294) );
  OR2_X1 U6533 ( .A1(n6363), .A2(n8448), .ZN(n6203) );
  NAND2_X1 U6534 ( .A1(n6071), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6027) );
  INV_X1 U6535 ( .A(n8598), .ZN(n10155) );
  INV_X1 U6536 ( .A(n8593), .ZN(n10146) );
  AND2_X1 U6537 ( .A1(n8039), .A2(n8036), .ZN(n7957) );
  INV_X1 U6538 ( .A(n10169), .ZN(n8800) );
  INV_X1 U6539 ( .A(n8636), .ZN(n8817) );
  INV_X1 U6540 ( .A(n8864), .ZN(n8875) );
  OR2_X1 U6541 ( .A1(n4522), .A2(n7963), .ZN(n8793) );
  INV_X1 U6542 ( .A(n10215), .ZN(n10213) );
  AND2_X1 U6543 ( .A1(n6629), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6725) );
  XNOR2_X1 U6544 ( .A(n6008), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8145) );
  INV_X1 U6545 ( .A(n5984), .ZN(n5985) );
  INV_X1 U6546 ( .A(n9926), .ZN(n9105) );
  OR2_X1 U6547 ( .A1(n9575), .A2(n4521), .ZN(n5933) );
  INV_X1 U6548 ( .A(n9528), .ZN(n9531) );
  INV_X1 U6549 ( .A(n9534), .ZN(n9507) );
  INV_X1 U6550 ( .A(n9503), .ZN(n9530) );
  NAND2_X1 U6551 ( .A1(n9953), .A2(n7154), .ZN(n10006) );
  INV_X1 U6552 ( .A(n10029), .ZN(n9950) );
  AND2_X1 U6553 ( .A1(n5947), .A2(n9897), .ZN(n6614) );
  NAND2_X1 U6554 ( .A1(n10084), .A2(n10009), .ZN(n10112) );
  INV_X1 U6555 ( .A(n10038), .ZN(n9897) );
  INV_X1 U6556 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5228) );
  INV_X1 U6557 ( .A(n8389), .ZN(n8399) );
  AND2_X1 U6558 ( .A1(n6921), .A2(n6920), .ZN(n8393) );
  NAND4_X1 U6559 ( .A1(n6206), .A2(n6205), .A3(n6204), .A4(n6203), .ZN(n8809)
         );
  INV_X1 U6560 ( .A(P2_U3893), .ZN(n8561) );
  INV_X1 U6561 ( .A(n10161), .ZN(n8571) );
  NAND2_X1 U6562 ( .A1(n7053), .A2(n10169), .ZN(n10174) );
  OR2_X1 U6563 ( .A1(n7053), .A2(n8815), .ZN(n10171) );
  NAND2_X1 U6564 ( .A1(n10233), .A2(n10196), .ZN(n8878) );
  INV_X1 U6565 ( .A(n10233), .ZN(n10231) );
  XOR2_X1 U6566 ( .A(n8691), .B(n8690), .Z(n8924) );
  OR2_X1 U6567 ( .A1(n10223), .A2(n10215), .ZN(n8951) );
  OR2_X1 U6568 ( .A1(n10223), .A2(n10217), .ZN(n8977) );
  AND2_X1 U6569 ( .A1(n6491), .A2(n6490), .ZN(n10223) );
  INV_X1 U6570 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7558) );
  INV_X1 U6571 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6833) );
  NOR2_X1 U6572 ( .A1(n5126), .A2(n5985), .ZN(n5986) );
  INV_X1 U6573 ( .A(n7694), .ZN(n7730) );
  OR2_X1 U6574 ( .A1(n5975), .A2(n5977), .ZN(n9919) );
  NAND2_X1 U6575 ( .A1(n5933), .A2(n5932), .ZN(n9362) );
  OR2_X1 U6576 ( .A1(n9939), .A2(n9397), .ZN(n9503) );
  OR2_X1 U6577 ( .A1(n9939), .A2(n6810), .ZN(n9528) );
  INV_X1 U6578 ( .A(n10006), .ZN(n9737) );
  NAND2_X1 U6579 ( .A1(n10141), .A2(n10095), .ZN(n9837) );
  INV_X1 U6580 ( .A(n10141), .ZN(n10139) );
  INV_X1 U6581 ( .A(n9669), .ZN(n9867) );
  INV_X1 U6582 ( .A(n10125), .ZN(n10123) );
  AND2_X2 U6583 ( .A1(n6620), .A2(n10036), .ZN(n10125) );
  INV_X1 U6584 ( .A(n10035), .ZN(n10034) );
  AND2_X1 U6585 ( .A1(n9897), .A2(n9896), .ZN(n10035) );
  INV_X1 U6586 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10588) );
  INV_X1 U6587 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10661) );
  INV_X1 U6588 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6768) );
  CLKBUF_X1 U6589 ( .A(n9906), .Z(n8152) );
  INV_X1 U6590 ( .A(SI_1_), .ZN(n5132) );
  AND2_X1 U6591 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5133) );
  NAND2_X1 U6592 ( .A1(n5911), .A2(n5133), .ZN(n5298) );
  AND2_X1 U6593 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5134) );
  NAND2_X1 U6594 ( .A1(n7931), .A2(n5134), .ZN(n6046) );
  NAND2_X1 U6595 ( .A1(n5135), .A2(SI_1_), .ZN(n5136) );
  NAND2_X1 U6596 ( .A1(n5137), .A2(n5136), .ZN(n5337) );
  INV_X1 U6597 ( .A(SI_2_), .ZN(n5138) );
  XNOR2_X1 U6598 ( .A(n5139), .B(n5138), .ZN(n5336) );
  NAND2_X1 U6599 ( .A1(n5337), .A2(n5336), .ZN(n5141) );
  NAND2_X1 U6600 ( .A1(n5139), .A2(SI_2_), .ZN(n5140) );
  NAND2_X1 U6601 ( .A1(n5141), .A2(n5140), .ZN(n5354) );
  INV_X1 U6602 ( .A(SI_3_), .ZN(n5144) );
  XNOR2_X1 U6603 ( .A(n5145), .B(n5144), .ZN(n5353) );
  NAND2_X1 U6604 ( .A1(n5354), .A2(n5353), .ZN(n5147) );
  NAND2_X1 U6605 ( .A1(n5145), .A2(SI_3_), .ZN(n5146) );
  MUX2_X1 U6606 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n6714), .Z(n5148) );
  INV_X1 U6607 ( .A(SI_4_), .ZN(n10587) );
  XNOR2_X1 U6608 ( .A(n5148), .B(n10587), .ZN(n5376) );
  NAND2_X1 U6609 ( .A1(n5148), .A2(SI_4_), .ZN(n5398) );
  MUX2_X1 U6610 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n5911), .Z(n5150) );
  NAND2_X1 U6611 ( .A1(n5150), .A2(SI_5_), .ZN(n5149) );
  AND2_X1 U6612 ( .A1(n5398), .A2(n5149), .ZN(n5152) );
  INV_X1 U6613 ( .A(n5149), .ZN(n5151) );
  INV_X1 U6614 ( .A(SI_5_), .ZN(n10421) );
  XNOR2_X1 U6615 ( .A(n5150), .B(n10421), .ZN(n5400) );
  MUX2_X1 U6616 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6714), .Z(n5153) );
  NAND2_X1 U6617 ( .A1(n5153), .A2(SI_6_), .ZN(n5154) );
  MUX2_X1 U6618 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6714), .Z(n5157) );
  XNOR2_X1 U6619 ( .A(n5157), .B(SI_7_), .ZN(n5421) );
  INV_X1 U6620 ( .A(n5421), .ZN(n5156) );
  NAND2_X1 U6621 ( .A1(n5157), .A2(SI_7_), .ZN(n5158) );
  MUX2_X1 U6622 ( .A(n6759), .B(n10655), .S(n6714), .Z(n5159) );
  NAND2_X1 U6623 ( .A1(n5159), .A2(n10617), .ZN(n5483) );
  INV_X1 U6624 ( .A(n5159), .ZN(n5160) );
  NAND2_X1 U6625 ( .A1(n5160), .A2(SI_8_), .ZN(n5161) );
  NAND2_X1 U6626 ( .A1(n5483), .A2(n5161), .ZN(n5468) );
  MUX2_X1 U6627 ( .A(n6766), .B(n6768), .S(n6714), .Z(n5163) );
  INV_X1 U6628 ( .A(SI_9_), .ZN(n5162) );
  NAND2_X1 U6629 ( .A1(n5163), .A2(n5162), .ZN(n5484) );
  AND2_X1 U6630 ( .A1(n5483), .A2(n5484), .ZN(n5528) );
  MUX2_X1 U6631 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n6714), .Z(n5167) );
  INV_X1 U6632 ( .A(n5532), .ZN(n5165) );
  INV_X1 U6633 ( .A(n5163), .ZN(n5164) );
  NAND2_X1 U6634 ( .A1(n5164), .A2(SI_9_), .ZN(n5530) );
  NAND2_X1 U6635 ( .A1(n5167), .A2(SI_10_), .ZN(n5168) );
  NAND2_X1 U6636 ( .A1(n5169), .A2(n5168), .ZN(n5557) );
  MUX2_X1 U6637 ( .A(n6833), .B(n5170), .S(n5911), .Z(n5171) );
  INV_X1 U6638 ( .A(n5171), .ZN(n5172) );
  NAND2_X1 U6639 ( .A1(n5172), .A2(SI_11_), .ZN(n5173) );
  NAND2_X1 U6640 ( .A1(n5174), .A2(n5173), .ZN(n5556) );
  MUX2_X1 U6641 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6714), .Z(n5176) );
  MUX2_X1 U6642 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6714), .Z(n5178) );
  XNOR2_X1 U6643 ( .A(n5178), .B(SI_13_), .ZN(n5602) );
  MUX2_X1 U6644 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6714), .Z(n5180) );
  XNOR2_X1 U6645 ( .A(n5180), .B(SI_14_), .ZN(n5622) );
  INV_X1 U6646 ( .A(n5622), .ZN(n5179) );
  NAND2_X1 U6647 ( .A1(n5180), .A2(SI_14_), .ZN(n5181) );
  MUX2_X1 U6648 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n5911), .Z(n5643) );
  NAND2_X1 U6649 ( .A1(n5182), .A2(n10564), .ZN(n5183) );
  NAND2_X1 U6650 ( .A1(n5184), .A2(n5183), .ZN(n5683) );
  MUX2_X1 U6651 ( .A(n7105), .B(n5185), .S(n6714), .Z(n5681) );
  NOR2_X1 U6652 ( .A1(n5187), .A2(SI_16_), .ZN(n5186) );
  NAND2_X1 U6653 ( .A1(n5187), .A2(SI_16_), .ZN(n5188) );
  INV_X1 U6654 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n5190) );
  MUX2_X1 U6655 ( .A(n5190), .B(n10561), .S(n6714), .Z(n5192) );
  INV_X1 U6656 ( .A(SI_17_), .ZN(n5191) );
  NAND2_X1 U6657 ( .A1(n5192), .A2(n5191), .ZN(n5195) );
  INV_X1 U6658 ( .A(n5192), .ZN(n5193) );
  NAND2_X1 U6659 ( .A1(n5193), .A2(SI_17_), .ZN(n5194) );
  NAND2_X1 U6660 ( .A1(n5195), .A2(n5194), .ZN(n5706) );
  MUX2_X1 U6661 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6714), .Z(n5197) );
  XNOR2_X1 U6662 ( .A(n5197), .B(n10423), .ZN(n5724) );
  INV_X1 U6663 ( .A(n5724), .ZN(n5196) );
  NAND2_X1 U6664 ( .A1(n5197), .A2(SI_18_), .ZN(n5198) );
  MUX2_X1 U6665 ( .A(n7283), .B(n10661), .S(n6714), .Z(n5200) );
  INV_X1 U6666 ( .A(SI_19_), .ZN(n5199) );
  NAND2_X1 U6667 ( .A1(n5200), .A2(n5199), .ZN(n5203) );
  INV_X1 U6668 ( .A(n5200), .ZN(n5201) );
  NAND2_X1 U6669 ( .A1(n5201), .A2(SI_19_), .ZN(n5202) );
  NAND2_X1 U6670 ( .A1(n5203), .A2(n5202), .ZN(n5282) );
  MUX2_X1 U6671 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n6714), .Z(n5741) );
  INV_X1 U6672 ( .A(n5741), .ZN(n5204) );
  MUX2_X1 U6673 ( .A(n7558), .B(n7559), .S(n6714), .Z(n5761) );
  MUX2_X1 U6674 ( .A(n7583), .B(n7580), .S(n6714), .Z(n5206) );
  INV_X1 U6675 ( .A(SI_22_), .ZN(n5205) );
  NAND2_X1 U6676 ( .A1(n5206), .A2(n5205), .ZN(n5780) );
  INV_X1 U6677 ( .A(n5206), .ZN(n5207) );
  NAND2_X1 U6678 ( .A1(n5207), .A2(SI_22_), .ZN(n5208) );
  NAND2_X1 U6679 ( .A1(n5780), .A2(n5208), .ZN(n5211) );
  INV_X1 U6680 ( .A(n5211), .ZN(n5209) );
  NAND2_X1 U6681 ( .A1(n5210), .A2(n5209), .ZN(n5781) );
  NAND2_X1 U6682 ( .A1(n5041), .A2(n5211), .ZN(n5212) );
  NAND2_X1 U6683 ( .A1(n5781), .A2(n5212), .ZN(n7579) );
  NOR2_X4 U6684 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5339) );
  INV_X2 U6685 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5402) );
  NAND2_X1 U6686 ( .A1(n5214), .A2(n5402), .ZN(n5215) );
  NOR2_X1 U6687 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5219) );
  NOR2_X1 U6688 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5218) );
  NOR2_X1 U6689 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5217) );
  NOR2_X1 U6690 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5216) );
  NOR2_X1 U6691 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n5223) );
  NOR2_X1 U6692 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5222) );
  NOR2_X1 U6693 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5221) );
  INV_X2 U6694 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5252) );
  NAND2_X1 U6695 ( .A1(n5685), .A2(n5252), .ZN(n5235) );
  INV_X1 U6696 ( .A(n5235), .ZN(n5225) );
  XNOR2_X2 U6697 ( .A(n5229), .B(n5228), .ZN(n9399) );
  INV_X2 U6698 ( .A(n6562), .ZN(n5441) );
  NAND2_X1 U6699 ( .A1(n7579), .A2(n5441), .ZN(n5232) );
  NAND2_X1 U6700 ( .A1(n8158), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5231) );
  NAND2_X1 U6701 ( .A1(n5234), .A2(n5253), .ZN(n5236) );
  INV_X1 U6702 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5237) );
  AND3_X1 U6703 ( .A1(n5942), .A2(n10335), .A3(n5945), .ZN(n5238) );
  OAI21_X1 U6704 ( .B1(n5242), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5239) );
  MUX2_X1 U6705 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5239), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n5241) );
  INV_X1 U6706 ( .A(n7770), .ZN(n5245) );
  NAND2_X1 U6707 ( .A1(n5240), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5244) );
  NAND2_X1 U6708 ( .A1(n5245), .A2(n5128), .ZN(n5292) );
  NAND2_X1 U6709 ( .A1(n4561), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5247) );
  NAND2_X1 U6710 ( .A1(n5964), .A2(n9292), .ZN(n5976) );
  INV_X1 U6711 ( .A(n5976), .ZN(n7152) );
  AND2_X2 U6712 ( .A1(n5292), .A2(n7152), .ZN(n5319) );
  INV_X2 U6713 ( .A(n5319), .ZN(n5389) );
  NAND2_X1 U6714 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), 
        .ZN(n5249) );
  INV_X1 U6715 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5250) );
  NAND2_X1 U6716 ( .A1(n5284), .A2(n9292), .ZN(n5962) );
  NAND2_X1 U6717 ( .A1(n5962), .A2(n5976), .ZN(n5258) );
  NAND2_X1 U6718 ( .A1(n5256), .A2(n10335), .ZN(n5257) );
  NAND2_X2 U6719 ( .A1(n5284), .A2(n9351), .ZN(n6567) );
  NAND2_X1 U6720 ( .A1(n5258), .A2(n6567), .ZN(n5260) );
  INV_X1 U6721 ( .A(n5292), .ZN(n5259) );
  INV_X2 U6722 ( .A(n5294), .ZN(n5900) );
  NAND2_X1 U6723 ( .A1(n5472), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5498) );
  INV_X1 U6724 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5628) );
  INV_X1 U6725 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n7590) );
  INV_X1 U6726 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9018) );
  INV_X1 U6727 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9025) );
  INV_X1 U6728 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5266) );
  NAND2_X1 U6729 ( .A1(n5767), .A2(n5266), .ZN(n5267) );
  NAND2_X1 U6730 ( .A1(n5790), .A2(n5267), .ZN(n9671) );
  NAND2_X1 U6731 ( .A1(n5271), .A2(n5272), .ZN(n9900) );
  XNOR2_X2 U6732 ( .A(n5270), .B(n5269), .ZN(n5275) );
  OR2_X1 U6733 ( .A1(n9671), .A2(n4520), .ZN(n5281) );
  INV_X1 U6734 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9670) );
  INV_X4 U6735 ( .A(n5691), .ZN(n6899) );
  NAND2_X1 U6736 ( .A1(n5928), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5278) );
  AND2_X2 U6737 ( .A1(n5275), .A2(n9909), .ZN(n5380) );
  NAND2_X1 U6738 ( .A1(n5792), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5277) );
  OAI211_X1 U6739 ( .C1(n9670), .C2(n6899), .A(n5278), .B(n5277), .ZN(n5279)
         );
  INV_X1 U6740 ( .A(n5279), .ZN(n5280) );
  NAND2_X1 U6741 ( .A1(n5281), .A2(n5280), .ZN(n9367) );
  AOI22_X1 U6742 ( .A1(n9669), .A2(n5319), .B1(n5900), .B2(n9367), .ZN(n9080)
         );
  XNOR2_X1 U6743 ( .A(n5283), .B(n5282), .ZN(n7282) );
  NAND2_X1 U6744 ( .A1(n7282), .A2(n5441), .ZN(n5287) );
  INV_X1 U6745 ( .A(n5284), .ZN(n5285) );
  AOI22_X1 U6746 ( .A1(n5285), .A2(n5727), .B1(n8158), .B2(
        P2_DATAO_REG_19__SCAN_IN), .ZN(n5286) );
  NAND2_X1 U6747 ( .A1(n5733), .A2(n9018), .ZN(n5288) );
  AND2_X1 U6748 ( .A1(n5747), .A2(n5288), .ZN(n9713) );
  INV_X1 U6749 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9522) );
  NAND2_X1 U6750 ( .A1(n5928), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5290) );
  NAND2_X1 U6751 ( .A1(n5792), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5289) );
  OAI211_X1 U6752 ( .C1(n9522), .C2(n6899), .A(n5290), .B(n5289), .ZN(n5291)
         );
  AOI21_X1 U6753 ( .B1(n9713), .B2(n5889), .A(n5291), .ZN(n9092) );
  OAI22_X1 U6754 ( .A1(n9879), .A2(n5389), .B1(n9092), .B2(n5294), .ZN(n5740)
         );
  OAI22_X1 U6755 ( .A1(n9879), .A2(n5496), .B1(n9092), .B2(n5389), .ZN(n5295)
         );
  XNOR2_X1 U6756 ( .A(n5295), .B(n5322), .ZN(n5739) );
  INV_X1 U6757 ( .A(SI_0_), .ZN(n5297) );
  INV_X1 U6758 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5296) );
  OAI21_X1 U6759 ( .B1(n7931), .B2(n5297), .A(n5296), .ZN(n5299) );
  AND2_X1 U6760 ( .A1(n5299), .A2(n5298), .ZN(n9910) );
  NAND2_X1 U6761 ( .A1(n5346), .A2(n10020), .ZN(n5305) );
  NAND2_X1 U6762 ( .A1(n5380), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5301) );
  INV_X1 U6763 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7330) );
  INV_X1 U6764 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6985) );
  INV_X1 U6765 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9929) );
  OR2_X1 U6766 ( .A1(n5360), .A2(n9929), .ZN(n5302) );
  AOI22_X1 U6767 ( .A1(n5319), .A2(n10020), .B1(n5259), .B2(n10534), .ZN(n5306) );
  NAND2_X1 U6768 ( .A1(n5307), .A2(n5306), .ZN(n6982) );
  NAND2_X1 U6769 ( .A1(n6983), .A2(n6982), .ZN(n6981) );
  NAND2_X1 U6770 ( .A1(n6981), .A2(n5308), .ZN(n6994) );
  NAND2_X1 U6771 ( .A1(n5355), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5313) );
  NAND2_X1 U6772 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n10534), .ZN(n5310) );
  MUX2_X1 U6773 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5310), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n5312) );
  INV_X1 U6774 ( .A(n5339), .ZN(n5311) );
  NAND2_X1 U6775 ( .A1(n5312), .A2(n5311), .ZN(n6795) );
  NAND2_X1 U6776 ( .A1(n5346), .A2(n10021), .ZN(n5321) );
  INV_X1 U6777 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6997) );
  INV_X1 U6778 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6794) );
  INV_X1 U6779 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5314) );
  NAND2_X1 U6780 ( .A1(n5380), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5315) );
  NAND2_X1 U6781 ( .A1(n6984), .A2(n5319), .ZN(n5320) );
  NAND2_X1 U6782 ( .A1(n5321), .A2(n5320), .ZN(n5323) );
  XNOR2_X1 U6783 ( .A(n5323), .B(n5898), .ZN(n5325) );
  INV_X1 U6784 ( .A(n10021), .ZN(n10041) );
  NOR2_X1 U6785 ( .A1(n10041), .A2(n5389), .ZN(n5324) );
  NAND2_X1 U6786 ( .A1(n5325), .A2(n5326), .ZN(n6991) );
  NAND2_X1 U6787 ( .A1(n6994), .A2(n6991), .ZN(n5329) );
  INV_X1 U6788 ( .A(n5325), .ZN(n5328) );
  INV_X1 U6789 ( .A(n5326), .ZN(n5327) );
  NAND2_X1 U6790 ( .A1(n5328), .A2(n5327), .ZN(n6992) );
  NAND2_X1 U6791 ( .A1(n5329), .A2(n6992), .ZN(n6888) );
  NAND2_X1 U6792 ( .A1(n5380), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5332) );
  INV_X1 U6793 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5330) );
  AND2_X1 U6794 ( .A1(n5332), .A2(n5331), .ZN(n5335) );
  INV_X1 U6795 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9405) );
  INV_X1 U6796 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6793) );
  OR2_X1 U6797 ( .A1(n5360), .A2(n6793), .ZN(n5333) );
  XNOR2_X1 U6798 ( .A(n5337), .B(n5336), .ZN(n6732) );
  NAND2_X1 U6799 ( .A1(n5355), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5344) );
  INV_X1 U6800 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9899) );
  NOR2_X1 U6801 ( .A1(n5339), .A2(n9899), .ZN(n5338) );
  MUX2_X1 U6802 ( .A(n9899), .B(n5338), .S(P1_IR_REG_2__SCAN_IN), .Z(n5342) );
  INV_X1 U6803 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5340) );
  NAND2_X1 U6804 ( .A1(n5339), .A2(n5340), .ZN(n5356) );
  INV_X1 U6805 ( .A(n5356), .ZN(n5341) );
  NOR2_X1 U6806 ( .A1(n5342), .A2(n5341), .ZN(n6796) );
  NAND2_X1 U6807 ( .A1(n5727), .A2(n6796), .ZN(n5343) );
  NOR2_X1 U6808 ( .A1(n10050), .A2(n5389), .ZN(n5345) );
  AOI21_X1 U6809 ( .B1(n5900), .B2(n4512), .A(n5345), .ZN(n5350) );
  NAND2_X1 U6810 ( .A1(n4512), .A2(n5319), .ZN(n5348) );
  NAND2_X1 U6811 ( .A1(n5346), .A2(n10005), .ZN(n5347) );
  NAND2_X1 U6812 ( .A1(n5348), .A2(n5347), .ZN(n5349) );
  XNOR2_X1 U6813 ( .A(n5350), .B(n5351), .ZN(n6889) );
  NAND2_X1 U6814 ( .A1(n5351), .A2(n5350), .ZN(n5352) );
  OAI21_X1 U6815 ( .B1(n6888), .B2(n6889), .A(n5352), .ZN(n7007) );
  XNOR2_X1 U6816 ( .A(n5354), .B(n5353), .ZN(n6717) );
  NAND2_X1 U6817 ( .A1(n8158), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5359) );
  NAND2_X1 U6818 ( .A1(n5356), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5357) );
  XNOR2_X1 U6819 ( .A(n5357), .B(P1_IR_REG_3__SCAN_IN), .ZN(n9426) );
  NAND2_X1 U6820 ( .A1(n5727), .A2(n9426), .ZN(n5358) );
  INV_X1 U6821 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6797) );
  INV_X1 U6822 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6775) );
  OR2_X1 U6823 ( .A1(n5361), .A2(n6775), .ZN(n5364) );
  NAND2_X1 U6824 ( .A1(n5380), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5363) );
  OR2_X1 U6825 ( .A1(n4521), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5362) );
  NAND2_X1 U6826 ( .A1(n9384), .A2(n5319), .ZN(n5366) );
  NAND2_X1 U6827 ( .A1(n5367), .A2(n5366), .ZN(n5368) );
  XNOR2_X1 U6828 ( .A(n5368), .B(n5322), .ZN(n5370) );
  INV_X1 U6829 ( .A(n7290), .ZN(n10055) );
  NOR2_X1 U6830 ( .A1(n10055), .A2(n5389), .ZN(n5369) );
  AOI21_X1 U6831 ( .B1(n5900), .B2(n9384), .A(n5369), .ZN(n5371) );
  XNOR2_X1 U6832 ( .A(n5370), .B(n5371), .ZN(n7008) );
  NAND2_X1 U6833 ( .A1(n7007), .A2(n7008), .ZN(n5374) );
  INV_X1 U6834 ( .A(n5370), .ZN(n5372) );
  NAND2_X1 U6835 ( .A1(n5372), .A2(n5371), .ZN(n5373) );
  NAND2_X1 U6836 ( .A1(n5374), .A2(n5373), .ZN(n7032) );
  INV_X1 U6837 ( .A(n7032), .ZN(n5394) );
  NAND2_X1 U6838 ( .A1(n5375), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5403) );
  XNOR2_X1 U6839 ( .A(n5403), .B(n5402), .ZN(n9437) );
  XNOR2_X1 U6840 ( .A(n5377), .B(n5376), .ZN(n6720) );
  OR2_X1 U6841 ( .A1(n6720), .A2(n6562), .ZN(n5379) );
  NAND2_X1 U6842 ( .A1(n5355), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5378) );
  OAI211_X1 U6843 ( .C1(n6783), .C2(n9437), .A(n5379), .B(n5378), .ZN(n9983)
         );
  NAND2_X1 U6844 ( .A1(n5921), .A2(n9983), .ZN(n5391) );
  NAND2_X1 U6845 ( .A1(n5928), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5388) );
  INV_X1 U6846 ( .A(n5380), .ZN(n5653) );
  INV_X1 U6847 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5381) );
  OR2_X1 U6848 ( .A1(n5653), .A2(n5381), .ZN(n5387) );
  INV_X1 U6849 ( .A(n5382), .ZN(n5409) );
  INV_X1 U6850 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7291) );
  INV_X1 U6851 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5383) );
  NAND2_X1 U6852 ( .A1(n7291), .A2(n5383), .ZN(n5384) );
  NAND2_X1 U6853 ( .A1(n5409), .A2(n5384), .ZN(n9977) );
  OR2_X1 U6854 ( .A1(n4521), .A2(n9977), .ZN(n5386) );
  INV_X1 U6855 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6777) );
  OR2_X1 U6856 ( .A1(n6899), .A2(n6777), .ZN(n5385) );
  NAND4_X1 U6857 ( .A1(n5388), .A2(n5387), .A3(n5386), .A4(n5385), .ZN(n6895)
         );
  NAND2_X1 U6858 ( .A1(n6895), .A2(n5754), .ZN(n5390) );
  NAND2_X1 U6859 ( .A1(n5391), .A2(n5390), .ZN(n5392) );
  XNOR2_X1 U6860 ( .A(n5392), .B(n5898), .ZN(n5396) );
  AOI22_X1 U6861 ( .A1(n5900), .A2(n6895), .B1(n5319), .B2(n9983), .ZN(n5395)
         );
  XNOR2_X1 U6862 ( .A(n5396), .B(n5395), .ZN(n7033) );
  OR2_X1 U6863 ( .A1(n5396), .A2(n5395), .ZN(n5397) );
  NAND2_X1 U6864 ( .A1(n5399), .A2(n5398), .ZN(n5401) );
  XNOR2_X1 U6865 ( .A(n5401), .B(n5400), .ZN(n6723) );
  OR2_X1 U6866 ( .A1(n6723), .A2(n6562), .ZN(n5407) );
  NAND2_X1 U6867 ( .A1(n5403), .A2(n5402), .ZN(n5404) );
  NAND2_X1 U6868 ( .A1(n5404), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5405) );
  XNOR2_X1 U6869 ( .A(n5405), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9454) );
  AOI22_X1 U6870 ( .A1(n8158), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n5727), .B2(
        n9454), .ZN(n5406) );
  NAND2_X1 U6871 ( .A1(n5921), .A2(n10067), .ZN(n5417) );
  NAND2_X1 U6872 ( .A1(n5928), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5415) );
  INV_X1 U6873 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5408) );
  OR2_X1 U6874 ( .A1(n5653), .A2(n5408), .ZN(n5414) );
  INV_X1 U6875 ( .A(n5447), .ZN(n5411) );
  INV_X1 U6876 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9446) );
  NAND2_X1 U6877 ( .A1(n5409), .A2(n9446), .ZN(n5410) );
  NAND2_X1 U6878 ( .A1(n5411), .A2(n5410), .ZN(n7218) );
  OR2_X1 U6879 ( .A1(n4521), .A2(n7218), .ZN(n5413) );
  INV_X1 U6880 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7159) );
  OR2_X1 U6881 ( .A1(n6899), .A2(n7159), .ZN(n5412) );
  NAND4_X1 U6882 ( .A1(n5415), .A2(n5414), .A3(n5413), .A4(n5412), .ZN(n9383)
         );
  NAND2_X1 U6883 ( .A1(n9383), .A2(n5754), .ZN(n5416) );
  NAND2_X1 U6884 ( .A1(n5417), .A2(n5416), .ZN(n5418) );
  XNOR2_X1 U6885 ( .A(n5418), .B(n5898), .ZN(n5439) );
  NAND2_X1 U6886 ( .A1(n5900), .A2(n9383), .ZN(n5420) );
  NAND2_X1 U6887 ( .A1(n10067), .A2(n5319), .ZN(n5419) );
  NAND2_X1 U6888 ( .A1(n5420), .A2(n5419), .ZN(n7216) );
  XNOR2_X1 U6889 ( .A(n5422), .B(n5421), .ZN(n6740) );
  NAND2_X1 U6890 ( .A1(n6740), .A2(n5441), .ZN(n5428) );
  BUF_X1 U6891 ( .A(n5423), .Z(n5424) );
  INV_X1 U6892 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5425) );
  NAND2_X1 U6893 ( .A1(n5424), .A2(n5425), .ZN(n5470) );
  NAND2_X1 U6894 ( .A1(n5470), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5426) );
  XNOR2_X1 U6895 ( .A(n5426), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6823) );
  AOI22_X1 U6896 ( .A1(n8158), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5727), .B2(
        n6823), .ZN(n5427) );
  NAND2_X1 U6897 ( .A1(n5428), .A2(n5427), .ZN(n10081) );
  NAND2_X1 U6898 ( .A1(n10081), .A2(n5921), .ZN(n5436) );
  NAND2_X1 U6899 ( .A1(n5928), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5434) );
  INV_X1 U6900 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n5429) );
  OR2_X1 U6901 ( .A1(n5653), .A2(n5429), .ZN(n5433) );
  AND2_X1 U6902 ( .A1(n5446), .A2(n6818), .ZN(n5430) );
  OR2_X1 U6903 ( .A1(n5430), .A2(n5472), .ZN(n7251) );
  OR2_X1 U6904 ( .A1(n4520), .A2(n7251), .ZN(n5432) );
  INV_X1 U6905 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7228) );
  OR2_X1 U6906 ( .A1(n6899), .A2(n7228), .ZN(n5431) );
  NAND4_X1 U6907 ( .A1(n5434), .A2(n5433), .A3(n5432), .A4(n5431), .ZN(n9381)
         );
  NAND2_X1 U6908 ( .A1(n9381), .A2(n5754), .ZN(n5435) );
  NAND2_X1 U6909 ( .A1(n5436), .A2(n5435), .ZN(n5437) );
  XNOR2_X1 U6910 ( .A(n5437), .B(n5322), .ZN(n5464) );
  AND2_X1 U6911 ( .A1(n5900), .A2(n9381), .ZN(n5438) );
  AOI21_X1 U6912 ( .B1(n10081), .B2(n5754), .A(n5438), .ZN(n5465) );
  XNOR2_X1 U6913 ( .A(n5464), .B(n5465), .ZN(n7248) );
  INV_X1 U6914 ( .A(n5439), .ZN(n5440) );
  NAND2_X1 U6915 ( .A1(n6736), .A2(n5441), .ZN(n5444) );
  OR2_X1 U6916 ( .A1(n5424), .A2(n9899), .ZN(n5442) );
  XNOR2_X1 U6917 ( .A(n5442), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6806) );
  AOI22_X1 U6918 ( .A1(n8158), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5727), .B2(
        n6806), .ZN(n5443) );
  NAND2_X1 U6919 ( .A1(n5444), .A2(n5443), .ZN(n10072) );
  NAND2_X1 U6920 ( .A1(n5921), .A2(n10072), .ZN(n5453) );
  NAND2_X1 U6921 ( .A1(n5928), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5451) );
  INV_X1 U6922 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5445) );
  OR2_X1 U6923 ( .A1(n5653), .A2(n5445), .ZN(n5450) );
  OAI21_X1 U6924 ( .B1(n5447), .B2(P1_REG3_REG_6__SCAN_IN), .A(n5446), .ZN(
        n7199) );
  OR2_X1 U6925 ( .A1(n4520), .A2(n7199), .ZN(n5449) );
  INV_X1 U6926 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7183) );
  OR2_X1 U6927 ( .A1(n6899), .A2(n7183), .ZN(n5448) );
  NAND4_X1 U6928 ( .A1(n5451), .A2(n5450), .A3(n5449), .A4(n5448), .ZN(n9382)
         );
  NAND2_X1 U6929 ( .A1(n9382), .A2(n5754), .ZN(n5452) );
  NAND2_X1 U6930 ( .A1(n5453), .A2(n5452), .ZN(n5454) );
  XNOR2_X1 U6931 ( .A(n5454), .B(n5322), .ZN(n5459) );
  NAND2_X1 U6932 ( .A1(n10072), .A2(n5754), .ZN(n5456) );
  NAND2_X1 U6933 ( .A1(n5900), .A2(n9382), .ZN(n5455) );
  NAND2_X1 U6934 ( .A1(n5456), .A2(n5455), .ZN(n5460) );
  XNOR2_X1 U6935 ( .A(n5459), .B(n5460), .ZN(n7196) );
  INV_X1 U6936 ( .A(n7196), .ZN(n5457) );
  NAND2_X1 U6937 ( .A1(n5458), .A2(n7193), .ZN(n5512) );
  INV_X1 U6938 ( .A(n7248), .ZN(n5463) );
  INV_X1 U6939 ( .A(n5459), .ZN(n5462) );
  INV_X1 U6940 ( .A(n5460), .ZN(n5461) );
  NAND2_X1 U6941 ( .A1(n5462), .A2(n5461), .ZN(n7245) );
  OR2_X1 U6942 ( .A1(n5463), .A2(n7245), .ZN(n5511) );
  INV_X1 U6943 ( .A(n5464), .ZN(n5466) );
  NAND2_X1 U6944 ( .A1(n5466), .A2(n5465), .ZN(n5517) );
  AND2_X1 U6945 ( .A1(n5511), .A2(n5517), .ZN(n5467) );
  NAND2_X1 U6946 ( .A1(n5537), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5491) );
  XNOR2_X1 U6947 ( .A(n5491), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6791) );
  AOI22_X1 U6948 ( .A1(n8158), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5727), .B2(
        n6791), .ZN(n5471) );
  NAND2_X1 U6949 ( .A1(n9962), .A2(n5921), .ZN(n5480) );
  NAND2_X1 U6950 ( .A1(n5380), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5478) );
  INV_X1 U6951 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6792) );
  OR2_X1 U6952 ( .A1(n5360), .A2(n6792), .ZN(n5477) );
  OR2_X1 U6953 ( .A1(n5472), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5473) );
  NAND2_X1 U6954 ( .A1(n5498), .A2(n5473), .ZN(n9963) );
  OR2_X1 U6955 ( .A1(n4520), .A2(n9963), .ZN(n5476) );
  INV_X1 U6956 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n5474) );
  OR2_X1 U6957 ( .A1(n6899), .A2(n5474), .ZN(n5475) );
  NAND4_X1 U6958 ( .A1(n5478), .A2(n5477), .A3(n5476), .A4(n5475), .ZN(n9380)
         );
  NAND2_X1 U6959 ( .A1(n9380), .A2(n5754), .ZN(n5479) );
  NAND2_X1 U6960 ( .A1(n5480), .A2(n5479), .ZN(n5481) );
  XNOR2_X1 U6961 ( .A(n5481), .B(n5322), .ZN(n5520) );
  XNOR2_X1 U6962 ( .A(n7444), .B(n5520), .ZN(n7384) );
  AND2_X1 U6963 ( .A1(n5900), .A2(n9380), .ZN(n5482) );
  AOI21_X1 U6964 ( .B1(n9962), .B2(n5754), .A(n5482), .ZN(n7385) );
  NAND2_X1 U6965 ( .A1(n5529), .A2(n5483), .ZN(n5485) );
  AND2_X1 U6966 ( .A1(n5484), .A2(n5530), .ZN(n5486) );
  NAND2_X1 U6967 ( .A1(n5485), .A2(n5486), .ZN(n5490) );
  INV_X1 U6968 ( .A(n5485), .ZN(n5488) );
  INV_X1 U6969 ( .A(n5486), .ZN(n5487) );
  NAND2_X1 U6970 ( .A1(n5490), .A2(n5489), .ZN(n6764) );
  NAND2_X1 U6971 ( .A1(n6764), .A2(n5441), .ZN(n5495) );
  INV_X1 U6972 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5535) );
  NAND2_X1 U6973 ( .A1(n5491), .A2(n5535), .ZN(n5492) );
  NAND2_X1 U6974 ( .A1(n5492), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5493) );
  XNOR2_X1 U6975 ( .A(n5493), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6876) );
  AOI22_X1 U6976 ( .A1(n8158), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5727), .B2(
        n6876), .ZN(n5494) );
  NAND2_X2 U6977 ( .A1(n5495), .A2(n5494), .ZN(n10096) );
  NAND2_X1 U6978 ( .A1(n10096), .A2(n5921), .ZN(n5506) );
  NAND2_X1 U6979 ( .A1(n5792), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5504) );
  INV_X1 U6980 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7404) );
  OR2_X1 U6981 ( .A1(n6899), .A2(n7404), .ZN(n5503) );
  NAND2_X1 U6982 ( .A1(n5498), .A2(n5497), .ZN(n5499) );
  NAND2_X1 U6983 ( .A1(n5542), .A2(n5499), .ZN(n7451) );
  OR2_X1 U6984 ( .A1(n4520), .A2(n7451), .ZN(n5502) );
  INV_X1 U6985 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5500) );
  OR2_X1 U6986 ( .A1(n5360), .A2(n5500), .ZN(n5501) );
  NAND4_X1 U6987 ( .A1(n5504), .A2(n5503), .A3(n5502), .A4(n5501), .ZN(n9379)
         );
  NAND2_X1 U6988 ( .A1(n9379), .A2(n5754), .ZN(n5505) );
  NAND2_X1 U6989 ( .A1(n5506), .A2(n5505), .ZN(n5507) );
  XNOR2_X1 U6990 ( .A(n5507), .B(n5322), .ZN(n5513) );
  NAND2_X1 U6991 ( .A1(n10096), .A2(n5754), .ZN(n5509) );
  NAND2_X1 U6992 ( .A1(n5900), .A2(n9379), .ZN(n5508) );
  NAND2_X1 U6993 ( .A1(n5509), .A2(n5508), .ZN(n5514) );
  NAND2_X1 U6994 ( .A1(n5513), .A2(n5514), .ZN(n7447) );
  AND2_X1 U6995 ( .A1(n7385), .A2(n7447), .ZN(n5510) );
  NAND2_X1 U6996 ( .A1(n7384), .A2(n5510), .ZN(n5527) );
  AND2_X1 U6997 ( .A1(n5512), .A2(n5511), .ZN(n5519) );
  INV_X1 U6998 ( .A(n5513), .ZN(n5516) );
  INV_X1 U6999 ( .A(n5514), .ZN(n5515) );
  NAND2_X1 U7000 ( .A1(n5516), .A2(n5515), .ZN(n7448) );
  AND2_X1 U7001 ( .A1(n5517), .A2(n7448), .ZN(n5518) );
  NAND2_X1 U7002 ( .A1(n5519), .A2(n5518), .ZN(n5525) );
  INV_X1 U7003 ( .A(n7448), .ZN(n5521) );
  INV_X1 U7004 ( .A(n5520), .ZN(n7443) );
  NOR2_X1 U7005 ( .A1(n5521), .A2(n7443), .ZN(n5523) );
  INV_X1 U7006 ( .A(n7447), .ZN(n5522) );
  NOR2_X1 U7007 ( .A1(n5523), .A2(n5522), .ZN(n5524) );
  NAND2_X1 U7008 ( .A1(n5525), .A2(n5524), .ZN(n5526) );
  NAND2_X1 U7009 ( .A1(n5527), .A2(n5526), .ZN(n5554) );
  INV_X1 U7010 ( .A(n5554), .ZN(n5552) );
  NAND2_X1 U7011 ( .A1(n5529), .A2(n5528), .ZN(n5531) );
  AND2_X1 U7012 ( .A1(n5531), .A2(n5530), .ZN(n5533) );
  XNOR2_X1 U7013 ( .A(n5533), .B(n5532), .ZN(n6761) );
  NAND2_X1 U7014 ( .A1(n6761), .A2(n5441), .ZN(n5540) );
  INV_X1 U7015 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5534) );
  NAND2_X1 U7016 ( .A1(n5535), .A2(n5534), .ZN(n5536) );
  OR2_X1 U7017 ( .A1(n5537), .A2(n5536), .ZN(n5558) );
  NAND2_X1 U7018 ( .A1(n5558), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5538) );
  XNOR2_X1 U7019 ( .A(n5538), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7073) );
  AOI22_X1 U7020 ( .A1(n8158), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5727), .B2(
        n7073), .ZN(n5539) );
  NAND2_X1 U7021 ( .A1(n5540), .A2(n5539), .ZN(n7545) );
  NAND2_X1 U7022 ( .A1(n7545), .A2(n5921), .ZN(n5549) );
  NAND2_X1 U7023 ( .A1(n5792), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5547) );
  INV_X1 U7024 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6879) );
  OR2_X1 U7025 ( .A1(n5360), .A2(n6879), .ZN(n5546) );
  AND2_X1 U7026 ( .A1(n5542), .A2(n5541), .ZN(n5543) );
  OR2_X1 U7027 ( .A1(n5543), .A2(n5562), .ZN(n7540) );
  OR2_X1 U7028 ( .A1(n4521), .A2(n7540), .ZN(n5545) );
  INV_X1 U7029 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6871) );
  OR2_X1 U7030 ( .A1(n6899), .A2(n6871), .ZN(n5544) );
  NAND4_X1 U7031 ( .A1(n5547), .A2(n5546), .A3(n5545), .A4(n5544), .ZN(n9378)
         );
  NAND2_X1 U7032 ( .A1(n9378), .A2(n5754), .ZN(n5548) );
  NAND2_X1 U7033 ( .A1(n5549), .A2(n5548), .ZN(n5550) );
  XNOR2_X1 U7034 ( .A(n5550), .B(n5898), .ZN(n5555) );
  INV_X1 U7035 ( .A(n5555), .ZN(n5551) );
  NAND2_X1 U7036 ( .A1(n5552), .A2(n5551), .ZN(n7537) );
  AND2_X1 U7037 ( .A1(n5900), .A2(n9378), .ZN(n5553) );
  AOI21_X1 U7038 ( .B1(n7545), .B2(n5319), .A(n5553), .ZN(n7538) );
  XNOR2_X1 U7039 ( .A(n5557), .B(n5556), .ZN(n6770) );
  NAND2_X1 U7040 ( .A1(n6770), .A2(n5441), .ZN(n5561) );
  NOR2_X1 U7041 ( .A1(n5558), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5580) );
  OR2_X1 U7042 ( .A1(n5580), .A2(n9899), .ZN(n5559) );
  XNOR2_X1 U7043 ( .A(n5559), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7078) );
  AOI22_X1 U7044 ( .A1(n8158), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5727), .B2(
        n7078), .ZN(n5560) );
  NAND2_X1 U7045 ( .A1(n7614), .A2(n5921), .ZN(n5569) );
  NAND2_X1 U7046 ( .A1(n5792), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5567) );
  INV_X1 U7047 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7079) );
  OR2_X1 U7048 ( .A1(n5360), .A2(n7079), .ZN(n5566) );
  NOR2_X1 U7049 ( .A1(n5562), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5563) );
  OR2_X1 U7050 ( .A1(n5584), .A2(n5563), .ZN(n7574) );
  OR2_X1 U7051 ( .A1(n4520), .A2(n7574), .ZN(n5565) );
  INV_X1 U7052 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7530) );
  OR2_X1 U7053 ( .A1(n6899), .A2(n7530), .ZN(n5564) );
  NAND4_X1 U7054 ( .A1(n5567), .A2(n5566), .A3(n5565), .A4(n5564), .ZN(n9377)
         );
  NAND2_X1 U7055 ( .A1(n9377), .A2(n5754), .ZN(n5568) );
  NAND2_X1 U7056 ( .A1(n5569), .A2(n5568), .ZN(n5570) );
  XNOR2_X1 U7057 ( .A(n5570), .B(n5898), .ZN(n5572) );
  AND2_X1 U7058 ( .A1(n5900), .A2(n9377), .ZN(n5571) );
  AOI21_X1 U7059 ( .B1(n7614), .B2(n5319), .A(n5571), .ZN(n5573) );
  NAND2_X1 U7060 ( .A1(n5572), .A2(n5573), .ZN(n9917) );
  INV_X1 U7061 ( .A(n5572), .ZN(n5575) );
  INV_X1 U7062 ( .A(n5573), .ZN(n5574) );
  NAND2_X1 U7063 ( .A1(n5575), .A2(n5574), .ZN(n5576) );
  AND2_X1 U7064 ( .A1(n9917), .A2(n5576), .ZN(n7572) );
  XNOR2_X1 U7065 ( .A(n5578), .B(n5577), .ZN(n6865) );
  NAND2_X1 U7066 ( .A1(n6865), .A2(n5441), .ZN(n5583) );
  INV_X1 U7067 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5579) );
  NAND2_X1 U7068 ( .A1(n5580), .A2(n5579), .ZN(n5581) );
  NAND2_X1 U7069 ( .A1(n5581), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5605) );
  XNOR2_X1 U7070 ( .A(n5605), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7373) );
  AOI22_X1 U7071 ( .A1(n8158), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5727), .B2(
        n7373), .ZN(n5582) );
  NAND2_X1 U7072 ( .A1(n10108), .A2(n5921), .ZN(n5593) );
  NAND2_X1 U7073 ( .A1(n5792), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5591) );
  INV_X1 U7074 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7071) );
  OR2_X1 U7075 ( .A1(n6899), .A2(n7071), .ZN(n5590) );
  INV_X1 U7076 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7077) );
  OR2_X1 U7077 ( .A1(n5360), .A2(n7077), .ZN(n5589) );
  INV_X1 U7078 ( .A(n5584), .ZN(n5586) );
  INV_X1 U7079 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5585) );
  NAND2_X1 U7080 ( .A1(n5586), .A2(n5585), .ZN(n5587) );
  NAND2_X1 U7081 ( .A1(n5611), .A2(n5587), .ZN(n9927) );
  OR2_X1 U7082 ( .A1(n4520), .A2(n9927), .ZN(n5588) );
  NAND4_X1 U7083 ( .A1(n5591), .A2(n5590), .A3(n5589), .A4(n5588), .ZN(n9376)
         );
  NAND2_X1 U7084 ( .A1(n9376), .A2(n5754), .ZN(n5592) );
  NAND2_X1 U7085 ( .A1(n5593), .A2(n5592), .ZN(n5594) );
  XNOR2_X1 U7086 ( .A(n5594), .B(n5898), .ZN(n5596) );
  AND2_X1 U7087 ( .A1(n5900), .A2(n9376), .ZN(n5595) );
  AOI21_X1 U7088 ( .B1(n10108), .B2(n5319), .A(n5595), .ZN(n5597) );
  NAND2_X1 U7089 ( .A1(n5596), .A2(n5597), .ZN(n5664) );
  INV_X1 U7090 ( .A(n5596), .ZN(n5599) );
  INV_X1 U7091 ( .A(n5597), .ZN(n5598) );
  NAND2_X1 U7092 ( .A1(n5599), .A2(n5598), .ZN(n5600) );
  AND2_X1 U7093 ( .A1(n5664), .A2(n5600), .ZN(n9915) );
  NAND2_X1 U7094 ( .A1(n9921), .A2(n5664), .ZN(n7722) );
  XNOR2_X1 U7095 ( .A(n5603), .B(n5602), .ZN(n6884) );
  NAND2_X1 U7096 ( .A1(n6884), .A2(n5441), .ZN(n5609) );
  INV_X1 U7097 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5604) );
  NAND2_X1 U7098 ( .A1(n5605), .A2(n5604), .ZN(n5606) );
  NAND2_X1 U7099 ( .A1(n5606), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5607) );
  XNOR2_X1 U7100 ( .A(n5607), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9496) );
  AOI22_X1 U7101 ( .A1(n9496), .A2(n5727), .B1(n8158), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n5608) );
  NAND2_X1 U7102 ( .A1(n7694), .A2(n5921), .ZN(n5619) );
  NAND2_X1 U7103 ( .A1(n5792), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5617) );
  NAND2_X1 U7104 ( .A1(n5611), .A2(n5610), .ZN(n5612) );
  NAND2_X1 U7105 ( .A1(n5629), .A2(n5612), .ZN(n7644) );
  OR2_X1 U7106 ( .A1(n4520), .A2(n7644), .ZN(n5616) );
  INV_X1 U7107 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n5613) );
  OR2_X1 U7108 ( .A1(n6899), .A2(n5613), .ZN(n5615) );
  INV_X1 U7109 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7362) );
  OR2_X1 U7110 ( .A1(n5360), .A2(n7362), .ZN(n5614) );
  NAND4_X1 U7111 ( .A1(n5617), .A2(n5616), .A3(n5615), .A4(n5614), .ZN(n9375)
         );
  NAND2_X1 U7112 ( .A1(n9375), .A2(n5754), .ZN(n5618) );
  NAND2_X1 U7113 ( .A1(n5619), .A2(n5618), .ZN(n5620) );
  XNOR2_X1 U7114 ( .A(n5620), .B(n5322), .ZN(n5639) );
  AND2_X1 U7115 ( .A1(n5900), .A2(n9375), .ZN(n5621) );
  AOI21_X1 U7116 ( .B1(n7694), .B2(n5319), .A(n5621), .ZN(n5640) );
  XNOR2_X1 U7117 ( .A(n5639), .B(n5640), .ZN(n7723) );
  NAND2_X1 U7118 ( .A1(n7722), .A2(n7723), .ZN(n7721) );
  XNOR2_X1 U7119 ( .A(n5623), .B(n5622), .ZN(n6978) );
  NAND2_X1 U7120 ( .A1(n6978), .A2(n5441), .ZN(n5627) );
  OR2_X1 U7121 ( .A1(n5624), .A2(n9899), .ZN(n5625) );
  XNOR2_X1 U7122 ( .A(n5625), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7377) );
  AOI22_X1 U7123 ( .A1(n8158), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5727), .B2(
        n7377), .ZN(n5626) );
  NAND2_X1 U7124 ( .A1(n9951), .A2(n5346), .ZN(n5637) );
  NAND2_X1 U7125 ( .A1(n5792), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5635) );
  INV_X1 U7126 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7376) );
  OR2_X1 U7127 ( .A1(n6899), .A2(n7376), .ZN(n5634) );
  NAND2_X1 U7128 ( .A1(n5629), .A2(n5628), .ZN(n5630) );
  NAND2_X1 U7129 ( .A1(n5649), .A2(n5630), .ZN(n9948) );
  OR2_X1 U7130 ( .A1(n4520), .A2(n9948), .ZN(n5633) );
  INV_X1 U7131 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n5631) );
  OR2_X1 U7132 ( .A1(n5360), .A2(n5631), .ZN(n5632) );
  NAND4_X1 U7133 ( .A1(n5635), .A2(n5634), .A3(n5633), .A4(n5632), .ZN(n9374)
         );
  NAND2_X1 U7134 ( .A1(n9374), .A2(n5754), .ZN(n5636) );
  NAND2_X1 U7135 ( .A1(n5637), .A2(n5636), .ZN(n5638) );
  XNOR2_X1 U7136 ( .A(n5638), .B(n5898), .ZN(n5667) );
  INV_X1 U7137 ( .A(n5667), .ZN(n5663) );
  INV_X1 U7138 ( .A(n5639), .ZN(n5641) );
  NAND2_X1 U7139 ( .A1(n5641), .A2(n5640), .ZN(n5662) );
  AND2_X1 U7140 ( .A1(n5663), .A2(n5662), .ZN(n5642) );
  NAND2_X1 U7141 ( .A1(n7721), .A2(n5642), .ZN(n8996) );
  XNOR2_X1 U7142 ( .A(n5643), .B(SI_15_), .ZN(n5644) );
  XNOR2_X1 U7143 ( .A(n5645), .B(n5644), .ZN(n7068) );
  NAND2_X1 U7144 ( .A1(n7068), .A2(n5441), .ZN(n5648) );
  XNOR2_X1 U7145 ( .A(n5646), .B(P1_IR_REG_15__SCAN_IN), .ZN(n7501) );
  AOI22_X1 U7146 ( .A1(n8158), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5727), .B2(
        n7501), .ZN(n5647) );
  NAND2_X1 U7147 ( .A1(n9121), .A2(n5921), .ZN(n5660) );
  INV_X1 U7148 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7369) );
  NAND2_X1 U7149 ( .A1(n5649), .A2(n7369), .ZN(n5650) );
  NAND2_X1 U7150 ( .A1(n5689), .A2(n5650), .ZN(n9119) );
  OR2_X1 U7151 ( .A1(n9119), .A2(n4521), .ZN(n5658) );
  INV_X1 U7152 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n5651) );
  OR2_X1 U7153 ( .A1(n5360), .A2(n5651), .ZN(n5657) );
  INV_X1 U7154 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n5652) );
  OR2_X1 U7155 ( .A1(n5653), .A2(n5652), .ZN(n5656) );
  INV_X1 U7156 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n5654) );
  OR2_X1 U7157 ( .A1(n6899), .A2(n5654), .ZN(n5655) );
  NAND4_X1 U7158 ( .A1(n5658), .A2(n5657), .A3(n5656), .A4(n5655), .ZN(n9373)
         );
  NAND2_X1 U7159 ( .A1(n9373), .A2(n5754), .ZN(n5659) );
  NAND2_X1 U7160 ( .A1(n5660), .A2(n5659), .ZN(n5661) );
  XNOR2_X1 U7161 ( .A(n5661), .B(n5898), .ZN(n5677) );
  OR2_X1 U7162 ( .A1(n5663), .A2(n5662), .ZN(n5666) );
  AND2_X1 U7163 ( .A1(n5664), .A2(n5666), .ZN(n5665) );
  NAND2_X1 U7164 ( .A1(n9921), .A2(n5665), .ZN(n5671) );
  INV_X1 U7165 ( .A(n5666), .ZN(n5669) );
  AND2_X1 U7166 ( .A1(n7723), .A2(n5667), .ZN(n5668) );
  OR2_X1 U7167 ( .A1(n5669), .A2(n5668), .ZN(n5670) );
  NAND2_X1 U7168 ( .A1(n5671), .A2(n5670), .ZN(n8997) );
  NAND2_X1 U7169 ( .A1(n9951), .A2(n5754), .ZN(n5673) );
  NAND2_X1 U7170 ( .A1(n5900), .A2(n9374), .ZN(n5672) );
  NAND2_X1 U7171 ( .A1(n5673), .A2(n5672), .ZN(n8999) );
  NAND2_X1 U7172 ( .A1(n8997), .A2(n8999), .ZN(n5676) );
  NAND3_X1 U7173 ( .A1(n8996), .A2(n5677), .A3(n5676), .ZN(n9112) );
  NAND2_X1 U7174 ( .A1(n9121), .A2(n5754), .ZN(n5675) );
  NAND2_X1 U7175 ( .A1(n5900), .A2(n9373), .ZN(n5674) );
  NAND2_X1 U7176 ( .A1(n5675), .A2(n5674), .ZN(n9115) );
  NAND2_X1 U7177 ( .A1(n9112), .A2(n9115), .ZN(n5680) );
  NAND2_X1 U7178 ( .A1(n8996), .A2(n5676), .ZN(n5679) );
  INV_X1 U7179 ( .A(n5677), .ZN(n5678) );
  NAND2_X1 U7180 ( .A1(n5679), .A2(n5678), .ZN(n9113) );
  NAND2_X1 U7181 ( .A1(n5680), .A2(n9113), .ZN(n9038) );
  INV_X1 U7182 ( .A(n9038), .ZN(n5701) );
  XNOR2_X1 U7183 ( .A(n5681), .B(SI_16_), .ZN(n5682) );
  XNOR2_X1 U7184 ( .A(n5683), .B(n5682), .ZN(n7102) );
  NAND2_X1 U7185 ( .A1(n7102), .A2(n5441), .ZN(n5687) );
  XNOR2_X1 U7186 ( .A(n5684), .B(n5685), .ZN(n7593) );
  AOI22_X1 U7187 ( .A1(n8158), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5727), .B2(
        n7593), .ZN(n5686) );
  NAND2_X1 U7188 ( .A1(n9045), .A2(n5346), .ZN(n5697) );
  INV_X1 U7189 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5688) );
  NAND2_X1 U7190 ( .A1(n5689), .A2(n5688), .ZN(n5690) );
  NAND2_X1 U7191 ( .A1(n5711), .A2(n5690), .ZN(n9043) );
  OR2_X1 U7192 ( .A1(n9043), .A2(n4521), .ZN(n5695) );
  NAND2_X1 U7193 ( .A1(n5928), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5694) );
  NAND2_X1 U7194 ( .A1(n5792), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5693) );
  NAND2_X1 U7195 ( .A1(n5691), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5692) );
  NAND4_X1 U7196 ( .A1(n5695), .A2(n5694), .A3(n5693), .A4(n5692), .ZN(n9372)
         );
  NAND2_X1 U7197 ( .A1(n9372), .A2(n5754), .ZN(n5696) );
  NAND2_X1 U7198 ( .A1(n5697), .A2(n5696), .ZN(n5698) );
  XNOR2_X1 U7199 ( .A(n5698), .B(n5322), .ZN(n5702) );
  NAND2_X1 U7200 ( .A1(n9045), .A2(n5754), .ZN(n5700) );
  NAND2_X1 U7201 ( .A1(n5900), .A2(n9372), .ZN(n5699) );
  NAND2_X1 U7202 ( .A1(n5700), .A2(n5699), .ZN(n5703) );
  NAND2_X2 U7203 ( .A1(n5701), .A2(n4599), .ZN(n9037) );
  INV_X1 U7204 ( .A(n5702), .ZN(n5705) );
  INV_X1 U7205 ( .A(n5703), .ZN(n5704) );
  NAND2_X1 U7206 ( .A1(n5705), .A2(n5704), .ZN(n9040) );
  XNOR2_X1 U7207 ( .A(n5707), .B(n5706), .ZN(n7130) );
  NAND2_X1 U7208 ( .A1(n7130), .A2(n5441), .ZN(n5710) );
  XNOR2_X1 U7209 ( .A(n5708), .B(P1_IR_REG_17__SCAN_IN), .ZN(n7752) );
  AOI22_X1 U7210 ( .A1(n8158), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5727), .B2(
        n7752), .ZN(n5709) );
  NAND2_X1 U7211 ( .A1(n9743), .A2(n5921), .ZN(n5717) );
  NAND2_X1 U7212 ( .A1(n5711), .A2(n7590), .ZN(n5712) );
  NAND2_X1 U7213 ( .A1(n5731), .A2(n5712), .ZN(n9741) );
  AOI22_X1 U7214 ( .A1(n5792), .A2(P1_REG0_REG_17__SCAN_IN), .B1(n5928), .B2(
        P1_REG1_REG_17__SCAN_IN), .ZN(n5715) );
  INV_X1 U7215 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n5713) );
  OR2_X1 U7216 ( .A1(n6899), .A2(n5713), .ZN(n5714) );
  OAI211_X1 U7217 ( .C1(n9741), .C2(n4521), .A(n5715), .B(n5714), .ZN(n9371)
         );
  NAND2_X1 U7218 ( .A1(n9371), .A2(n5319), .ZN(n5716) );
  NAND2_X1 U7219 ( .A1(n5717), .A2(n5716), .ZN(n5718) );
  XNOR2_X1 U7220 ( .A(n5718), .B(n5322), .ZN(n5720) );
  AND2_X1 U7221 ( .A1(n9371), .A2(n5900), .ZN(n5719) );
  AOI21_X1 U7222 ( .B1(n9743), .B2(n5319), .A(n5719), .ZN(n5721) );
  XNOR2_X1 U7223 ( .A(n5720), .B(n5721), .ZN(n9050) );
  INV_X1 U7224 ( .A(n5720), .ZN(n5722) );
  NAND2_X1 U7225 ( .A1(n5722), .A2(n5721), .ZN(n5723) );
  XNOR2_X1 U7226 ( .A(n5725), .B(n5724), .ZN(n7213) );
  NAND2_X1 U7227 ( .A1(n7213), .A2(n5441), .ZN(n5729) );
  XNOR2_X1 U7228 ( .A(n5726), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9524) );
  AOI22_X1 U7229 ( .A1(n8158), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9524), .B2(
        n5727), .ZN(n5728) );
  NAND2_X1 U7230 ( .A1(n9816), .A2(n5346), .ZN(n5737) );
  INV_X1 U7231 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n7744) );
  INV_X1 U7232 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5730) );
  NAND2_X1 U7233 ( .A1(n5731), .A2(n5730), .ZN(n5732) );
  NAND2_X1 U7234 ( .A1(n5733), .A2(n5732), .ZN(n9729) );
  OR2_X1 U7235 ( .A1(n9729), .A2(n4521), .ZN(n5735) );
  AOI22_X1 U7236 ( .A1(n5792), .A2(P1_REG0_REG_18__SCAN_IN), .B1(n5928), .B2(
        P1_REG1_REG_18__SCAN_IN), .ZN(n5734) );
  OAI211_X1 U7237 ( .C1(n6899), .C2(n7744), .A(n5735), .B(n5734), .ZN(n9370)
         );
  NAND2_X1 U7238 ( .A1(n9370), .A2(n5319), .ZN(n5736) );
  NAND2_X1 U7239 ( .A1(n5737), .A2(n5736), .ZN(n5738) );
  AOI22_X1 U7240 ( .A1(n9816), .A2(n5319), .B1(n5900), .B2(n9370), .ZN(n9087)
         );
  XOR2_X1 U7241 ( .A(n5740), .B(n5739), .Z(n9015) );
  XNOR2_X1 U7242 ( .A(n5741), .B(n10419), .ZN(n5742) );
  XNOR2_X1 U7243 ( .A(n5743), .B(n5742), .ZN(n7431) );
  NAND2_X1 U7244 ( .A1(n7431), .A2(n5441), .ZN(n5745) );
  NAND2_X1 U7245 ( .A1(n8158), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5744) );
  NAND2_X1 U7246 ( .A1(n9698), .A2(n5346), .ZN(n5756) );
  INV_X1 U7247 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5746) );
  NAND2_X1 U7248 ( .A1(n5747), .A2(n5746), .ZN(n5748) );
  NAND2_X1 U7249 ( .A1(n5765), .A2(n5748), .ZN(n9700) );
  OR2_X1 U7250 ( .A1(n9700), .A2(n4521), .ZN(n5753) );
  INV_X1 U7251 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9701) );
  NAND2_X1 U7252 ( .A1(n5792), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5750) );
  NAND2_X1 U7253 ( .A1(n5928), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5749) );
  OAI211_X1 U7254 ( .C1(n9701), .C2(n6899), .A(n5750), .B(n5749), .ZN(n5751)
         );
  INV_X1 U7255 ( .A(n5751), .ZN(n5752) );
  NAND2_X1 U7256 ( .A1(n5753), .A2(n5752), .ZN(n9024) );
  NAND2_X1 U7257 ( .A1(n9024), .A2(n5754), .ZN(n5755) );
  NAND2_X1 U7258 ( .A1(n5756), .A2(n5755), .ZN(n5757) );
  XNOR2_X1 U7259 ( .A(n5757), .B(n5898), .ZN(n9072) );
  AND2_X1 U7260 ( .A1(n9024), .A2(n5900), .ZN(n5758) );
  AOI21_X1 U7261 ( .B1(n9698), .B2(n5319), .A(n5758), .ZN(n9071) );
  INV_X1 U7262 ( .A(n9071), .ZN(n5760) );
  INV_X1 U7263 ( .A(n9072), .ZN(n5759) );
  XNOR2_X1 U7264 ( .A(n5761), .B(SI_21_), .ZN(n5762) );
  XNOR2_X1 U7265 ( .A(n4714), .B(n5762), .ZN(n7557) );
  NAND2_X1 U7266 ( .A1(n7557), .A2(n5441), .ZN(n5764) );
  NAND2_X1 U7267 ( .A1(n8158), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5763) );
  NAND2_X1 U7268 ( .A1(n5765), .A2(n9025), .ZN(n5766) );
  AND2_X1 U7269 ( .A1(n5767), .A2(n5766), .ZN(n9684) );
  NAND2_X1 U7270 ( .A1(n9684), .A2(n5889), .ZN(n5773) );
  INV_X1 U7271 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n5770) );
  NAND2_X1 U7272 ( .A1(n5380), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5769) );
  NAND2_X1 U7273 ( .A1(n5928), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5768) );
  OAI211_X1 U7274 ( .C1(n5770), .C2(n6899), .A(n5769), .B(n5768), .ZN(n5771)
         );
  INV_X1 U7275 ( .A(n5771), .ZN(n5772) );
  NAND2_X1 U7276 ( .A1(n5773), .A2(n5772), .ZN(n9368) );
  AOI22_X1 U7277 ( .A1(n9683), .A2(n5319), .B1(n5900), .B2(n9368), .ZN(n5778)
         );
  NAND2_X1 U7278 ( .A1(n9683), .A2(n5921), .ZN(n5775) );
  NAND2_X1 U7279 ( .A1(n9368), .A2(n5319), .ZN(n5774) );
  NAND2_X1 U7280 ( .A1(n5775), .A2(n5774), .ZN(n5776) );
  XNOR2_X1 U7281 ( .A(n5776), .B(n5322), .ZN(n5777) );
  XOR2_X1 U7282 ( .A(n5778), .B(n5777), .Z(n9022) );
  AOI22_X1 U7283 ( .A1(n9669), .A2(n5346), .B1(n5754), .B2(n9367), .ZN(n5779)
         );
  NAND2_X1 U7284 ( .A1(n5781), .A2(n5780), .ZN(n5804) );
  MUX2_X1 U7285 ( .A(n7639), .B(n10567), .S(n6714), .Z(n5783) );
  INV_X1 U7286 ( .A(SI_23_), .ZN(n5782) );
  NAND2_X1 U7287 ( .A1(n5783), .A2(n5782), .ZN(n5805) );
  INV_X1 U7288 ( .A(n5783), .ZN(n5784) );
  NAND2_X1 U7289 ( .A1(n5784), .A2(SI_23_), .ZN(n5785) );
  XNOR2_X1 U7290 ( .A(n5804), .B(n5803), .ZN(n7636) );
  NAND2_X1 U7291 ( .A1(n7636), .A2(n5441), .ZN(n5787) );
  NAND2_X1 U7292 ( .A1(n8158), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5786) );
  INV_X1 U7293 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5789) );
  NAND2_X1 U7294 ( .A1(n5790), .A2(n5789), .ZN(n5791) );
  NAND2_X1 U7295 ( .A1(n5837), .A2(n5791), .ZN(n9009) );
  OR2_X1 U7296 ( .A1(n9009), .A2(n4521), .ZN(n5798) );
  INV_X1 U7297 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n5795) );
  NAND2_X1 U7298 ( .A1(n5928), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5794) );
  NAND2_X1 U7299 ( .A1(n5792), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5793) );
  OAI211_X1 U7300 ( .C1(n5795), .C2(n6899), .A(n5794), .B(n5793), .ZN(n5796)
         );
  INV_X1 U7301 ( .A(n5796), .ZN(n5797) );
  NAND2_X1 U7302 ( .A1(n5798), .A2(n5797), .ZN(n9366) );
  AOI22_X1 U7303 ( .A1(n9862), .A2(n5921), .B1(n5319), .B2(n9366), .ZN(n5799)
         );
  XNOR2_X1 U7304 ( .A(n5799), .B(n5322), .ZN(n5801) );
  AOI22_X1 U7305 ( .A1(n9862), .A2(n5319), .B1(n5900), .B2(n9366), .ZN(n5800)
         );
  NAND2_X1 U7306 ( .A1(n5801), .A2(n5800), .ZN(n5802) );
  OAI21_X1 U7307 ( .B1(n5801), .B2(n5800), .A(n5802), .ZN(n9006) );
  INV_X1 U7308 ( .A(n5802), .ZN(n9060) );
  INV_X1 U7309 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7766) );
  MUX2_X1 U7310 ( .A(n7766), .B(n10588), .S(n5911), .Z(n5806) );
  NAND2_X1 U7311 ( .A1(n5806), .A2(n10577), .ZN(n5829) );
  INV_X1 U7312 ( .A(n5806), .ZN(n5807) );
  NAND2_X1 U7313 ( .A1(n5807), .A2(SI_24_), .ZN(n5808) );
  XNOR2_X1 U7314 ( .A(n5828), .B(n5827), .ZN(n7731) );
  NAND2_X1 U7315 ( .A1(n7731), .A2(n5441), .ZN(n5810) );
  NAND2_X1 U7316 ( .A1(n8158), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5809) );
  NAND2_X1 U7317 ( .A1(n9782), .A2(n5346), .ZN(n5818) );
  XNOR2_X1 U7318 ( .A(n5837), .B(P1_REG3_REG_24__SCAN_IN), .ZN(n9640) );
  NAND2_X1 U7319 ( .A1(n9640), .A2(n5889), .ZN(n5816) );
  INV_X1 U7320 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n5813) );
  NAND2_X1 U7321 ( .A1(n5928), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5812) );
  NAND2_X1 U7322 ( .A1(n5792), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5811) );
  OAI211_X1 U7323 ( .C1(n5813), .C2(n6899), .A(n5812), .B(n5811), .ZN(n5814)
         );
  INV_X1 U7324 ( .A(n5814), .ZN(n5815) );
  NAND2_X1 U7325 ( .A1(n5816), .A2(n5815), .ZN(n9365) );
  NAND2_X1 U7326 ( .A1(n9365), .A2(n5319), .ZN(n5817) );
  NAND2_X1 U7327 ( .A1(n5818), .A2(n5817), .ZN(n5819) );
  XNOR2_X1 U7328 ( .A(n5819), .B(n5898), .ZN(n5821) );
  AND2_X1 U7329 ( .A1(n9365), .A2(n5900), .ZN(n5820) );
  AOI21_X1 U7330 ( .B1(n9782), .B2(n5319), .A(n5820), .ZN(n5822) );
  NAND2_X1 U7331 ( .A1(n5821), .A2(n5822), .ZN(n5826) );
  INV_X1 U7332 ( .A(n5821), .ZN(n5824) );
  INV_X1 U7333 ( .A(n5822), .ZN(n5823) );
  NAND2_X1 U7334 ( .A1(n5824), .A2(n5823), .ZN(n5825) );
  AND2_X1 U7335 ( .A1(n5826), .A2(n5825), .ZN(n9059) );
  INV_X1 U7336 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8149) );
  INV_X1 U7337 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7772) );
  MUX2_X1 U7338 ( .A(n8149), .B(n7772), .S(n6714), .Z(n5831) );
  INV_X1 U7339 ( .A(SI_25_), .ZN(n5830) );
  NAND2_X1 U7340 ( .A1(n5831), .A2(n5830), .ZN(n5851) );
  INV_X1 U7341 ( .A(n5831), .ZN(n5832) );
  NAND2_X1 U7342 ( .A1(n5832), .A2(SI_25_), .ZN(n5833) );
  XNOR2_X1 U7343 ( .A(n5850), .B(n5849), .ZN(n7769) );
  NAND2_X1 U7344 ( .A1(n7769), .A2(n5441), .ZN(n5835) );
  NAND2_X1 U7345 ( .A1(n8158), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5834) );
  INV_X1 U7346 ( .A(n9857), .ZN(n5845) );
  INV_X1 U7347 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9065) );
  INV_X1 U7348 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5836) );
  OAI21_X1 U7349 ( .B1(n5837), .B2(n9065), .A(n5836), .ZN(n5838) );
  AND2_X1 U7350 ( .A1(n5838), .A2(n5860), .ZN(n9625) );
  NAND2_X1 U7351 ( .A1(n9625), .A2(n5889), .ZN(n5844) );
  INV_X1 U7352 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n5841) );
  NAND2_X1 U7353 ( .A1(n5928), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5840) );
  NAND2_X1 U7354 ( .A1(n5792), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5839) );
  OAI211_X1 U7355 ( .C1(n5841), .C2(n6899), .A(n5840), .B(n5839), .ZN(n5842)
         );
  INV_X1 U7356 ( .A(n5842), .ZN(n5843) );
  NAND2_X1 U7357 ( .A1(n5844), .A2(n5843), .ZN(n9364) );
  INV_X1 U7358 ( .A(n9364), .ZN(n9064) );
  OAI22_X1 U7359 ( .A1(n5845), .A2(n5389), .B1(n9064), .B2(n5294), .ZN(n5872)
         );
  NAND2_X1 U7360 ( .A1(n9857), .A2(n5921), .ZN(n5847) );
  NAND2_X1 U7361 ( .A1(n9364), .A2(n5319), .ZN(n5846) );
  NAND2_X1 U7362 ( .A1(n5847), .A2(n5846), .ZN(n5848) );
  XNOR2_X1 U7363 ( .A(n5848), .B(n5322), .ZN(n5871) );
  XOR2_X1 U7364 ( .A(n5872), .B(n5871), .Z(n9031) );
  NAND2_X1 U7365 ( .A1(n5850), .A2(n5849), .ZN(n5852) );
  NAND2_X1 U7366 ( .A1(n5852), .A2(n5851), .ZN(n5877) );
  INV_X1 U7367 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7817) );
  INV_X1 U7368 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10439) );
  MUX2_X1 U7369 ( .A(n7817), .B(n10439), .S(n6714), .Z(n5853) );
  INV_X1 U7370 ( .A(SI_26_), .ZN(n10578) );
  NAND2_X1 U7371 ( .A1(n5853), .A2(n10578), .ZN(n5878) );
  INV_X1 U7372 ( .A(n5853), .ZN(n5854) );
  NAND2_X1 U7373 ( .A1(n5854), .A2(SI_26_), .ZN(n5855) );
  XNOR2_X1 U7374 ( .A(n5877), .B(n5876), .ZN(n7816) );
  NAND2_X1 U7375 ( .A1(n7816), .A2(n5441), .ZN(n5857) );
  NAND2_X1 U7376 ( .A1(n8158), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5856) );
  NAND2_X1 U7377 ( .A1(n9853), .A2(n5346), .ZN(n5868) );
  INV_X1 U7378 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5859) );
  NAND2_X1 U7379 ( .A1(n5860), .A2(n5859), .ZN(n5861) );
  NAND2_X1 U7380 ( .A1(n5924), .A2(n5861), .ZN(n9610) );
  OR2_X1 U7381 ( .A1(n9610), .A2(n4520), .ZN(n5866) );
  INV_X1 U7382 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9609) );
  NAND2_X1 U7383 ( .A1(n5928), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5863) );
  NAND2_X1 U7384 ( .A1(n5792), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5862) );
  OAI211_X1 U7385 ( .C1(n9609), .C2(n6899), .A(n5863), .B(n5862), .ZN(n5864)
         );
  INV_X1 U7386 ( .A(n5864), .ZN(n5865) );
  NAND2_X1 U7387 ( .A1(n9363), .A2(n5319), .ZN(n5867) );
  NAND2_X1 U7388 ( .A1(n5868), .A2(n5867), .ZN(n5869) );
  XNOR2_X1 U7389 ( .A(n5869), .B(n5322), .ZN(n5908) );
  AND2_X1 U7390 ( .A1(n9363), .A2(n5900), .ZN(n5870) );
  AOI21_X1 U7391 ( .B1(n9853), .B2(n5319), .A(n5870), .ZN(n5906) );
  XNOR2_X1 U7392 ( .A(n5908), .B(n5906), .ZN(n9098) );
  INV_X1 U7393 ( .A(n5871), .ZN(n5874) );
  INV_X1 U7394 ( .A(n5872), .ZN(n5873) );
  NAND2_X1 U7395 ( .A1(n5874), .A2(n5873), .ZN(n9099) );
  NAND2_X1 U7396 ( .A1(n5877), .A2(n5876), .ZN(n5879) );
  NAND2_X1 U7397 ( .A1(n5879), .A2(n5878), .ZN(n5885) );
  INV_X1 U7398 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n6343) );
  INV_X1 U7399 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5880) );
  MUX2_X1 U7400 ( .A(n6343), .B(n5880), .S(n6714), .Z(n5881) );
  INV_X1 U7401 ( .A(SI_27_), .ZN(n10657) );
  NAND2_X1 U7402 ( .A1(n5881), .A2(n10657), .ZN(n5909) );
  INV_X1 U7403 ( .A(n5881), .ZN(n5882) );
  NAND2_X1 U7404 ( .A1(n5882), .A2(SI_27_), .ZN(n5883) );
  NAND2_X1 U7405 ( .A1(n5885), .A2(n5884), .ZN(n5910) );
  OR2_X1 U7406 ( .A1(n5885), .A2(n5884), .ZN(n5886) );
  NAND2_X1 U7407 ( .A1(n5910), .A2(n5886), .ZN(n7857) );
  NAND2_X1 U7408 ( .A1(n7857), .A2(n5441), .ZN(n5888) );
  NAND2_X1 U7409 ( .A1(n8158), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5887) );
  NAND2_X1 U7410 ( .A1(n9849), .A2(n5921), .ZN(n5897) );
  XNOR2_X1 U7411 ( .A(n5924), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9595) );
  NAND2_X1 U7412 ( .A1(n9595), .A2(n5889), .ZN(n5895) );
  INV_X1 U7413 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n5892) );
  NAND2_X1 U7414 ( .A1(n5928), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5891) );
  NAND2_X1 U7415 ( .A1(n5792), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5890) );
  OAI211_X1 U7416 ( .C1(n5892), .C2(n6899), .A(n5891), .B(n5890), .ZN(n5893)
         );
  INV_X1 U7417 ( .A(n5893), .ZN(n5894) );
  NAND2_X1 U7418 ( .A1(n9104), .A2(n5319), .ZN(n5896) );
  NAND2_X1 U7419 ( .A1(n5897), .A2(n5896), .ZN(n5899) );
  XNOR2_X1 U7420 ( .A(n5899), .B(n5898), .ZN(n5903) );
  INV_X1 U7421 ( .A(n5903), .ZN(n5905) );
  AND2_X1 U7422 ( .A1(n9104), .A2(n5900), .ZN(n5901) );
  AOI21_X1 U7423 ( .B1(n9849), .B2(n5319), .A(n5901), .ZN(n5902) );
  INV_X1 U7424 ( .A(n5902), .ZN(n5904) );
  AOI21_X1 U7425 ( .B1(n5905), .B2(n5904), .A(n5965), .ZN(n8990) );
  INV_X1 U7426 ( .A(n5906), .ZN(n5907) );
  NAND2_X1 U7427 ( .A1(n5908), .A2(n5907), .ZN(n8991) );
  NAND2_X1 U7428 ( .A1(n5910), .A2(n5909), .ZN(n5917) );
  INV_X1 U7429 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n6354) );
  INV_X1 U7430 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n5912) );
  MUX2_X1 U7431 ( .A(n6354), .B(n5912), .S(n6714), .Z(n5913) );
  INV_X1 U7432 ( .A(SI_28_), .ZN(n10435) );
  NAND2_X1 U7433 ( .A1(n5913), .A2(n10435), .ZN(n6369) );
  INV_X1 U7434 ( .A(n5913), .ZN(n5914) );
  NAND2_X1 U7435 ( .A1(n5914), .A2(SI_28_), .ZN(n5915) );
  NAND2_X1 U7436 ( .A1(n5917), .A2(n5916), .ZN(n6370) );
  OR2_X1 U7437 ( .A1(n5917), .A2(n5916), .ZN(n5918) );
  NAND2_X1 U7438 ( .A1(n6370), .A2(n5918), .ZN(n7884) );
  NAND2_X1 U7439 ( .A1(n7884), .A2(n5441), .ZN(n5920) );
  NAND2_X1 U7440 ( .A1(n8158), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5919) );
  NAND2_X1 U7441 ( .A1(n9760), .A2(n5921), .ZN(n5935) );
  INV_X1 U7442 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5923) );
  INV_X1 U7443 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5922) );
  OAI21_X1 U7444 ( .B1(n5924), .B2(n5923), .A(n5922), .ZN(n5927) );
  INV_X1 U7445 ( .A(n5924), .ZN(n5926) );
  AND2_X1 U7446 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P1_REG3_REG_27__SCAN_IN), 
        .ZN(n5925) );
  NAND2_X1 U7447 ( .A1(n5926), .A2(n5925), .ZN(n9558) );
  NAND2_X1 U7448 ( .A1(n5927), .A2(n9558), .ZN(n9575) );
  INV_X1 U7449 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9574) );
  NAND2_X1 U7450 ( .A1(n5792), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5930) );
  NAND2_X1 U7451 ( .A1(n5928), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5929) );
  OAI211_X1 U7452 ( .C1(n9574), .C2(n6899), .A(n5930), .B(n5929), .ZN(n5931)
         );
  INV_X1 U7453 ( .A(n5931), .ZN(n5932) );
  NAND2_X1 U7454 ( .A1(n9362), .A2(n5319), .ZN(n5934) );
  NAND2_X1 U7455 ( .A1(n5935), .A2(n5934), .ZN(n5936) );
  XNOR2_X1 U7456 ( .A(n5936), .B(n5322), .ZN(n5938) );
  AOI22_X1 U7457 ( .A1(n9760), .A2(n5319), .B1(n5900), .B2(n9362), .ZN(n5937)
         );
  XNOR2_X1 U7458 ( .A(n5938), .B(n5937), .ZN(n5966) );
  NAND2_X1 U7459 ( .A1(n7770), .A2(P1_B_REG_SCAN_IN), .ZN(n5940) );
  MUX2_X1 U7460 ( .A(n5940), .B(P1_B_REG_SCAN_IN), .S(n5939), .Z(n5941) );
  NAND2_X1 U7461 ( .A1(n5941), .A2(n5959), .ZN(n9896) );
  OAI22_X1 U7462 ( .A1(n9896), .A2(P1_D_REG_0__SCAN_IN), .B1(n5959), .B2(n5939), .ZN(n6619) );
  INV_X1 U7463 ( .A(n6619), .ZN(n5947) );
  NAND2_X1 U7464 ( .A1(n5943), .A2(n5942), .ZN(n5944) );
  NAND2_X1 U7465 ( .A1(n5944), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5946) );
  NAND3_X1 U7466 ( .A1(n5292), .A2(n9352), .A3(P1_STATE_REG_SCAN_IN), .ZN(
        n10038) );
  INV_X1 U7467 ( .A(n9896), .ZN(n6610) );
  NOR4_X1 U7468 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5951) );
  NOR4_X1 U7469 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n5950) );
  NOR4_X1 U7470 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5949) );
  NOR4_X1 U7471 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5948) );
  NAND4_X1 U7472 ( .A1(n5951), .A2(n5950), .A3(n5949), .A4(n5948), .ZN(n5957)
         );
  NOR2_X1 U7473 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .ZN(
        n5955) );
  NOR4_X1 U7474 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5954) );
  NOR4_X1 U7475 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5953) );
  NOR4_X1 U7476 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5952) );
  NAND4_X1 U7477 ( .A1(n5955), .A2(n5954), .A3(n5953), .A4(n5952), .ZN(n5956)
         );
  NOR2_X1 U7478 ( .A1(n5957), .A2(n5956), .ZN(n6608) );
  NAND2_X1 U7479 ( .A1(n6608), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5958) );
  NAND2_X1 U7480 ( .A1(n6610), .A2(n5958), .ZN(n5960) );
  INV_X1 U7481 ( .A(n5959), .ZN(n7831) );
  NAND2_X1 U7482 ( .A1(n7770), .A2(n7831), .ZN(n9898) );
  NAND2_X1 U7483 ( .A1(n5960), .A2(n9898), .ZN(n7149) );
  INV_X1 U7484 ( .A(n7149), .ZN(n5961) );
  NAND2_X1 U7485 ( .A1(n6614), .A2(n5961), .ZN(n5975) );
  INV_X1 U7486 ( .A(n5964), .ZN(n9350) );
  NAND2_X1 U7487 ( .A1(n9351), .A2(n5964), .ZN(n9289) );
  NAND2_X1 U7488 ( .A1(n10116), .A2(n9289), .ZN(n5977) );
  NAND3_X1 U7489 ( .A1(n8992), .A2(n9097), .A3(n5966), .ZN(n5987) );
  INV_X1 U7490 ( .A(n6605), .ZN(n7324) );
  OR2_X1 U7491 ( .A1(n7324), .A2(n9292), .ZN(n7161) );
  OR2_X1 U7492 ( .A1(n5975), .A2(n7161), .ZN(n5968) );
  NOR2_X1 U7493 ( .A1(n10038), .A2(n5964), .ZN(n5967) );
  AND2_X2 U7494 ( .A1(n5285), .A2(n5963), .ZN(n9222) );
  INV_X1 U7495 ( .A(n9399), .ZN(n9397) );
  OR2_X1 U7496 ( .A1(n9558), .A2(n4520), .ZN(n5974) );
  INV_X1 U7497 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9557) );
  NAND2_X1 U7498 ( .A1(n5792), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5971) );
  INV_X1 U7499 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6615) );
  OR2_X1 U7500 ( .A1(n5360), .A2(n6615), .ZN(n5970) );
  OAI211_X1 U7501 ( .C1(n9557), .C2(n6899), .A(n5971), .B(n5970), .ZN(n5972)
         );
  INV_X1 U7502 ( .A(n5972), .ZN(n5973) );
  NAND2_X1 U7503 ( .A1(n5974), .A2(n5973), .ZN(n9361) );
  AOI22_X1 U7504 ( .A1(n9104), .A2(n9101), .B1(n9103), .B2(n9361), .ZN(n9569)
         );
  INV_X1 U7505 ( .A(n9575), .ZN(n5981) );
  INV_X1 U7506 ( .A(n9292), .ZN(n9294) );
  NAND2_X1 U7507 ( .A1(n9294), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9349) );
  OR2_X1 U7508 ( .A1(n6567), .A2(n5976), .ZN(n7323) );
  NAND3_X1 U7509 ( .A1(n5977), .A2(n9349), .A3(n7323), .ZN(n5978) );
  OAI21_X1 U7510 ( .B1(n6619), .B2(n7149), .A(n5978), .ZN(n5980) );
  NAND2_X1 U7511 ( .A1(n5962), .A2(n6782), .ZN(n7147) );
  AND3_X1 U7512 ( .A1(n7147), .A2(n9352), .A3(n5292), .ZN(n5979) );
  NAND2_X1 U7513 ( .A1(n5980), .A2(n5979), .ZN(n6890) );
  AOI22_X1 U7514 ( .A1(n5981), .A2(n9105), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n5982) );
  OAI21_X1 U7515 ( .B1(n9569), .B2(n9914), .A(n5982), .ZN(n5983) );
  AOI21_X1 U7516 ( .B1(n9760), .B2(n9924), .A(n5983), .ZN(n5984) );
  NAND3_X1 U7517 ( .A1(n5988), .A2(n5987), .A3(n5986), .ZN(P1_U3220) );
  INV_X1 U7518 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6492) );
  INV_X1 U7519 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5991) );
  NAND2_X1 U7520 ( .A1(n6185), .A2(n5991), .ZN(n6195) );
  NAND2_X1 U7521 ( .A1(n6218), .A2(n6004), .ZN(n6229) );
  INV_X1 U7522 ( .A(n6229), .ZN(n5995) );
  INV_X1 U7523 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5994) );
  NAND3_X1 U7524 ( .A1(n5995), .A2(n6232), .A3(n5994), .ZN(n5996) );
  OR2_X1 U7525 ( .A1(n5997), .A2(n6003), .ZN(n5998) );
  NAND2_X1 U7526 ( .A1(n6257), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5999) );
  XNOR2_X2 U7527 ( .A(n5999), .B(n4763), .ZN(n8597) );
  INV_X1 U7528 ( .A(n7307), .ZN(n6009) );
  NOR2_X1 U7529 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n6002) );
  NOR2_X1 U7530 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n6001) );
  NOR2_X1 U7531 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n6000) );
  NAND4_X1 U7532 ( .A1(n6002), .A2(n6001), .A3(n6000), .A4(n6218), .ZN(n6007)
         );
  NAND4_X1 U7533 ( .A1(n6232), .A2(n6005), .A3(n6004), .A4(n6003), .ZN(n6006)
         );
  NAND2_X1 U7534 ( .A1(n6010), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6008) );
  INV_X1 U7535 ( .A(n10208), .ZN(n10184) );
  NOR2_X1 U7536 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n6012) );
  INV_X1 U7537 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6014) );
  NOR2_X1 U7538 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n6015) );
  NAND2_X2 U7539 ( .A1(n6018), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6032) );
  NAND2_X1 U7540 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), 
        .ZN(n6019) );
  XNOR2_X2 U7541 ( .A(n6020), .B(P2_IR_REG_29__SCAN_IN), .ZN(n6023) );
  INV_X2 U7542 ( .A(n6023), .ZN(n6024) );
  INV_X1 U7543 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6021) );
  OR2_X1 U7544 ( .A1(n7471), .A2(n6021), .ZN(n6030) );
  BUF_X2 U7545 ( .A(n6023), .Z(n8245) );
  NAND2_X4 U7546 ( .A1(n6025), .A2(n8245), .ZN(n7474) );
  OR2_X1 U7547 ( .A1(n7474), .A2(n6692), .ZN(n6029) );
  INV_X1 U7548 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6026) );
  OR2_X1 U7549 ( .A1(n6375), .A2(n6026), .ZN(n6028) );
  NAND4_X2 U7550 ( .A1(n6030), .A2(n6029), .A3(n6028), .A4(n6027), .ZN(n8419)
         );
  XNOR2_X2 U7551 ( .A(n6032), .B(n6031), .ZN(n6444) );
  XNOR2_X2 U7552 ( .A(n6033), .B(n6014), .ZN(n6445) );
  NAND2_X4 U7553 ( .A1(n6444), .A2(n6445), .ZN(n6627) );
  INV_X1 U7554 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8981) );
  OR2_X1 U7555 ( .A1(n6632), .A2(n8981), .ZN(n6035) );
  INV_X1 U7556 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6037) );
  OR2_X1 U7557 ( .A1(n6066), .A2(n6037), .ZN(n6039) );
  OR2_X1 U7558 ( .A1(n6065), .A2(n6732), .ZN(n6038) );
  INV_X1 U7559 ( .A(n7306), .ZN(n6384) );
  NAND2_X1 U7560 ( .A1(n8419), .A2(n6384), .ZN(n7989) );
  NAND2_X1 U7561 ( .A1(n6071), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6043) );
  NAND2_X1 U7562 ( .A1(n6070), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6042) );
  INV_X1 U7563 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7050) );
  OR2_X1 U7564 ( .A1(n6375), .A2(n7050), .ZN(n6041) );
  INV_X1 U7565 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7055) );
  NAND2_X1 U7566 ( .A1(n4506), .A2(SI_0_), .ZN(n6045) );
  INV_X1 U7567 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6044) );
  NAND2_X1 U7568 ( .A1(n6045), .A2(n6044), .ZN(n6047) );
  NAND2_X1 U7569 ( .A1(n6047), .A2(n6046), .ZN(n8987) );
  MUX2_X1 U7570 ( .A(n6929), .B(n8987), .S(n6627), .Z(n7057) );
  OR2_X1 U7571 ( .A1(n6381), .A2(n7057), .ZN(n7311) );
  NAND2_X1 U7572 ( .A1(n6071), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6051) );
  INV_X1 U7573 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6661) );
  INV_X1 U7574 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7319) );
  INV_X1 U7575 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6660) );
  NAND2_X1 U7576 ( .A1(n7311), .A2(n7987), .ZN(n7296) );
  NAND2_X1 U7577 ( .A1(n7297), .A2(n6056), .ZN(n7980) );
  NAND2_X1 U7578 ( .A1(n7469), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6062) );
  INV_X1 U7579 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6057) );
  OR2_X1 U7580 ( .A1(n7471), .A2(n6057), .ZN(n6061) );
  OR2_X1 U7581 ( .A1(n6375), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6060) );
  INV_X1 U7582 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6058) );
  NAND2_X1 U7583 ( .A1(n6063), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6064) );
  XNOR2_X1 U7584 ( .A(n6064), .B(n5989), .ZN(n6716) );
  OR2_X1 U7585 ( .A1(n6065), .A2(n6717), .ZN(n6068) );
  OR2_X1 U7586 ( .A1(n6066), .A2(n5143), .ZN(n6067) );
  OAI211_X1 U7587 ( .C1(n6627), .C2(n6716), .A(n6068), .B(n6067), .ZN(n7137)
         );
  NAND2_X1 U7588 ( .A1(n8418), .A2(n10186), .ZN(n7995) );
  NAND2_X1 U7589 ( .A1(n8003), .A2(n7995), .ZN(n7424) );
  INV_X1 U7590 ( .A(n7424), .ZN(n7948) );
  NAND2_X1 U7591 ( .A1(n7980), .A2(n7948), .ZN(n6069) );
  NAND2_X1 U7592 ( .A1(n6069), .A2(n8003), .ZN(n7204) );
  NAND2_X1 U7593 ( .A1(n6070), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6078) );
  INV_X1 U7594 ( .A(n6071), .ZN(n6237) );
  INV_X1 U7595 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n6072) );
  OR2_X1 U7596 ( .A1(n6237), .A2(n6072), .ZN(n6077) );
  NAND2_X1 U7597 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6073) );
  AND2_X1 U7598 ( .A1(n6088), .A2(n6073), .ZN(n10168) );
  OR2_X1 U7599 ( .A1(n6375), .A2(n10168), .ZN(n6076) );
  INV_X1 U7600 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6074) );
  OR2_X1 U7601 ( .A1(n7474), .A2(n6074), .ZN(n6075) );
  NAND4_X1 U7602 ( .A1(n6078), .A2(n6077), .A3(n6076), .A4(n6075), .ZN(n8417)
         );
  NAND2_X1 U7603 ( .A1(n6080), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6082) );
  INV_X1 U7604 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6081) );
  INV_X1 U7605 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6083) );
  OR2_X1 U7606 ( .A1(n6066), .A2(n6083), .ZN(n6085) );
  OR2_X1 U7607 ( .A1(n6065), .A2(n6720), .ZN(n6084) );
  OAI211_X1 U7608 ( .C1(n6627), .C2(n6974), .A(n6085), .B(n6084), .ZN(n7210)
         );
  XNOR2_X1 U7609 ( .A(n8417), .B(n10170), .ZN(n6388) );
  NAND2_X1 U7610 ( .A1(n7204), .A2(n7993), .ZN(n7203) );
  INV_X1 U7611 ( .A(n8417), .ZN(n7427) );
  NAND2_X1 U7612 ( .A1(n7427), .A2(n7210), .ZN(n7996) );
  NAND2_X1 U7613 ( .A1(n7203), .A2(n7996), .ZN(n7433) );
  NAND2_X1 U7614 ( .A1(n7469), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6093) );
  INV_X1 U7615 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7436) );
  OR2_X1 U7616 ( .A1(n6363), .A2(n7436), .ZN(n6092) );
  NAND2_X1 U7617 ( .A1(n6088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6089) );
  AND2_X1 U7618 ( .A1(n6099), .A2(n6089), .ZN(n7437) );
  OR2_X1 U7619 ( .A1(n6375), .A2(n7437), .ZN(n6091) );
  INV_X1 U7620 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6659) );
  OR2_X1 U7621 ( .A1(n7471), .A2(n6659), .ZN(n6090) );
  NAND4_X1 U7622 ( .A1(n6093), .A2(n6092), .A3(n6091), .A4(n6090), .ZN(n8416)
         );
  NAND2_X1 U7623 ( .A1(n6105), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6095) );
  INV_X1 U7624 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6094) );
  XNOR2_X1 U7625 ( .A(n6095), .B(n6094), .ZN(n7101) );
  OR2_X1 U7626 ( .A1(n6065), .A2(n6723), .ZN(n6097) );
  INV_X1 U7627 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6721) );
  OR2_X1 U7628 ( .A1(n7936), .A2(n6721), .ZN(n6096) );
  OAI211_X1 U7629 ( .C1(n6627), .C2(n7101), .A(n6097), .B(n6096), .ZN(n7439)
         );
  INV_X1 U7630 ( .A(n7439), .ZN(n10193) );
  NAND2_X1 U7631 ( .A1(n8416), .A2(n10193), .ZN(n8004) );
  NAND2_X1 U7632 ( .A1(n7433), .A2(n8004), .ZN(n7460) );
  OR2_X1 U7633 ( .A1(n8416), .A2(n10193), .ZN(n7997) );
  NAND2_X1 U7634 ( .A1(n6070), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6104) );
  INV_X1 U7635 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n6098) );
  OR2_X1 U7636 ( .A1(n6237), .A2(n6098), .ZN(n6103) );
  NAND2_X1 U7637 ( .A1(n6099), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6100) );
  AND2_X1 U7638 ( .A1(n6120), .A2(n6100), .ZN(n7276) );
  OR2_X1 U7639 ( .A1(n6375), .A2(n7276), .ZN(n6102) );
  INV_X1 U7640 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7464) );
  OR2_X1 U7641 ( .A1(n7474), .A2(n7464), .ZN(n6101) );
  NAND4_X1 U7642 ( .A1(n6104), .A2(n6103), .A3(n6102), .A4(n6101), .ZN(n8415)
         );
  INV_X1 U7643 ( .A(n8415), .ZN(n7513) );
  INV_X1 U7644 ( .A(n6112), .ZN(n6106) );
  NAND2_X1 U7645 ( .A1(n6106), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6107) );
  AOI22_X1 U7646 ( .A1(n6270), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6269), .B2(
        n7127), .ZN(n6109) );
  INV_X2 U7647 ( .A(n6065), .ZN(n6139) );
  NAND2_X1 U7648 ( .A1(n6736), .A2(n6139), .ZN(n6108) );
  NAND2_X1 U7649 ( .A1(n6109), .A2(n6108), .ZN(n7466) );
  NAND2_X1 U7650 ( .A1(n7513), .A2(n7466), .ZN(n7999) );
  AND2_X1 U7651 ( .A1(n7997), .A2(n7999), .ZN(n8010) );
  NAND2_X1 U7652 ( .A1(n7460), .A2(n8010), .ZN(n6110) );
  INV_X1 U7653 ( .A(n7466), .ZN(n7484) );
  NAND2_X1 U7654 ( .A1(n7484), .A2(n8415), .ZN(n8008) );
  NAND2_X1 U7655 ( .A1(n6110), .A2(n8008), .ZN(n7511) );
  NAND2_X1 U7656 ( .A1(n6740), .A2(n6139), .ZN(n6117) );
  NAND2_X1 U7657 ( .A1(n6112), .A2(n6111), .ZN(n6140) );
  NAND2_X1 U7658 ( .A1(n6140), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6114) );
  INV_X1 U7659 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6113) );
  NAND2_X1 U7660 ( .A1(n6114), .A2(n6113), .ZN(n6127) );
  OR2_X1 U7661 ( .A1(n6114), .A2(n6113), .ZN(n6115) );
  AOI22_X1 U7662 ( .A1(n6270), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6269), .B2(
        n7266), .ZN(n6116) );
  NAND2_X1 U7663 ( .A1(n7469), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6125) );
  INV_X1 U7664 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6676) );
  OR2_X1 U7665 ( .A1(n6363), .A2(n6676), .ZN(n6124) );
  NAND2_X1 U7666 ( .A1(n6120), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6121) );
  AND2_X1 U7667 ( .A1(n6132), .A2(n6121), .ZN(n7517) );
  OR2_X1 U7668 ( .A1(n6375), .A2(n7517), .ZN(n6123) );
  INV_X1 U7669 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6675) );
  OR2_X1 U7670 ( .A1(n7471), .A2(n6675), .ZN(n6122) );
  NAND4_X1 U7671 ( .A1(n6125), .A2(n6124), .A3(n6123), .A4(n6122), .ZN(n8414)
         );
  XNOR2_X1 U7672 ( .A(n10201), .B(n8414), .ZN(n8017) );
  NAND2_X1 U7673 ( .A1(n7511), .A2(n8017), .ZN(n6126) );
  INV_X1 U7674 ( .A(n8414), .ZN(n8020) );
  OR2_X1 U7675 ( .A1(n8020), .A2(n10201), .ZN(n8026) );
  NAND2_X1 U7676 ( .A1(n6757), .A2(n6139), .ZN(n6131) );
  NAND2_X1 U7677 ( .A1(n6127), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6129) );
  INV_X1 U7678 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6128) );
  INV_X1 U7679 ( .A(n6758), .ZN(n7345) );
  AOI22_X1 U7680 ( .A1(n6270), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6269), .B2(
        n7345), .ZN(n6130) );
  NAND2_X1 U7681 ( .A1(n6131), .A2(n6130), .ZN(n7568) );
  NAND2_X1 U7682 ( .A1(n7469), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6138) );
  INV_X1 U7683 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7566) );
  OR2_X1 U7684 ( .A1(n7474), .A2(n7566), .ZN(n6137) );
  NAND2_X1 U7685 ( .A1(n6132), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6133) );
  AND2_X1 U7686 ( .A1(n6151), .A2(n6133), .ZN(n7565) );
  OR2_X1 U7687 ( .A1(n6375), .A2(n7565), .ZN(n6136) );
  INV_X1 U7688 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6134) );
  OR2_X1 U7689 ( .A1(n7471), .A2(n6134), .ZN(n6135) );
  NAND4_X1 U7690 ( .A1(n6138), .A2(n6137), .A3(n6136), .A4(n6135), .ZN(n8413)
         );
  NOR2_X1 U7691 ( .A1(n7568), .A2(n6398), .ZN(n8027) );
  NAND2_X1 U7692 ( .A1(n7568), .A2(n6398), .ZN(n8022) );
  NAND2_X1 U7693 ( .A1(n6764), .A2(n6139), .ZN(n6149) );
  INV_X1 U7694 ( .A(n6140), .ZN(n6142) );
  NOR2_X1 U7695 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n6141) );
  INV_X1 U7696 ( .A(n6146), .ZN(n6143) );
  NAND2_X1 U7697 ( .A1(n6143), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6144) );
  MUX2_X1 U7698 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6144), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n6147) );
  INV_X1 U7699 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6145) );
  NAND2_X1 U7700 ( .A1(n6146), .A2(n6145), .ZN(n6158) );
  NAND2_X1 U7701 ( .A1(n6147), .A2(n6158), .ZN(n6765) );
  INV_X1 U7702 ( .A(n6765), .ZN(n7630) );
  AOI22_X1 U7703 ( .A1(n6270), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6269), .B2(
        n7630), .ZN(n6148) );
  NAND2_X1 U7704 ( .A1(n7469), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6157) );
  INV_X1 U7705 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7668) );
  OR2_X1 U7706 ( .A1(n6363), .A2(n7668), .ZN(n6156) );
  NAND2_X1 U7707 ( .A1(n6151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6152) );
  AND2_X1 U7708 ( .A1(n6165), .A2(n6152), .ZN(n7679) );
  OR2_X1 U7709 ( .A1(n6375), .A2(n7679), .ZN(n6155) );
  INV_X1 U7710 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6153) );
  OR2_X1 U7711 ( .A1(n7471), .A2(n6153), .ZN(n6154) );
  NAND4_X1 U7712 ( .A1(n6157), .A2(n6156), .A3(n6155), .A4(n6154), .ZN(n8412)
         );
  NAND2_X1 U7713 ( .A1(n7718), .A2(n7775), .ZN(n8023) );
  NAND2_X1 U7714 ( .A1(n8014), .A2(n8023), .ZN(n7955) );
  NAND2_X1 U7715 ( .A1(n6761), .A2(n6139), .ZN(n6164) );
  NAND2_X1 U7716 ( .A1(n6158), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6159) );
  MUX2_X1 U7717 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6159), .S(
        P2_IR_REG_10__SCAN_IN), .Z(n6162) );
  INV_X1 U7718 ( .A(n6160), .ZN(n6161) );
  NAND2_X1 U7719 ( .A1(n6162), .A2(n6161), .ZN(n6763) );
  INV_X1 U7720 ( .A(n6763), .ZN(n7712) );
  AOI22_X1 U7721 ( .A1(n6270), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6269), .B2(
        n7712), .ZN(n6163) );
  NAND2_X1 U7722 ( .A1(n7469), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6171) );
  INV_X1 U7723 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7740) );
  OR2_X1 U7724 ( .A1(n7474), .A2(n7740), .ZN(n6170) );
  NAND2_X1 U7725 ( .A1(n6165), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6166) );
  AND2_X1 U7726 ( .A1(n6177), .A2(n6166), .ZN(n7779) );
  OR2_X1 U7727 ( .A1(n6375), .A2(n7779), .ZN(n6169) );
  INV_X1 U7728 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6167) );
  OR2_X1 U7729 ( .A1(n7471), .A2(n6167), .ZN(n6168) );
  NAND4_X1 U7730 ( .A1(n6171), .A2(n6170), .A3(n6169), .A4(n6168), .ZN(n8411)
         );
  OR2_X1 U7731 ( .A1(n10212), .A2(n7820), .ZN(n8039) );
  AND2_X1 U7732 ( .A1(n8039), .A2(n8014), .ZN(n8028) );
  NAND2_X1 U7733 ( .A1(n10212), .A2(n7820), .ZN(n8036) );
  NAND2_X1 U7734 ( .A1(n6172), .A2(n8036), .ZN(n7783) );
  NAND2_X1 U7735 ( .A1(n6770), .A2(n6139), .ZN(n6175) );
  OR2_X1 U7736 ( .A1(n6160), .A2(n8981), .ZN(n6173) );
  XNOR2_X1 U7737 ( .A(n6173), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7796) );
  AOI22_X1 U7738 ( .A1(n6270), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6269), .B2(
        n7796), .ZN(n6174) );
  NAND2_X1 U7739 ( .A1(n6175), .A2(n6174), .ZN(n7819) );
  NAND2_X1 U7740 ( .A1(n7469), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6183) );
  INV_X1 U7741 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6176) );
  OR2_X1 U7742 ( .A1(n7471), .A2(n6176), .ZN(n6182) );
  NAND2_X1 U7743 ( .A1(n6177), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6178) );
  AND2_X1 U7744 ( .A1(n6189), .A2(n6178), .ZN(n7824) );
  OR2_X1 U7745 ( .A1(n6375), .A2(n7824), .ZN(n6181) );
  INV_X1 U7746 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6179) );
  OR2_X1 U7747 ( .A1(n6363), .A2(n6179), .ZN(n6180) );
  NAND2_X1 U7748 ( .A1(n7819), .A2(n7879), .ZN(n8041) );
  INV_X1 U7749 ( .A(n7959), .ZN(n6184) );
  NAND2_X1 U7750 ( .A1(n6865), .A2(n6139), .ZN(n6188) );
  OR2_X1 U7751 ( .A1(n6185), .A2(n8981), .ZN(n6186) );
  XNOR2_X1 U7752 ( .A(n6186), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7813) );
  AOI22_X1 U7753 ( .A1(n6270), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6269), .B2(
        n7813), .ZN(n6187) );
  NAND2_X1 U7754 ( .A1(n7469), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6194) );
  INV_X1 U7755 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7792) );
  OR2_X1 U7756 ( .A1(n7471), .A2(n7792), .ZN(n6193) );
  NAND2_X1 U7757 ( .A1(n6189), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6190) );
  AND2_X1 U7758 ( .A1(n6201), .A2(n6190), .ZN(n7876) );
  OR2_X1 U7759 ( .A1(n6375), .A2(n7876), .ZN(n6192) );
  INV_X1 U7760 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7840) );
  OR2_X1 U7761 ( .A1(n7474), .A2(n7840), .ZN(n6191) );
  NAND4_X1 U7762 ( .A1(n6194), .A2(n6193), .A3(n6192), .A4(n6191), .ZN(n8409)
         );
  INV_X1 U7763 ( .A(n8409), .ZN(n7907) );
  NAND2_X1 U7764 ( .A1(n7873), .A2(n7907), .ZN(n8044) );
  NAND2_X1 U7765 ( .A1(n8045), .A2(n8044), .ZN(n8047) );
  NAND2_X1 U7766 ( .A1(n7835), .A2(n8045), .ZN(n7861) );
  NAND2_X1 U7767 ( .A1(n6884), .A2(n6139), .ZN(n6198) );
  NAND2_X1 U7768 ( .A1(n6195), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6196) );
  XNOR2_X1 U7769 ( .A(n6196), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8473) );
  AOI22_X1 U7770 ( .A1(n6270), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6269), .B2(
        n8473), .ZN(n6197) );
  NAND2_X1 U7771 ( .A1(n7469), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6206) );
  INV_X1 U7772 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8440) );
  OR2_X1 U7773 ( .A1(n7471), .A2(n8440), .ZN(n6205) );
  NAND2_X1 U7774 ( .A1(n6201), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6202) );
  AND2_X1 U7775 ( .A1(n6211), .A2(n6202), .ZN(n7910) );
  OR2_X1 U7776 ( .A1(n6375), .A2(n7910), .ZN(n6204) );
  INV_X1 U7777 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8448) );
  INV_X1 U7778 ( .A(n8809), .ZN(n7905) );
  NOR2_X1 U7779 ( .A1(n8048), .A2(n7905), .ZN(n6207) );
  INV_X1 U7780 ( .A(n8048), .ZN(n7917) );
  NAND2_X1 U7781 ( .A1(n6978), .A2(n6139), .ZN(n6210) );
  NAND2_X1 U7782 ( .A1(n6208), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6231) );
  XNOR2_X1 U7783 ( .A(n6231), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8482) );
  AOI22_X1 U7784 ( .A1(n6270), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6269), .B2(
        n8482), .ZN(n6209) );
  NAND2_X1 U7785 ( .A1(n7469), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6217) );
  INV_X1 U7786 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8874) );
  OR2_X1 U7787 ( .A1(n7471), .A2(n8874), .ZN(n6216) );
  NAND2_X1 U7788 ( .A1(n6211), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6212) );
  AND2_X1 U7789 ( .A1(n6223), .A2(n6212), .ZN(n8814) );
  OR2_X1 U7790 ( .A1(n6375), .A2(n8814), .ZN(n6215) );
  INV_X1 U7791 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6213) );
  OR2_X1 U7792 ( .A1(n7474), .A2(n6213), .ZN(n6214) );
  NAND4_X1 U7793 ( .A1(n6217), .A2(n6216), .A3(n6215), .A4(n6214), .ZN(n8794)
         );
  INV_X1 U7794 ( .A(n8794), .ZN(n8173) );
  OR2_X1 U7795 ( .A1(n8974), .A2(n8173), .ZN(n8057) );
  NAND2_X1 U7796 ( .A1(n8974), .A2(n8173), .ZN(n8056) );
  NAND2_X1 U7797 ( .A1(n7068), .A2(n6139), .ZN(n6222) );
  NAND2_X1 U7798 ( .A1(n6231), .A2(n6218), .ZN(n6219) );
  NAND2_X1 U7799 ( .A1(n6219), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6220) );
  XNOR2_X1 U7800 ( .A(n6220), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8519) );
  AOI22_X1 U7801 ( .A1(n6270), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6269), .B2(
        n8519), .ZN(n6221) );
  NAND2_X1 U7802 ( .A1(n7469), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6228) );
  INV_X1 U7803 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8797) );
  OR2_X1 U7804 ( .A1(n6363), .A2(n8797), .ZN(n6227) );
  NAND2_X1 U7805 ( .A1(n6223), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6224) );
  AND2_X1 U7806 ( .A1(n6235), .A2(n6224), .ZN(n8798) );
  OR2_X1 U7807 ( .A1(n6375), .A2(n8798), .ZN(n6226) );
  INV_X1 U7808 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8871) );
  OR2_X1 U7809 ( .A1(n7471), .A2(n8871), .ZN(n6225) );
  NAND4_X1 U7810 ( .A1(n6228), .A2(n6227), .A3(n6226), .A4(n6225), .ZN(n8811)
         );
  INV_X1 U7811 ( .A(n8811), .ZN(n8262) );
  AND2_X1 U7812 ( .A1(n8967), .A2(n8262), .ZN(n8068) );
  OR2_X1 U7813 ( .A1(n8967), .A2(n8262), .ZN(n8063) );
  NAND2_X1 U7814 ( .A1(n7102), .A2(n6139), .ZN(n6234) );
  NAND2_X1 U7815 ( .A1(n6229), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6230) );
  NAND2_X1 U7816 ( .A1(n6231), .A2(n6230), .ZN(n6243) );
  XNOR2_X1 U7817 ( .A(n6243), .B(n6232), .ZN(n8527) );
  AOI22_X1 U7818 ( .A1(n6270), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6269), .B2(
        n8527), .ZN(n6233) );
  NAND2_X1 U7819 ( .A1(n6235), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U7820 ( .A1(n6248), .A2(n6236), .ZN(n8788) );
  NAND2_X1 U7821 ( .A1(n6360), .A2(n8788), .ZN(n6241) );
  INV_X1 U7822 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8868) );
  OR2_X1 U7823 ( .A1(n7471), .A2(n8868), .ZN(n6240) );
  INV_X1 U7824 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8959) );
  OR2_X1 U7825 ( .A1(n6237), .A2(n8959), .ZN(n6239) );
  INV_X1 U7826 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8787) );
  OR2_X1 U7827 ( .A1(n6363), .A2(n8787), .ZN(n6238) );
  NAND4_X1 U7828 ( .A1(n6241), .A2(n6240), .A3(n6239), .A4(n6238), .ZN(n8795)
         );
  NAND2_X1 U7829 ( .A1(n8961), .A2(n8769), .ZN(n8072) );
  NAND2_X1 U7830 ( .A1(n8780), .A2(n8072), .ZN(n6242) );
  NAND2_X1 U7831 ( .A1(n7130), .A2(n6139), .ZN(n6246) );
  OAI21_X1 U7832 ( .B1(n6243), .B2(P2_IR_REG_16__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6244) );
  XNOR2_X1 U7833 ( .A(n6244), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8567) );
  AOI22_X1 U7834 ( .A1(n6270), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6269), .B2(
        n8567), .ZN(n6245) );
  NAND2_X1 U7835 ( .A1(n6248), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6249) );
  NAND2_X1 U7836 ( .A1(n6262), .A2(n6249), .ZN(n8776) );
  NAND2_X1 U7837 ( .A1(n8776), .A2(n6360), .ZN(n6253) );
  NAND2_X1 U7838 ( .A1(n7469), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6252) );
  INV_X1 U7839 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8865) );
  OR2_X1 U7840 ( .A1(n7471), .A2(n8865), .ZN(n6251) );
  INV_X1 U7841 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8775) );
  OR2_X1 U7842 ( .A1(n7474), .A2(n8775), .ZN(n6250) );
  INV_X1 U7843 ( .A(n8080), .ZN(n6254) );
  NAND2_X1 U7844 ( .A1(n8955), .A2(n8753), .ZN(n8066) );
  NAND2_X1 U7845 ( .A1(n7213), .A2(n6139), .ZN(n6261) );
  NAND2_X1 U7846 ( .A1(n4591), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6255) );
  MUX2_X1 U7847 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6255), .S(
        P2_IR_REG_18__SCAN_IN), .Z(n6256) );
  INV_X1 U7848 ( .A(n6256), .ZN(n6259) );
  INV_X1 U7849 ( .A(n6257), .ZN(n6258) );
  NOR2_X1 U7850 ( .A1(n6259), .A2(n6258), .ZN(n8574) );
  AOI22_X1 U7851 ( .A1(n6270), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6269), .B2(
        n8574), .ZN(n6260) );
  NAND2_X1 U7852 ( .A1(n6262), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6263) );
  NAND2_X1 U7853 ( .A1(n6273), .A2(n6263), .ZN(n8758) );
  NAND2_X1 U7854 ( .A1(n8758), .A2(n6360), .ZN(n6268) );
  NAND2_X1 U7855 ( .A1(n6070), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6265) );
  NAND2_X1 U7856 ( .A1(n7469), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6264) );
  AND2_X1 U7857 ( .A1(n6265), .A2(n6264), .ZN(n6267) );
  INV_X1 U7858 ( .A(n7474), .ZN(n6275) );
  NAND2_X1 U7859 ( .A1(n6275), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6266) );
  NAND2_X1 U7860 ( .A1(n8365), .A2(n8771), .ZN(n8079) );
  NAND2_X1 U7861 ( .A1(n8081), .A2(n8079), .ZN(n8755) );
  NAND2_X1 U7862 ( .A1(n8860), .A2(n8081), .ZN(n8741) );
  NAND2_X1 U7863 ( .A1(n7282), .A2(n6139), .ZN(n6272) );
  AOI22_X1 U7864 ( .A1(n6270), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6438), .B2(
        n6269), .ZN(n6271) );
  NAND2_X1 U7865 ( .A1(n6273), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6274) );
  NAND2_X1 U7866 ( .A1(n6282), .A2(n6274), .ZN(n8748) );
  NAND2_X1 U7867 ( .A1(n8748), .A2(n6360), .ZN(n6278) );
  AOI22_X1 U7868 ( .A1(n6070), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n7469), .B2(
        P2_REG0_REG_19__SCAN_IN), .ZN(n6277) );
  NAND2_X1 U7869 ( .A1(n6275), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6276) );
  NAND2_X1 U7870 ( .A1(n8944), .A2(n8754), .ZN(n8086) );
  NAND2_X1 U7871 ( .A1(n8085), .A2(n8086), .ZN(n6416) );
  NAND2_X1 U7872 ( .A1(n8741), .A2(n8743), .ZN(n8740) );
  NAND2_X1 U7873 ( .A1(n7431), .A2(n6139), .ZN(n6281) );
  INV_X1 U7874 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6279) );
  OR2_X1 U7875 ( .A1(n7936), .A2(n6279), .ZN(n6280) );
  NAND2_X1 U7876 ( .A1(n6282), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6283) );
  NAND2_X1 U7877 ( .A1(n6293), .A2(n6283), .ZN(n8736) );
  NAND2_X1 U7878 ( .A1(n8736), .A2(n6360), .ZN(n6288) );
  INV_X1 U7879 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8735) );
  NAND2_X1 U7880 ( .A1(n6070), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6285) );
  NAND2_X1 U7881 ( .A1(n7469), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6284) );
  OAI211_X1 U7882 ( .C1(n8735), .C2(n7474), .A(n6285), .B(n6284), .ZN(n6286)
         );
  INV_X1 U7883 ( .A(n6286), .ZN(n6287) );
  NAND2_X1 U7884 ( .A1(n7557), .A2(n6139), .ZN(n6290) );
  OR2_X1 U7885 ( .A1(n7936), .A2(n7558), .ZN(n6289) );
  INV_X1 U7886 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n6291) );
  NAND2_X1 U7887 ( .A1(n6293), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6294) );
  NAND2_X1 U7888 ( .A1(n6300), .A2(n6294), .ZN(n8726) );
  INV_X1 U7889 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8725) );
  NAND2_X1 U7890 ( .A1(n6070), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6296) );
  NAND2_X1 U7891 ( .A1(n7469), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6295) );
  OAI211_X1 U7892 ( .C1(n8725), .C2(n6363), .A(n6296), .B(n6295), .ZN(n6297)
         );
  AND2_X1 U7893 ( .A1(n8713), .A2(n8094), .ZN(n8699) );
  NAND2_X1 U7894 ( .A1(n7579), .A2(n6139), .ZN(n6299) );
  OR2_X1 U7895 ( .A1(n7936), .A2(n7583), .ZN(n6298) );
  OR2_X2 U7896 ( .A1(n6300), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6307) );
  NAND2_X1 U7897 ( .A1(n6300), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6301) );
  NAND2_X1 U7898 ( .A1(n6307), .A2(n6301), .ZN(n8710) );
  INV_X1 U7899 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8709) );
  NAND2_X1 U7900 ( .A1(n6070), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6303) );
  NAND2_X1 U7901 ( .A1(n7469), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6302) );
  OAI211_X1 U7902 ( .C1(n8709), .C2(n7474), .A(n6303), .B(n6302), .ZN(n6304)
         );
  AND2_X1 U7903 ( .A1(n8699), .A2(n7979), .ZN(n8687) );
  NAND2_X1 U7904 ( .A1(n7636), .A2(n6139), .ZN(n6306) );
  OR2_X1 U7905 ( .A1(n7936), .A2(n7639), .ZN(n6305) );
  NAND2_X1 U7906 ( .A1(n6307), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6308) );
  NAND2_X1 U7907 ( .A1(n6319), .A2(n6308), .ZN(n8696) );
  NAND2_X1 U7908 ( .A1(n8696), .A2(n6360), .ZN(n6313) );
  INV_X1 U7909 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8695) );
  NAND2_X1 U7910 ( .A1(n6070), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6310) );
  NAND2_X1 U7911 ( .A1(n7469), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6309) );
  OAI211_X1 U7912 ( .C1(n8695), .C2(n6363), .A(n6310), .B(n6309), .ZN(n6311)
         );
  INV_X1 U7913 ( .A(n6311), .ZN(n6312) );
  INV_X1 U7914 ( .A(n8102), .ZN(n8098) );
  AND2_X1 U7915 ( .A1(n8687), .A2(n8098), .ZN(n6316) );
  INV_X1 U7916 ( .A(n7979), .ZN(n6315) );
  NAND2_X1 U7917 ( .A1(n8927), .A2(n8294), .ZN(n7977) );
  NAND2_X1 U7918 ( .A1(n8737), .A2(n8282), .ZN(n8714) );
  AND2_X1 U7919 ( .A1(n7977), .A2(n8700), .ZN(n6314) );
  NAND2_X1 U7920 ( .A1(n7731), .A2(n6139), .ZN(n6318) );
  OR2_X1 U7921 ( .A1(n7936), .A2(n7766), .ZN(n6317) );
  INV_X1 U7922 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10413) );
  NAND2_X1 U7923 ( .A1(n6319), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6320) );
  NAND2_X1 U7924 ( .A1(n6329), .A2(n6320), .ZN(n8683) );
  NAND2_X1 U7925 ( .A1(n8683), .A2(n6360), .ZN(n6326) );
  INV_X1 U7926 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6323) );
  NAND2_X1 U7927 ( .A1(n7469), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6322) );
  NAND2_X1 U7928 ( .A1(n6070), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6321) );
  OAI211_X1 U7929 ( .C1(n6323), .C2(n7474), .A(n6322), .B(n6321), .ZN(n6324)
         );
  INV_X1 U7930 ( .A(n6324), .ZN(n6325) );
  NAND2_X1 U7931 ( .A1(n8915), .A2(n8305), .ZN(n8099) );
  AND2_X1 U7932 ( .A1(n8099), .A2(n8674), .ZN(n8101) );
  NAND2_X1 U7933 ( .A1(n7769), .A2(n6139), .ZN(n6328) );
  OR2_X1 U7934 ( .A1(n6066), .A2(n8149), .ZN(n6327) );
  NAND2_X1 U7935 ( .A1(n6329), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6330) );
  NAND2_X1 U7936 ( .A1(n6347), .A2(n6330), .ZN(n8666) );
  NAND2_X1 U7937 ( .A1(n8666), .A2(n6360), .ZN(n6335) );
  INV_X1 U7938 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8671) );
  NAND2_X1 U7939 ( .A1(n7469), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6332) );
  NAND2_X1 U7940 ( .A1(n6070), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6331) );
  OAI211_X1 U7941 ( .C1(n6363), .C2(n8671), .A(n6332), .B(n6331), .ZN(n6333)
         );
  INV_X1 U7942 ( .A(n6333), .ZN(n6334) );
  NAND2_X1 U7943 ( .A1(n8909), .A2(n8385), .ZN(n8109) );
  NAND2_X1 U7944 ( .A1(n7816), .A2(n6139), .ZN(n6337) );
  OR2_X1 U7945 ( .A1(n7936), .A2(n7817), .ZN(n6336) );
  NAND2_X1 U7946 ( .A1(n8648), .A2(n6360), .ZN(n6342) );
  INV_X1 U7947 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8647) );
  NAND2_X1 U7948 ( .A1(n6070), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6339) );
  NAND2_X1 U7949 ( .A1(n7469), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6338) );
  OAI211_X1 U7950 ( .C1(n8647), .C2(n6363), .A(n6339), .B(n6338), .ZN(n6340)
         );
  INV_X1 U7951 ( .A(n6340), .ZN(n6341) );
  NOR2_X1 U7952 ( .A1(n8903), .A2(n8306), .ZN(n8112) );
  NAND2_X1 U7953 ( .A1(n8903), .A2(n8306), .ZN(n7968) );
  NAND2_X1 U7954 ( .A1(n7857), .A2(n6139), .ZN(n6345) );
  OR2_X1 U7955 ( .A1(n7936), .A2(n6343), .ZN(n6344) );
  OAI21_X1 U7956 ( .B1(n6347), .B2(P2_REG3_REG_26__SCAN_IN), .A(
        P2_REG3_REG_27__SCAN_IN), .ZN(n6348) );
  INV_X1 U7957 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10448) );
  INV_X1 U7958 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n10607) );
  NAND2_X1 U7959 ( .A1(n10448), .A2(n10607), .ZN(n6346) );
  NAND2_X1 U7960 ( .A1(n6348), .A2(n6358), .ZN(n8638) );
  NAND2_X1 U7961 ( .A1(n8638), .A2(n6360), .ZN(n6353) );
  INV_X1 U7962 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8637) );
  NAND2_X1 U7963 ( .A1(n6070), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6350) );
  NAND2_X1 U7964 ( .A1(n7469), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6349) );
  OAI211_X1 U7965 ( .C1(n8637), .C2(n7474), .A(n6350), .B(n6349), .ZN(n6351)
         );
  INV_X1 U7966 ( .A(n6351), .ZN(n6352) );
  OR2_X1 U7967 ( .A1(n8897), .A2(n8386), .ZN(n8117) );
  OAI21_X1 U7968 ( .B1(n8628), .B2(n8629), .A(n8117), .ZN(n8620) );
  NAND2_X1 U7969 ( .A1(n7884), .A2(n6139), .ZN(n6356) );
  OR2_X1 U7970 ( .A1(n7936), .A2(n6354), .ZN(n6355) );
  INV_X1 U7971 ( .A(n6358), .ZN(n6357) );
  NAND2_X1 U7972 ( .A1(n6357), .A2(n10599), .ZN(n8604) );
  NAND2_X1 U7973 ( .A1(n6358), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6359) );
  NAND2_X1 U7974 ( .A1(n8604), .A2(n6359), .ZN(n8625) );
  NAND2_X1 U7975 ( .A1(n8625), .A2(n6360), .ZN(n6366) );
  INV_X1 U7976 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8624) );
  NAND2_X1 U7977 ( .A1(n7469), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6362) );
  NAND2_X1 U7978 ( .A1(n6070), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6361) );
  OAI211_X1 U7979 ( .C1(n8624), .C2(n6363), .A(n6362), .B(n6361), .ZN(n6364)
         );
  INV_X1 U7980 ( .A(n6364), .ZN(n6365) );
  NAND2_X1 U7981 ( .A1(n8620), .A2(n8622), .ZN(n6368) );
  INV_X1 U7982 ( .A(n8633), .ZN(n8252) );
  OR2_X1 U7983 ( .A1(n8891), .A2(n8252), .ZN(n6367) );
  NAND2_X1 U7984 ( .A1(n6368), .A2(n6367), .ZN(n7939) );
  NAND2_X1 U7985 ( .A1(n6370), .A2(n6369), .ZN(n7923) );
  MUX2_X1 U7986 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n7931), .Z(n7921) );
  NAND2_X1 U7987 ( .A1(n7925), .A2(n6372), .ZN(n9907) );
  OR2_X1 U7988 ( .A1(n9907), .A2(n6065), .ZN(n6374) );
  INV_X1 U7989 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8244) );
  OR2_X1 U7990 ( .A1(n6066), .A2(n8244), .ZN(n6373) );
  OR2_X1 U7991 ( .A1(n8604), .A2(n6375), .ZN(n7478) );
  INV_X1 U7992 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8613) );
  NAND2_X1 U7993 ( .A1(n7469), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6377) );
  NAND2_X1 U7994 ( .A1(n6070), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6376) );
  OAI211_X1 U7995 ( .C1(n8613), .C2(n7474), .A(n6377), .B(n6376), .ZN(n6378)
         );
  INV_X1 U7996 ( .A(n6378), .ZN(n6379) );
  NAND2_X1 U7997 ( .A1(n7478), .A2(n6379), .ZN(n8623) );
  INV_X1 U7998 ( .A(n8623), .ZN(n6380) );
  NAND2_X1 U7999 ( .A1(n8615), .A2(n6380), .ZN(n7940) );
  INV_X1 U8000 ( .A(n8619), .ZN(n6457) );
  INV_X1 U8001 ( .A(n7057), .ZN(n7021) );
  NAND2_X1 U8002 ( .A1(n6381), .A2(n7021), .ZN(n7314) );
  OR2_X1 U8003 ( .A1(n8420), .A2(n7020), .ZN(n7301) );
  NAND2_X1 U8004 ( .A1(n7312), .A2(n7301), .ZN(n6383) );
  NAND2_X1 U8005 ( .A1(n4796), .A2(n6384), .ZN(n6385) );
  NAND2_X1 U8006 ( .A1(n8418), .A2(n7137), .ZN(n6386) );
  INV_X1 U8007 ( .A(n8418), .ZN(n7207) );
  NAND2_X1 U8008 ( .A1(n7207), .A2(n10186), .ZN(n6387) );
  NAND2_X1 U8009 ( .A1(n7205), .A2(n6388), .ZN(n6390) );
  NAND2_X1 U8010 ( .A1(n7427), .A2(n10170), .ZN(n6389) );
  INV_X1 U8011 ( .A(n8416), .ZN(n7271) );
  NAND2_X1 U8012 ( .A1(n7434), .A2(n7271), .ZN(n6391) );
  NAND2_X1 U8013 ( .A1(n6391), .A2(n7439), .ZN(n6393) );
  OR2_X1 U8014 ( .A1(n7434), .A2(n7271), .ZN(n6392) );
  AND2_X1 U8015 ( .A1(n7466), .A2(n8415), .ZN(n6394) );
  NOR2_X1 U8016 ( .A1(n10201), .A2(n8414), .ZN(n6396) );
  NAND2_X1 U8017 ( .A1(n10201), .A2(n8414), .ZN(n6395) );
  INV_X1 U8018 ( .A(n7568), .ZN(n10203) );
  NAND2_X1 U8019 ( .A1(n6397), .A2(n10203), .ZN(n6401) );
  INV_X1 U8020 ( .A(n7563), .ZN(n6399) );
  INV_X1 U8021 ( .A(n8413), .ZN(n6398) );
  NAND2_X1 U8022 ( .A1(n6399), .A2(n6398), .ZN(n6400) );
  OR2_X1 U8023 ( .A1(n7718), .A2(n8412), .ZN(n6402) );
  NAND2_X1 U8024 ( .A1(n10212), .A2(n8411), .ZN(n6403) );
  NAND2_X1 U8025 ( .A1(n7784), .A2(n7959), .ZN(n6405) );
  INV_X1 U8026 ( .A(n7879), .ZN(n8410) );
  NAND2_X1 U8027 ( .A1(n7819), .A2(n8410), .ZN(n6404) );
  AND2_X1 U8028 ( .A1(n7873), .A2(n8409), .ZN(n6406) );
  OR2_X1 U8029 ( .A1(n8048), .A2(n8809), .ZN(n8049) );
  NAND2_X1 U8030 ( .A1(n8048), .A2(n8809), .ZN(n8051) );
  NAND2_X1 U8031 ( .A1(n8049), .A2(n8051), .ZN(n7961) );
  NAND2_X1 U8032 ( .A1(n8974), .A2(n8794), .ZN(n6407) );
  NAND2_X1 U8033 ( .A1(n6408), .A2(n6407), .ZN(n8792) );
  AND2_X1 U8034 ( .A1(n8967), .A2(n8811), .ZN(n7963) );
  NAND2_X1 U8035 ( .A1(n8069), .A2(n8072), .ZN(n8782) );
  NAND2_X1 U8036 ( .A1(n8961), .A2(n8795), .ZN(n6411) );
  NAND2_X1 U8037 ( .A1(n8781), .A2(n6411), .ZN(n8764) );
  NAND2_X1 U8038 ( .A1(n8080), .A2(n8066), .ZN(n8065) );
  INV_X1 U8039 ( .A(n8753), .ZN(n8784) );
  NAND2_X1 U8040 ( .A1(n8955), .A2(n8784), .ZN(n6412) );
  OR2_X1 U8041 ( .A1(n8365), .A2(n8744), .ZN(n6413) );
  NAND2_X1 U8042 ( .A1(n8751), .A2(n6413), .ZN(n6415) );
  NAND2_X1 U8043 ( .A1(n8365), .A2(n8744), .ZN(n6414) );
  NAND2_X1 U8044 ( .A1(n6415), .A2(n6414), .ZN(n8742) );
  NAND2_X1 U8045 ( .A1(n8742), .A2(n6416), .ZN(n6418) );
  INV_X1 U8046 ( .A(n8754), .ZN(n8408) );
  NAND2_X1 U8047 ( .A1(n8944), .A2(n8408), .ZN(n6417) );
  NAND2_X1 U8048 ( .A1(n8094), .A2(n8093), .ZN(n8718) );
  INV_X1 U8049 ( .A(n8733), .ZN(n8707) );
  NAND2_X1 U8050 ( .A1(n7979), .A2(n7977), .ZN(n8651) );
  NOR2_X1 U8051 ( .A1(n8915), .A2(n8693), .ZN(n8657) );
  NOR2_X1 U8052 ( .A1(n8657), .A2(n5125), .ZN(n6419) );
  OR2_X1 U8053 ( .A1(n8921), .A2(n8706), .ZN(n8655) );
  AND2_X1 U8054 ( .A1(n6419), .A2(n8655), .ZN(n6425) );
  INV_X1 U8055 ( .A(n6425), .ZN(n6420) );
  NAND2_X1 U8056 ( .A1(n8921), .A2(n8706), .ZN(n8654) );
  OR2_X1 U8057 ( .A1(n6420), .A2(n8654), .ZN(n6424) );
  AND2_X1 U8058 ( .A1(n8651), .A2(n6424), .ZN(n6422) );
  NAND2_X1 U8059 ( .A1(n8915), .A2(n8693), .ZN(n8658) );
  NOR2_X1 U8060 ( .A1(n5125), .A2(n8659), .ZN(n6429) );
  INV_X1 U8061 ( .A(n6429), .ZN(n6421) );
  AND2_X1 U8062 ( .A1(n6422), .A2(n6421), .ZN(n6423) );
  NAND2_X1 U8063 ( .A1(n8652), .A2(n6423), .ZN(n6431) );
  INV_X1 U8064 ( .A(n6424), .ZN(n6427) );
  INV_X1 U8065 ( .A(n8294), .ZN(n8723) );
  OR2_X1 U8066 ( .A1(n8927), .A2(n8723), .ZN(n8653) );
  AND2_X1 U8067 ( .A1(n8653), .A2(n6425), .ZN(n6426) );
  NAND2_X1 U8068 ( .A1(n8903), .A2(n8664), .ZN(n6433) );
  NOR2_X1 U8069 ( .A1(n8903), .A2(n8664), .ZN(n6432) );
  NOR2_X1 U8070 ( .A1(n8891), .A2(n8633), .ZN(n6434) );
  INV_X1 U8071 ( .A(n8891), .ZN(n8127) );
  OAI22_X1 U8072 ( .A1(n8621), .A2(n6434), .B1(n8127), .B2(n8252), .ZN(n6435)
         );
  XNOR2_X1 U8073 ( .A(n6435), .B(n4758), .ZN(n6440) );
  NAND2_X1 U8074 ( .A1(n6438), .A2(n8145), .ZN(n6487) );
  NAND2_X1 U8075 ( .A1(n6440), .A2(n8813), .ZN(n6456) );
  INV_X1 U8076 ( .A(n8145), .ZN(n7581) );
  OAI21_X1 U8077 ( .B1(n8141), .B2(n8145), .A(n8597), .ZN(n6441) );
  INV_X1 U8078 ( .A(n6441), .ZN(n6442) );
  AND2_X1 U8079 ( .A1(n10215), .A2(n6442), .ZN(n6443) );
  NAND2_X1 U8080 ( .A1(n8141), .A2(n8597), .ZN(n7018) );
  INV_X1 U8081 ( .A(n6444), .ZN(n8142) );
  INV_X1 U8082 ( .A(n8555), .ZN(n8588) );
  NAND2_X1 U8083 ( .A1(n8142), .A2(n8588), .ZN(n6446) );
  AND2_X1 U8084 ( .A1(n6627), .A2(n6446), .ZN(n7023) );
  INV_X1 U8085 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n6450) );
  NAND2_X1 U8086 ( .A1(n7469), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6449) );
  INV_X1 U8087 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n6447) );
  OR2_X1 U8088 ( .A1(n7471), .A2(n6447), .ZN(n6448) );
  OAI211_X1 U8089 ( .C1(n6450), .C2(n6363), .A(n6449), .B(n6448), .ZN(n6451)
         );
  INV_X1 U8090 ( .A(n6451), .ZN(n6452) );
  NAND2_X1 U8091 ( .A1(n7478), .A2(n6452), .ZN(n8407) );
  AOI21_X1 U8092 ( .B1(P2_B_REG_SCAN_IN), .B2(n6627), .A(n8770), .ZN(n8606) );
  AOI22_X1 U8093 ( .A1(n8633), .A2(n8808), .B1(n8407), .B2(n8606), .ZN(n6453)
         );
  NAND2_X1 U8094 ( .A1(n6456), .A2(n6455), .ZN(n8611) );
  NAND2_X1 U8095 ( .A1(n6458), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6461) );
  INV_X1 U8096 ( .A(n6461), .ZN(n6459) );
  NAND2_X1 U8097 ( .A1(n6459), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n6462) );
  INV_X1 U8098 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6460) );
  NAND2_X1 U8099 ( .A1(n6461), .A2(n6460), .ZN(n6463) );
  XNOR2_X1 U8100 ( .A(n7767), .B(P2_B_REG_SCAN_IN), .ZN(n6466) );
  NAND2_X1 U8101 ( .A1(n6463), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6465) );
  INV_X1 U8102 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6464) );
  NAND2_X1 U8103 ( .A1(n6466), .A2(n8150), .ZN(n6469) );
  NAND2_X1 U8104 ( .A1(n6467), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6468) );
  NAND2_X1 U8105 ( .A1(n6469), .A2(n6727), .ZN(n6724) );
  OR2_X1 U8106 ( .A1(n6724), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6471) );
  INV_X1 U8107 ( .A(n6727), .ZN(n7818) );
  NAND2_X1 U8108 ( .A1(n8150), .A2(n7818), .ZN(n6470) );
  NAND2_X1 U8109 ( .A1(n6471), .A2(n6470), .ZN(n7041) );
  NAND2_X1 U8110 ( .A1(n7818), .A2(n7767), .ZN(n6472) );
  OAI21_X2 U8111 ( .B1(n6724), .B2(P2_D_REG_0__SCAN_IN), .A(n6472), .ZN(n7040)
         );
  NOR2_X1 U8112 ( .A1(n7041), .A2(n7040), .ZN(n6497) );
  NOR2_X1 U8113 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6476) );
  NOR4_X1 U8114 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6475) );
  NOR4_X1 U8115 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6474) );
  NOR4_X1 U8116 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n6473) );
  NAND4_X1 U8117 ( .A1(n6476), .A2(n6475), .A3(n6474), .A4(n6473), .ZN(n6482)
         );
  NOR4_X1 U8118 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6480) );
  NOR4_X1 U8119 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n6479) );
  NOR4_X1 U8120 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6478) );
  NOR4_X1 U8121 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6477) );
  NAND4_X1 U8122 ( .A1(n6480), .A2(n6479), .A3(n6478), .A4(n6477), .ZN(n6481)
         );
  NOR2_X1 U8123 ( .A1(n6482), .A2(n6481), .ZN(n6483) );
  OR2_X1 U8124 ( .A1(n6724), .A2(n6483), .ZN(n6495) );
  NAND2_X1 U8125 ( .A1(n6497), .A2(n6495), .ZN(n6905) );
  INV_X1 U8126 ( .A(n6905), .ZN(n6486) );
  INV_X1 U8127 ( .A(n8150), .ZN(n6484) );
  INV_X1 U8128 ( .A(n7767), .ZN(n6726) );
  NAND3_X1 U8129 ( .A1(n6484), .A2(n6727), .A3(n6726), .ZN(n6630) );
  NAND2_X1 U8130 ( .A1(n4600), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6485) );
  XNOR2_X1 U8131 ( .A(n6485), .B(n6011), .ZN(n6629) );
  NOR2_X1 U8132 ( .A1(n6487), .A2(n8141), .ZN(n6488) );
  NAND2_X1 U8133 ( .A1(n7013), .A2(n6488), .ZN(n6918) );
  NAND2_X1 U8134 ( .A1(n7048), .A2(n6918), .ZN(n6489) );
  NAND2_X1 U8135 ( .A1(n6922), .A2(n6489), .ZN(n6491) );
  NAND3_X1 U8136 ( .A1(n8133), .A2(n6918), .A3(n10215), .ZN(n6916) );
  NAND2_X1 U8137 ( .A1(n6916), .A2(n8815), .ZN(n6906) );
  NAND2_X1 U8138 ( .A1(n6906), .A2(n7025), .ZN(n6490) );
  MUX2_X1 U8139 ( .A(n6492), .B(n6504), .S(n10221), .Z(n6493) );
  INV_X1 U8140 ( .A(n8615), .ZN(n6506) );
  NAND2_X1 U8141 ( .A1(n6493), .A2(n5123), .ZN(P2_U3456) );
  INV_X1 U8142 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6505) );
  INV_X1 U8143 ( .A(n6630), .ZN(n6494) );
  AOI21_X1 U8144 ( .B1(n8124), .B2(n7018), .A(n6494), .ZN(n6907) );
  NAND2_X1 U8145 ( .A1(n6495), .A2(n6725), .ZN(n6496) );
  NOR2_X1 U8146 ( .A1(n6497), .A2(n6496), .ZN(n6498) );
  NAND3_X1 U8147 ( .A1(n7014), .A2(n8145), .A3(n8597), .ZN(n6499) );
  OAI21_X1 U8148 ( .B1(n6924), .B2(n7040), .A(n7044), .ZN(n6502) );
  INV_X1 U8149 ( .A(n7044), .ZN(n6500) );
  NAND2_X1 U8150 ( .A1(n6500), .A2(n7041), .ZN(n6501) );
  AND2_X1 U8151 ( .A1(n6502), .A2(n6501), .ZN(n6503) );
  MUX2_X1 U8152 ( .A(n6505), .B(n6504), .S(n10233), .Z(n6507) );
  NAND2_X1 U8153 ( .A1(n10233), .A2(n10213), .ZN(n8864) );
  NAND2_X1 U8154 ( .A1(n6507), .A2(n5122), .ZN(P2_U3488) );
  INV_X1 U8155 ( .A(n6509), .ZN(n6508) );
  NAND2_X1 U8156 ( .A1(n6508), .A2(n10021), .ZN(n6571) );
  NAND2_X1 U8157 ( .A1(n6509), .A2(n10041), .ZN(n9298) );
  NAND2_X1 U8158 ( .A1(n9386), .A2(n10020), .ZN(n10010) );
  NAND2_X1 U8159 ( .A1(n6569), .A2(n10010), .ZN(n6511) );
  NAND2_X1 U8160 ( .A1(n4513), .A2(n10041), .ZN(n6510) );
  NAND2_X1 U8161 ( .A1(n6511), .A2(n6510), .ZN(n10000) );
  OR2_X1 U8162 ( .A1(n6512), .A2(n10050), .ZN(n6572) );
  NAND2_X1 U8163 ( .A1(n6512), .A2(n10050), .ZN(n9299) );
  NAND2_X1 U8164 ( .A1(n10000), .A2(n10001), .ZN(n6514) );
  INV_X1 U8165 ( .A(n6512), .ZN(n7009) );
  NAND2_X1 U8166 ( .A1(n7009), .A2(n10050), .ZN(n6513) );
  NAND2_X1 U8167 ( .A1(n6514), .A2(n6513), .ZN(n7287) );
  XNOR2_X2 U8168 ( .A(n9384), .B(n7290), .ZN(n9230) );
  INV_X1 U8169 ( .A(n9230), .ZN(n7288) );
  NAND2_X1 U8170 ( .A1(n7287), .A2(n7288), .ZN(n6516) );
  INV_X1 U8171 ( .A(n9384), .ZN(n7036) );
  NAND2_X1 U8172 ( .A1(n7036), .A2(n10055), .ZN(n6515) );
  NAND2_X1 U8173 ( .A1(n6516), .A2(n6515), .ZN(n9981) );
  OR2_X1 U8174 ( .A1(n6895), .A2(n10063), .ZN(n9127) );
  NAND2_X1 U8175 ( .A1(n6895), .A2(n10063), .ZN(n9300) );
  NAND2_X1 U8176 ( .A1(n9127), .A2(n9300), .ZN(n9982) );
  NAND2_X1 U8177 ( .A1(n9981), .A2(n9982), .ZN(n6518) );
  INV_X1 U8178 ( .A(n6895), .ZN(n7157) );
  NAND2_X1 U8179 ( .A1(n7157), .A2(n10063), .ZN(n6517) );
  NAND2_X1 U8180 ( .A1(n6518), .A2(n6517), .ZN(n7155) );
  INV_X1 U8181 ( .A(n9383), .ZN(n7181) );
  NAND2_X1 U8182 ( .A1(n7181), .A2(n10067), .ZN(n9128) );
  NAND2_X1 U8183 ( .A1(n9139), .A2(n9383), .ZN(n9302) );
  NAND2_X1 U8184 ( .A1(n9128), .A2(n9302), .ZN(n9232) );
  NAND2_X1 U8185 ( .A1(n7155), .A2(n9232), .ZN(n6520) );
  NAND2_X1 U8186 ( .A1(n7181), .A2(n9139), .ZN(n6519) );
  NAND2_X1 U8187 ( .A1(n6520), .A2(n6519), .ZN(n7178) );
  NOR2_X1 U8188 ( .A1(n10072), .A2(n9132), .ZN(n9125) );
  NAND2_X1 U8189 ( .A1(n10072), .A2(n9132), .ZN(n9129) );
  INV_X1 U8190 ( .A(n9129), .ZN(n9233) );
  OR2_X1 U8191 ( .A1(n9125), .A2(n9233), .ZN(n7179) );
  NAND2_X1 U8192 ( .A1(n7178), .A2(n7179), .ZN(n6522) );
  OR2_X1 U8193 ( .A1(n10072), .A2(n9382), .ZN(n6521) );
  NAND2_X1 U8194 ( .A1(n6522), .A2(n6521), .ZN(n7223) );
  INV_X1 U8195 ( .A(n9381), .ZN(n7180) );
  OR2_X1 U8196 ( .A1(n10081), .A2(n7180), .ZN(n9147) );
  NAND2_X1 U8197 ( .A1(n10081), .A2(n7180), .ZN(n7395) );
  NAND2_X1 U8198 ( .A1(n9147), .A2(n7395), .ZN(n9145) );
  OR2_X1 U8199 ( .A1(n10081), .A2(n9381), .ZN(n6523) );
  INV_X1 U8200 ( .A(n9380), .ZN(n7226) );
  INV_X1 U8201 ( .A(n9148), .ZN(n6524) );
  AND2_X1 U8202 ( .A1(n9962), .A2(n7226), .ZN(n9151) );
  OR2_X1 U8203 ( .A1(n9962), .A2(n9380), .ZN(n6525) );
  INV_X1 U8204 ( .A(n9379), .ZN(n6526) );
  OR2_X1 U8205 ( .A1(n10096), .A2(n6526), .ZN(n9161) );
  NAND2_X1 U8206 ( .A1(n10096), .A2(n6526), .ZN(n9162) );
  NAND2_X1 U8207 ( .A1(n9161), .A2(n9162), .ZN(n7397) );
  INV_X1 U8208 ( .A(n9378), .ZN(n6527) );
  NOR2_X1 U8209 ( .A1(n7545), .A2(n6527), .ZN(n9157) );
  INV_X1 U8210 ( .A(n9157), .ZN(n9305) );
  NAND2_X1 U8211 ( .A1(n7545), .A2(n6527), .ZN(n9163) );
  NAND2_X1 U8212 ( .A1(n7349), .A2(n7350), .ZN(n6529) );
  OR2_X1 U8213 ( .A1(n7545), .A2(n9378), .ZN(n6528) );
  NOR2_X1 U8214 ( .A1(n7614), .A2(n9377), .ZN(n6531) );
  INV_X1 U8215 ( .A(n7614), .ZN(n7611) );
  INV_X1 U8216 ( .A(n9377), .ZN(n6530) );
  OR2_X1 U8217 ( .A1(n7614), .A2(n6530), .ZN(n9164) );
  NAND2_X1 U8218 ( .A1(n7614), .A2(n6530), .ZN(n9165) );
  NAND2_X1 U8219 ( .A1(n9164), .A2(n9165), .ZN(n9240) );
  INV_X1 U8220 ( .A(n9376), .ZN(n6532) );
  OR2_X1 U8221 ( .A1(n10108), .A2(n6532), .ZN(n9167) );
  NAND2_X1 U8222 ( .A1(n10108), .A2(n6532), .ZN(n9312) );
  NAND2_X1 U8223 ( .A1(n9167), .A2(n9312), .ZN(n9241) );
  NAND2_X1 U8224 ( .A1(n7650), .A2(n9241), .ZN(n6534) );
  NAND2_X1 U8225 ( .A1(n10108), .A2(n9376), .ZN(n6533) );
  NAND2_X1 U8226 ( .A1(n6534), .A2(n6533), .ZN(n7640) );
  INV_X1 U8227 ( .A(n9375), .ZN(n9000) );
  OR2_X1 U8228 ( .A1(n7694), .A2(n9000), .ZN(n9175) );
  AND2_X1 U8229 ( .A1(n7694), .A2(n9000), .ZN(n9171) );
  NAND2_X1 U8230 ( .A1(n9175), .A2(n9316), .ZN(n9242) );
  NAND2_X1 U8231 ( .A1(n7640), .A2(n9242), .ZN(n6536) );
  NAND2_X1 U8232 ( .A1(n7694), .A2(n9375), .ZN(n6535) );
  NOR2_X1 U8233 ( .A1(n9121), .A2(n9373), .ZN(n6537) );
  INV_X1 U8234 ( .A(n9372), .ZN(n7848) );
  OR2_X1 U8235 ( .A1(n9045), .A2(n7848), .ZN(n9181) );
  NAND2_X1 U8236 ( .A1(n9045), .A2(n7848), .ZN(n9296) );
  NAND2_X1 U8237 ( .A1(n9045), .A2(n9372), .ZN(n6538) );
  NAND2_X1 U8238 ( .A1(n6539), .A2(n6538), .ZN(n9738) );
  AND2_X1 U8239 ( .A1(n9743), .A2(n9371), .ZN(n6540) );
  NOR2_X1 U8240 ( .A1(n9816), .A2(n9370), .ZN(n6541) );
  NAND2_X1 U8241 ( .A1(n9816), .A2(n9370), .ZN(n6542) );
  NAND2_X1 U8242 ( .A1(n6543), .A2(n6542), .ZN(n9718) );
  INV_X1 U8243 ( .A(n9718), .ZN(n6544) );
  NAND2_X1 U8244 ( .A1(n9879), .A2(n9092), .ZN(n6545) );
  NAND2_X1 U8245 ( .A1(n9698), .A2(n9024), .ZN(n6546) );
  NAND2_X1 U8246 ( .A1(n6547), .A2(n6546), .ZN(n9681) );
  OR2_X1 U8247 ( .A1(n9683), .A2(n9368), .ZN(n6548) );
  NAND2_X1 U8248 ( .A1(n9669), .A2(n9367), .ZN(n6550) );
  OR2_X1 U8249 ( .A1(n9862), .A2(n9366), .ZN(n6552) );
  INV_X1 U8250 ( .A(n9630), .ZN(n6553) );
  NAND2_X1 U8251 ( .A1(n9782), .A2(n9365), .ZN(n6554) );
  AND2_X1 U8252 ( .A1(n9857), .A2(n9364), .ZN(n6556) );
  NOR2_X1 U8253 ( .A1(n9853), .A2(n9363), .ZN(n6557) );
  INV_X1 U8254 ( .A(n9104), .ZN(n6558) );
  NOR2_X1 U8255 ( .A1(n9849), .A2(n6558), .ZN(n9213) );
  INV_X1 U8256 ( .A(n9213), .ZN(n9259) );
  NAND2_X1 U8257 ( .A1(n9849), .A2(n6558), .ZN(n9215) );
  NAND2_X1 U8258 ( .A1(n9592), .A2(n9591), .ZN(n9590) );
  OR2_X1 U8259 ( .A1(n9104), .A2(n9849), .ZN(n6559) );
  NAND2_X1 U8260 ( .A1(n9590), .A2(n6559), .ZN(n9573) );
  NAND2_X1 U8261 ( .A1(n9760), .A2(n9362), .ZN(n6560) );
  OR2_X1 U8262 ( .A1(n9760), .A2(n9362), .ZN(n6561) );
  NAND2_X1 U8263 ( .A1(n8158), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6563) );
  INV_X1 U8264 ( .A(n9361), .ZN(n6565) );
  NAND2_X1 U8265 ( .A1(n9560), .A2(n6565), .ZN(n9257) );
  NAND2_X1 U8266 ( .A1(n9283), .A2(n9257), .ZN(n9254) );
  INV_X1 U8267 ( .A(n10122), .ZN(n10084) );
  NAND2_X1 U8268 ( .A1(n5962), .A2(n6567), .ZN(n6568) );
  NAND3_X1 U8269 ( .A1(n7323), .A2(n7324), .A3(n6568), .ZN(n10009) );
  INV_X1 U8270 ( .A(n6569), .ZN(n6570) );
  INV_X1 U8271 ( .A(n10020), .ZN(n7004) );
  NOR2_X1 U8272 ( .A1(n9386), .A2(n7004), .ZN(n7002) );
  NAND2_X1 U8273 ( .A1(n10011), .A2(n6571), .ZN(n9992) );
  INV_X1 U8274 ( .A(n10001), .ZN(n9993) );
  NAND2_X1 U8275 ( .A1(n9992), .A2(n9993), .ZN(n9991) );
  NAND2_X1 U8276 ( .A1(n9384), .A2(n10055), .ZN(n9301) );
  NAND2_X1 U8277 ( .A1(n7284), .A2(n9301), .ZN(n6574) );
  NAND2_X1 U8278 ( .A1(n7036), .A2(n7290), .ZN(n6573) );
  NAND2_X1 U8279 ( .A1(n6574), .A2(n6573), .ZN(n9974) );
  NAND2_X1 U8280 ( .A1(n9126), .A2(n9128), .ZN(n7224) );
  INV_X1 U8281 ( .A(n7224), .ZN(n6578) );
  INV_X1 U8282 ( .A(n9152), .ZN(n6576) );
  INV_X1 U8283 ( .A(n9151), .ZN(n6575) );
  NAND2_X1 U8284 ( .A1(n6575), .A2(n7395), .ZN(n9150) );
  NAND2_X1 U8285 ( .A1(n6576), .A2(n9150), .ZN(n6577) );
  NAND3_X1 U8286 ( .A1(n6578), .A2(n9238), .A3(n9129), .ZN(n9307) );
  NAND2_X1 U8287 ( .A1(n9147), .A2(n4802), .ZN(n6579) );
  INV_X1 U8288 ( .A(n9236), .ZN(n6580) );
  NAND2_X1 U8289 ( .A1(n9238), .A2(n6580), .ZN(n9304) );
  NAND2_X1 U8290 ( .A1(n9307), .A2(n9304), .ZN(n7351) );
  INV_X1 U8291 ( .A(n9241), .ZN(n7660) );
  NAND2_X1 U8292 ( .A1(n6581), .A2(n9316), .ZN(n9941) );
  INV_X1 U8293 ( .A(n9374), .ZN(n7847) );
  NOR2_X1 U8294 ( .A1(n9951), .A2(n7847), .ZN(n9173) );
  INV_X1 U8295 ( .A(n9173), .ZN(n9319) );
  NAND2_X1 U8296 ( .A1(n9319), .A2(n9177), .ZN(n9943) );
  INV_X1 U8297 ( .A(n9943), .ZN(n9942) );
  INV_X1 U8298 ( .A(n9373), .ZN(n9001) );
  NOR2_X1 U8299 ( .A1(n9121), .A2(n9001), .ZN(n9321) );
  INV_X1 U8300 ( .A(n9321), .ZN(n9179) );
  NAND2_X1 U8301 ( .A1(n9121), .A2(n9001), .ZN(n9178) );
  INV_X1 U8302 ( .A(n9371), .ZN(n9090) );
  OR2_X1 U8303 ( .A1(n9743), .A2(n9090), .ZN(n9183) );
  NAND2_X1 U8304 ( .A1(n9743), .A2(n9090), .ZN(n9191) );
  NAND2_X1 U8305 ( .A1(n9183), .A2(n9191), .ZN(n9182) );
  INV_X1 U8306 ( .A(n9370), .ZN(n6583) );
  OR2_X1 U8307 ( .A1(n9816), .A2(n6583), .ZN(n9194) );
  NAND2_X1 U8308 ( .A1(n9816), .A2(n6583), .ZN(n9192) );
  NAND2_X1 U8309 ( .A1(n9194), .A2(n9192), .ZN(n9723) );
  INV_X1 U8310 ( .A(n9092), .ZN(n9369) );
  OR2_X1 U8311 ( .A1(n9879), .A2(n9369), .ZN(n9184) );
  NAND2_X1 U8312 ( .A1(n9184), .A2(n6584), .ZN(n9717) );
  XNOR2_X1 U8313 ( .A(n9698), .B(n9024), .ZN(n9691) );
  INV_X1 U8314 ( .A(n9024), .ZN(n9187) );
  AND2_X1 U8315 ( .A1(n9698), .A2(n9187), .ZN(n9124) );
  INV_X1 U8316 ( .A(n9124), .ZN(n9188) );
  NAND2_X1 U8317 ( .A1(n6585), .A2(n9188), .ZN(n9677) );
  XNOR2_X1 U8318 ( .A(n9683), .B(n9368), .ZN(n9680) );
  NAND2_X1 U8319 ( .A1(n9677), .A2(n9680), .ZN(n6586) );
  INV_X1 U8320 ( .A(n9368), .ZN(n9196) );
  NAND2_X1 U8321 ( .A1(n9683), .A2(n9196), .ZN(n9199) );
  INV_X1 U8322 ( .A(n9367), .ZN(n6587) );
  OR2_X1 U8323 ( .A1(n9669), .A2(n6587), .ZN(n9200) );
  NAND2_X1 U8324 ( .A1(n9669), .A2(n6587), .ZN(n9202) );
  NAND2_X1 U8325 ( .A1(n9663), .A2(n9662), .ZN(n6588) );
  INV_X1 U8326 ( .A(n9366), .ZN(n9082) );
  OR2_X1 U8327 ( .A1(n9862), .A2(n9082), .ZN(n9203) );
  NAND2_X1 U8328 ( .A1(n9862), .A2(n9082), .ZN(n9632) );
  NAND2_X1 U8329 ( .A1(n9203), .A2(n9632), .ZN(n9250) );
  INV_X1 U8330 ( .A(n9365), .ZN(n6589) );
  NAND2_X1 U8331 ( .A1(n9782), .A2(n6589), .ZN(n9269) );
  AND2_X1 U8332 ( .A1(n9631), .A2(n9632), .ZN(n6590) );
  OR2_X1 U8333 ( .A1(n9857), .A2(n9064), .ZN(n9264) );
  INV_X1 U8334 ( .A(n9264), .ZN(n9211) );
  NAND2_X1 U8335 ( .A1(n9857), .A2(n9064), .ZN(n9207) );
  XNOR2_X1 U8336 ( .A(n9853), .B(n9363), .ZN(n9604) );
  NAND2_X1 U8337 ( .A1(n9600), .A2(n9604), .ZN(n9584) );
  INV_X1 U8338 ( .A(n9363), .ZN(n9210) );
  NAND2_X1 U8339 ( .A1(n9853), .A2(n9210), .ZN(n9583) );
  NAND2_X1 U8340 ( .A1(n9584), .A2(n9583), .ZN(n6591) );
  NAND2_X1 U8341 ( .A1(n6591), .A2(n9252), .ZN(n9586) );
  INV_X1 U8342 ( .A(n9362), .ZN(n6592) );
  NAND2_X1 U8343 ( .A1(n9760), .A2(n6592), .ZN(n9216) );
  INV_X1 U8344 ( .A(n9254), .ZN(n6593) );
  NAND2_X1 U8345 ( .A1(n5285), .A2(n9351), .ZN(n6595) );
  NAND2_X1 U8346 ( .A1(n5964), .A2(n9294), .ZN(n6594) );
  INV_X1 U8347 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9552) );
  INV_X1 U8348 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n6596) );
  OR2_X1 U8349 ( .A1(n5360), .A2(n6596), .ZN(n6598) );
  NAND2_X1 U8350 ( .A1(n5792), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6597) );
  OAI211_X1 U8351 ( .C1(n6899), .C2(n9552), .A(n6598), .B(n6597), .ZN(n9360)
         );
  INV_X1 U8352 ( .A(n9360), .ZN(n9336) );
  INV_X1 U8353 ( .A(P1_B_REG_SCAN_IN), .ZN(n6599) );
  OR2_X1 U8354 ( .A1(n4519), .A2(n6599), .ZN(n6600) );
  NAND2_X1 U8355 ( .A1(n9103), .A2(n6600), .ZN(n8163) );
  NAND2_X1 U8356 ( .A1(n9362), .A2(n9101), .ZN(n6601) );
  OAI21_X1 U8357 ( .B1(n9336), .B2(n8163), .A(n6601), .ZN(n6602) );
  INV_X1 U8358 ( .A(n9853), .ZN(n9608) );
  INV_X1 U8359 ( .A(n9951), .ZN(n10117) );
  NAND2_X1 U8360 ( .A1(n10024), .A2(n10050), .ZN(n7289) );
  AND2_X1 U8361 ( .A1(n9987), .A2(n9139), .ZN(n7184) );
  INV_X1 U8362 ( .A(n10072), .ZN(n9135) );
  NAND2_X1 U8363 ( .A1(n7184), .A2(n9135), .ZN(n7229) );
  INV_X1 U8364 ( .A(n7545), .ZN(n10103) );
  OR2_X2 U8365 ( .A1(n7529), .A2(n7614), .ZN(n7651) );
  NAND2_X1 U8366 ( .A1(n9887), .A2(n9740), .ZN(n9739) );
  NOR2_X2 U8367 ( .A1(n9816), .A2(n9739), .ZN(n9728) );
  NOR2_X1 U8368 ( .A1(n9857), .A2(n9638), .ZN(n9624) );
  NAND2_X1 U8369 ( .A1(n9608), .A2(n9624), .ZN(n9607) );
  NAND2_X1 U8370 ( .A1(n6605), .A2(n9292), .ZN(n10003) );
  AOI21_X1 U8371 ( .B1(n9560), .B2(n9577), .A(n10003), .ZN(n6606) );
  NAND2_X1 U8372 ( .A1(n6606), .A2(n9550), .ZN(n9562) );
  NAND2_X1 U8373 ( .A1(n9566), .A2(n9562), .ZN(n6607) );
  AOI21_X1 U8374 ( .B1(n9564), .B2(n10112), .A(n6607), .ZN(n6621) );
  INV_X1 U8375 ( .A(n6608), .ZN(n6609) );
  NAND2_X1 U8376 ( .A1(n6610), .A2(n6609), .ZN(n6613) );
  OAI21_X1 U8377 ( .B1(n9896), .B2(P1_D_REG_1__SCAN_IN), .A(n9898), .ZN(n6612)
         );
  NAND2_X1 U8378 ( .A1(n10122), .A2(n9350), .ZN(n6611) );
  MUX2_X1 U8379 ( .A(n6615), .B(n6621), .S(n10141), .Z(n6618) );
  NAND2_X1 U8380 ( .A1(n9560), .A2(n6616), .ZN(n6617) );
  NAND2_X1 U8381 ( .A1(n6618), .A2(n6617), .ZN(P1_U3551) );
  INV_X1 U8382 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6622) );
  MUX2_X1 U8383 ( .A(n6622), .B(n6621), .S(n10125), .Z(n6625) );
  NAND2_X1 U8384 ( .A1(n9560), .A2(n6623), .ZN(n6624) );
  NAND2_X1 U8385 ( .A1(n6625), .A2(n6624), .ZN(P1_U3519) );
  NAND2_X1 U8386 ( .A1(n5259), .A2(n9352), .ZN(n6781) );
  NAND2_X1 U8387 ( .A1(n8133), .A2(n6630), .ZN(n6626) );
  NAND2_X1 U8388 ( .A1(n6626), .A2(n6629), .ZN(n6655) );
  NAND2_X1 U8389 ( .A1(n6655), .A2(n6627), .ZN(n6628) );
  NAND2_X1 U8390 ( .A1(n6628), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U8391 ( .A(n6629), .ZN(n7132) );
  OR2_X1 U8392 ( .A1(n6630), .A2(n7132), .ZN(n6686) );
  MUX2_X1 U8393 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6021), .S(n6036), .Z(n8423)
         );
  AND2_X1 U8394 ( .A1(n6929), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6633) );
  NAND2_X1 U8395 ( .A1(n6632), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6634) );
  OAI21_X1 U8396 ( .B1(n6718), .B2(n6633), .A(n6634), .ZN(n10144) );
  OR2_X1 U8397 ( .A1(n10144), .A2(n6660), .ZN(n10142) );
  NAND2_X1 U8398 ( .A1(n10142), .A2(n6634), .ZN(n8422) );
  NAND2_X1 U8399 ( .A1(n8423), .A2(n8422), .ZN(n8421) );
  NAND2_X1 U8400 ( .A1(n6036), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6635) );
  NAND2_X1 U8401 ( .A1(n8421), .A2(n6635), .ZN(n6636) );
  NAND2_X1 U8402 ( .A1(n6636), .A2(n6716), .ZN(n6956) );
  INV_X1 U8403 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6637) );
  MUX2_X1 U8404 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6637), .S(n6974), .Z(n6955)
         );
  NAND2_X1 U8405 ( .A1(n6974), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6638) );
  NAND2_X1 U8406 ( .A1(n6960), .A2(n6638), .ZN(n6639) );
  NAND2_X1 U8407 ( .A1(n6639), .A2(n7101), .ZN(n7116) );
  NAND2_X1 U8408 ( .A1(n7118), .A2(n7116), .ZN(n6640) );
  XNOR2_X1 U8409 ( .A(n7127), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n7115) );
  NAND2_X1 U8410 ( .A1(n6640), .A2(n7115), .ZN(n7120) );
  INV_X1 U8411 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6641) );
  OR2_X1 U8412 ( .A1(n7127), .A2(n6641), .ZN(n6642) );
  NAND2_X1 U8413 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n6758), .ZN(n6645) );
  OAI21_X1 U8414 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n6758), .A(n6645), .ZN(
        n7340) );
  NOR2_X1 U8415 ( .A1(n7341), .A2(n7340), .ZN(n7339) );
  AND2_X1 U8416 ( .A1(n6758), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6646) );
  NAND2_X1 U8417 ( .A1(n6648), .A2(n6765), .ZN(n6647) );
  INV_X1 U8418 ( .A(n6647), .ZN(n6649) );
  NAND2_X1 U8419 ( .A1(n6763), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6650) );
  OAI21_X1 U8420 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n6763), .A(n6650), .ZN(
        n7708) );
  INV_X1 U8421 ( .A(n6650), .ZN(n6651) );
  INV_X1 U8422 ( .A(n7796), .ZN(n7802) );
  NAND2_X1 U8423 ( .A1(n6652), .A2(n7802), .ZN(n7789) );
  OAI21_X1 U8424 ( .B1(n6652), .B2(n7802), .A(n7789), .ZN(n6653) );
  NOR2_X1 U8425 ( .A1(n6176), .A2(n6653), .ZN(n7790) );
  AOI21_X1 U8426 ( .B1(n6653), .B2(n6176), .A(n7790), .ZN(n6654) );
  NOR2_X1 U8427 ( .A1(n6444), .A2(P2_U3151), .ZN(n7885) );
  AND2_X1 U8428 ( .A1(n6655), .A2(n7885), .ZN(n6688) );
  INV_X1 U8429 ( .A(n6688), .ZN(n6932) );
  NOR2_X1 U8430 ( .A1(n6654), .A2(n10152), .ZN(n6713) );
  NOR2_X1 U8431 ( .A1(n8555), .A2(P2_U3151), .ZN(n7858) );
  NAND2_X1 U8432 ( .A1(n6655), .A2(n7858), .ZN(n6656) );
  MUX2_X1 U8433 ( .A(n8561), .B(n6656), .S(n6444), .Z(n8598) );
  NOR2_X1 U8434 ( .A1(n8598), .A2(n7802), .ZN(n6712) );
  MUX2_X1 U8435 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8555), .Z(n7803) );
  XNOR2_X1 U8436 ( .A(n7803), .B(n7796), .ZN(n6684) );
  MUX2_X1 U8437 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8555), .Z(n6657) );
  OR2_X1 U8438 ( .A1(n6657), .A2(n6763), .ZN(n6682) );
  XNOR2_X1 U8439 ( .A(n6657), .B(n7712), .ZN(n7702) );
  MUX2_X1 U8440 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8555), .Z(n6658) );
  OR2_X1 U8441 ( .A1(n6658), .A2(n6765), .ZN(n6681) );
  XNOR2_X1 U8442 ( .A(n6658), .B(n7630), .ZN(n7621) );
  MUX2_X1 U8443 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8555), .Z(n6679) );
  OR2_X1 U8444 ( .A1(n6679), .A2(n6758), .ZN(n6680) );
  MUX2_X1 U8445 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8555), .Z(n6673) );
  INV_X1 U8446 ( .A(n6673), .ZN(n6674) );
  INV_X1 U8447 ( .A(n7101), .ZN(n6672) );
  MUX2_X1 U8448 ( .A(n7436), .B(n6659), .S(n8555), .Z(n6671) );
  INV_X1 U8449 ( .A(n6974), .ZN(n6670) );
  MUX2_X1 U8450 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8555), .Z(n6668) );
  INV_X1 U8451 ( .A(n6668), .ZN(n6669) );
  MUX2_X1 U8452 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8555), .Z(n6666) );
  INV_X1 U8453 ( .A(n6666), .ZN(n6667) );
  INV_X1 U8454 ( .A(n6036), .ZN(n8433) );
  MUX2_X1 U8455 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8555), .Z(n6664) );
  INV_X1 U8456 ( .A(n6664), .ZN(n6665) );
  INV_X1 U8457 ( .A(n6718), .ZN(n10156) );
  MUX2_X1 U8458 ( .A(n6661), .B(n6660), .S(n6445), .Z(n6663) );
  XNOR2_X1 U8459 ( .A(n6663), .B(n6718), .ZN(n10149) );
  INV_X1 U8460 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6662) );
  MUX2_X1 U8461 ( .A(n7055), .B(n6662), .S(n8555), .Z(n6930) );
  NAND2_X1 U8462 ( .A1(n10149), .A2(n10148), .ZN(n10147) );
  OAI21_X1 U8463 ( .B1(n10156), .B2(n6663), .A(n10147), .ZN(n8432) );
  XOR2_X1 U8464 ( .A(n6036), .B(n6664), .Z(n8431) );
  NAND2_X1 U8465 ( .A1(n8432), .A2(n8431), .ZN(n8430) );
  OAI21_X1 U8466 ( .B1(n8433), .B2(n6665), .A(n8430), .ZN(n6938) );
  XNOR2_X1 U8467 ( .A(n6666), .B(n6716), .ZN(n6939) );
  NOR2_X1 U8468 ( .A1(n6938), .A2(n6939), .ZN(n6937) );
  XOR2_X1 U8469 ( .A(n6974), .B(n6668), .Z(n6953) );
  NAND2_X1 U8470 ( .A1(n6954), .A2(n6953), .ZN(n6952) );
  OAI21_X1 U8471 ( .B1(n6670), .B2(n6669), .A(n6952), .ZN(n7091) );
  XNOR2_X1 U8472 ( .A(n6671), .B(n7101), .ZN(n7090) );
  NAND2_X1 U8473 ( .A1(n7091), .A2(n7090), .ZN(n7089) );
  OAI21_X1 U8474 ( .B1(n6672), .B2(n6671), .A(n7089), .ZN(n7107) );
  XOR2_X1 U8475 ( .A(n7127), .B(n6673), .Z(n7108) );
  NOR2_X1 U8476 ( .A1(n7107), .A2(n7108), .ZN(n7106) );
  MUX2_X1 U8477 ( .A(n6676), .B(n6675), .S(n8555), .Z(n6677) );
  XNOR2_X1 U8478 ( .A(n6677), .B(n7266), .ZN(n7257) );
  INV_X1 U8479 ( .A(n6677), .ZN(n6678) );
  OAI22_X1 U8480 ( .A1(n7258), .A2(n7257), .B1(n6678), .B2(n6741), .ZN(n7335)
         );
  XNOR2_X1 U8481 ( .A(n6679), .B(n7345), .ZN(n7334) );
  NAND2_X1 U8482 ( .A1(n7335), .A2(n7334), .ZN(n7333) );
  NAND2_X1 U8483 ( .A1(n6680), .A2(n7333), .ZN(n7620) );
  NAND2_X1 U8484 ( .A1(n7621), .A2(n7620), .ZN(n7619) );
  NAND2_X1 U8485 ( .A1(n6681), .A2(n7619), .ZN(n7701) );
  NAND2_X1 U8486 ( .A1(n7702), .A2(n7701), .ZN(n7700) );
  NAND2_X1 U8487 ( .A1(n6682), .A2(n7700), .ZN(n6683) );
  OR2_X1 U8488 ( .A1(n6684), .A2(n6683), .ZN(n6685) );
  NAND2_X1 U8489 ( .A1(n6684), .A2(n6683), .ZN(n7804) );
  NAND2_X1 U8490 ( .A1(P2_U3893), .A2(n6444), .ZN(n8593) );
  AOI21_X1 U8491 ( .B1(n6685), .B2(n7804), .A(n8593), .ZN(n6711) );
  INV_X1 U8492 ( .A(n6686), .ZN(n6687) );
  INV_X1 U8493 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n10262) );
  AND2_X1 U8494 ( .A1(n6688), .A2(n8588), .ZN(n10161) );
  NAND2_X1 U8495 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n6763), .ZN(n6705) );
  AND2_X1 U8496 ( .A1(n6929), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6689) );
  NAND2_X1 U8497 ( .A1(n6632), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6690) );
  OAI21_X1 U8498 ( .B1(n6718), .B2(n6689), .A(n6690), .ZN(n10157) );
  OR2_X1 U8499 ( .A1(n10157), .A2(n6661), .ZN(n10158) );
  NAND2_X1 U8500 ( .A1(n10158), .A2(n6690), .ZN(n8427) );
  NAND2_X1 U8501 ( .A1(n6036), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6693) );
  NAND2_X1 U8502 ( .A1(n8426), .A2(n6693), .ZN(n6694) );
  NAND2_X1 U8503 ( .A1(n6974), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6696) );
  XNOR2_X1 U8504 ( .A(n7127), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n7109) );
  NAND2_X1 U8505 ( .A1(n6698), .A2(n7109), .ZN(n7114) );
  OR2_X1 U8506 ( .A1(n7127), .A2(n7464), .ZN(n6699) );
  NAND2_X1 U8507 ( .A1(n7114), .A2(n6699), .ZN(n6700) );
  NAND2_X1 U8508 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n6758), .ZN(n6702) );
  OAI21_X1 U8509 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n6758), .A(n6702), .ZN(
        n7332) );
  INV_X1 U8510 ( .A(n6703), .ZN(n6704) );
  OAI21_X1 U8511 ( .B1(n6763), .B2(P2_REG2_REG_10__SCAN_IN), .A(n6705), .ZN(
        n7698) );
  OAI21_X1 U8512 ( .B1(n6706), .B2(P2_REG2_REG_11__SCAN_IN), .A(n7798), .ZN(
        n6707) );
  NAND2_X1 U8513 ( .A1(n10161), .A2(n6707), .ZN(n6709) );
  AND2_X1 U8514 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7825) );
  INV_X1 U8515 ( .A(n7825), .ZN(n6708) );
  OAI211_X1 U8516 ( .C1(n8565), .C2(n10262), .A(n6709), .B(n6708), .ZN(n6710)
         );
  OR4_X1 U8517 ( .A1(n6713), .A2(n6712), .A3(n6711), .A4(n6710), .ZN(P2_U3193)
         );
  NAND2_X1 U8518 ( .A1(n6714), .A2(P1_U3086), .ZN(n9908) );
  NAND2_X1 U8519 ( .A1(n4507), .A2(P1_U3086), .ZN(n9906) );
  INV_X1 U8520 ( .A(n9906), .ZN(n9902) );
  AOI22_X1 U8521 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9426), .B1(n9902), .B2(
        P2_DATAO_REG_3__SCAN_IN), .ZN(n6715) );
  OAI21_X1 U8522 ( .B1(n6717), .B2(n9908), .A(n6715), .ZN(P1_U3352) );
  NOR2_X1 U8523 ( .A1(n7931), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8984) );
  INV_X1 U8524 ( .A(n8984), .ZN(n8243) );
  AND2_X1 U8525 ( .A1(n4506), .A2(P2_U3151), .ZN(n7635) );
  INV_X2 U8526 ( .A(n7635), .ZN(n8986) );
  OAI222_X1 U8527 ( .A1(n8243), .A2(n5143), .B1(n8986), .B2(n6717), .C1(
        P2_U3151), .C2(n6716), .ZN(P2_U3292) );
  OAI222_X1 U8528 ( .A1(n6718), .A2(P2_U3151), .B1(n8986), .B2(n6730), .C1(
        n8243), .C2(n5131), .ZN(P2_U3294) );
  OAI222_X1 U8529 ( .A1(n6036), .A2(P2_U3151), .B1(n8986), .B2(n6732), .C1(
        n8243), .C2(n6037), .ZN(P2_U3293) );
  OAI222_X1 U8530 ( .A1(n6974), .A2(P2_U3151), .B1(n8986), .B2(n6720), .C1(
        n8243), .C2(n6083), .ZN(P2_U3291) );
  INV_X1 U8531 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6719) );
  OAI222_X1 U8532 ( .A1(n9437), .A2(P1_U3086), .B1(n9908), .B2(n6720), .C1(
        n6719), .C2(n8152), .ZN(P1_U3351) );
  OAI222_X1 U8533 ( .A1(n8243), .A2(n6721), .B1(n8986), .B2(n6723), .C1(
        P2_U3151), .C2(n7101), .ZN(P2_U3290) );
  INV_X1 U8534 ( .A(n9454), .ZN(n9447) );
  INV_X1 U8535 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6722) );
  OAI222_X1 U8536 ( .A1(n9447), .A2(P1_U3086), .B1(n9908), .B2(n6723), .C1(
        n6722), .C2(n9906), .ZN(P1_U3350) );
  NAND2_X1 U8537 ( .A1(n6923), .A2(n6724), .ZN(n6744) );
  INV_X1 U8538 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6729) );
  INV_X1 U8539 ( .A(n6725), .ZN(n6915) );
  NOR3_X1 U8540 ( .A1(n6727), .A2(n6915), .A3(n6726), .ZN(n6728) );
  AOI21_X1 U8541 ( .B1(n6744), .B2(n6729), .A(n6728), .ZN(P2_U3376) );
  INV_X1 U8542 ( .A(n9908), .ZN(n7633) );
  INV_X1 U8543 ( .A(n7633), .ZN(n7771) );
  OAI222_X1 U8544 ( .A1(n6795), .A2(P1_U3086), .B1(n7771), .B2(n6730), .C1(
        n5043), .C2(n8152), .ZN(P1_U3354) );
  INV_X1 U8545 ( .A(n6796), .ZN(n9408) );
  INV_X1 U8546 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6731) );
  OAI222_X1 U8547 ( .A1(n9408), .A2(P1_U3086), .B1(n7771), .B2(n6732), .C1(
        n6731), .C2(n9906), .ZN(P1_U3353) );
  INV_X1 U8548 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6735) );
  INV_X1 U8549 ( .A(n7041), .ZN(n6733) );
  NAND2_X1 U8550 ( .A1(n6733), .A2(n6923), .ZN(n6734) );
  OAI21_X1 U8551 ( .B1(n6923), .B2(n6735), .A(n6734), .ZN(P2_U3377) );
  INV_X1 U8552 ( .A(n6736), .ZN(n6739) );
  AOI22_X1 U8553 ( .A1(n7127), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n8984), .ZN(n6737) );
  OAI21_X1 U8554 ( .B1(n6739), .B2(n8986), .A(n6737), .ZN(P2_U3289) );
  INV_X1 U8555 ( .A(n6806), .ZN(n9462) );
  INV_X1 U8556 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6738) );
  OAI222_X1 U8557 ( .A1(n9462), .A2(P1_U3086), .B1(n9908), .B2(n6739), .C1(
        n6738), .C2(n9906), .ZN(P1_U3349) );
  INV_X1 U8558 ( .A(n6823), .ZN(n6819) );
  INV_X1 U8559 ( .A(n6740), .ZN(n6742) );
  INV_X1 U8560 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10409) );
  OAI222_X1 U8561 ( .A1(n6819), .A2(P1_U3086), .B1(n7771), .B2(n6742), .C1(
        n10409), .C2(n9906), .ZN(P1_U3348) );
  INV_X1 U8562 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6743) );
  OAI222_X1 U8563 ( .A1(n8243), .A2(n6743), .B1(n8986), .B2(n6742), .C1(
        P2_U3151), .C2(n6741), .ZN(P2_U3288) );
  INV_X1 U8564 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n6745) );
  NOR2_X1 U8565 ( .A1(n6834), .A2(n6745), .ZN(P2_U3256) );
  INV_X1 U8566 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n6746) );
  NOR2_X1 U8567 ( .A1(n6834), .A2(n6746), .ZN(P2_U3253) );
  INV_X1 U8568 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n6747) );
  NOR2_X1 U8569 ( .A1(n6834), .A2(n6747), .ZN(P2_U3254) );
  INV_X1 U8570 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n6748) );
  NOR2_X1 U8571 ( .A1(n6834), .A2(n6748), .ZN(P2_U3252) );
  INV_X1 U8572 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n6749) );
  NOR2_X1 U8573 ( .A1(n6834), .A2(n6749), .ZN(P2_U3257) );
  INV_X1 U8574 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n6750) );
  NOR2_X1 U8575 ( .A1(n6834), .A2(n6750), .ZN(P2_U3248) );
  INV_X1 U8576 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n6751) );
  NOR2_X1 U8577 ( .A1(n6834), .A2(n6751), .ZN(P2_U3246) );
  INV_X1 U8578 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n6752) );
  NOR2_X1 U8579 ( .A1(n6834), .A2(n6752), .ZN(P2_U3247) );
  INV_X1 U8580 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n6753) );
  NOR2_X1 U8581 ( .A1(n6834), .A2(n6753), .ZN(P2_U3255) );
  INV_X1 U8582 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n6754) );
  NOR2_X1 U8583 ( .A1(n6834), .A2(n6754), .ZN(P2_U3250) );
  INV_X1 U8584 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n6755) );
  NOR2_X1 U8585 ( .A1(n6834), .A2(n6755), .ZN(P2_U3249) );
  INV_X1 U8586 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n6756) );
  NOR2_X1 U8587 ( .A1(n6834), .A2(n6756), .ZN(P2_U3251) );
  INV_X1 U8588 ( .A(n6757), .ZN(n6760) );
  OAI222_X1 U8589 ( .A1(n8243), .A2(n6759), .B1(n8986), .B2(n6760), .C1(
        P2_U3151), .C2(n6758), .ZN(P2_U3287) );
  INV_X1 U8590 ( .A(n6791), .ZN(n6859) );
  OAI222_X1 U8591 ( .A1(n6859), .A2(P1_U3086), .B1(n7771), .B2(n6760), .C1(
        n10655), .C2(n9906), .ZN(P1_U3347) );
  INV_X1 U8592 ( .A(n6761), .ZN(n6769) );
  INV_X1 U8593 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6762) );
  OAI222_X1 U8594 ( .A1(n8986), .A2(n6769), .B1(n6763), .B2(P2_U3151), .C1(
        n6762), .C2(n8243), .ZN(P2_U3285) );
  INV_X1 U8595 ( .A(n6764), .ZN(n6767) );
  OAI222_X1 U8596 ( .A1(n8243), .A2(n6766), .B1(n8986), .B2(n6767), .C1(
        P2_U3151), .C2(n6765), .ZN(P2_U3286) );
  INV_X1 U8597 ( .A(n6876), .ZN(n6790) );
  OAI222_X1 U8598 ( .A1(n8152), .A2(n6768), .B1(n7771), .B2(n6767), .C1(n6790), 
        .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U8599 ( .A(n7073), .ZN(n7081) );
  INV_X1 U8600 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10635) );
  OAI222_X1 U8601 ( .A1(P1_U3086), .A2(n7081), .B1(n7771), .B2(n6769), .C1(
        n10635), .C2(n9906), .ZN(P1_U3345) );
  INV_X1 U8602 ( .A(n6770), .ZN(n6832) );
  AOI22_X1 U8603 ( .A1(n7078), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9902), .ZN(n6771) );
  OAI21_X1 U8604 ( .B1(n6832), .B2(n9908), .A(n6771), .ZN(P1_U3344) );
  NOR2_X1 U8605 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(n6876), .ZN(n6772) );
  AOI21_X1 U8606 ( .B1(n6876), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6772), .ZN(
        n6780) );
  MUX2_X1 U8607 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n5330), .S(n6796), .Z(n9414)
         );
  MUX2_X1 U8608 ( .A(n5314), .B(P1_REG2_REG_1__SCAN_IN), .S(n6795), .Z(n9391)
         );
  AND2_X1 U8609 ( .A1(n10534), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9401) );
  NAND2_X1 U8610 ( .A1(n9391), .A2(n9401), .ZN(n9390) );
  INV_X1 U8611 ( .A(n6795), .ZN(n9392) );
  NAND2_X1 U8612 ( .A1(n9392), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6773) );
  NAND2_X1 U8613 ( .A1(n9390), .A2(n6773), .ZN(n9413) );
  NAND2_X1 U8614 ( .A1(n9414), .A2(n9413), .ZN(n9412) );
  NAND2_X1 U8615 ( .A1(n6796), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6774) );
  NAND2_X1 U8616 ( .A1(n9412), .A2(n6774), .ZN(n9419) );
  XNOR2_X1 U8617 ( .A(n9426), .B(n6775), .ZN(n9420) );
  NAND2_X1 U8618 ( .A1(n9419), .A2(n9420), .ZN(n9418) );
  NAND2_X1 U8619 ( .A1(n9426), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6776) );
  NAND2_X1 U8620 ( .A1(n9418), .A2(n6776), .ZN(n9435) );
  MUX2_X1 U8621 ( .A(n6777), .B(P1_REG2_REG_4__SCAN_IN), .S(n9437), .Z(n9436)
         );
  NAND2_X1 U8622 ( .A1(n9435), .A2(n9436), .ZN(n9434) );
  OAI21_X1 U8623 ( .B1(n9437), .B2(n6777), .A(n9434), .ZN(n9451) );
  MUX2_X1 U8624 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n7159), .S(n9454), .Z(n9452)
         );
  NAND2_X1 U8625 ( .A1(n9451), .A2(n9452), .ZN(n9450) );
  OAI21_X1 U8626 ( .B1(n9447), .B2(n7159), .A(n9450), .ZN(n9466) );
  MUX2_X1 U8627 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n7183), .S(n6806), .Z(n9467)
         );
  NAND2_X1 U8628 ( .A1(n9466), .A2(n9467), .ZN(n9465) );
  OAI21_X1 U8629 ( .B1(n9462), .B2(n7183), .A(n9465), .ZN(n6816) );
  MUX2_X1 U8630 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n7228), .S(n6823), .Z(n6817)
         );
  AND2_X1 U8631 ( .A1(n6816), .A2(n6817), .ZN(n6831) );
  AOI21_X1 U8632 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n6823), .A(n6831), .ZN(
        n6862) );
  MUX2_X1 U8633 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n5474), .S(n6791), .Z(n6778)
         );
  INV_X1 U8634 ( .A(n6778), .ZN(n6861) );
  NOR2_X1 U8635 ( .A1(n6862), .A2(n6861), .ZN(n6860) );
  AOI21_X1 U8636 ( .B1(n6791), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6860), .ZN(
        n6779) );
  NAND2_X1 U8637 ( .A1(n6780), .A2(n6779), .ZN(n6870) );
  OAI21_X1 U8638 ( .B1(n6780), .B2(n6779), .A(n6870), .ZN(n6814) );
  AND2_X1 U8639 ( .A1(n6781), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6788) );
  NAND2_X1 U8640 ( .A1(n6782), .A2(n9352), .ZN(n6784) );
  NAND2_X1 U8641 ( .A1(n6784), .A2(n6783), .ZN(n6787) );
  INV_X1 U8642 ( .A(n6787), .ZN(n6785) );
  NAND2_X1 U8643 ( .A1(n6788), .A2(n6785), .ZN(n9939) );
  NOR2_X1 U8644 ( .A1(n9399), .A2(n4519), .ZN(n9402) );
  INV_X1 U8645 ( .A(n9402), .ZN(n6786) );
  OR2_X1 U8646 ( .A1(n9939), .A2(n6786), .ZN(n9534) );
  NAND2_X1 U8647 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7454) );
  AND2_X1 U8648 ( .A1(n6788), .A2(n6787), .ZN(n9936) );
  NAND2_X1 U8649 ( .A1(n9936), .A2(P1_ADDR_REG_9__SCAN_IN), .ZN(n6789) );
  OAI211_X1 U8650 ( .C1(n9503), .C2(n6790), .A(n7454), .B(n6789), .ZN(n6813)
         );
  AOI22_X1 U8651 ( .A1(P1_REG1_REG_9__SCAN_IN), .A2(n6790), .B1(n6876), .B2(
        n5500), .ZN(n6809) );
  MUX2_X1 U8652 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n6792), .S(n6791), .Z(n6855)
         );
  INV_X1 U8653 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10133) );
  MUX2_X1 U8654 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6793), .S(n6796), .Z(n9411)
         );
  MUX2_X1 U8655 ( .A(n6794), .B(P1_REG1_REG_1__SCAN_IN), .S(n6795), .Z(n9388)
         );
  AND2_X1 U8656 ( .A1(n10534), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9389) );
  NAND2_X1 U8657 ( .A1(n9388), .A2(n9389), .ZN(n9387) );
  OAI21_X1 U8658 ( .B1(n6794), .B2(n6795), .A(n9387), .ZN(n9410) );
  NAND2_X1 U8659 ( .A1(n9411), .A2(n9410), .ZN(n9423) );
  NAND2_X1 U8660 ( .A1(n6796), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9422) );
  NAND2_X1 U8661 ( .A1(n9423), .A2(n9422), .ZN(n6799) );
  MUX2_X1 U8662 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6797), .S(n9426), .Z(n6798)
         );
  NAND2_X1 U8663 ( .A1(n6799), .A2(n6798), .ZN(n9440) );
  NAND2_X1 U8664 ( .A1(n9426), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9439) );
  NAND2_X1 U8665 ( .A1(n9440), .A2(n9439), .ZN(n6802) );
  INV_X1 U8666 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6800) );
  MUX2_X1 U8667 ( .A(n6800), .B(P1_REG1_REG_4__SCAN_IN), .S(n9437), .Z(n6801)
         );
  NAND2_X1 U8668 ( .A1(n6802), .A2(n6801), .ZN(n9457) );
  INV_X1 U8669 ( .A(n9457), .ZN(n6805) );
  NOR2_X1 U8670 ( .A1(n9437), .A2(n6800), .ZN(n9453) );
  INV_X1 U8671 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6803) );
  MUX2_X1 U8672 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6803), .S(n9454), .Z(n6804)
         );
  OAI21_X1 U8673 ( .B1(n6805), .B2(n9453), .A(n6804), .ZN(n9471) );
  NAND2_X1 U8674 ( .A1(n9454), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9470) );
  INV_X1 U8675 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10131) );
  MUX2_X1 U8676 ( .A(n10131), .B(P1_REG1_REG_6__SCAN_IN), .S(n6806), .Z(n9469)
         );
  AOI21_X1 U8677 ( .B1(n9471), .B2(n9470), .A(n9469), .ZN(n9468) );
  NOR2_X1 U8678 ( .A1(n9462), .A2(n10131), .ZN(n6822) );
  MUX2_X1 U8679 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n10133), .S(n6823), .Z(n6807)
         );
  OAI21_X1 U8680 ( .B1(n9468), .B2(n6822), .A(n6807), .ZN(n6826) );
  OAI21_X1 U8681 ( .B1(n10133), .B2(n6819), .A(n6826), .ZN(n6854) );
  NAND2_X1 U8682 ( .A1(n6855), .A2(n6854), .ZN(n6853) );
  OAI21_X1 U8683 ( .B1(n6859), .B2(n6792), .A(n6853), .ZN(n6808) );
  NOR2_X1 U8684 ( .A1(n6809), .A2(n6808), .ZN(n6877) );
  AOI21_X1 U8685 ( .B1(n6809), .B2(n6808), .A(n6877), .ZN(n6811) );
  INV_X1 U8686 ( .A(n4519), .ZN(n6810) );
  NOR2_X1 U8687 ( .A1(n6811), .A2(n9528), .ZN(n6812) );
  AOI211_X1 U8688 ( .C1(n6814), .C2(n9507), .A(n6813), .B(n6812), .ZN(n6815)
         );
  INV_X1 U8689 ( .A(n6815), .ZN(P1_U3252) );
  OAI21_X1 U8690 ( .B1(n6817), .B2(n6816), .A(n9507), .ZN(n6830) );
  NOR2_X1 U8691 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6818), .ZN(n6821) );
  NOR2_X1 U8692 ( .A1(n9503), .A2(n6819), .ZN(n6820) );
  AOI211_X1 U8693 ( .C1(n9936), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n6821), .B(
        n6820), .ZN(n6829) );
  INV_X1 U8694 ( .A(n6822), .ZN(n6825) );
  MUX2_X1 U8695 ( .A(n10133), .B(P1_REG1_REG_7__SCAN_IN), .S(n6823), .Z(n6824)
         );
  NAND2_X1 U8696 ( .A1(n6825), .A2(n6824), .ZN(n6827) );
  OAI211_X1 U8697 ( .C1(n9468), .C2(n6827), .A(n9531), .B(n6826), .ZN(n6828)
         );
  OAI211_X1 U8698 ( .C1(n6831), .C2(n6830), .A(n6829), .B(n6828), .ZN(P1_U3250) );
  OAI222_X1 U8699 ( .A1(n8243), .A2(n6833), .B1(n8986), .B2(n6832), .C1(
        P2_U3151), .C2(n7802), .ZN(P2_U3284) );
  INV_X1 U8700 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n6835) );
  NOR2_X1 U8701 ( .A1(n6834), .A2(n6835), .ZN(P2_U3262) );
  INV_X1 U8702 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n6836) );
  NOR2_X1 U8703 ( .A1(n6834), .A2(n6836), .ZN(P2_U3234) );
  INV_X1 U8704 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n6837) );
  NOR2_X1 U8705 ( .A1(n6834), .A2(n6837), .ZN(P2_U3263) );
  INV_X1 U8706 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n6838) );
  NOR2_X1 U8707 ( .A1(n6834), .A2(n6838), .ZN(P2_U3258) );
  INV_X1 U8708 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n6839) );
  NOR2_X1 U8709 ( .A1(n6834), .A2(n6839), .ZN(P2_U3261) );
  INV_X1 U8710 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n6840) );
  NOR2_X1 U8711 ( .A1(n6834), .A2(n6840), .ZN(P2_U3260) );
  INV_X1 U8712 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n6841) );
  NOR2_X1 U8713 ( .A1(n6834), .A2(n6841), .ZN(P2_U3259) );
  INV_X1 U8714 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n6842) );
  NOR2_X1 U8715 ( .A1(n6834), .A2(n6842), .ZN(P2_U3243) );
  INV_X1 U8716 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n6843) );
  NOR2_X1 U8717 ( .A1(n6834), .A2(n6843), .ZN(P2_U3242) );
  INV_X1 U8718 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n6844) );
  NOR2_X1 U8719 ( .A1(n6834), .A2(n6844), .ZN(P2_U3241) );
  INV_X1 U8720 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n6845) );
  NOR2_X1 U8721 ( .A1(n6834), .A2(n6845), .ZN(P2_U3240) );
  INV_X1 U8722 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n6846) );
  NOR2_X1 U8723 ( .A1(n6834), .A2(n6846), .ZN(P2_U3239) );
  INV_X1 U8724 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n6847) );
  NOR2_X1 U8725 ( .A1(n6834), .A2(n6847), .ZN(P2_U3238) );
  INV_X1 U8726 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n6848) );
  NOR2_X1 U8727 ( .A1(n6834), .A2(n6848), .ZN(P2_U3237) );
  INV_X1 U8728 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n6849) );
  NOR2_X1 U8729 ( .A1(n6834), .A2(n6849), .ZN(P2_U3236) );
  INV_X1 U8730 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n6850) );
  NOR2_X1 U8731 ( .A1(n6834), .A2(n6850), .ZN(P2_U3235) );
  INV_X1 U8732 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n6851) );
  NOR2_X1 U8733 ( .A1(n6834), .A2(n6851), .ZN(P2_U3245) );
  INV_X1 U8734 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n6852) );
  NOR2_X1 U8735 ( .A1(n6834), .A2(n6852), .ZN(P2_U3244) );
  OAI211_X1 U8736 ( .C1(n6855), .C2(n6854), .A(n9531), .B(n6853), .ZN(n6858)
         );
  AND2_X1 U8737 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6856) );
  AOI21_X1 U8738 ( .B1(n9936), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n6856), .ZN(
        n6857) );
  OAI211_X1 U8739 ( .C1(n9503), .C2(n6859), .A(n6858), .B(n6857), .ZN(n6864)
         );
  AOI211_X1 U8740 ( .C1(n6862), .C2(n6861), .A(n6860), .B(n9534), .ZN(n6863)
         );
  OR2_X1 U8741 ( .A1(n6864), .A2(n6863), .ZN(P1_U3251) );
  INV_X1 U8742 ( .A(n6865), .ZN(n6867) );
  INV_X1 U8743 ( .A(n7813), .ZN(n8447) );
  INV_X1 U8744 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6866) );
  OAI222_X1 U8745 ( .A1(n8986), .A2(n6867), .B1(n8447), .B2(P2_U3151), .C1(
        n6866), .C2(n8243), .ZN(P2_U3283) );
  INV_X1 U8746 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10645) );
  INV_X1 U8747 ( .A(n7373), .ZN(n7364) );
  OAI222_X1 U8748 ( .A1(n8152), .A2(n10645), .B1(n7771), .B2(n6867), .C1(
        P1_U3086), .C2(n7364), .ZN(P1_U3343) );
  CLKBUF_X2 U8749 ( .A(P1_U3973), .Z(n9385) );
  NOR2_X1 U8750 ( .A1(n9936), .A2(n9385), .ZN(P1_U3085) );
  AND2_X1 U8751 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6868) );
  AOI21_X1 U8752 ( .B1(n9936), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n6868), .ZN(
        n6869) );
  INV_X1 U8753 ( .A(n6869), .ZN(n6875) );
  OAI21_X1 U8754 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n6876), .A(n6870), .ZN(
        n6873) );
  MUX2_X1 U8755 ( .A(n6871), .B(P1_REG2_REG_10__SCAN_IN), .S(n7073), .Z(n6872)
         );
  NOR2_X1 U8756 ( .A1(n6872), .A2(n6873), .ZN(n7072) );
  AOI211_X1 U8757 ( .C1(n6873), .C2(n6872), .A(n7072), .B(n9534), .ZN(n6874)
         );
  AOI211_X1 U8758 ( .C1(n9530), .C2(n7073), .A(n6875), .B(n6874), .ZN(n6883)
         );
  NOR2_X1 U8759 ( .A1(P1_REG1_REG_9__SCAN_IN), .A2(n6876), .ZN(n6878) );
  NOR2_X1 U8760 ( .A1(n6878), .A2(n6877), .ZN(n6881) );
  MUX2_X1 U8761 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6879), .S(n7073), .Z(n6880)
         );
  NAND2_X1 U8762 ( .A1(n6880), .A2(n6881), .ZN(n7080) );
  OAI211_X1 U8763 ( .C1(n6881), .C2(n6880), .A(n9531), .B(n7080), .ZN(n6882)
         );
  NAND2_X1 U8764 ( .A1(n6883), .A2(n6882), .ZN(P1_U3253) );
  INV_X1 U8765 ( .A(n6884), .ZN(n6887) );
  AOI22_X1 U8766 ( .A1(n9496), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9902), .ZN(n6885) );
  OAI21_X1 U8767 ( .B1(n6887), .B2(n7771), .A(n6885), .ZN(P1_U3342) );
  AOI22_X1 U8768 ( .A1(n8473), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n8984), .ZN(n6886) );
  OAI21_X1 U8769 ( .B1(n6887), .B2(n8986), .A(n6886), .ZN(P2_U3282) );
  XOR2_X1 U8770 ( .A(n6888), .B(n6889), .Z(n6893) );
  NOR2_X1 U8771 ( .A1(n6890), .A2(P1_U3086), .ZN(n6998) );
  AOI22_X1 U8772 ( .A1(n9103), .A2(n9384), .B1(n6984), .B2(n9101), .ZN(n9994)
         );
  OAI22_X1 U8773 ( .A1(n6998), .A2(n9405), .B1(n9914), .B2(n9994), .ZN(n6891)
         );
  AOI21_X1 U8774 ( .B1(n10005), .B2(n9924), .A(n6891), .ZN(n6892) );
  OAI21_X1 U8775 ( .B1(n6893), .B2(n9919), .A(n6892), .ZN(P1_U3237) );
  NAND2_X1 U8776 ( .A1(n9385), .A2(n4512), .ZN(n6894) );
  OAI21_X1 U8777 ( .B1(n9385), .B2(n6037), .A(n6894), .ZN(P1_U3556) );
  NAND2_X1 U8778 ( .A1(n9385), .A2(n6895), .ZN(n6896) );
  OAI21_X1 U8779 ( .B1(n9385), .B2(n6083), .A(n6896), .ZN(P1_U3558) );
  NAND2_X1 U8780 ( .A1(n9385), .A2(n6984), .ZN(n6897) );
  OAI21_X1 U8781 ( .B1(n9385), .B2(n5131), .A(n6897), .ZN(P1_U3555) );
  NAND2_X1 U8782 ( .A1(n9024), .A2(n9385), .ZN(n6898) );
  OAI21_X1 U8783 ( .B1(n6279), .B2(n9385), .A(n6898), .ZN(P1_U3574) );
  INV_X1 U8784 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6904) );
  NAND2_X1 U8785 ( .A1(n5792), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6902) );
  INV_X1 U8786 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n8164) );
  OR2_X1 U8787 ( .A1(n5360), .A2(n8164), .ZN(n6901) );
  INV_X1 U8788 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9543) );
  OR2_X1 U8789 ( .A1(n6899), .A2(n9543), .ZN(n6900) );
  AND3_X1 U8790 ( .A1(n6902), .A2(n6901), .A3(n6900), .ZN(n9225) );
  INV_X1 U8791 ( .A(n9225), .ZN(n9286) );
  NAND2_X1 U8792 ( .A1(n9286), .A2(n9385), .ZN(n6903) );
  OAI21_X1 U8793 ( .B1(n9385), .B2(n6904), .A(n6903), .ZN(P1_U3585) );
  NAND2_X1 U8794 ( .A1(n6906), .A2(n6905), .ZN(n6908) );
  OAI211_X1 U8795 ( .C1(n6911), .C2(n6918), .A(n6908), .B(n6907), .ZN(n6909)
         );
  NAND2_X1 U8796 ( .A1(n6909), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6914) );
  INV_X1 U8797 ( .A(n6923), .ZN(n6910) );
  NOR2_X1 U8798 ( .A1(n7048), .A2(n6910), .ZN(n8143) );
  INV_X1 U8799 ( .A(n6911), .ZN(n6912) );
  NAND2_X1 U8800 ( .A1(n8143), .A2(n6912), .ZN(n6913) );
  NAND2_X1 U8801 ( .A1(n6914), .A2(n6913), .ZN(n7133) );
  NOR2_X1 U8802 ( .A1(n7133), .A2(n6915), .ZN(n7063) );
  NAND2_X1 U8803 ( .A1(n6381), .A2(n7057), .ZN(n7981) );
  NAND2_X1 U8804 ( .A1(n7311), .A2(n7981), .ZN(n7946) );
  INV_X1 U8805 ( .A(n6916), .ZN(n6917) );
  NAND2_X1 U8806 ( .A1(n6922), .A2(n6917), .ZN(n6921) );
  INV_X1 U8807 ( .A(n6918), .ZN(n6919) );
  NAND2_X1 U8808 ( .A1(n7025), .A2(n6919), .ZN(n6920) );
  NAND2_X1 U8809 ( .A1(n6922), .A2(n10213), .ZN(n6925) );
  INV_X1 U8810 ( .A(n8324), .ZN(n8405) );
  NOR2_X1 U8811 ( .A1(n7048), .A2(n7023), .ZN(n6926) );
  OAI22_X1 U8812 ( .A1(n8405), .A2(n7057), .B1(n6055), .B2(n8398), .ZN(n6927)
         );
  AOI21_X1 U8813 ( .B1(n7946), .B2(n8381), .A(n6927), .ZN(n6928) );
  OAI21_X1 U8814 ( .B1(n7063), .B2(n7050), .A(n6928), .ZN(P2_U3172) );
  INV_X1 U8815 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6936) );
  XNOR2_X1 U8816 ( .A(n6930), .B(n6929), .ZN(n6931) );
  AOI21_X1 U8817 ( .B1(n6932), .B2(n8593), .A(n6931), .ZN(n6933) );
  AOI21_X1 U8818 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .A(n6933), .ZN(
        n6935) );
  OAI211_X1 U8819 ( .C1(n8565), .C2(n6936), .A(n6935), .B(n6934), .ZN(P2_U3182) );
  AOI21_X1 U8820 ( .B1(n6939), .B2(n6938), .A(n6937), .ZN(n6951) );
  INV_X1 U8821 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6943) );
  INV_X1 U8822 ( .A(n6958), .ZN(n6940) );
  AOI21_X1 U8823 ( .B1(n6057), .B2(n6941), .A(n6940), .ZN(n6942) );
  OAI22_X1 U8824 ( .A1(n8565), .A2(n6943), .B1(n10152), .B2(n6942), .ZN(n6949)
         );
  INV_X1 U8825 ( .A(n6966), .ZN(n6944) );
  AOI21_X1 U8826 ( .B1(n6058), .B2(n6945), .A(n6944), .ZN(n6947) );
  NOR2_X1 U8827 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10634), .ZN(n7135) );
  INV_X1 U8828 ( .A(n7135), .ZN(n6946) );
  OAI21_X1 U8829 ( .B1(n8571), .B2(n6947), .A(n6946), .ZN(n6948) );
  AOI211_X1 U8830 ( .C1(n4895), .C2(n10155), .A(n6949), .B(n6948), .ZN(n6950)
         );
  OAI21_X1 U8831 ( .B1(n6951), .B2(n8593), .A(n6950), .ZN(P2_U3185) );
  OAI211_X1 U8832 ( .C1(n6954), .C2(n6953), .A(n6952), .B(n10146), .ZN(n6973)
         );
  INV_X1 U8833 ( .A(n8565), .ZN(n10145) );
  INV_X1 U8834 ( .A(n6955), .ZN(n6957) );
  NAND3_X1 U8835 ( .A1(n6958), .A2(n6957), .A3(n6956), .ZN(n6959) );
  AOI21_X1 U8836 ( .B1(n6960), .B2(n6959), .A(n10152), .ZN(n6971) );
  INV_X1 U8837 ( .A(n6961), .ZN(n6963) );
  NOR2_X1 U8838 ( .A1(n6963), .A2(n6962), .ZN(n6967) );
  INV_X1 U8839 ( .A(n6964), .ZN(n6965) );
  AOI21_X1 U8840 ( .B1(n6967), .B2(n6966), .A(n6965), .ZN(n6969) );
  NOR2_X1 U8841 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10440), .ZN(n7173) );
  INV_X1 U8842 ( .A(n7173), .ZN(n6968) );
  OAI21_X1 U8843 ( .B1(n8571), .B2(n6969), .A(n6968), .ZN(n6970) );
  AOI211_X1 U8844 ( .C1(n10145), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n6971), .B(
        n6970), .ZN(n6972) );
  OAI211_X1 U8845 ( .C1(n8598), .C2(n6974), .A(n6973), .B(n6972), .ZN(P2_U3186) );
  OAI21_X1 U8846 ( .B1(n8813), .B2(n10196), .A(n7946), .ZN(n6975) );
  NAND2_X1 U8847 ( .A1(n8420), .A2(n8810), .ZN(n7049) );
  OAI211_X1 U8848 ( .C1(n10215), .C2(n7057), .A(n6975), .B(n7049), .ZN(n6988)
         );
  NAND2_X1 U8849 ( .A1(n6988), .A2(n10233), .ZN(n6976) );
  OAI21_X1 U8850 ( .B1(n10233), .B2(n6662), .A(n6976), .ZN(P2_U3459) );
  INV_X1 U8851 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n10568) );
  NAND2_X1 U8852 ( .A1(n8745), .A2(P2_U3893), .ZN(n6977) );
  OAI21_X1 U8853 ( .B1(P2_U3893), .B2(n10568), .A(n6977), .ZN(P2_U3511) );
  INV_X1 U8854 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10638) );
  INV_X1 U8855 ( .A(n6978), .ZN(n6979) );
  INV_X1 U8856 ( .A(n7377), .ZN(n9514) );
  OAI222_X1 U8857 ( .A1(n8152), .A2(n10638), .B1(n7771), .B2(n6979), .C1(n9514), .C2(P1_U3086), .ZN(P1_U3341) );
  INV_X1 U8858 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6980) );
  INV_X1 U8859 ( .A(n8482), .ZN(n8492) );
  OAI222_X1 U8860 ( .A1(n8243), .A2(n6980), .B1(n8986), .B2(n6979), .C1(
        P2_U3151), .C2(n8492), .ZN(P2_U3281) );
  OAI21_X1 U8861 ( .B1(n6983), .B2(n6982), .A(n6981), .ZN(n9398) );
  NAND2_X1 U8862 ( .A1(n6984), .A2(n9103), .ZN(n7326) );
  OAI22_X1 U8863 ( .A1(n6998), .A2(n6985), .B1(n9914), .B2(n7326), .ZN(n6986)
         );
  AOI21_X1 U8864 ( .B1(n10020), .B2(n9924), .A(n6986), .ZN(n6987) );
  OAI21_X1 U8865 ( .B1(n9919), .B2(n9398), .A(n6987), .ZN(P1_U3232) );
  INV_X1 U8866 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6990) );
  NAND2_X1 U8867 ( .A1(n6988), .A2(n10221), .ZN(n6989) );
  OAI21_X1 U8868 ( .B1(n6990), .B2(n10221), .A(n6989), .ZN(P2_U3390) );
  NAND2_X1 U8869 ( .A1(n6992), .A2(n6991), .ZN(n6993) );
  XOR2_X1 U8870 ( .A(n6994), .B(n6993), .Z(n7001) );
  NAND2_X1 U8871 ( .A1(n9386), .A2(n9101), .ZN(n6996) );
  NAND2_X1 U8872 ( .A1(n4512), .A2(n9103), .ZN(n6995) );
  AND2_X1 U8873 ( .A1(n6996), .A2(n6995), .ZN(n10015) );
  OAI22_X1 U8874 ( .A1(n6998), .A2(n6997), .B1(n9914), .B2(n10015), .ZN(n6999)
         );
  AOI21_X1 U8875 ( .B1(n10021), .B2(n9924), .A(n6999), .ZN(n7000) );
  OAI21_X1 U8876 ( .B1(n7001), .B2(n9919), .A(n7000), .ZN(P1_U3222) );
  INV_X1 U8877 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7006) );
  INV_X1 U8878 ( .A(n7002), .ZN(n10013) );
  NAND2_X1 U8879 ( .A1(n9386), .A2(n7004), .ZN(n9297) );
  NAND2_X1 U8880 ( .A1(n10013), .A2(n9297), .ZN(n9229) );
  OAI21_X1 U8881 ( .B1(n10112), .B2(n9996), .A(n9229), .ZN(n7003) );
  OAI211_X1 U8882 ( .C1(n7324), .C2(n7004), .A(n7003), .B(n7326), .ZN(n9838)
         );
  NAND2_X1 U8883 ( .A1(n10125), .A2(n9838), .ZN(n7005) );
  OAI21_X1 U8884 ( .B1(n10125), .B2(n7006), .A(n7005), .ZN(P1_U3453) );
  XOR2_X1 U8885 ( .A(n7008), .B(n7007), .Z(n7012) );
  OAI22_X1 U8886 ( .A1(n7009), .A2(n9089), .B1(n7157), .B2(n9091), .ZN(n7285)
         );
  AOI22_X1 U8887 ( .A1(n9117), .A2(n7285), .B1(n9924), .B2(n7290), .ZN(n7011)
         );
  MUX2_X1 U8888 ( .A(n9926), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n7010) );
  OAI211_X1 U8889 ( .C1(n7012), .C2(n9919), .A(n7011), .B(n7010), .ZN(P1_U3218) );
  OR2_X1 U8890 ( .A1(n7169), .A2(n7021), .ZN(n7022) );
  NAND2_X1 U8891 ( .A1(n7022), .A2(n7311), .ZN(n7061) );
  XOR2_X1 U8892 ( .A(n7062), .B(n7061), .Z(n7031) );
  INV_X1 U8893 ( .A(n6381), .ZN(n7027) );
  INV_X1 U8894 ( .A(n7023), .ZN(n7024) );
  NOR2_X1 U8895 ( .A1(n7048), .A2(n7024), .ZN(n7026) );
  NAND2_X1 U8896 ( .A1(n7026), .A2(n7025), .ZN(n8384) );
  OAI22_X1 U8897 ( .A1(n8398), .A2(n4796), .B1(n7027), .B2(n8384), .ZN(n7029)
         );
  NOR2_X1 U8898 ( .A1(n7063), .A2(n7319), .ZN(n7028) );
  AOI211_X1 U8899 ( .C1(n7020), .C2(n8324), .A(n7029), .B(n7028), .ZN(n7030)
         );
  OAI21_X1 U8900 ( .B1(n8393), .B2(n7031), .A(n7030), .ZN(P2_U3162) );
  AOI21_X1 U8901 ( .B1(n7032), .B2(n7033), .A(n9919), .ZN(n7035) );
  NAND2_X1 U8902 ( .A1(n7035), .A2(n7034), .ZN(n7039) );
  OAI22_X1 U8903 ( .A1(n7036), .A2(n9089), .B1(n7181), .B2(n9091), .ZN(n9975)
         );
  AND2_X1 U8904 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9431) );
  INV_X1 U8905 ( .A(n9924), .ZN(n9070) );
  OAI22_X1 U8906 ( .A1(n9070), .A2(n10063), .B1(n9977), .B2(n9926), .ZN(n7037)
         );
  AOI211_X1 U8907 ( .C1(n9117), .C2(n9975), .A(n9431), .B(n7037), .ZN(n7038)
         );
  NAND2_X1 U8908 ( .A1(n7039), .A2(n7038), .ZN(P1_U3230) );
  INV_X1 U8909 ( .A(n7040), .ZN(n7043) );
  NAND2_X1 U8910 ( .A1(n7044), .A2(n7041), .ZN(n7042) );
  OAI21_X1 U8911 ( .B1(n7044), .B2(n7043), .A(n7042), .ZN(n7045) );
  INV_X1 U8912 ( .A(n7045), .ZN(n7046) );
  NAND2_X1 U8913 ( .A1(n7047), .A2(n7046), .ZN(n7053) );
  AND2_X1 U8914 ( .A1(n7048), .A2(n10215), .ZN(n7052) );
  OAI21_X1 U8915 ( .B1(n10169), .B2(n7050), .A(n7049), .ZN(n7051) );
  AOI21_X1 U8916 ( .B1(n7052), .B2(n7946), .A(n7051), .ZN(n7054) );
  MUX2_X1 U8917 ( .A(n7055), .B(n7054), .S(n10174), .Z(n7056) );
  OAI21_X1 U8918 ( .B1(n10171), .B2(n7057), .A(n7056), .ZN(P2_U3233) );
  INV_X1 U8919 ( .A(n7058), .ZN(n7059) );
  NOR2_X1 U8920 ( .A1(n7059), .A2(n8420), .ZN(n7060) );
  AOI21_X1 U8921 ( .B1(n7062), .B2(n7061), .A(n7060), .ZN(n7141) );
  XNOR2_X1 U8922 ( .A(n7306), .B(n7169), .ZN(n7138) );
  XOR2_X1 U8923 ( .A(n8419), .B(n7138), .Z(n7140) );
  XOR2_X1 U8924 ( .A(n7141), .B(n7140), .Z(n7067) );
  OAI22_X1 U8925 ( .A1(n8398), .A2(n7207), .B1(n6055), .B2(n8384), .ZN(n7065)
         );
  NOR2_X1 U8926 ( .A1(n7063), .A2(n6026), .ZN(n7064) );
  AOI211_X1 U8927 ( .C1(n7306), .C2(n8324), .A(n7065), .B(n7064), .ZN(n7066)
         );
  OAI21_X1 U8928 ( .B1(n7067), .B2(n8393), .A(n7066), .ZN(P2_U3177) );
  INV_X1 U8929 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7069) );
  INV_X1 U8930 ( .A(n7068), .ZN(n7070) );
  INV_X1 U8931 ( .A(n8519), .ZN(n8509) );
  OAI222_X1 U8932 ( .A1(n8243), .A2(n7069), .B1(n8986), .B2(n7070), .C1(
        P2_U3151), .C2(n8509), .ZN(P2_U3280) );
  INV_X1 U8933 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10463) );
  INV_X1 U8934 ( .A(n7501), .ZN(n7379) );
  OAI222_X1 U8935 ( .A1(n9906), .A2(n10463), .B1(n7771), .B2(n7070), .C1(n7379), .C2(P1_U3086), .ZN(P1_U3340) );
  MUX2_X1 U8936 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n7071), .S(n7373), .Z(n7076)
         );
  AOI21_X1 U8937 ( .B1(n7073), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7072), .ZN(
        n9485) );
  NAND2_X1 U8938 ( .A1(n7078), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7074) );
  OAI21_X1 U8939 ( .B1(n7078), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7074), .ZN(
        n9484) );
  NOR2_X1 U8940 ( .A1(n9485), .A2(n9484), .ZN(n9483) );
  AOI21_X1 U8941 ( .B1(n7078), .B2(P1_REG2_REG_11__SCAN_IN), .A(n9483), .ZN(
        n7075) );
  NAND2_X1 U8942 ( .A1(n7076), .A2(n7075), .ZN(n7372) );
  OAI21_X1 U8943 ( .B1(n7076), .B2(n7075), .A(n7372), .ZN(n7086) );
  MUX2_X1 U8944 ( .A(n7077), .B(P1_REG1_REG_12__SCAN_IN), .S(n7373), .Z(n7083)
         );
  INV_X1 U8945 ( .A(n7078), .ZN(n9477) );
  MUX2_X1 U8946 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n7079), .S(n7078), .Z(n9481)
         );
  OAI21_X1 U8947 ( .B1(n7081), .B2(n6879), .A(n7080), .ZN(n9482) );
  NAND2_X1 U8948 ( .A1(n9481), .A2(n9482), .ZN(n9480) );
  OAI21_X1 U8949 ( .B1(n9477), .B2(n7079), .A(n9480), .ZN(n7082) );
  NOR2_X1 U8950 ( .A1(n7082), .A2(n7083), .ZN(n7363) );
  AOI21_X1 U8951 ( .B1(n7083), .B2(n7082), .A(n7363), .ZN(n7084) );
  NOR2_X1 U8952 ( .A1(n9528), .A2(n7084), .ZN(n7085) );
  AOI21_X1 U8953 ( .B1(n9507), .B2(n7086), .A(n7085), .ZN(n7088) );
  AND2_X1 U8954 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9911) );
  AOI21_X1 U8955 ( .B1(n9936), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n9911), .ZN(
        n7087) );
  OAI211_X1 U8956 ( .C1(n7364), .C2(n9503), .A(n7088), .B(n7087), .ZN(P1_U3255) );
  OAI211_X1 U8957 ( .C1(n7091), .C2(n7090), .A(n7089), .B(n10146), .ZN(n7100)
         );
  AOI21_X1 U8958 ( .B1(n7118), .B2(n7092), .A(n10152), .ZN(n7098) );
  INV_X1 U8959 ( .A(n7112), .ZN(n7093) );
  AOI21_X1 U8960 ( .B1(n7436), .B2(n7094), .A(n7093), .ZN(n7096) );
  NOR2_X1 U8961 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6086), .ZN(n7240) );
  INV_X1 U8962 ( .A(n7240), .ZN(n7095) );
  OAI21_X1 U8963 ( .B1(n8571), .B2(n7096), .A(n7095), .ZN(n7097) );
  AOI211_X1 U8964 ( .C1(n10145), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n7098), .B(
        n7097), .ZN(n7099) );
  OAI211_X1 U8965 ( .C1(n8598), .C2(n7101), .A(n7100), .B(n7099), .ZN(P2_U3187) );
  INV_X1 U8966 ( .A(n7102), .ZN(n7104) );
  AOI22_X1 U8967 ( .A1(n7593), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n9902), .ZN(n7103) );
  OAI21_X1 U8968 ( .B1(n7104), .B2(n9908), .A(n7103), .ZN(P1_U3339) );
  INV_X1 U8969 ( .A(n8527), .ZN(n8537) );
  OAI222_X1 U8970 ( .A1(n8243), .A2(n7105), .B1(P2_U3151), .B2(n8537), .C1(
        n7104), .C2(n8986), .ZN(P2_U3279) );
  AOI21_X1 U8971 ( .B1(n7108), .B2(n7107), .A(n7106), .ZN(n7129) );
  INV_X1 U8972 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7125) );
  INV_X1 U8973 ( .A(n7109), .ZN(n7111) );
  NAND3_X1 U8974 ( .A1(n7112), .A2(n7111), .A3(n7110), .ZN(n7113) );
  AOI21_X1 U8975 ( .B1(n7114), .B2(n7113), .A(n8571), .ZN(n7122) );
  INV_X1 U8976 ( .A(n7115), .ZN(n7117) );
  NAND3_X1 U8977 ( .A1(n7118), .A2(n7117), .A3(n7116), .ZN(n7119) );
  AOI21_X1 U8978 ( .B1(n7120), .B2(n7119), .A(n10152), .ZN(n7121) );
  NOR2_X1 U8979 ( .A1(n7122), .A2(n7121), .ZN(n7124) );
  INV_X1 U8980 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10398) );
  NOR2_X1 U8981 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10398), .ZN(n7277) );
  INV_X1 U8982 ( .A(n7277), .ZN(n7123) );
  OAI211_X1 U8983 ( .C1(n8565), .C2(n7125), .A(n7124), .B(n7123), .ZN(n7126)
         );
  AOI21_X1 U8984 ( .B1(n7127), .B2(n10155), .A(n7126), .ZN(n7128) );
  OAI21_X1 U8985 ( .B1(n7129), .B2(n8593), .A(n7128), .ZN(P2_U3188) );
  INV_X1 U8986 ( .A(n7130), .ZN(n7166) );
  AOI22_X1 U8987 ( .A1(n8567), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n8984), .ZN(n7131) );
  OAI21_X1 U8988 ( .B1(n7166), .B2(n8986), .A(n7131), .ZN(P2_U3278) );
  AND2_X1 U8989 ( .A1(n7132), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7637) );
  NOR2_X1 U8990 ( .A1(n4796), .A2(n8384), .ZN(n7134) );
  AOI211_X1 U8991 ( .C1(n8337), .C2(n8417), .A(n7135), .B(n7134), .ZN(n7136)
         );
  OAI21_X1 U8992 ( .B1(n10186), .B2(n8405), .A(n7136), .ZN(n7145) );
  XNOR2_X1 U8993 ( .A(n8235), .B(n7137), .ZN(n7168) );
  XNOR2_X1 U8994 ( .A(n7168), .B(n8418), .ZN(n7143) );
  INV_X1 U8995 ( .A(n7138), .ZN(n7139) );
  OAI22_X1 U8996 ( .A1(n7141), .A2(n7140), .B1(n7139), .B2(n8419), .ZN(n7142)
         );
  NOR2_X1 U8997 ( .A1(n7142), .A2(n7143), .ZN(n7167) );
  AOI211_X1 U8998 ( .C1(n7143), .C2(n7142), .A(n8393), .B(n7167), .ZN(n7144)
         );
  AOI211_X1 U8999 ( .C1(n10634), .C2(n8389), .A(n7145), .B(n7144), .ZN(n7146)
         );
  INV_X1 U9000 ( .A(n7146), .ZN(P2_U3158) );
  INV_X1 U9001 ( .A(n7147), .ZN(n7148) );
  NOR2_X1 U9002 ( .A1(n7149), .A2(n7148), .ZN(n7150) );
  NAND2_X1 U9003 ( .A1(n10036), .A2(n7150), .ZN(n7151) );
  NAND2_X1 U9004 ( .A1(n5285), .A2(n7152), .ZN(n7153) );
  OR2_X1 U9005 ( .A1(n10033), .A2(n7153), .ZN(n9953) );
  OR2_X1 U9006 ( .A1(n10033), .A2(n10009), .ZN(n7154) );
  XOR2_X1 U9007 ( .A(n9232), .B(n7155), .Z(n10070) );
  XOR2_X1 U9008 ( .A(n9232), .B(n7156), .Z(n7158) );
  OAI22_X1 U9009 ( .A1(n9132), .A2(n9091), .B1(n7157), .B2(n9089), .ZN(n7217)
         );
  AOI21_X1 U9010 ( .B1(n7158), .B2(n9996), .A(n7217), .ZN(n10069) );
  MUX2_X1 U9011 ( .A(n7159), .B(n10069), .S(n9734), .Z(n7164) );
  INV_X1 U9012 ( .A(n9987), .ZN(n7160) );
  AOI211_X1 U9013 ( .C1(n10067), .C2(n7160), .A(n10003), .B(n7184), .ZN(n10066) );
  OAI22_X1 U9014 ( .A1(n10029), .A2(n9139), .B1(n7218), .B2(n9699), .ZN(n7162)
         );
  AOI21_X1 U9015 ( .B1(n10066), .B2(n10025), .A(n7162), .ZN(n7163) );
  OAI211_X1 U9016 ( .C1(n9737), .C2(n10070), .A(n7164), .B(n7163), .ZN(
        P1_U3288) );
  INV_X1 U9017 ( .A(n7752), .ZN(n7165) );
  OAI222_X1 U9018 ( .A1(n8152), .A2(n10561), .B1(n7771), .B2(n7166), .C1(n7165), .C2(P1_U3086), .ZN(P1_U3338) );
  AOI21_X1 U9019 ( .B1(n7168), .B2(n8418), .A(n7167), .ZN(n7171) );
  XNOR2_X1 U9020 ( .A(n8228), .B(n7210), .ZN(n7236) );
  XNOR2_X1 U9021 ( .A(n7236), .B(n8417), .ZN(n7170) );
  NAND2_X1 U9022 ( .A1(n7171), .A2(n7170), .ZN(n7237) );
  OAI21_X1 U9023 ( .B1(n7171), .B2(n7170), .A(n7237), .ZN(n7172) );
  NAND2_X1 U9024 ( .A1(n7172), .A2(n8381), .ZN(n7177) );
  AOI21_X1 U9025 ( .B1(n8402), .B2(n8418), .A(n7173), .ZN(n7174) );
  OAI21_X1 U9026 ( .B1(n7271), .B2(n8398), .A(n7174), .ZN(n7175) );
  AOI21_X1 U9027 ( .B1(n7210), .B2(n8324), .A(n7175), .ZN(n7176) );
  OAI211_X1 U9028 ( .C1(n10168), .C2(n8399), .A(n7177), .B(n7176), .ZN(
        P2_U3170) );
  XOR2_X1 U9029 ( .A(n4518), .B(n7179), .Z(n10077) );
  XOR2_X1 U9030 ( .A(n7179), .B(n7224), .Z(n7182) );
  OAI22_X1 U9031 ( .A1(n7181), .A2(n9089), .B1(n7180), .B2(n9091), .ZN(n7197)
         );
  AOI21_X1 U9032 ( .B1(n7182), .B2(n9996), .A(n7197), .ZN(n10076) );
  MUX2_X1 U9033 ( .A(n7183), .B(n10076), .S(n9734), .Z(n7189) );
  INV_X1 U9034 ( .A(n7184), .ZN(n7186) );
  INV_X1 U9035 ( .A(n7229), .ZN(n7185) );
  AOI21_X1 U9036 ( .B1(n10072), .B2(n7186), .A(n7185), .ZN(n10074) );
  NOR2_X1 U9037 ( .A1(n9746), .A2(n10003), .ZN(n9639) );
  OAI22_X1 U9038 ( .A1(n10029), .A2(n9135), .B1(n7199), .B2(n9699), .ZN(n7187)
         );
  AOI21_X1 U9039 ( .B1(n10074), .B2(n9639), .A(n7187), .ZN(n7188) );
  OAI211_X1 U9040 ( .C1(n9737), .C2(n10077), .A(n7189), .B(n7188), .ZN(
        P1_U3287) );
  NAND2_X1 U9041 ( .A1(n9104), .A2(n9385), .ZN(n7190) );
  OAI21_X1 U9042 ( .B1(n9385), .B2(n6343), .A(n7190), .ZN(P1_U3581) );
  NAND2_X1 U9043 ( .A1(n7191), .A2(n7192), .ZN(n7195) );
  NAND2_X1 U9044 ( .A1(n7191), .A2(n7193), .ZN(n7246) );
  INV_X1 U9045 ( .A(n7246), .ZN(n7194) );
  AOI21_X1 U9046 ( .B1(n7196), .B2(n7195), .A(n7194), .ZN(n7202) );
  AOI22_X1 U9047 ( .A1(n9117), .A2(n7197), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3086), .ZN(n7198) );
  OAI21_X1 U9048 ( .B1(n7199), .B2(n9926), .A(n7198), .ZN(n7200) );
  AOI21_X1 U9049 ( .B1(n10072), .B2(n9924), .A(n7200), .ZN(n7201) );
  OAI21_X1 U9050 ( .B1(n7202), .B2(n9919), .A(n7201), .ZN(P1_U3239) );
  OAI21_X1 U9051 ( .B1(n7204), .B2(n7993), .A(n7203), .ZN(n10165) );
  XNOR2_X1 U9052 ( .A(n7205), .B(n7993), .ZN(n7206) );
  OAI222_X1 U9053 ( .A1(n8768), .A2(n7207), .B1(n8770), .B2(n7271), .C1(n7206), 
        .C2(n8765), .ZN(n10164) );
  AOI21_X1 U9054 ( .B1(n10196), .B2(n10165), .A(n10164), .ZN(n7212) );
  OAI22_X1 U9055 ( .A1(n10170), .A2(n8951), .B1(n10221), .B2(n6072), .ZN(n7208) );
  INV_X1 U9056 ( .A(n7208), .ZN(n7209) );
  OAI21_X1 U9057 ( .B1(n7212), .B2(n10223), .A(n7209), .ZN(P2_U3402) );
  AOI22_X1 U9058 ( .A1(n8875), .A2(n7210), .B1(n10231), .B2(
        P2_REG1_REG_4__SCAN_IN), .ZN(n7211) );
  OAI21_X1 U9059 ( .B1(n7212), .B2(n10231), .A(n7211), .ZN(P2_U3463) );
  INV_X1 U9060 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10606) );
  INV_X1 U9061 ( .A(n7213), .ZN(n7234) );
  INV_X1 U9062 ( .A(n9524), .ZN(n7762) );
  OAI222_X1 U9063 ( .A1(n8152), .A2(n10606), .B1(n7771), .B2(n7234), .C1(
        P1_U3086), .C2(n7762), .ZN(P1_U3337) );
  NAND2_X1 U9064 ( .A1(n7214), .A2(n7192), .ZN(n7215) );
  XOR2_X1 U9065 ( .A(n7216), .B(n7215), .Z(n7222) );
  AOI22_X1 U9066 ( .A1(n9117), .A2(n7217), .B1(P1_REG3_REG_5__SCAN_IN), .B2(
        P1_U3086), .ZN(n7221) );
  INV_X1 U9067 ( .A(n7218), .ZN(n7219) );
  AOI22_X1 U9068 ( .A1(n7219), .A2(n9105), .B1(n9924), .B2(n10067), .ZN(n7220)
         );
  OAI211_X1 U9069 ( .C1(n7222), .C2(n9919), .A(n7221), .B(n7220), .ZN(P1_U3227) );
  XNOR2_X1 U9070 ( .A(n7223), .B(n4612), .ZN(n10085) );
  NAND2_X1 U9071 ( .A1(n7224), .A2(n4802), .ZN(n7225) );
  NAND2_X1 U9072 ( .A1(n7225), .A2(n9129), .ZN(n7394) );
  XNOR2_X1 U9073 ( .A(n7394), .B(n4612), .ZN(n7227) );
  OAI22_X1 U9074 ( .A1(n9132), .A2(n9089), .B1(n7226), .B2(n9091), .ZN(n7249)
         );
  AOI21_X1 U9075 ( .B1(n7227), .B2(n9996), .A(n7249), .ZN(n10083) );
  MUX2_X1 U9076 ( .A(n7228), .B(n10083), .S(n9734), .Z(n7233) );
  AOI211_X1 U9077 ( .C1(n10081), .C2(n7229), .A(n10003), .B(n4920), .ZN(n10080) );
  INV_X1 U9078 ( .A(n10081), .ZN(n7230) );
  OAI22_X1 U9079 ( .A1(n10029), .A2(n7230), .B1(n9699), .B2(n7251), .ZN(n7231)
         );
  AOI21_X1 U9080 ( .B1(n10080), .B2(n10025), .A(n7231), .ZN(n7232) );
  OAI211_X1 U9081 ( .C1(n9737), .C2(n10085), .A(n7233), .B(n7232), .ZN(
        P1_U3286) );
  INV_X1 U9082 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7235) );
  INV_X1 U9083 ( .A(n8574), .ZN(n8586) );
  OAI222_X1 U9084 ( .A1(n8243), .A2(n7235), .B1(n8586), .B2(P2_U3151), .C1(
        n8986), .C2(n7234), .ZN(P2_U3277) );
  XNOR2_X1 U9085 ( .A(n8228), .B(n7439), .ZN(n7270) );
  XNOR2_X1 U9086 ( .A(n7270), .B(n8416), .ZN(n7272) );
  INV_X1 U9087 ( .A(n7236), .ZN(n7238) );
  OAI21_X1 U9088 ( .B1(n7238), .B2(n8417), .A(n7237), .ZN(n7273) );
  XOR2_X1 U9089 ( .A(n7272), .B(n7273), .Z(n7244) );
  NOR2_X1 U9090 ( .A1(n7427), .A2(n8384), .ZN(n7239) );
  AOI211_X1 U9091 ( .C1(n8337), .C2(n8415), .A(n7240), .B(n7239), .ZN(n7241)
         );
  OAI21_X1 U9092 ( .B1(n7437), .B2(n8399), .A(n7241), .ZN(n7242) );
  AOI21_X1 U9093 ( .B1(n7439), .B2(n8324), .A(n7242), .ZN(n7243) );
  OAI21_X1 U9094 ( .B1(n7244), .B2(n8393), .A(n7243), .ZN(P2_U3167) );
  NAND2_X1 U9095 ( .A1(n7246), .A2(n7245), .ZN(n7247) );
  XOR2_X1 U9096 ( .A(n7248), .B(n7247), .Z(n7254) );
  AOI22_X1 U9097 ( .A1(n9117), .A2(n7249), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3086), .ZN(n7250) );
  OAI21_X1 U9098 ( .B1(n7251), .B2(n9926), .A(n7250), .ZN(n7252) );
  AOI21_X1 U9099 ( .B1(n10081), .B2(n9924), .A(n7252), .ZN(n7253) );
  OAI21_X1 U9100 ( .B1(n7254), .B2(n9919), .A(n7253), .ZN(P1_U3213) );
  AOI21_X1 U9101 ( .B1(n7256), .B2(n6675), .A(n7255), .ZN(n7269) );
  XNOR2_X1 U9102 ( .A(n7258), .B(n7257), .ZN(n7259) );
  NAND2_X1 U9103 ( .A1(n7259), .A2(n10146), .ZN(n7268) );
  INV_X1 U9104 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7260) );
  NAND2_X1 U9105 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7415) );
  OAI21_X1 U9106 ( .B1(n8565), .B2(n7260), .A(n7415), .ZN(n7265) );
  AOI21_X1 U9107 ( .B1(n7262), .B2(n6676), .A(n7261), .ZN(n7263) );
  NOR2_X1 U9108 ( .A1(n7263), .A2(n8571), .ZN(n7264) );
  AOI211_X1 U9109 ( .C1(n10155), .C2(n7266), .A(n7265), .B(n7264), .ZN(n7267)
         );
  OAI211_X1 U9110 ( .C1(n7269), .C2(n10152), .A(n7268), .B(n7267), .ZN(
        P2_U3189) );
  XNOR2_X1 U9111 ( .A(n8228), .B(n7466), .ZN(n7410) );
  XNOR2_X1 U9112 ( .A(n7410), .B(n8415), .ZN(n7274) );
  OAI211_X1 U9113 ( .C1(n7275), .C2(n7274), .A(n7411), .B(n8381), .ZN(n7281)
         );
  INV_X1 U9114 ( .A(n7276), .ZN(n7465) );
  AOI21_X1 U9115 ( .B1(n8402), .B2(n8416), .A(n7277), .ZN(n7278) );
  OAI21_X1 U9116 ( .B1(n8020), .B2(n8398), .A(n7278), .ZN(n7279) );
  AOI21_X1 U9117 ( .B1(n7465), .B2(n8389), .A(n7279), .ZN(n7280) );
  OAI211_X1 U9118 ( .C1(n7484), .C2(n8405), .A(n7281), .B(n7280), .ZN(P2_U3179) );
  INV_X1 U9119 ( .A(n7282), .ZN(n8166) );
  OAI222_X1 U9120 ( .A1(n8243), .A2(n7283), .B1(n8986), .B2(n8166), .C1(n8597), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  XNOR2_X1 U9121 ( .A(n9230), .B(n7284), .ZN(n7286) );
  AOI21_X1 U9122 ( .B1(n7286), .B2(n9996), .A(n7285), .ZN(n10056) );
  XNOR2_X1 U9123 ( .A(n7288), .B(n7287), .ZN(n10059) );
  INV_X1 U9124 ( .A(n7289), .ZN(n10002) );
  OAI211_X1 U9125 ( .C1(n10002), .C2(n10055), .A(n10073), .B(n9984), .ZN(
        n10054) );
  NAND2_X1 U9126 ( .A1(n9950), .A2(n7290), .ZN(n7293) );
  AOI22_X1 U9127 ( .A1(n10033), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n10019), .B2(
        n7291), .ZN(n7292) );
  OAI211_X1 U9128 ( .C1(n10054), .C2(n9746), .A(n7293), .B(n7292), .ZN(n7294)
         );
  AOI21_X1 U9129 ( .B1(n10059), .B2(n10006), .A(n7294), .ZN(n7295) );
  OAI21_X1 U9130 ( .B1(n10056), .B2(n10033), .A(n7295), .ZN(P1_U3290) );
  AOI21_X1 U9131 ( .B1(n7296), .B2(n7982), .A(n7988), .ZN(n7299) );
  INV_X1 U9132 ( .A(n7297), .ZN(n7298) );
  NOR2_X1 U9133 ( .A1(n7299), .A2(n7298), .ZN(n10179) );
  NAND2_X1 U9134 ( .A1(n8817), .A2(n7423), .ZN(n8618) );
  AOI22_X1 U9135 ( .A1(n8808), .A2(n8420), .B1(n8418), .B2(n8810), .ZN(n7305)
         );
  INV_X1 U9136 ( .A(n7300), .ZN(n7303) );
  AND3_X1 U9137 ( .A1(n7312), .A2(n7988), .A3(n7301), .ZN(n7302) );
  OAI21_X1 U9138 ( .B1(n7303), .B2(n7302), .A(n8813), .ZN(n7304) );
  OAI211_X1 U9139 ( .C1(n10179), .C2(n7739), .A(n7305), .B(n7304), .ZN(n10181)
         );
  NAND2_X1 U9140 ( .A1(n7306), .A2(n10213), .ZN(n10180) );
  OAI22_X1 U9141 ( .A1(n10180), .A2(n7307), .B1(n10169), .B2(n6026), .ZN(n7308) );
  NOR2_X1 U9142 ( .A1(n10181), .A2(n7308), .ZN(n7309) );
  MUX2_X1 U9143 ( .A(n6692), .B(n7309), .S(n10174), .Z(n7310) );
  OAI21_X1 U9144 ( .B1(n10179), .B2(n8618), .A(n7310), .ZN(P2_U3231) );
  INV_X1 U9145 ( .A(n7313), .ZN(n7949) );
  XNOR2_X1 U9146 ( .A(n7311), .B(n7949), .ZN(n10175) );
  AOI22_X1 U9147 ( .A1(n8808), .A2(n6381), .B1(n8419), .B2(n8810), .ZN(n7317)
         );
  OAI21_X1 U9148 ( .B1(n7314), .B2(n7313), .A(n7312), .ZN(n7315) );
  NAND2_X1 U9149 ( .A1(n7315), .A2(n8813), .ZN(n7316) );
  OAI211_X1 U9150 ( .C1(n10175), .C2(n7739), .A(n7317), .B(n7316), .ZN(n10177)
         );
  NAND2_X1 U9151 ( .A1(n10177), .A2(n10174), .ZN(n7322) );
  OAI22_X1 U9152 ( .A1(n10171), .A2(n7318), .B1(n10169), .B2(n7319), .ZN(n7320) );
  AOI21_X1 U9153 ( .B1(n8636), .B2(P2_REG2_REG_1__SCAN_IN), .A(n7320), .ZN(
        n7321) );
  OAI211_X1 U9154 ( .C1(n10175), .C2(n8618), .A(n7322), .B(n7321), .ZN(
        P2_U3232) );
  INV_X2 U9155 ( .A(n10033), .ZN(n9734) );
  OAI21_X1 U9156 ( .B1(n9639), .B2(n9950), .A(n10020), .ZN(n7329) );
  NAND3_X1 U9157 ( .A1(n9229), .A2(n7324), .A3(n7323), .ZN(n7325) );
  AOI21_X1 U9158 ( .B1(n7326), .B2(n7325), .A(n10033), .ZN(n7327) );
  AOI21_X1 U9159 ( .B1(n10019), .B2(P1_REG3_REG_0__SCAN_IN), .A(n7327), .ZN(
        n7328) );
  OAI211_X1 U9160 ( .C1(n9734), .C2(n7330), .A(n7329), .B(n7328), .ZN(P1_U3293) );
  AOI21_X1 U9161 ( .B1(n4605), .B2(n7332), .A(n7331), .ZN(n7348) );
  OAI21_X1 U9162 ( .B1(n7335), .B2(n7334), .A(n7333), .ZN(n7336) );
  NAND2_X1 U9163 ( .A1(n7336), .A2(n10146), .ZN(n7347) );
  INV_X1 U9164 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7338) );
  NOR2_X1 U9165 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n4616), .ZN(n7552) );
  INV_X1 U9166 ( .A(n7552), .ZN(n7337) );
  OAI21_X1 U9167 ( .B1(n8565), .B2(n7338), .A(n7337), .ZN(n7344) );
  AOI21_X1 U9168 ( .B1(n7341), .B2(n7340), .A(n7339), .ZN(n7342) );
  NOR2_X1 U9169 ( .A1(n7342), .A2(n10152), .ZN(n7343) );
  AOI211_X1 U9170 ( .C1(n10155), .C2(n7345), .A(n7344), .B(n7343), .ZN(n7346)
         );
  OAI211_X1 U9171 ( .C1(n7348), .C2(n8571), .A(n7347), .B(n7346), .ZN(P2_U3190) );
  XNOR2_X1 U9172 ( .A(n7349), .B(n7350), .ZN(n10106) );
  INV_X1 U9173 ( .A(n10106), .ZN(n7360) );
  XNOR2_X1 U9174 ( .A(n7351), .B(n9237), .ZN(n7354) );
  NAND2_X1 U9175 ( .A1(n9379), .A2(n9101), .ZN(n7353) );
  NAND2_X1 U9176 ( .A1(n9377), .A2(n9103), .ZN(n7352) );
  AND2_X1 U9177 ( .A1(n7353), .A2(n7352), .ZN(n7543) );
  OAI21_X1 U9178 ( .B1(n7354), .B2(n10016), .A(n7543), .ZN(n10104) );
  OAI211_X1 U9179 ( .C1(n7355), .C2(n10103), .A(n7529), .B(n10073), .ZN(n10102) );
  OAI22_X1 U9180 ( .A1(n9734), .A2(n6871), .B1(n7540), .B2(n9699), .ZN(n7356)
         );
  AOI21_X1 U9181 ( .B1(n9950), .B2(n7545), .A(n7356), .ZN(n7357) );
  OAI21_X1 U9182 ( .B1(n10102), .B2(n9746), .A(n7357), .ZN(n7358) );
  AOI21_X1 U9183 ( .B1(n10104), .B2(n9734), .A(n7358), .ZN(n7359) );
  OAI21_X1 U9184 ( .B1(n7360), .B2(n9737), .A(n7359), .ZN(P1_U3283) );
  NAND2_X1 U9185 ( .A1(n8645), .A2(P2_U3893), .ZN(n7361) );
  OAI21_X1 U9186 ( .B1(P2_U3893), .B2(n5880), .A(n7361), .ZN(P2_U3518) );
  NAND2_X1 U9187 ( .A1(n9496), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n9513) );
  MUX2_X1 U9188 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n7362), .S(n9496), .Z(n9497)
         );
  AOI21_X1 U9189 ( .B1(n7364), .B2(n7077), .A(n7363), .ZN(n9498) );
  NAND2_X1 U9190 ( .A1(n9497), .A2(n9498), .ZN(n9510) );
  NAND2_X1 U9191 ( .A1(n9513), .A2(n9510), .ZN(n7367) );
  NAND2_X1 U9192 ( .A1(n7377), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7368) );
  OAI21_X1 U9193 ( .B1(n7377), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7368), .ZN(
        n7365) );
  INV_X1 U9194 ( .A(n7365), .ZN(n7366) );
  NAND2_X1 U9195 ( .A1(n7367), .A2(n7366), .ZN(n9516) );
  NAND2_X1 U9196 ( .A1(n9516), .A2(n7368), .ZN(n7490) );
  XNOR2_X1 U9197 ( .A(n7490), .B(n7379), .ZN(n7489) );
  XNOR2_X1 U9198 ( .A(n7489), .B(P1_REG1_REG_15__SCAN_IN), .ZN(n7383) );
  NOR2_X1 U9199 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7369), .ZN(n7371) );
  NOR2_X1 U9200 ( .A1(n9503), .A2(n7379), .ZN(n7370) );
  AOI211_X1 U9201 ( .C1(n9936), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n7371), .B(
        n7370), .ZN(n7382) );
  NAND2_X1 U9202 ( .A1(n9496), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7375) );
  OAI21_X1 U9203 ( .B1(n9496), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7375), .ZN(
        n9491) );
  OAI21_X1 U9204 ( .B1(n7373), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7372), .ZN(
        n9492) );
  NOR2_X1 U9205 ( .A1(n9491), .A2(n9492), .ZN(n9490) );
  INV_X1 U9206 ( .A(n9490), .ZN(n7374) );
  NAND2_X1 U9207 ( .A1(n7375), .A2(n7374), .ZN(n9508) );
  XNOR2_X1 U9208 ( .A(n7377), .B(n7376), .ZN(n9509) );
  NAND2_X1 U9209 ( .A1(n9508), .A2(n9509), .ZN(n9506) );
  NAND2_X1 U9210 ( .A1(n7377), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7378) );
  NAND2_X1 U9211 ( .A1(n9506), .A2(n7378), .ZN(n7502) );
  XNOR2_X1 U9212 ( .A(n7502), .B(n7379), .ZN(n7380) );
  NAND2_X1 U9213 ( .A1(n7380), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n7504) );
  OAI211_X1 U9214 ( .C1(n7380), .C2(P1_REG2_REG_15__SCAN_IN), .A(n9507), .B(
        n7504), .ZN(n7381) );
  OAI211_X1 U9215 ( .C1(n7383), .C2(n9528), .A(n7382), .B(n7381), .ZN(P1_U3258) );
  NAND2_X1 U9216 ( .A1(n7384), .A2(n7385), .ZN(n7446) );
  OAI21_X1 U9217 ( .B1(n7385), .B2(n7384), .A(n7446), .ZN(n7391) );
  NAND2_X1 U9218 ( .A1(n9379), .A2(n9103), .ZN(n7387) );
  NAND2_X1 U9219 ( .A1(n9381), .A2(n9101), .ZN(n7386) );
  NAND2_X1 U9220 ( .A1(n7387), .A2(n7386), .ZN(n9959) );
  AOI22_X1 U9221 ( .A1(n9117), .A2(n9959), .B1(P1_REG3_REG_8__SCAN_IN), .B2(
        P1_U3086), .ZN(n7389) );
  NAND2_X1 U9222 ( .A1(n9924), .A2(n9962), .ZN(n7388) );
  OAI211_X1 U9223 ( .C1(n9926), .C2(n9963), .A(n7389), .B(n7388), .ZN(n7390)
         );
  AOI21_X1 U9224 ( .B1(n7391), .B2(n9097), .A(n7390), .ZN(n7392) );
  INV_X1 U9225 ( .A(n7392), .ZN(P1_U3221) );
  XNOR2_X1 U9226 ( .A(n7393), .B(n7397), .ZN(n10094) );
  INV_X1 U9227 ( .A(n10094), .ZN(n7409) );
  NAND2_X1 U9228 ( .A1(n7394), .A2(n4612), .ZN(n7396) );
  NAND2_X1 U9229 ( .A1(n7396), .A2(n7395), .ZN(n9958) );
  OR2_X1 U9230 ( .A1(n9958), .A2(n9968), .ZN(n9960) );
  NAND2_X1 U9231 ( .A1(n9960), .A2(n9148), .ZN(n7398) );
  XNOR2_X1 U9232 ( .A(n7398), .B(n7397), .ZN(n7399) );
  NAND2_X1 U9233 ( .A1(n7399), .A2(n9996), .ZN(n7400) );
  NAND2_X1 U9234 ( .A1(n9380), .A2(n9101), .ZN(n7452) );
  NAND2_X1 U9235 ( .A1(n7400), .A2(n7452), .ZN(n10100) );
  NAND2_X1 U9236 ( .A1(n10100), .A2(n9734), .ZN(n7408) );
  INV_X1 U9237 ( .A(n10096), .ZN(n7403) );
  XNOR2_X1 U9238 ( .A(n9969), .B(n7403), .ZN(n7401) );
  NAND2_X1 U9239 ( .A1(n7401), .A2(n10073), .ZN(n7402) );
  NAND2_X1 U9240 ( .A1(n9378), .A2(n9103), .ZN(n7453) );
  NAND2_X1 U9241 ( .A1(n7402), .A2(n7453), .ZN(n10097) );
  NOR2_X1 U9242 ( .A1(n7403), .A2(n10029), .ZN(n7406) );
  OAI22_X1 U9243 ( .A1(n9734), .A2(n7404), .B1(n7451), .B2(n9699), .ZN(n7405)
         );
  AOI211_X1 U9244 ( .C1(n10097), .C2(n10025), .A(n7406), .B(n7405), .ZN(n7407)
         );
  OAI211_X1 U9245 ( .C1(n9737), .C2(n7409), .A(n7408), .B(n7407), .ZN(P1_U3284) );
  XNOR2_X1 U9246 ( .A(n8235), .B(n10201), .ZN(n7548) );
  XNOR2_X1 U9247 ( .A(n7548), .B(n8414), .ZN(n7414) );
  OR2_X1 U9248 ( .A1(n7513), .A2(n7410), .ZN(n7412) );
  AOI21_X1 U9249 ( .B1(n7414), .B2(n7413), .A(n7549), .ZN(n7421) );
  INV_X1 U9250 ( .A(n7415), .ZN(n7417) );
  NOR2_X1 U9251 ( .A1(n7513), .A2(n8384), .ZN(n7416) );
  AOI211_X1 U9252 ( .C1(n8337), .C2(n8413), .A(n7417), .B(n7416), .ZN(n7418)
         );
  OAI21_X1 U9253 ( .B1(n7517), .B2(n8399), .A(n7418), .ZN(n7419) );
  AOI21_X1 U9254 ( .B1(n10201), .B2(n8324), .A(n7419), .ZN(n7420) );
  OAI21_X1 U9255 ( .B1(n7421), .B2(n8393), .A(n7420), .ZN(P2_U3153) );
  NAND2_X1 U9256 ( .A1(n7431), .A2(n7633), .ZN(n7422) );
  OAI211_X1 U9257 ( .C1(n10568), .C2(n8152), .A(n7422), .B(n9349), .ZN(
        P1_U3335) );
  NAND2_X1 U9258 ( .A1(n7739), .A2(n4725), .ZN(n10166) );
  XNOR2_X1 U9259 ( .A(n7980), .B(n7424), .ZN(n10187) );
  XNOR2_X1 U9260 ( .A(n7948), .B(n7425), .ZN(n7426) );
  OAI222_X1 U9261 ( .A1(n8770), .A2(n7427), .B1(n8768), .B2(n4796), .C1(n8765), 
        .C2(n7426), .ZN(n10189) );
  NAND2_X1 U9262 ( .A1(n10189), .A2(n8817), .ZN(n7430) );
  OAI22_X1 U9263 ( .A1(n10171), .A2(n10186), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n10169), .ZN(n7428) );
  AOI21_X1 U9264 ( .B1(n8636), .B2(P2_REG2_REG_3__SCAN_IN), .A(n7428), .ZN(
        n7429) );
  OAI211_X1 U9265 ( .C1(n8822), .C2(n10187), .A(n7430), .B(n7429), .ZN(
        P2_U3230) );
  INV_X1 U9266 ( .A(n7431), .ZN(n7432) );
  OAI222_X1 U9267 ( .A1(n8986), .A2(n7432), .B1(n8243), .B2(n6279), .C1(n8141), 
        .C2(P2_U3151), .ZN(P2_U3275) );
  XNOR2_X1 U9268 ( .A(n8416), .B(n7439), .ZN(n7950) );
  XOR2_X1 U9269 ( .A(n7433), .B(n7950), .Z(n10191) );
  XOR2_X1 U9270 ( .A(n7434), .B(n7950), .Z(n7435) );
  AOI222_X1 U9271 ( .A1(n8813), .A2(n7435), .B1(n8415), .B2(n8810), .C1(n8417), 
        .C2(n8808), .ZN(n10192) );
  MUX2_X1 U9272 ( .A(n7436), .B(n10192), .S(n10174), .Z(n7441) );
  INV_X1 U9273 ( .A(n7437), .ZN(n7438) );
  AOI22_X1 U9274 ( .A1(n8801), .A2(n7439), .B1(n8800), .B2(n7438), .ZN(n7440)
         );
  OAI211_X1 U9275 ( .C1(n10191), .C2(n8822), .A(n7441), .B(n7440), .ZN(
        P2_U3228) );
  NAND2_X1 U9276 ( .A1(n8633), .A2(P2_U3893), .ZN(n7442) );
  OAI21_X1 U9277 ( .B1(P2_U3893), .B2(n5912), .A(n7442), .ZN(P2_U3519) );
  NAND2_X1 U9278 ( .A1(n7444), .A2(n7443), .ZN(n7445) );
  NAND2_X1 U9279 ( .A1(n7446), .A2(n7445), .ZN(n7450) );
  NAND2_X1 U9280 ( .A1(n7448), .A2(n7447), .ZN(n7449) );
  XNOR2_X1 U9281 ( .A(n7450), .B(n7449), .ZN(n7459) );
  NOR2_X1 U9282 ( .A1(n9926), .A2(n7451), .ZN(n7457) );
  AND2_X1 U9283 ( .A1(n7453), .A2(n7452), .ZN(n7455) );
  OAI21_X1 U9284 ( .B1(n9914), .B2(n7455), .A(n7454), .ZN(n7456) );
  AOI211_X1 U9285 ( .C1(n10096), .C2(n9924), .A(n7457), .B(n7456), .ZN(n7458)
         );
  OAI21_X1 U9286 ( .B1(n7459), .B2(n9919), .A(n7458), .ZN(P1_U3231) );
  XNOR2_X1 U9287 ( .A(n8415), .B(n7466), .ZN(n7951) );
  NAND2_X1 U9288 ( .A1(n7460), .A2(n7997), .ZN(n7461) );
  XOR2_X1 U9289 ( .A(n7951), .B(n7461), .Z(n7481) );
  XNOR2_X1 U9290 ( .A(n7462), .B(n7951), .ZN(n7463) );
  AOI222_X1 U9291 ( .A1(n8813), .A2(n7463), .B1(n8414), .B2(n8810), .C1(n8416), 
        .C2(n8808), .ZN(n7480) );
  MUX2_X1 U9292 ( .A(n7464), .B(n7480), .S(n10174), .Z(n7468) );
  AOI22_X1 U9293 ( .A1(n8801), .A2(n7466), .B1(n8800), .B2(n7465), .ZN(n7467)
         );
  OAI211_X1 U9294 ( .C1(n7481), .C2(n8822), .A(n7468), .B(n7467), .ZN(P2_U3227) );
  INV_X1 U9295 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10437) );
  INV_X1 U9296 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n7475) );
  NAND2_X1 U9297 ( .A1(n7469), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7473) );
  INV_X1 U9298 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n7470) );
  OR2_X1 U9299 ( .A1(n7471), .A2(n7470), .ZN(n7472) );
  OAI211_X1 U9300 ( .C1(n7475), .C2(n7474), .A(n7473), .B(n7472), .ZN(n7476)
         );
  INV_X1 U9301 ( .A(n7476), .ZN(n7477) );
  NAND2_X1 U9302 ( .A1(n8607), .A2(P2_U3893), .ZN(n7479) );
  OAI21_X1 U9303 ( .B1(P2_U3893), .B2(n10437), .A(n7479), .ZN(P2_U3522) );
  INV_X1 U9304 ( .A(n10196), .ZN(n10217) );
  OAI21_X1 U9305 ( .B1(n10217), .B2(n7481), .A(n7480), .ZN(n7486) );
  OAI22_X1 U9306 ( .A1(n7484), .A2(n8951), .B1(n10221), .B2(n6098), .ZN(n7482)
         );
  AOI21_X1 U9307 ( .B1(n7486), .B2(n10221), .A(n7482), .ZN(n7483) );
  INV_X1 U9308 ( .A(n7483), .ZN(P2_U3408) );
  OAI22_X1 U9309 ( .A1(n8864), .A2(n7484), .B1(n10233), .B2(n6641), .ZN(n7485)
         );
  AOI21_X1 U9310 ( .B1(n7486), .B2(n10233), .A(n7485), .ZN(n7487) );
  INV_X1 U9311 ( .A(n7487), .ZN(P2_U3465) );
  INV_X1 U9312 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9831) );
  NOR2_X1 U9313 ( .A1(n7593), .A2(n9831), .ZN(n7488) );
  AOI21_X1 U9314 ( .B1(n9831), .B2(n7593), .A(n7488), .ZN(n7497) );
  NAND2_X1 U9315 ( .A1(n7489), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n7492) );
  NAND2_X1 U9316 ( .A1(n7490), .A2(n7501), .ZN(n7491) );
  NAND2_X1 U9317 ( .A1(n7492), .A2(n7491), .ZN(n7496) );
  AND2_X1 U9318 ( .A1(n7593), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n7494) );
  NOR2_X1 U9319 ( .A1(n7593), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n7493) );
  INV_X1 U9320 ( .A(n7601), .ZN(n7495) );
  AOI21_X1 U9321 ( .B1(n7497), .B2(n7496), .A(n7495), .ZN(n7510) );
  AND2_X1 U9322 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7500) );
  INV_X1 U9323 ( .A(n7593), .ZN(n7498) );
  NOR2_X1 U9324 ( .A1(n9503), .A2(n7498), .ZN(n7499) );
  AOI211_X1 U9325 ( .C1(n9936), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n7500), .B(
        n7499), .ZN(n7509) );
  NAND2_X1 U9326 ( .A1(n7502), .A2(n7501), .ZN(n7503) );
  NAND2_X1 U9327 ( .A1(n7504), .A2(n7503), .ZN(n7507) );
  INV_X1 U9328 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7505) );
  XNOR2_X1 U9329 ( .A(n7593), .B(n7505), .ZN(n7506) );
  NAND2_X1 U9330 ( .A1(n7507), .A2(n7506), .ZN(n7586) );
  OAI211_X1 U9331 ( .C1(n7507), .C2(n7506), .A(n7586), .B(n9507), .ZN(n7508)
         );
  OAI211_X1 U9332 ( .C1(n7510), .C2(n9528), .A(n7509), .B(n7508), .ZN(P1_U3259) );
  XNOR2_X1 U9333 ( .A(n7511), .B(n8017), .ZN(n10198) );
  XOR2_X1 U9334 ( .A(n7512), .B(n8017), .Z(n7515) );
  OAI22_X1 U9335 ( .A1(n7513), .A2(n8768), .B1(n6398), .B2(n8770), .ZN(n7514)
         );
  AOI21_X1 U9336 ( .B1(n7515), .B2(n8813), .A(n7514), .ZN(n7516) );
  OAI21_X1 U9337 ( .B1(n7739), .B2(n10198), .A(n7516), .ZN(n10199) );
  NAND2_X1 U9338 ( .A1(n10199), .A2(n8817), .ZN(n7520) );
  OAI22_X1 U9339 ( .A1(n10174), .A2(n6676), .B1(n7517), .B2(n10169), .ZN(n7518) );
  AOI21_X1 U9340 ( .B1(n8801), .B2(n10201), .A(n7518), .ZN(n7519) );
  OAI211_X1 U9341 ( .C1(n10198), .C2(n8618), .A(n7520), .B(n7519), .ZN(
        P2_U3226) );
  XNOR2_X1 U9342 ( .A(n7521), .B(n9240), .ZN(n7609) );
  INV_X1 U9343 ( .A(n7609), .ZN(n7535) );
  INV_X1 U9344 ( .A(n7522), .ZN(n7523) );
  AOI211_X1 U9345 ( .C1(n9240), .C2(n7524), .A(n10016), .B(n7523), .ZN(n7527)
         );
  NAND2_X1 U9346 ( .A1(n9376), .A2(n9103), .ZN(n7526) );
  NAND2_X1 U9347 ( .A1(n9378), .A2(n9101), .ZN(n7525) );
  NAND2_X1 U9348 ( .A1(n7526), .A2(n7525), .ZN(n7576) );
  OR2_X1 U9349 ( .A1(n7527), .A2(n7576), .ZN(n7607) );
  NAND2_X1 U9350 ( .A1(n7607), .A2(n9734), .ZN(n7534) );
  INV_X1 U9351 ( .A(n7651), .ZN(n7528) );
  AOI211_X1 U9352 ( .C1(n7614), .C2(n7529), .A(n10003), .B(n7528), .ZN(n7608)
         );
  NOR2_X1 U9353 ( .A1(n7611), .A2(n10029), .ZN(n7532) );
  OAI22_X1 U9354 ( .A1(n9734), .A2(n7530), .B1(n7574), .B2(n9699), .ZN(n7531)
         );
  AOI211_X1 U9355 ( .C1(n7608), .C2(n10025), .A(n7532), .B(n7531), .ZN(n7533)
         );
  OAI211_X1 U9356 ( .C1(n9737), .C2(n7535), .A(n7534), .B(n7533), .ZN(P1_U3282) );
  NAND2_X1 U9357 ( .A1(n7537), .A2(n7536), .ZN(n7539) );
  XNOR2_X1 U9358 ( .A(n7539), .B(n7538), .ZN(n7547) );
  OR2_X1 U9359 ( .A1(n9926), .A2(n7540), .ZN(n7542) );
  NAND2_X1 U9360 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7541) );
  OAI211_X1 U9361 ( .C1(n9914), .C2(n7543), .A(n7542), .B(n7541), .ZN(n7544)
         );
  AOI21_X1 U9362 ( .B1(n7545), .B2(n9924), .A(n7544), .ZN(n7546) );
  OAI21_X1 U9363 ( .B1(n7547), .B2(n9919), .A(n7546), .ZN(P1_U3217) );
  XNOR2_X1 U9364 ( .A(n7568), .B(n8235), .ZN(n7680) );
  XNOR2_X1 U9365 ( .A(n7680), .B(n8413), .ZN(n7681) );
  INV_X1 U9366 ( .A(n7548), .ZN(n7550) );
  XOR2_X1 U9367 ( .A(n7681), .B(n7682), .Z(n7556) );
  NOR2_X1 U9368 ( .A1(n8020), .A2(n8384), .ZN(n7551) );
  AOI211_X1 U9369 ( .C1(n8337), .C2(n8412), .A(n7552), .B(n7551), .ZN(n7553)
         );
  OAI21_X1 U9370 ( .B1(n7565), .B2(n8399), .A(n7553), .ZN(n7554) );
  AOI21_X1 U9371 ( .B1(n7568), .B2(n8324), .A(n7554), .ZN(n7555) );
  OAI21_X1 U9372 ( .B1(n7556), .B2(n8393), .A(n7555), .ZN(P2_U3161) );
  INV_X1 U9373 ( .A(n7557), .ZN(n7560) );
  OAI222_X1 U9374 ( .A1(n8986), .A2(n7560), .B1(P2_U3151), .B2(n7013), .C1(
        n7558), .C2(n8243), .ZN(P2_U3274) );
  OAI222_X1 U9375 ( .A1(P1_U3086), .A2(n9350), .B1(n9908), .B2(n7560), .C1(
        n7559), .C2(n9906), .ZN(P1_U3334) );
  INV_X1 U9376 ( .A(n8022), .ZN(n7561) );
  OR2_X1 U9377 ( .A1(n8027), .A2(n7561), .ZN(n7954) );
  XOR2_X1 U9378 ( .A(n7954), .B(n7562), .Z(n10204) );
  XNOR2_X1 U9379 ( .A(n7563), .B(n7954), .ZN(n7564) );
  OAI222_X1 U9380 ( .A1(n8770), .A2(n7775), .B1(n8768), .B2(n8020), .C1(n7564), 
        .C2(n8765), .ZN(n10206) );
  NAND2_X1 U9381 ( .A1(n10206), .A2(n8817), .ZN(n7570) );
  OAI22_X1 U9382 ( .A1(n8817), .A2(n7566), .B1(n7565), .B2(n10169), .ZN(n7567)
         );
  AOI21_X1 U9383 ( .B1(n8801), .B2(n7568), .A(n7567), .ZN(n7569) );
  OAI211_X1 U9384 ( .C1(n10204), .C2(n8822), .A(n7570), .B(n7569), .ZN(
        P2_U3225) );
  OAI21_X1 U9385 ( .B1(n7572), .B2(n7571), .A(n9918), .ZN(n7573) );
  NAND2_X1 U9386 ( .A1(n7573), .A2(n9097), .ZN(n7578) );
  AND2_X1 U9387 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9479) );
  NOR2_X1 U9388 ( .A1(n9926), .A2(n7574), .ZN(n7575) );
  AOI211_X1 U9389 ( .C1(n9117), .C2(n7576), .A(n9479), .B(n7575), .ZN(n7577)
         );
  OAI211_X1 U9390 ( .C1(n7611), .C2(n9070), .A(n7578), .B(n7577), .ZN(P1_U3236) );
  INV_X1 U9391 ( .A(n7579), .ZN(n7582) );
  OAI222_X1 U9392 ( .A1(n5963), .A2(P1_U3086), .B1(n7771), .B2(n7582), .C1(
        n7580), .C2(n8152), .ZN(P1_U3333) );
  OAI222_X1 U9393 ( .A1(n8243), .A2(n7583), .B1(n8986), .B2(n7582), .C1(n7581), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  OR2_X1 U9394 ( .A1(n7752), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7747) );
  NAND2_X1 U9395 ( .A1(n7752), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7584) );
  NAND2_X1 U9396 ( .A1(n7747), .A2(n7584), .ZN(n7589) );
  NAND2_X1 U9397 ( .A1(n7593), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7585) );
  NAND2_X1 U9398 ( .A1(n7586), .A2(n7585), .ZN(n7588) );
  INV_X1 U9399 ( .A(n7748), .ZN(n7587) );
  AOI21_X1 U9400 ( .B1(n7589), .B2(n7588), .A(n7587), .ZN(n7606) );
  INV_X1 U9401 ( .A(n9936), .ZN(n9541) );
  INV_X1 U9402 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n7592) );
  NOR2_X1 U9403 ( .A1(n7590), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9055) );
  INV_X1 U9404 ( .A(n9055), .ZN(n7591) );
  OAI21_X1 U9405 ( .B1(n9541), .B2(n7592), .A(n7591), .ZN(n7604) );
  OR2_X1 U9406 ( .A1(n7593), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n7599) );
  NAND2_X1 U9407 ( .A1(n7601), .A2(n7599), .ZN(n7597) );
  INV_X1 U9408 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n7594) );
  OR2_X1 U9409 ( .A1(n7752), .A2(n7594), .ZN(n7596) );
  NAND2_X1 U9410 ( .A1(n7752), .A2(n7594), .ZN(n7595) );
  NAND2_X1 U9411 ( .A1(n7596), .A2(n7595), .ZN(n7598) );
  NAND2_X1 U9412 ( .A1(n7597), .A2(n7598), .ZN(n7754) );
  INV_X1 U9413 ( .A(n7598), .ZN(n7600) );
  NAND3_X1 U9414 ( .A1(n7601), .A2(n7600), .A3(n7599), .ZN(n7602) );
  AOI21_X1 U9415 ( .B1(n7754), .B2(n7602), .A(n9528), .ZN(n7603) );
  AOI211_X1 U9416 ( .C1(n9530), .C2(n7752), .A(n7604), .B(n7603), .ZN(n7605)
         );
  OAI21_X1 U9417 ( .B1(n7606), .B2(n9534), .A(n7605), .ZN(P1_U3260) );
  AOI211_X1 U9418 ( .C1(n10112), .C2(n7609), .A(n7608), .B(n7607), .ZN(n7616)
         );
  INV_X1 U9419 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7610) );
  OAI22_X1 U9420 ( .A1(n7611), .A2(n9894), .B1(n10125), .B2(n7610), .ZN(n7612)
         );
  INV_X1 U9421 ( .A(n7612), .ZN(n7613) );
  OAI21_X1 U9422 ( .B1(n7616), .B2(n10123), .A(n7613), .ZN(P1_U3486) );
  AOI22_X1 U9423 ( .A1(n7614), .A2(n6616), .B1(n10139), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n7615) );
  OAI21_X1 U9424 ( .B1(n7616), .B2(n10139), .A(n7615), .ZN(P1_U3533) );
  AOI21_X1 U9425 ( .B1(n7668), .B2(n7618), .A(n7617), .ZN(n7632) );
  INV_X1 U9426 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10254) );
  OAI21_X1 U9427 ( .B1(n7621), .B2(n7620), .A(n7619), .ZN(n7622) );
  NAND2_X1 U9428 ( .A1(n7622), .A2(n10146), .ZN(n7624) );
  NOR2_X1 U9429 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6150), .ZN(n7677) );
  INV_X1 U9430 ( .A(n7677), .ZN(n7623) );
  OAI211_X1 U9431 ( .C1(n8565), .C2(n10254), .A(n7624), .B(n7623), .ZN(n7629)
         );
  AOI21_X1 U9432 ( .B1(n7626), .B2(n6153), .A(n7625), .ZN(n7627) );
  NOR2_X1 U9433 ( .A1(n7627), .A2(n10152), .ZN(n7628) );
  AOI211_X1 U9434 ( .C1(n10155), .C2(n7630), .A(n7629), .B(n7628), .ZN(n7631)
         );
  OAI21_X1 U9435 ( .B1(n7632), .B2(n8571), .A(n7631), .ZN(P2_U3191) );
  NAND2_X1 U9436 ( .A1(n7636), .A2(n7633), .ZN(n7634) );
  OR2_X1 U9437 ( .A1(n9352), .A2(P1_U3086), .ZN(n9358) );
  OAI211_X1 U9438 ( .C1(n10567), .C2(n9906), .A(n7634), .B(n9358), .ZN(
        P1_U3332) );
  NAND2_X1 U9439 ( .A1(n7636), .A2(n7635), .ZN(n7638) );
  INV_X1 U9440 ( .A(n7637), .ZN(n8147) );
  OAI211_X1 U9441 ( .C1(n7639), .C2(n8243), .A(n7638), .B(n8147), .ZN(P2_U3272) );
  XOR2_X1 U9442 ( .A(n7640), .B(n9242), .Z(n7690) );
  INV_X1 U9443 ( .A(n7690), .ZN(n7649) );
  XNOR2_X1 U9444 ( .A(n7641), .B(n9242), .ZN(n7642) );
  AOI22_X1 U9445 ( .A1(n9103), .A2(n9374), .B1(n9376), .B2(n9101), .ZN(n7725)
         );
  OAI21_X1 U9446 ( .B1(n7642), .B2(n10016), .A(n7725), .ZN(n7688) );
  OAI21_X1 U9447 ( .B1(n7730), .B2(n7653), .A(n10073), .ZN(n7643) );
  NOR2_X1 U9448 ( .A1(n7643), .A2(n9954), .ZN(n7689) );
  NAND2_X1 U9449 ( .A1(n7689), .A2(n10025), .ZN(n7646) );
  INV_X1 U9450 ( .A(n7644), .ZN(n7727) );
  AOI22_X1 U9451 ( .A1(n10033), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7727), .B2(
        n10019), .ZN(n7645) );
  OAI211_X1 U9452 ( .C1(n7730), .C2(n10029), .A(n7646), .B(n7645), .ZN(n7647)
         );
  AOI21_X1 U9453 ( .B1(n7688), .B2(n9734), .A(n7647), .ZN(n7648) );
  OAI21_X1 U9454 ( .B1(n7649), .B2(n9737), .A(n7648), .ZN(P1_U3280) );
  XNOR2_X1 U9455 ( .A(n7650), .B(n7660), .ZN(n10113) );
  NAND2_X1 U9456 ( .A1(n7651), .A2(n10108), .ZN(n7652) );
  NAND2_X1 U9457 ( .A1(n7652), .A2(n10073), .ZN(n7654) );
  OR2_X1 U9458 ( .A1(n7654), .A2(n7653), .ZN(n10109) );
  INV_X1 U9459 ( .A(n9927), .ZN(n7655) );
  AOI22_X1 U9460 ( .A1(n10033), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7655), .B2(
        n10019), .ZN(n7657) );
  NAND2_X1 U9461 ( .A1(n10108), .A2(n9950), .ZN(n7656) );
  OAI211_X1 U9462 ( .C1(n10109), .C2(n9746), .A(n7657), .B(n7656), .ZN(n7664)
         );
  OAI21_X1 U9463 ( .B1(n7660), .B2(n7659), .A(n7658), .ZN(n7662) );
  AOI22_X1 U9464 ( .A1(n9101), .A2(n9377), .B1(n9375), .B2(n9103), .ZN(n9913)
         );
  INV_X1 U9465 ( .A(n9913), .ZN(n7661) );
  AOI21_X1 U9466 ( .B1(n7662), .B2(n9996), .A(n7661), .ZN(n10110) );
  NOR2_X1 U9467 ( .A1(n10110), .A2(n10033), .ZN(n7663) );
  AOI211_X1 U9468 ( .C1(n10113), .C2(n10006), .A(n7664), .B(n7663), .ZN(n7665)
         );
  INV_X1 U9469 ( .A(n7665), .ZN(P1_U3281) );
  XOR2_X1 U9470 ( .A(n7666), .B(n7955), .Z(n7667) );
  OAI222_X1 U9471 ( .A1(n8770), .A2(n7820), .B1(n8768), .B2(n6398), .C1(n8765), 
        .C2(n7667), .ZN(n7715) );
  INV_X1 U9472 ( .A(n7715), .ZN(n7675) );
  OAI22_X1 U9473 ( .A1(n8817), .A2(n7668), .B1(n7679), .B2(n10169), .ZN(n7669)
         );
  AOI21_X1 U9474 ( .B1(n8801), .B2(n7718), .A(n7669), .ZN(n7674) );
  NAND2_X1 U9475 ( .A1(n7670), .A2(n7955), .ZN(n7671) );
  AND2_X1 U9476 ( .A1(n7733), .A2(n7671), .ZN(n7716) );
  INV_X1 U9477 ( .A(n8822), .ZN(n7672) );
  NAND2_X1 U9478 ( .A1(n7716), .A2(n7672), .ZN(n7673) );
  OAI211_X1 U9479 ( .C1(n7675), .C2(n8636), .A(n7674), .B(n7673), .ZN(P2_U3224) );
  NOR2_X1 U9480 ( .A1(n6398), .A2(n8384), .ZN(n7676) );
  AOI211_X1 U9481 ( .C1(n8337), .C2(n8411), .A(n7677), .B(n7676), .ZN(n7678)
         );
  OAI21_X1 U9482 ( .B1(n7679), .B2(n8399), .A(n7678), .ZN(n7686) );
  XNOR2_X1 U9483 ( .A(n7718), .B(n8235), .ZN(n7774) );
  XNOR2_X1 U9484 ( .A(n7774), .B(n8412), .ZN(n7684) );
  AOI211_X1 U9485 ( .C1(n7684), .C2(n7683), .A(n8393), .B(n7773), .ZN(n7685)
         );
  AOI211_X1 U9486 ( .C1(n7718), .C2(n8324), .A(n7686), .B(n7685), .ZN(n7687)
         );
  INV_X1 U9487 ( .A(n7687), .ZN(P2_U3171) );
  AOI211_X1 U9488 ( .C1(n7690), .C2(n10112), .A(n7689), .B(n7688), .ZN(n7696)
         );
  INV_X1 U9489 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n7691) );
  OAI22_X1 U9490 ( .A1(n7730), .A2(n9894), .B1(n10125), .B2(n7691), .ZN(n7692)
         );
  INV_X1 U9491 ( .A(n7692), .ZN(n7693) );
  OAI21_X1 U9492 ( .B1(n7696), .B2(n10123), .A(n7693), .ZN(P1_U3492) );
  AOI22_X1 U9493 ( .A1(n7694), .A2(n6616), .B1(n10139), .B2(
        P1_REG1_REG_13__SCAN_IN), .ZN(n7695) );
  OAI21_X1 U9494 ( .B1(n7696), .B2(n10139), .A(n7695), .ZN(P1_U3535) );
  AOI21_X1 U9495 ( .B1(n7699), .B2(n7698), .A(n7697), .ZN(n7714) );
  INV_X1 U9496 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n10258) );
  OAI21_X1 U9497 ( .B1(n7702), .B2(n7701), .A(n7700), .ZN(n7703) );
  NAND2_X1 U9498 ( .A1(n7703), .A2(n10146), .ZN(n7706) );
  INV_X1 U9499 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7704) );
  NOR2_X1 U9500 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7704), .ZN(n7777) );
  INV_X1 U9501 ( .A(n7777), .ZN(n7705) );
  OAI211_X1 U9502 ( .C1(n8565), .C2(n10258), .A(n7706), .B(n7705), .ZN(n7711)
         );
  AOI21_X1 U9503 ( .B1(n4598), .B2(n7708), .A(n7707), .ZN(n7709) );
  NOR2_X1 U9504 ( .A1(n7709), .A2(n10152), .ZN(n7710) );
  AOI211_X1 U9505 ( .C1(n10155), .C2(n7712), .A(n7711), .B(n7710), .ZN(n7713)
         );
  OAI21_X1 U9506 ( .B1(n7714), .B2(n8571), .A(n7713), .ZN(P2_U3192) );
  AOI21_X1 U9507 ( .B1(n7716), .B2(n10196), .A(n7715), .ZN(n7720) );
  AOI22_X1 U9508 ( .A1(n8875), .A2(n7718), .B1(n10231), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n7717) );
  OAI21_X1 U9509 ( .B1(n7720), .B2(n10231), .A(n7717), .ZN(P2_U3468) );
  AOI22_X1 U9510 ( .A1(n8973), .A2(n7718), .B1(n10223), .B2(
        P2_REG0_REG_9__SCAN_IN), .ZN(n7719) );
  OAI21_X1 U9511 ( .B1(n7720), .B2(n10223), .A(n7719), .ZN(P2_U3417) );
  OAI21_X1 U9512 ( .B1(n7723), .B2(n7722), .A(n7721), .ZN(n7724) );
  NAND2_X1 U9513 ( .A1(n7724), .A2(n9097), .ZN(n7729) );
  NAND2_X1 U9514 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n9494) );
  OAI21_X1 U9515 ( .B1(n9914), .B2(n7725), .A(n9494), .ZN(n7726) );
  AOI21_X1 U9516 ( .B1(n7727), .B2(n9105), .A(n7726), .ZN(n7728) );
  OAI211_X1 U9517 ( .C1(n7730), .C2(n9070), .A(n7729), .B(n7728), .ZN(P1_U3234) );
  INV_X1 U9518 ( .A(n7731), .ZN(n7768) );
  INV_X1 U9519 ( .A(n5939), .ZN(n7732) );
  OAI222_X1 U9520 ( .A1(n9906), .A2(n10588), .B1(n9908), .B2(n7768), .C1(
        P1_U3086), .C2(n7732), .ZN(P1_U3331) );
  NAND2_X1 U9521 ( .A1(n7733), .A2(n8014), .ZN(n7734) );
  XNOR2_X1 U9522 ( .A(n7734), .B(n7957), .ZN(n10209) );
  XOR2_X1 U9523 ( .A(n7957), .B(n7735), .Z(n7736) );
  NAND2_X1 U9524 ( .A1(n7736), .A2(n8813), .ZN(n7738) );
  AOI22_X1 U9525 ( .A1(n8410), .A2(n8810), .B1(n8808), .B2(n8412), .ZN(n7737)
         );
  OAI211_X1 U9526 ( .C1(n10209), .C2(n7739), .A(n7738), .B(n7737), .ZN(n10210)
         );
  NAND2_X1 U9527 ( .A1(n10210), .A2(n10174), .ZN(n7743) );
  OAI22_X1 U9528 ( .A1(n10174), .A2(n7740), .B1(n7779), .B2(n10169), .ZN(n7741) );
  AOI21_X1 U9529 ( .B1(n10212), .B2(n8801), .A(n7741), .ZN(n7742) );
  OAI211_X1 U9530 ( .C1(n10209), .C2(n8618), .A(n7743), .B(n7742), .ZN(
        P2_U3223) );
  OR2_X1 U9531 ( .A1(n9524), .A2(n7744), .ZN(n7746) );
  NAND2_X1 U9532 ( .A1(n9524), .A2(n7744), .ZN(n7745) );
  AND2_X1 U9533 ( .A1(n7746), .A2(n7745), .ZN(n7751) );
  NAND2_X1 U9534 ( .A1(n7748), .A2(n7747), .ZN(n7750) );
  INV_X1 U9535 ( .A(n9521), .ZN(n7749) );
  AOI211_X1 U9536 ( .C1(n7751), .C2(n7750), .A(n9534), .B(n7749), .ZN(n7765)
         );
  INV_X1 U9537 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9821) );
  MUX2_X1 U9538 ( .A(n9821), .B(P1_REG1_REG_18__SCAN_IN), .S(n9524), .Z(n7759)
         );
  OR2_X1 U9539 ( .A1(n7752), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n7753) );
  NAND2_X1 U9540 ( .A1(n7754), .A2(n7753), .ZN(n7758) );
  NOR2_X1 U9541 ( .A1(n9524), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n7756) );
  AND2_X1 U9542 ( .A1(n9524), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n7755) );
  INV_X1 U9543 ( .A(n9526), .ZN(n7757) );
  AOI211_X1 U9544 ( .C1(n7759), .C2(n7758), .A(n9528), .B(n7757), .ZN(n7764)
         );
  AND2_X1 U9545 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n7760) );
  AOI21_X1 U9546 ( .B1(n9936), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n7760), .ZN(
        n7761) );
  OAI21_X1 U9547 ( .B1(n9503), .B2(n7762), .A(n7761), .ZN(n7763) );
  OR3_X1 U9548 ( .A1(n7765), .A2(n7764), .A3(n7763), .ZN(P1_U3261) );
  OAI222_X1 U9549 ( .A1(n8986), .A2(n7768), .B1(P2_U3151), .B2(n7767), .C1(
        n7766), .C2(n8243), .ZN(P2_U3271) );
  INV_X1 U9550 ( .A(n7769), .ZN(n8151) );
  OAI222_X1 U9551 ( .A1(n8152), .A2(n7772), .B1(n7771), .B2(n8151), .C1(
        P1_U3086), .C2(n7770), .ZN(P1_U3330) );
  XOR2_X1 U9552 ( .A(n8235), .B(n10212), .Z(n7821) );
  XOR2_X1 U9553 ( .A(n7822), .B(n7821), .Z(n7782) );
  NOR2_X1 U9554 ( .A1(n7775), .A2(n8384), .ZN(n7776) );
  AOI211_X1 U9555 ( .C1(n8337), .C2(n8410), .A(n7777), .B(n7776), .ZN(n7778)
         );
  OAI21_X1 U9556 ( .B1(n7779), .B2(n8399), .A(n7778), .ZN(n7780) );
  AOI21_X1 U9557 ( .B1(n10212), .B2(n8324), .A(n7780), .ZN(n7781) );
  OAI21_X1 U9558 ( .B1(n7782), .B2(n8393), .A(n7781), .ZN(P2_U3157) );
  XNOR2_X1 U9559 ( .A(n7783), .B(n7959), .ZN(n10218) );
  XNOR2_X1 U9560 ( .A(n7784), .B(n7959), .ZN(n7785) );
  OAI222_X1 U9561 ( .A1(n8770), .A2(n7907), .B1(n8768), .B2(n7820), .C1(n7785), 
        .C2(n8765), .ZN(n10220) );
  NAND2_X1 U9562 ( .A1(n10220), .A2(n8817), .ZN(n7788) );
  OAI22_X1 U9563 ( .A1(n8817), .A2(n6179), .B1(n7824), .B2(n10169), .ZN(n7786)
         );
  AOI21_X1 U9564 ( .B1(n7819), .B2(n8801), .A(n7786), .ZN(n7787) );
  OAI211_X1 U9565 ( .C1(n8822), .C2(n10218), .A(n7788), .B(n7787), .ZN(
        P2_U3222) );
  INV_X1 U9566 ( .A(n7789), .ZN(n7791) );
  NOR2_X1 U9567 ( .A1(n7791), .A2(n7790), .ZN(n7794) );
  AOI22_X1 U9568 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n7813), .B1(n8447), .B2(
        n7792), .ZN(n7793) );
  NOR2_X1 U9569 ( .A1(n7794), .A2(n7793), .ZN(n8438) );
  AOI21_X1 U9570 ( .B1(n7794), .B2(n7793), .A(n8438), .ZN(n7815) );
  INV_X1 U9571 ( .A(n7795), .ZN(n7797) );
  MUX2_X1 U9572 ( .A(n7840), .B(P2_REG2_REG_12__SCAN_IN), .S(n7813), .Z(n7799)
         );
  INV_X1 U9573 ( .A(n7799), .ZN(n7800) );
  AOI21_X1 U9574 ( .B1(n7801), .B2(n7800), .A(n8446), .ZN(n7811) );
  NOR2_X1 U9575 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10459), .ZN(n7877) );
  AOI21_X1 U9576 ( .B1(n10145), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n7877), .ZN(
        n7810) );
  MUX2_X1 U9577 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8555), .Z(n8441) );
  XNOR2_X1 U9578 ( .A(n8441), .B(n7813), .ZN(n7807) );
  OR2_X1 U9579 ( .A1(n7803), .A2(n7802), .ZN(n7805) );
  NAND2_X1 U9580 ( .A1(n7805), .A2(n7804), .ZN(n7806) );
  NAND2_X1 U9581 ( .A1(n7807), .A2(n7806), .ZN(n8442) );
  OAI21_X1 U9582 ( .B1(n7807), .B2(n7806), .A(n8442), .ZN(n7808) );
  NAND2_X1 U9583 ( .A1(n7808), .A2(n10146), .ZN(n7809) );
  OAI211_X1 U9584 ( .C1(n7811), .C2(n8571), .A(n7810), .B(n7809), .ZN(n7812)
         );
  AOI21_X1 U9585 ( .B1(n7813), .B2(n10155), .A(n7812), .ZN(n7814) );
  OAI21_X1 U9586 ( .B1(n7815), .B2(n10152), .A(n7814), .ZN(P2_U3194) );
  INV_X1 U9587 ( .A(n7816), .ZN(n7832) );
  OAI222_X1 U9588 ( .A1(n8986), .A2(n7832), .B1(P2_U3151), .B2(n7818), .C1(
        n7817), .C2(n8243), .ZN(P2_U3269) );
  INV_X1 U9589 ( .A(n7819), .ZN(n10216) );
  XNOR2_X1 U9590 ( .A(n7959), .B(n8235), .ZN(n7870) );
  OAI211_X1 U9591 ( .C1(n7823), .C2(n7870), .A(n7872), .B(n8381), .ZN(n7830)
         );
  INV_X1 U9592 ( .A(n7824), .ZN(n7828) );
  AOI21_X1 U9593 ( .B1(n8402), .B2(n8411), .A(n7825), .ZN(n7826) );
  OAI21_X1 U9594 ( .B1(n7907), .B2(n8398), .A(n7826), .ZN(n7827) );
  AOI21_X1 U9595 ( .B1(n7828), .B2(n8389), .A(n7827), .ZN(n7829) );
  OAI211_X1 U9596 ( .C1(n10216), .C2(n8405), .A(n7830), .B(n7829), .ZN(
        P2_U3176) );
  OAI222_X1 U9597 ( .A1(n9906), .A2(n10439), .B1(n9908), .B2(n7832), .C1(
        P1_U3086), .C2(n7831), .ZN(P1_U3329) );
  NAND2_X1 U9598 ( .A1(n7833), .A2(n8047), .ZN(n7834) );
  NAND2_X1 U9599 ( .A1(n7835), .A2(n7834), .ZN(n8880) );
  XNOR2_X1 U9600 ( .A(n7836), .B(n4774), .ZN(n7837) );
  NAND2_X1 U9601 ( .A1(n7837), .A2(n8813), .ZN(n7839) );
  AOI22_X1 U9602 ( .A1(n8410), .A2(n8808), .B1(n8810), .B2(n8809), .ZN(n7838)
         );
  NAND2_X1 U9603 ( .A1(n7839), .A2(n7838), .ZN(n8882) );
  NAND2_X1 U9604 ( .A1(n8882), .A2(n8817), .ZN(n7843) );
  OAI22_X1 U9605 ( .A1(n8817), .A2(n7840), .B1(n7876), .B2(n10169), .ZN(n7841)
         );
  AOI21_X1 U9606 ( .B1(n7873), .B2(n8801), .A(n7841), .ZN(n7842) );
  OAI211_X1 U9607 ( .C1(n8880), .C2(n8822), .A(n7843), .B(n7842), .ZN(P2_U3221) );
  XNOR2_X1 U9608 ( .A(n7844), .B(n7846), .ZN(n9835) );
  INV_X1 U9609 ( .A(n9835), .ZN(n7856) );
  AOI211_X1 U9610 ( .C1(n7846), .C2(n7845), .A(n10016), .B(n4587), .ZN(n7849)
         );
  OAI22_X1 U9611 ( .A1(n7848), .A2(n9091), .B1(n7847), .B2(n9089), .ZN(n9116)
         );
  OR2_X1 U9612 ( .A1(n7849), .A2(n9116), .ZN(n9833) );
  INV_X1 U9613 ( .A(n9121), .ZN(n9895) );
  AOI21_X1 U9614 ( .B1(n4597), .B2(n9121), .A(n10003), .ZN(n7850) );
  AND2_X1 U9615 ( .A1(n7850), .A2(n4533), .ZN(n9834) );
  NAND2_X1 U9616 ( .A1(n9834), .A2(n10025), .ZN(n7853) );
  INV_X1 U9617 ( .A(n9119), .ZN(n7851) );
  AOI22_X1 U9618 ( .A1(n10033), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n7851), .B2(
        n10019), .ZN(n7852) );
  OAI211_X1 U9619 ( .C1(n9895), .C2(n10029), .A(n7853), .B(n7852), .ZN(n7854)
         );
  AOI21_X1 U9620 ( .B1(n9833), .B2(n9734), .A(n7854), .ZN(n7855) );
  OAI21_X1 U9621 ( .B1(n9737), .B2(n7856), .A(n7855), .ZN(P1_U3278) );
  INV_X1 U9622 ( .A(n7857), .ZN(n7860) );
  AOI21_X1 U9623 ( .B1(n8984), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n7858), .ZN(
        n7859) );
  OAI21_X1 U9624 ( .B1(n7860), .B2(n8986), .A(n7859), .ZN(P2_U3268) );
  OAI222_X1 U9625 ( .A1(n4519), .A2(P1_U3086), .B1(n9908), .B2(n7860), .C1(
        n9906), .C2(n5880), .ZN(P1_U3328) );
  XNOR2_X1 U9626 ( .A(n7861), .B(n7961), .ZN(n7918) );
  NAND2_X1 U9627 ( .A1(n7862), .A2(n7961), .ZN(n7863) );
  NAND3_X1 U9628 ( .A1(n7864), .A2(n8813), .A3(n7863), .ZN(n7866) );
  AOI22_X1 U9629 ( .A1(n8808), .A2(n8409), .B1(n8794), .B2(n8810), .ZN(n7865)
         );
  NAND2_X1 U9630 ( .A1(n7866), .A2(n7865), .ZN(n7916) );
  OAI22_X1 U9631 ( .A1(n7917), .A2(n8815), .B1(n7910), .B2(n10169), .ZN(n7867)
         );
  OAI21_X1 U9632 ( .B1(n7916), .B2(n7867), .A(n8817), .ZN(n7869) );
  NAND2_X1 U9633 ( .A1(n8636), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7868) );
  OAI211_X1 U9634 ( .C1(n7918), .C2(n8822), .A(n7869), .B(n7868), .ZN(P2_U3220) );
  INV_X1 U9635 ( .A(n7873), .ZN(n8879) );
  OR2_X1 U9636 ( .A1(n7870), .A2(n7879), .ZN(n7871) );
  NAND2_X1 U9637 ( .A1(n7872), .A2(n7871), .ZN(n7874) );
  XNOR2_X1 U9638 ( .A(n7873), .B(n8235), .ZN(n7902) );
  XOR2_X1 U9639 ( .A(n8409), .B(n7902), .Z(n7875) );
  OAI211_X1 U9640 ( .C1(n7874), .C2(n7875), .A(n7904), .B(n8381), .ZN(n7883)
         );
  INV_X1 U9641 ( .A(n7876), .ZN(n7881) );
  AOI21_X1 U9642 ( .B1(n8337), .B2(n8809), .A(n7877), .ZN(n7878) );
  OAI21_X1 U9643 ( .B1(n7879), .B2(n8384), .A(n7878), .ZN(n7880) );
  AOI21_X1 U9644 ( .B1(n8389), .B2(n7881), .A(n7880), .ZN(n7882) );
  OAI211_X1 U9645 ( .C1(n8879), .C2(n8405), .A(n7883), .B(n7882), .ZN(P2_U3164) );
  INV_X1 U9646 ( .A(n7884), .ZN(n8153) );
  AOI21_X1 U9647 ( .B1(n8984), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n7885), .ZN(
        n7886) );
  OAI21_X1 U9648 ( .B1(n8153), .B2(n8986), .A(n7886), .ZN(P2_U3267) );
  XNOR2_X1 U9649 ( .A(n7887), .B(n9245), .ZN(n9830) );
  INV_X1 U9650 ( .A(n9830), .ZN(n7901) );
  INV_X1 U9651 ( .A(n7888), .ZN(n7889) );
  AOI21_X1 U9652 ( .B1(n7891), .B2(n7890), .A(n7889), .ZN(n7893) );
  OAI22_X1 U9653 ( .A1(n9090), .A2(n9091), .B1(n9001), .B2(n9089), .ZN(n9041)
         );
  INV_X1 U9654 ( .A(n9041), .ZN(n7892) );
  OAI21_X1 U9655 ( .B1(n7893), .B2(n10016), .A(n7892), .ZN(n9828) );
  INV_X1 U9656 ( .A(n9045), .ZN(n9891) );
  NAND2_X1 U9657 ( .A1(n9045), .A2(n4533), .ZN(n7894) );
  NAND2_X1 U9658 ( .A1(n7894), .A2(n10073), .ZN(n7895) );
  NOR2_X1 U9659 ( .A1(n9740), .A2(n7895), .ZN(n9829) );
  NAND2_X1 U9660 ( .A1(n9829), .A2(n10025), .ZN(n7898) );
  INV_X1 U9661 ( .A(n9043), .ZN(n7896) );
  AOI22_X1 U9662 ( .A1(n10033), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n7896), .B2(
        n10019), .ZN(n7897) );
  OAI211_X1 U9663 ( .C1(n9891), .C2(n10029), .A(n7898), .B(n7897), .ZN(n7899)
         );
  AOI21_X1 U9664 ( .B1(n9828), .B2(n9734), .A(n7899), .ZN(n7900) );
  OAI21_X1 U9665 ( .B1(n9737), .B2(n7901), .A(n7900), .ZN(P1_U3277) );
  NAND2_X1 U9666 ( .A1(n7902), .A2(n8409), .ZN(n7903) );
  XNOR2_X1 U9667 ( .A(n8048), .B(n8235), .ZN(n8169) );
  XNOR2_X1 U9668 ( .A(n8169), .B(n7905), .ZN(n7906) );
  XNOR2_X1 U9669 ( .A(n8168), .B(n7906), .ZN(n7913) );
  NOR2_X1 U9670 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6199), .ZN(n8450) );
  NOR2_X1 U9671 ( .A1(n7907), .A2(n8384), .ZN(n7908) );
  AOI211_X1 U9672 ( .C1(n8337), .C2(n8794), .A(n8450), .B(n7908), .ZN(n7909)
         );
  OAI21_X1 U9673 ( .B1(n7910), .B2(n8399), .A(n7909), .ZN(n7911) );
  AOI21_X1 U9674 ( .B1(n8048), .B2(n8324), .A(n7911), .ZN(n7912) );
  OAI21_X1 U9675 ( .B1(n7913), .B2(n8393), .A(n7912), .ZN(P2_U3174) );
  MUX2_X1 U9676 ( .A(n7916), .B(P2_REG0_REG_13__SCAN_IN), .S(n10223), .Z(n7915) );
  OAI22_X1 U9677 ( .A1(n7918), .A2(n8977), .B1(n7917), .B2(n8951), .ZN(n7914)
         );
  OR2_X1 U9678 ( .A1(n7915), .A2(n7914), .ZN(P2_U3429) );
  MUX2_X1 U9679 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n7916), .S(n10233), .Z(n7920) );
  OAI22_X1 U9680 ( .A1(n7918), .A2(n8878), .B1(n7917), .B2(n8864), .ZN(n7919)
         );
  OR2_X1 U9681 ( .A1(n7920), .A2(n7919), .ZN(P2_U3472) );
  INV_X1 U9682 ( .A(n7921), .ZN(n7922) );
  MUX2_X1 U9683 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n4507), .Z(n7928) );
  XNOR2_X1 U9684 ( .A(n7928), .B(SI_30_), .ZN(n7929) );
  INV_X1 U9685 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8154) );
  NOR2_X1 U9686 ( .A1(n7936), .A2(n8154), .ZN(n7926) );
  INV_X1 U9687 ( .A(n8888), .ZN(n8826) );
  INV_X1 U9688 ( .A(n8407), .ZN(n7927) );
  OR2_X1 U9689 ( .A1(n8826), .A2(n7927), .ZN(n8132) );
  INV_X1 U9690 ( .A(n8132), .ZN(n8126) );
  MUX2_X1 U9691 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n4506), .Z(n7933) );
  INV_X1 U9692 ( .A(SI_31_), .ZN(n7932) );
  XNOR2_X1 U9693 ( .A(n7933), .B(n7932), .ZN(n7934) );
  NAND2_X1 U9694 ( .A1(n8980), .A2(n6139), .ZN(n7938) );
  OR2_X1 U9695 ( .A1(n7936), .A2(n6904), .ZN(n7937) );
  INV_X1 U9696 ( .A(n7939), .ZN(n7943) );
  NOR2_X1 U9697 ( .A1(n8888), .A2(n8407), .ZN(n8131) );
  INV_X1 U9698 ( .A(n8131), .ZN(n7941) );
  NAND2_X1 U9699 ( .A1(n7941), .A2(n7940), .ZN(n8128) );
  INV_X1 U9700 ( .A(n8130), .ZN(n8136) );
  OAI21_X1 U9701 ( .B1(n8888), .B2(n8823), .A(n8136), .ZN(n7942) );
  INV_X1 U9702 ( .A(n8674), .ZN(n7945) );
  INV_X1 U9703 ( .A(n8065), .ZN(n8766) );
  INV_X1 U9704 ( .A(n8782), .ZN(n8779) );
  INV_X1 U9705 ( .A(n8806), .ZN(n8804) );
  INV_X1 U9706 ( .A(n7946), .ZN(n7947) );
  AND4_X1 U9707 ( .A1(n7988), .A2(n7949), .A3(n7948), .A4(n7947), .ZN(n7952)
         );
  NAND4_X1 U9708 ( .A1(n7952), .A2(n7993), .A3(n7951), .A4(n7950), .ZN(n7953)
         );
  NOR3_X1 U9709 ( .A1(n7955), .A2(n7954), .A3(n7953), .ZN(n7956) );
  NAND3_X1 U9710 ( .A1(n7957), .A2(n7956), .A3(n8017), .ZN(n7958) );
  NOR2_X1 U9711 ( .A1(n7959), .A2(n7958), .ZN(n7960) );
  NAND3_X1 U9712 ( .A1(n7961), .A2(n4774), .A3(n7960), .ZN(n7962) );
  NOR2_X1 U9713 ( .A1(n8804), .A2(n7962), .ZN(n7964) );
  NAND4_X1 U9714 ( .A1(n8766), .A2(n8779), .A3(n7964), .A4(n8793), .ZN(n7965)
         );
  NOR2_X1 U9715 ( .A1(n8755), .A2(n7965), .ZN(n7966) );
  NAND3_X1 U9716 ( .A1(n8731), .A2(n8743), .A3(n7966), .ZN(n7967) );
  OR4_X1 U9717 ( .A1(n8691), .A2(n8651), .A3(n8718), .A4(n7967), .ZN(n7969) );
  INV_X1 U9718 ( .A(n7968), .ZN(n8113) );
  NAND2_X1 U9719 ( .A1(n8104), .A2(n8099), .ZN(n8677) );
  OR4_X1 U9720 ( .A1(n7969), .A2(n8643), .A3(n8662), .A4(n8677), .ZN(n7971) );
  INV_X1 U9721 ( .A(n8622), .ZN(n7970) );
  MUX2_X1 U9722 ( .A(n8252), .B(n8127), .S(n8133), .Z(n8122) );
  AND2_X1 U9723 ( .A1(n8674), .A2(n7977), .ZN(n7978) );
  MUX2_X1 U9724 ( .A(n7979), .B(n7978), .S(n8133), .Z(n8097) );
  INV_X1 U9725 ( .A(n7980), .ZN(n7984) );
  AND2_X1 U9726 ( .A1(n7982), .A2(n7981), .ZN(n7985) );
  NAND3_X1 U9727 ( .A1(n7984), .A2(n8003), .A3(n7983), .ZN(n7992) );
  INV_X1 U9728 ( .A(n7985), .ZN(n7986) );
  NAND3_X1 U9729 ( .A1(n7988), .A2(n7987), .A3(n7986), .ZN(n7990) );
  NAND3_X1 U9730 ( .A1(n7990), .A2(n7995), .A3(n7989), .ZN(n7991) );
  MUX2_X1 U9731 ( .A(n7992), .B(n7991), .S(n8124), .Z(n7994) );
  NAND2_X1 U9732 ( .A1(n7994), .A2(n7993), .ZN(n8007) );
  INV_X1 U9733 ( .A(n7995), .ZN(n7998) );
  OAI211_X1 U9734 ( .C1(n8007), .C2(n7998), .A(n7997), .B(n7996), .ZN(n8002)
         );
  AND2_X1 U9735 ( .A1(n8008), .A2(n8004), .ZN(n8001) );
  INV_X1 U9736 ( .A(n7999), .ZN(n8000) );
  AOI21_X1 U9737 ( .B1(n8002), .B2(n8001), .A(n8000), .ZN(n8013) );
  INV_X1 U9738 ( .A(n8003), .ZN(n8006) );
  NAND2_X1 U9739 ( .A1(n8417), .A2(n10170), .ZN(n8005) );
  OAI211_X1 U9740 ( .C1(n8007), .C2(n8006), .A(n8005), .B(n8004), .ZN(n8011)
         );
  INV_X1 U9741 ( .A(n8008), .ZN(n8009) );
  AOI21_X1 U9742 ( .B1(n8011), .B2(n8010), .A(n8009), .ZN(n8012) );
  MUX2_X1 U9743 ( .A(n8013), .B(n8012), .S(n8124), .Z(n8019) );
  NAND2_X1 U9744 ( .A1(n8023), .A2(n8022), .ZN(n8029) );
  INV_X1 U9745 ( .A(n8027), .ZN(n8015) );
  NAND2_X1 U9746 ( .A1(n8015), .A2(n8014), .ZN(n8016) );
  MUX2_X1 U9747 ( .A(n8029), .B(n8016), .S(n8124), .Z(n8025) );
  INV_X1 U9748 ( .A(n8025), .ZN(n8018) );
  NAND3_X1 U9749 ( .A1(n8019), .A2(n8018), .A3(n8017), .ZN(n8035) );
  NAND2_X1 U9750 ( .A1(n10201), .A2(n8020), .ZN(n8021) );
  AND2_X1 U9751 ( .A1(n8022), .A2(n8021), .ZN(n8024) );
  OAI211_X1 U9752 ( .C1(n8025), .C2(n8024), .A(n8023), .B(n8036), .ZN(n8032)
         );
  NOR2_X1 U9753 ( .A1(n8027), .A2(n4794), .ZN(n8030) );
  OAI21_X1 U9754 ( .B1(n8030), .B2(n8029), .A(n8028), .ZN(n8031) );
  MUX2_X1 U9755 ( .A(n8032), .B(n8031), .S(n8133), .Z(n8033) );
  INV_X1 U9756 ( .A(n8033), .ZN(n8034) );
  NAND2_X1 U9757 ( .A1(n8035), .A2(n8034), .ZN(n8043) );
  AND2_X1 U9758 ( .A1(n8041), .A2(n8036), .ZN(n8038) );
  INV_X1 U9759 ( .A(n8040), .ZN(n8037) );
  INV_X1 U9760 ( .A(n8041), .ZN(n8042) );
  MUX2_X1 U9761 ( .A(n8045), .B(n8044), .S(n8124), .Z(n8046) );
  MUX2_X1 U9762 ( .A(n8809), .B(n8048), .S(n8124), .Z(n8052) );
  INV_X1 U9763 ( .A(n8049), .ZN(n8050) );
  NAND2_X1 U9764 ( .A1(n8052), .A2(n8051), .ZN(n8053) );
  NAND2_X1 U9765 ( .A1(n8054), .A2(n8053), .ZN(n8055) );
  NAND2_X1 U9766 ( .A1(n8055), .A2(n8806), .ZN(n8062) );
  INV_X1 U9767 ( .A(n8056), .ZN(n8059) );
  NAND2_X1 U9768 ( .A1(n8063), .A2(n8057), .ZN(n8058) );
  MUX2_X1 U9769 ( .A(n8059), .B(n8058), .S(n8133), .Z(n8060) );
  NOR2_X1 U9770 ( .A1(n8060), .A2(n8068), .ZN(n8061) );
  NAND2_X1 U9771 ( .A1(n8062), .A2(n8061), .ZN(n8071) );
  NAND2_X1 U9772 ( .A1(n8071), .A2(n8063), .ZN(n8064) );
  AOI21_X1 U9773 ( .B1(n8079), .B2(n8066), .A(n8133), .ZN(n8067) );
  INV_X1 U9774 ( .A(n8068), .ZN(n8070) );
  AOI21_X1 U9775 ( .B1(n8071), .B2(n8070), .A(n4736), .ZN(n8074) );
  INV_X1 U9776 ( .A(n8072), .ZN(n8073) );
  OAI21_X1 U9777 ( .B1(n8074), .B2(n8073), .A(n8133), .ZN(n8075) );
  NAND2_X1 U9778 ( .A1(n8076), .A2(n8075), .ZN(n8084) );
  NAND2_X1 U9779 ( .A1(n8085), .A2(n8081), .ZN(n8077) );
  NOR2_X1 U9780 ( .A1(n8084), .A2(n8077), .ZN(n8078) );
  MUX2_X1 U9781 ( .A(n8079), .B(n8078), .S(n8124), .Z(n8091) );
  AND2_X1 U9782 ( .A1(n8081), .A2(n8080), .ZN(n8083) );
  INV_X1 U9783 ( .A(n8086), .ZN(n8082) );
  AOI21_X1 U9784 ( .B1(n8084), .B2(n8083), .A(n8082), .ZN(n8090) );
  NAND2_X1 U9785 ( .A1(n8731), .A2(n8085), .ZN(n8088) );
  NAND2_X1 U9786 ( .A1(n8714), .A2(n8086), .ZN(n8087) );
  MUX2_X1 U9787 ( .A(n8088), .B(n8087), .S(n8124), .Z(n8089) );
  NAND2_X1 U9788 ( .A1(n8094), .A2(n8713), .ZN(n8092) );
  MUX2_X1 U9789 ( .A(n8092), .B(n4703), .S(n8133), .Z(n8096) );
  INV_X1 U9790 ( .A(n8651), .ZN(n8703) );
  MUX2_X1 U9791 ( .A(n8094), .B(n8093), .S(n8124), .Z(n8095) );
  NAND3_X1 U9792 ( .A1(n8103), .A2(n8104), .A3(n8098), .ZN(n8100) );
  NAND2_X1 U9793 ( .A1(n8100), .A2(n8099), .ZN(n8107) );
  NAND2_X1 U9794 ( .A1(n8105), .A2(n8104), .ZN(n8106) );
  MUX2_X1 U9795 ( .A(n8107), .B(n8106), .S(n8124), .Z(n8111) );
  MUX2_X1 U9796 ( .A(n8109), .B(n8108), .S(n8133), .Z(n8110) );
  OAI211_X1 U9797 ( .C1(n8111), .C2(n8662), .A(n8641), .B(n8110), .ZN(n8116)
         );
  MUX2_X1 U9798 ( .A(n8113), .B(n8112), .S(n8124), .Z(n8114) );
  NOR2_X1 U9799 ( .A1(n8629), .A2(n8114), .ZN(n8115) );
  NAND2_X1 U9800 ( .A1(n8897), .A2(n8386), .ZN(n8118) );
  MUX2_X1 U9801 ( .A(n8118), .B(n8117), .S(n8133), .Z(n8119) );
  INV_X1 U9802 ( .A(n8119), .ZN(n8120) );
  NAND3_X1 U9803 ( .A1(n4753), .A2(n8124), .A3(n8123), .ZN(n8125) );
  AOI211_X1 U9804 ( .C1(n8127), .C2(n8129), .A(n8126), .B(n8125), .ZN(n8140)
         );
  AOI211_X1 U9805 ( .C1(n8133), .C2(n8132), .A(n8131), .B(n8130), .ZN(n8134)
         );
  AOI211_X1 U9806 ( .C1(n8137), .C2(n8136), .A(n8135), .B(n8134), .ZN(n8138)
         );
  NAND3_X1 U9807 ( .A1(n8143), .A2(n8142), .A3(n8555), .ZN(n8144) );
  OAI211_X1 U9808 ( .C1(n8145), .C2(n8147), .A(n8144), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8146) );
  OAI21_X1 U9809 ( .B1(n8148), .B2(n8147), .A(n8146), .ZN(P2_U3296) );
  OAI222_X1 U9810 ( .A1(n8986), .A2(n8151), .B1(P2_U3151), .B2(n8150), .C1(
        n8149), .C2(n8243), .ZN(P2_U3270) );
  OAI222_X1 U9811 ( .A1(n9399), .A2(P1_U3086), .B1(n9908), .B2(n8153), .C1(
        n8152), .C2(n5912), .ZN(P1_U3327) );
  INV_X1 U9812 ( .A(n8157), .ZN(n9905) );
  OAI222_X1 U9813 ( .A1(n8243), .A2(n8154), .B1(n8986), .B2(n9905), .C1(
        P2_U3151), .C2(n4505), .ZN(P2_U3265) );
  NAND2_X1 U9814 ( .A1(n8980), .A2(n5441), .ZN(n8156) );
  NAND2_X1 U9815 ( .A1(n8158), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8155) );
  INV_X1 U9816 ( .A(n9545), .ZN(n9842) );
  NAND2_X1 U9817 ( .A1(n8157), .A2(n5441), .ZN(n8160) );
  NAND2_X1 U9818 ( .A1(n8158), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8159) );
  OR2_X1 U9819 ( .A1(n9225), .A2(n8163), .ZN(n9542) );
  MUX2_X1 U9820 ( .A(n8164), .B(n9840), .S(n10141), .Z(n8165) );
  OAI21_X1 U9821 ( .B1(n9842), .B2(n9837), .A(n8165), .ZN(P1_U3553) );
  OAI222_X1 U9822 ( .A1(n5284), .A2(P1_U3086), .B1(n9908), .B2(n8166), .C1(
        n10661), .C2(n9906), .ZN(P1_U3336) );
  INV_X1 U9823 ( .A(n8257), .ZN(n8171) );
  XNOR2_X1 U9824 ( .A(n8974), .B(n8235), .ZN(n8172) );
  XNOR2_X1 U9825 ( .A(n8172), .B(n8794), .ZN(n8261) );
  INV_X1 U9826 ( .A(n8172), .ZN(n8174) );
  NAND2_X1 U9827 ( .A1(n8174), .A2(n8173), .ZN(n8175) );
  XNOR2_X1 U9828 ( .A(n8967), .B(n8235), .ZN(n8176) );
  XNOR2_X1 U9829 ( .A(n8176), .B(n8811), .ZN(n8394) );
  NAND2_X1 U9830 ( .A1(n8176), .A2(n8811), .ZN(n8177) );
  XNOR2_X1 U9831 ( .A(n8961), .B(n8235), .ZN(n8178) );
  XOR2_X1 U9832 ( .A(n8795), .B(n8178), .Z(n8312) );
  NAND2_X1 U9833 ( .A1(n8178), .A2(n8795), .ZN(n8179) );
  XNOR2_X1 U9834 ( .A(n8955), .B(n8228), .ZN(n8181) );
  NAND2_X1 U9835 ( .A1(n8181), .A2(n8753), .ZN(n8366) );
  OAI21_X1 U9836 ( .B1(n8181), .B2(n8753), .A(n8366), .ZN(n8321) );
  XNOR2_X1 U9837 ( .A(n8365), .B(n8228), .ZN(n8182) );
  NAND2_X1 U9838 ( .A1(n8182), .A2(n8771), .ZN(n8276) );
  INV_X1 U9839 ( .A(n8182), .ZN(n8183) );
  NAND2_X1 U9840 ( .A1(n8183), .A2(n8744), .ZN(n8184) );
  NAND2_X1 U9841 ( .A1(n8185), .A2(n8367), .ZN(n8275) );
  NAND2_X1 U9842 ( .A1(n8275), .A2(n8276), .ZN(n8210) );
  XNOR2_X1 U9843 ( .A(n8944), .B(n8228), .ZN(n8186) );
  NAND2_X1 U9844 ( .A1(n8186), .A2(n8754), .ZN(n8340) );
  INV_X1 U9845 ( .A(n8186), .ZN(n8187) );
  NAND2_X1 U9846 ( .A1(n8187), .A2(n8408), .ZN(n8188) );
  NAND2_X1 U9847 ( .A1(n8210), .A2(n8277), .ZN(n8279) );
  NAND2_X1 U9848 ( .A1(n8279), .A2(n8340), .ZN(n8287) );
  XNOR2_X1 U9849 ( .A(n8228), .B(n8737), .ZN(n8189) );
  NAND2_X1 U9850 ( .A1(n8189), .A2(n8282), .ZN(n8289) );
  INV_X1 U9851 ( .A(n8189), .ZN(n8190) );
  NAND2_X1 U9852 ( .A1(n8190), .A2(n8745), .ZN(n8191) );
  XNOR2_X1 U9853 ( .A(n8927), .B(n8235), .ZN(n8193) );
  INV_X1 U9854 ( .A(n8193), .ZN(n8192) );
  NAND2_X1 U9855 ( .A1(n8192), .A2(n8294), .ZN(n8203) );
  INV_X1 U9856 ( .A(n8203), .ZN(n8200) );
  XNOR2_X1 U9857 ( .A(n8193), .B(n8294), .ZN(n8351) );
  INV_X1 U9858 ( .A(n8351), .ZN(n8194) );
  XNOR2_X1 U9859 ( .A(n8933), .B(n8228), .ZN(n8195) );
  NAND2_X1 U9860 ( .A1(n8195), .A2(n8733), .ZN(n8350) );
  OR2_X1 U9861 ( .A1(n8194), .A2(n8350), .ZN(n8202) );
  INV_X1 U9862 ( .A(n8202), .ZN(n8199) );
  INV_X1 U9863 ( .A(n8195), .ZN(n8196) );
  NAND2_X1 U9864 ( .A1(n8196), .A2(n8707), .ZN(n8197) );
  AND2_X1 U9865 ( .A1(n8290), .A2(n8351), .ZN(n8198) );
  NAND2_X1 U9866 ( .A1(n8287), .A2(n8211), .ZN(n8208) );
  XOR2_X1 U9867 ( .A(n8235), .B(n8921), .Z(n8217) );
  INV_X1 U9868 ( .A(n8217), .ZN(n8206) );
  INV_X1 U9869 ( .A(n8201), .ZN(n8205) );
  AND2_X1 U9870 ( .A1(n8289), .A2(n8202), .ZN(n8354) );
  AND2_X1 U9871 ( .A1(n8354), .A2(n8203), .ZN(n8204) );
  AND2_X1 U9872 ( .A1(n8206), .A2(n8213), .ZN(n8207) );
  AND2_X1 U9873 ( .A1(n8277), .A2(n8211), .ZN(n8209) );
  INV_X1 U9874 ( .A(n8211), .ZN(n8212) );
  XNOR2_X1 U9875 ( .A(n8915), .B(n8228), .ZN(n8220) );
  NAND2_X1 U9876 ( .A1(n8220), .A2(n8305), .ZN(n8300) );
  INV_X1 U9877 ( .A(n8220), .ZN(n8221) );
  NAND2_X1 U9878 ( .A1(n8221), .A2(n8693), .ZN(n8222) );
  NAND2_X1 U9879 ( .A1(n8223), .A2(n8329), .ZN(n8299) );
  NAND2_X1 U9880 ( .A1(n8299), .A2(n8300), .ZN(n8227) );
  XNOR2_X1 U9881 ( .A(n8909), .B(n8228), .ZN(n8224) );
  NAND2_X1 U9882 ( .A1(n8224), .A2(n8385), .ZN(n8376) );
  INV_X1 U9883 ( .A(n8224), .ZN(n8225) );
  NAND2_X1 U9884 ( .A1(n8225), .A2(n8679), .ZN(n8226) );
  NAND2_X1 U9885 ( .A1(n8227), .A2(n8301), .ZN(n8303) );
  NAND2_X1 U9886 ( .A1(n8303), .A2(n8376), .ZN(n8229) );
  XNOR2_X1 U9887 ( .A(n8903), .B(n8228), .ZN(n8230) );
  XNOR2_X1 U9888 ( .A(n8230), .B(n8664), .ZN(n8377) );
  NAND2_X1 U9889 ( .A1(n8230), .A2(n8306), .ZN(n8231) );
  XNOR2_X1 U9890 ( .A(n8897), .B(n8235), .ZN(n8233) );
  XNOR2_X1 U9891 ( .A(n8233), .B(n8645), .ZN(n8246) );
  INV_X1 U9892 ( .A(n8233), .ZN(n8234) );
  NAND2_X1 U9893 ( .A1(n8248), .A2(n5121), .ZN(n8237) );
  XOR2_X1 U9894 ( .A(n8235), .B(n8622), .Z(n8236) );
  XNOR2_X1 U9895 ( .A(n8237), .B(n8236), .ZN(n8242) );
  NAND2_X1 U9896 ( .A1(n8623), .A2(n8337), .ZN(n8239) );
  AOI22_X1 U9897 ( .A1(n8625), .A2(n8389), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8238) );
  OAI211_X1 U9898 ( .C1(n8386), .C2(n8384), .A(n8239), .B(n8238), .ZN(n8240)
         );
  AOI21_X1 U9899 ( .B1(n8891), .B2(n8324), .A(n8240), .ZN(n8241) );
  OAI21_X1 U9900 ( .B1(n8242), .B2(n8393), .A(n8241), .ZN(P2_U3160) );
  OAI222_X1 U9901 ( .A1(n8986), .A2(n9907), .B1(P2_U3151), .B2(n8245), .C1(
        n8244), .C2(n8243), .ZN(P2_U3266) );
  INV_X1 U9902 ( .A(n8897), .ZN(n8256) );
  AOI21_X1 U9903 ( .B1(n8247), .B2(n8246), .A(n8393), .ZN(n8250) );
  NAND2_X1 U9904 ( .A1(n8250), .A2(n8249), .ZN(n8255) );
  AOI22_X1 U9905 ( .A1(n8638), .A2(n8389), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8251) );
  OAI21_X1 U9906 ( .B1(n8252), .B2(n8398), .A(n8251), .ZN(n8253) );
  AOI21_X1 U9907 ( .B1(n8402), .B2(n8664), .A(n8253), .ZN(n8254) );
  OAI211_X1 U9908 ( .C1(n8256), .C2(n8405), .A(n8255), .B(n8254), .ZN(P2_U3154) );
  INV_X1 U9909 ( .A(n8259), .ZN(n8260) );
  AOI21_X1 U9910 ( .B1(n8261), .B2(n8257), .A(n8260), .ZN(n8267) );
  NAND2_X1 U9911 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8470) );
  OAI21_X1 U9912 ( .B1(n8398), .B2(n8262), .A(n8470), .ZN(n8263) );
  AOI21_X1 U9913 ( .B1(n8402), .B2(n8809), .A(n8263), .ZN(n8264) );
  OAI21_X1 U9914 ( .B1(n8399), .B2(n8814), .A(n8264), .ZN(n8265) );
  AOI21_X1 U9915 ( .B1(n8974), .B2(n8324), .A(n8265), .ZN(n8266) );
  OAI21_X1 U9916 ( .B1(n8267), .B2(n8393), .A(n8266), .ZN(P2_U3155) );
  INV_X1 U9917 ( .A(n8269), .ZN(n8331) );
  AOI21_X1 U9918 ( .B1(n8706), .B2(n8268), .A(n8331), .ZN(n8274) );
  AOI22_X1 U9919 ( .A1(n8723), .A2(n8402), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8271) );
  NAND2_X1 U9920 ( .A1(n8696), .A2(n8389), .ZN(n8270) );
  OAI211_X1 U9921 ( .C1(n8305), .C2(n8398), .A(n8271), .B(n8270), .ZN(n8272)
         );
  AOI21_X1 U9922 ( .B1(n8921), .B2(n8324), .A(n8272), .ZN(n8273) );
  OAI21_X1 U9923 ( .B1(n8274), .B2(n8393), .A(n8273), .ZN(P2_U3156) );
  INV_X1 U9924 ( .A(n8944), .ZN(n8286) );
  INV_X1 U9925 ( .A(n8275), .ZN(n8370) );
  INV_X1 U9926 ( .A(n8276), .ZN(n8278) );
  NOR3_X1 U9927 ( .A1(n8370), .A2(n8278), .A3(n8277), .ZN(n8280) );
  INV_X1 U9928 ( .A(n8279), .ZN(n8343) );
  OAI21_X1 U9929 ( .B1(n8280), .B2(n8343), .A(n8381), .ZN(n8285) );
  NAND2_X1 U9930 ( .A1(n8744), .A2(n8402), .ZN(n8281) );
  NAND2_X1 U9931 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8595) );
  OAI211_X1 U9932 ( .C1(n8282), .C2(n8398), .A(n8281), .B(n8595), .ZN(n8283)
         );
  AOI21_X1 U9933 ( .B1(n8748), .B2(n8389), .A(n8283), .ZN(n8284) );
  OAI211_X1 U9934 ( .C1(n8286), .C2(n8405), .A(n8285), .B(n8284), .ZN(P2_U3159) );
  INV_X1 U9935 ( .A(n8933), .ZN(n8298) );
  NAND2_X1 U9936 ( .A1(n8287), .A2(n8341), .ZN(n8355) );
  INV_X1 U9937 ( .A(n8355), .ZN(n8344) );
  INV_X1 U9938 ( .A(n8289), .ZN(n8288) );
  NOR3_X1 U9939 ( .A1(n8344), .A2(n8288), .A3(n8290), .ZN(n8292) );
  NAND2_X1 U9940 ( .A1(n8355), .A2(n8289), .ZN(n8291) );
  OAI21_X1 U9941 ( .B1(n8292), .B2(n8353), .A(n8381), .ZN(n8297) );
  AOI22_X1 U9942 ( .A1(n8745), .A2(n8402), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8293) );
  OAI21_X1 U9943 ( .B1(n8294), .B2(n8398), .A(n8293), .ZN(n8295) );
  AOI21_X1 U9944 ( .B1(n8726), .B2(n8389), .A(n8295), .ZN(n8296) );
  OAI211_X1 U9945 ( .C1(n8298), .C2(n8405), .A(n8297), .B(n8296), .ZN(P2_U3163) );
  INV_X1 U9946 ( .A(n8909), .ZN(n8311) );
  INV_X1 U9947 ( .A(n8299), .ZN(n8332) );
  INV_X1 U9948 ( .A(n8300), .ZN(n8302) );
  NOR3_X1 U9949 ( .A1(n8332), .A2(n8302), .A3(n8301), .ZN(n8304) );
  INV_X1 U9950 ( .A(n8303), .ZN(n8379) );
  OAI21_X1 U9951 ( .B1(n8304), .B2(n8379), .A(n8381), .ZN(n8310) );
  INV_X1 U9952 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n10622) );
  OAI22_X1 U9953 ( .A1(n8305), .A2(n8384), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10622), .ZN(n8308) );
  NOR2_X1 U9954 ( .A1(n8306), .A2(n8398), .ZN(n8307) );
  AOI211_X1 U9955 ( .C1(n8666), .C2(n8389), .A(n8308), .B(n8307), .ZN(n8309)
         );
  OAI211_X1 U9956 ( .C1(n8311), .C2(n8405), .A(n8310), .B(n8309), .ZN(P2_U3165) );
  XNOR2_X1 U9957 ( .A(n8313), .B(n8312), .ZN(n8318) );
  NAND2_X1 U9958 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8516) );
  NAND2_X1 U9959 ( .A1(n8402), .A2(n8811), .ZN(n8314) );
  OAI211_X1 U9960 ( .C1(n8398), .C2(n8753), .A(n8516), .B(n8314), .ZN(n8315)
         );
  AOI21_X1 U9961 ( .B1(n8389), .B2(n8788), .A(n8315), .ZN(n8317) );
  NAND2_X1 U9962 ( .A1(n8961), .A2(n8324), .ZN(n8316) );
  OAI211_X1 U9963 ( .C1(n8318), .C2(n8393), .A(n8317), .B(n8316), .ZN(P2_U3166) );
  INV_X1 U9964 ( .A(n8320), .ZN(n8369) );
  AOI21_X1 U9965 ( .B1(n8321), .B2(n8319), .A(n8369), .ZN(n8327) );
  NAND2_X1 U9966 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8540) );
  NAND2_X1 U9967 ( .A1(n8402), .A2(n8795), .ZN(n8322) );
  OAI211_X1 U9968 ( .C1(n8398), .C2(n8771), .A(n8540), .B(n8322), .ZN(n8323)
         );
  AOI21_X1 U9969 ( .B1(n8776), .B2(n8389), .A(n8323), .ZN(n8326) );
  NAND2_X1 U9970 ( .A1(n8955), .A2(n8324), .ZN(n8325) );
  OAI211_X1 U9971 ( .C1(n8327), .C2(n8393), .A(n8326), .B(n8325), .ZN(P2_U3168) );
  INV_X1 U9972 ( .A(n8915), .ZN(n8681) );
  INV_X1 U9973 ( .A(n8328), .ZN(n8330) );
  NOR3_X1 U9974 ( .A1(n8331), .A2(n8330), .A3(n8329), .ZN(n8333) );
  OAI21_X1 U9975 ( .B1(n8333), .B2(n8332), .A(n8381), .ZN(n8339) );
  INV_X1 U9976 ( .A(n8683), .ZN(n8335) );
  AOI22_X1 U9977 ( .A1(n8706), .A2(n8402), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8334) );
  OAI21_X1 U9978 ( .B1(n8335), .B2(n8399), .A(n8334), .ZN(n8336) );
  AOI21_X1 U9979 ( .B1(n8679), .B2(n8337), .A(n8336), .ZN(n8338) );
  OAI211_X1 U9980 ( .C1(n8681), .C2(n8405), .A(n8339), .B(n8338), .ZN(P2_U3169) );
  INV_X1 U9981 ( .A(n8737), .ZN(n8938) );
  INV_X1 U9982 ( .A(n8340), .ZN(n8342) );
  NOR3_X1 U9983 ( .A1(n8343), .A2(n8342), .A3(n8341), .ZN(n8345) );
  OAI21_X1 U9984 ( .B1(n8345), .B2(n8344), .A(n8381), .ZN(n8349) );
  NOR2_X1 U9985 ( .A1(n8754), .A2(n8384), .ZN(n8347) );
  INV_X1 U9986 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10658) );
  OAI22_X1 U9987 ( .A1(n8733), .A2(n8398), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10658), .ZN(n8346) );
  AOI211_X1 U9988 ( .C1(n8736), .C2(n8389), .A(n8347), .B(n8346), .ZN(n8348)
         );
  OAI211_X1 U9989 ( .C1(n8938), .C2(n8405), .A(n8349), .B(n8348), .ZN(P2_U3173) );
  INV_X1 U9990 ( .A(n8927), .ZN(n8364) );
  INV_X1 U9991 ( .A(n8350), .ZN(n8352) );
  NOR3_X1 U9992 ( .A1(n8353), .A2(n8352), .A3(n8351), .ZN(n8359) );
  NAND2_X1 U9993 ( .A1(n8355), .A2(n8354), .ZN(n8357) );
  AND2_X1 U9994 ( .A1(n8357), .A2(n8356), .ZN(n8358) );
  OAI21_X1 U9995 ( .B1(n8359), .B2(n8358), .A(n8381), .ZN(n8363) );
  AOI22_X1 U9996 ( .A1(n8707), .A2(n8402), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8360) );
  OAI21_X1 U9997 ( .B1(n8219), .B2(n8398), .A(n8360), .ZN(n8361) );
  AOI21_X1 U9998 ( .B1(n8710), .B2(n8389), .A(n8361), .ZN(n8362) );
  OAI211_X1 U9999 ( .C1(n8364), .C2(n8405), .A(n8363), .B(n8362), .ZN(P2_U3175) );
  INV_X1 U10000 ( .A(n8365), .ZN(n8952) );
  INV_X1 U10001 ( .A(n8366), .ZN(n8368) );
  NOR3_X1 U10002 ( .A1(n8369), .A2(n8368), .A3(n8367), .ZN(n8371) );
  OAI21_X1 U10003 ( .B1(n8371), .B2(n8370), .A(n8381), .ZN(n8375) );
  NOR2_X1 U10004 ( .A1(n8753), .A2(n8384), .ZN(n8373) );
  NAND2_X1 U10005 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8564) );
  OAI21_X1 U10006 ( .B1(n8754), .B2(n8398), .A(n8564), .ZN(n8372) );
  AOI211_X1 U10007 ( .C1(n8758), .C2(n8389), .A(n8373), .B(n8372), .ZN(n8374)
         );
  OAI211_X1 U10008 ( .C1(n8952), .C2(n8405), .A(n8375), .B(n8374), .ZN(
        P2_U3178) );
  INV_X1 U10009 ( .A(n8903), .ZN(n8392) );
  INV_X1 U10010 ( .A(n8376), .ZN(n8378) );
  NOR3_X1 U10011 ( .A1(n8379), .A2(n8378), .A3(n8377), .ZN(n8383) );
  INV_X1 U10012 ( .A(n8380), .ZN(n8382) );
  OAI21_X1 U10013 ( .B1(n8383), .B2(n8382), .A(n8381), .ZN(n8391) );
  OAI22_X1 U10014 ( .A1(n8385), .A2(n8384), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10448), .ZN(n8388) );
  NOR2_X1 U10015 ( .A1(n8386), .A2(n8398), .ZN(n8387) );
  AOI211_X1 U10016 ( .C1(n8648), .C2(n8389), .A(n8388), .B(n8387), .ZN(n8390)
         );
  OAI211_X1 U10017 ( .C1(n8392), .C2(n8405), .A(n8391), .B(n8390), .ZN(
        P2_U3180) );
  INV_X1 U10018 ( .A(n8967), .ZN(n8406) );
  AOI21_X1 U10019 ( .B1(n8395), .B2(n8394), .A(n8393), .ZN(n8397) );
  NAND2_X1 U10020 ( .A1(n8397), .A2(n8396), .ZN(n8404) );
  NAND2_X1 U10021 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8496) );
  OAI21_X1 U10022 ( .B1(n8398), .B2(n8769), .A(n8496), .ZN(n8401) );
  NOR2_X1 U10023 ( .A1(n8399), .A2(n8798), .ZN(n8400) );
  AOI211_X1 U10024 ( .C1(n8402), .C2(n8794), .A(n8401), .B(n8400), .ZN(n8403)
         );
  OAI211_X1 U10025 ( .C1(n8406), .C2(n8405), .A(n8404), .B(n8403), .ZN(
        P2_U3181) );
  MUX2_X1 U10026 ( .A(n8407), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8561), .Z(
        P2_U3521) );
  MUX2_X1 U10027 ( .A(n8623), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8561), .Z(
        P2_U3520) );
  MUX2_X1 U10028 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8664), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10029 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8679), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10030 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8693), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10031 ( .A(n8706), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8561), .Z(
        P2_U3514) );
  MUX2_X1 U10032 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8723), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10033 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8707), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10034 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8408), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10035 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8744), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10036 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8784), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10037 ( .A(n8795), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8561), .Z(
        P2_U3507) );
  MUX2_X1 U10038 ( .A(n8811), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8561), .Z(
        P2_U3506) );
  MUX2_X1 U10039 ( .A(n8794), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8561), .Z(
        P2_U3505) );
  MUX2_X1 U10040 ( .A(n8809), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8561), .Z(
        P2_U3504) );
  MUX2_X1 U10041 ( .A(n8409), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8561), .Z(
        P2_U3503) );
  MUX2_X1 U10042 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8410), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U10043 ( .A(n8411), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8561), .Z(
        P2_U3501) );
  MUX2_X1 U10044 ( .A(n8412), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8561), .Z(
        P2_U3500) );
  MUX2_X1 U10045 ( .A(n8413), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8561), .Z(
        P2_U3499) );
  MUX2_X1 U10046 ( .A(n8414), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8561), .Z(
        P2_U3498) );
  MUX2_X1 U10047 ( .A(n8415), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8561), .Z(
        P2_U3497) );
  MUX2_X1 U10048 ( .A(n8416), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8561), .Z(
        P2_U3496) );
  MUX2_X1 U10049 ( .A(n8417), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8561), .Z(
        P2_U3495) );
  MUX2_X1 U10050 ( .A(n8418), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8561), .Z(
        P2_U3494) );
  MUX2_X1 U10051 ( .A(n8419), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8561), .Z(
        P2_U3493) );
  MUX2_X1 U10052 ( .A(n8420), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8561), .Z(
        P2_U3492) );
  MUX2_X1 U10053 ( .A(n6381), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8561), .Z(
        P2_U3491) );
  INV_X1 U10054 ( .A(n10152), .ZN(n8425) );
  OAI21_X1 U10055 ( .B1(n8423), .B2(n8422), .A(n8421), .ZN(n8424) );
  AOI22_X1 U10056 ( .A1(n10145), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(n8425), .B2(
        n8424), .ZN(n8437) );
  OAI21_X1 U10057 ( .B1(n8428), .B2(n8427), .A(n8426), .ZN(n8429) );
  AOI22_X1 U10058 ( .A1(n10161), .A2(n8429), .B1(P2_U3151), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n8436) );
  OAI211_X1 U10059 ( .C1(n8432), .C2(n8431), .A(n8430), .B(n10146), .ZN(n8435)
         );
  NAND2_X1 U10060 ( .A1(n10155), .A2(n8433), .ZN(n8434) );
  NAND4_X1 U10061 ( .A1(n8437), .A2(n8436), .A3(n8435), .A4(n8434), .ZN(
        P2_U3184) );
  AOI21_X1 U10062 ( .B1(n8440), .B2(n8439), .A(n8460), .ZN(n8458) );
  MUX2_X1 U10063 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8555), .Z(n8463) );
  XNOR2_X1 U10064 ( .A(n8463), .B(n8473), .ZN(n8445) );
  OR2_X1 U10065 ( .A1(n8441), .A2(n8447), .ZN(n8443) );
  NAND2_X1 U10066 ( .A1(n8443), .A2(n8442), .ZN(n8444) );
  NAND2_X1 U10067 ( .A1(n8445), .A2(n8444), .ZN(n8465) );
  OAI21_X1 U10068 ( .B1(n8445), .B2(n8444), .A(n8465), .ZN(n8455) );
  INV_X1 U10069 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n10270) );
  NOR2_X1 U10070 ( .A1(n8565), .A2(n10270), .ZN(n8454) );
  XNOR2_X1 U10071 ( .A(n8473), .B(n8472), .ZN(n8449) );
  NOR2_X1 U10072 ( .A1(n8448), .A2(n8449), .ZN(n8474) );
  AOI21_X1 U10073 ( .B1(n8449), .B2(n8448), .A(n8474), .ZN(n8452) );
  INV_X1 U10074 ( .A(n8450), .ZN(n8451) );
  OAI21_X1 U10075 ( .B1(n8571), .B2(n8452), .A(n8451), .ZN(n8453) );
  AOI211_X1 U10076 ( .C1(n10146), .C2(n8455), .A(n8454), .B(n8453), .ZN(n8457)
         );
  NAND2_X1 U10077 ( .A1(n10155), .A2(n8473), .ZN(n8456) );
  OAI211_X1 U10078 ( .C1(n8458), .C2(n10152), .A(n8457), .B(n8456), .ZN(
        P2_U3195) );
  NOR2_X1 U10079 ( .A1(n8473), .A2(n8459), .ZN(n8461) );
  AOI22_X1 U10080 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8482), .B1(n8492), .B2(
        n8874), .ZN(n8462) );
  AOI21_X1 U10081 ( .B1(n4590), .B2(n8462), .A(n8485), .ZN(n8484) );
  INV_X1 U10082 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n10274) );
  MUX2_X1 U10083 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8555), .Z(n8487) );
  XNOR2_X1 U10084 ( .A(n8487), .B(n8482), .ZN(n8468) );
  INV_X1 U10085 ( .A(n8463), .ZN(n8464) );
  NAND2_X1 U10086 ( .A1(n8473), .A2(n8464), .ZN(n8466) );
  NAND2_X1 U10087 ( .A1(n8466), .A2(n8465), .ZN(n8467) );
  NAND2_X1 U10088 ( .A1(n8468), .A2(n8467), .ZN(n8488) );
  OAI21_X1 U10089 ( .B1(n8468), .B2(n8467), .A(n8488), .ZN(n8469) );
  NAND2_X1 U10090 ( .A1(n8469), .A2(n10146), .ZN(n8471) );
  OAI211_X1 U10091 ( .C1(n8565), .C2(n10274), .A(n8471), .B(n8470), .ZN(n8481)
         );
  NOR2_X1 U10092 ( .A1(n8473), .A2(n8472), .ZN(n8475) );
  NOR2_X1 U10093 ( .A1(n8475), .A2(n8474), .ZN(n8478) );
  MUX2_X1 U10094 ( .A(n6213), .B(P2_REG2_REG_14__SCAN_IN), .S(n8482), .Z(n8476) );
  INV_X1 U10095 ( .A(n8476), .ZN(n8477) );
  AOI21_X1 U10096 ( .B1(n8478), .B2(n8477), .A(n8494), .ZN(n8479) );
  NOR2_X1 U10097 ( .A1(n8479), .A2(n8571), .ZN(n8480) );
  AOI211_X1 U10098 ( .C1(n10155), .C2(n8482), .A(n8481), .B(n8480), .ZN(n8483)
         );
  OAI21_X1 U10099 ( .B1(n8484), .B2(n10152), .A(n8483), .ZN(P2_U3196) );
  XOR2_X1 U10100 ( .A(n8504), .B(n8509), .Z(n8486) );
  NOR2_X1 U10101 ( .A1(n8871), .A2(n8486), .ZN(n8505) );
  AOI21_X1 U10102 ( .B1(n8871), .B2(n8486), .A(n8505), .ZN(n8503) );
  MUX2_X1 U10103 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8555), .Z(n8510) );
  XNOR2_X1 U10104 ( .A(n8510), .B(n8519), .ZN(n8491) );
  OR2_X1 U10105 ( .A1(n8487), .A2(n8492), .ZN(n8489) );
  NAND2_X1 U10106 ( .A1(n8489), .A2(n8488), .ZN(n8490) );
  NAND2_X1 U10107 ( .A1(n8491), .A2(n8490), .ZN(n8511) );
  OAI21_X1 U10108 ( .B1(n8491), .B2(n8490), .A(n8511), .ZN(n8500) );
  INV_X1 U10109 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n10278) );
  NOR2_X1 U10110 ( .A1(n8565), .A2(n10278), .ZN(n8499) );
  XNOR2_X1 U10111 ( .A(n8519), .B(n8518), .ZN(n8495) );
  AOI21_X1 U10112 ( .B1(n8495), .B2(n8797), .A(n8520), .ZN(n8497) );
  OAI21_X1 U10113 ( .B1(n8571), .B2(n8497), .A(n8496), .ZN(n8498) );
  AOI211_X1 U10114 ( .C1(n10146), .C2(n8500), .A(n8499), .B(n8498), .ZN(n8502)
         );
  NAND2_X1 U10115 ( .A1(n10155), .A2(n8519), .ZN(n8501) );
  OAI211_X1 U10116 ( .C1(n8503), .C2(n10152), .A(n8502), .B(n8501), .ZN(
        P2_U3197) );
  NOR2_X1 U10117 ( .A1(n8519), .A2(n8504), .ZN(n8506) );
  NOR2_X1 U10118 ( .A1(n8506), .A2(n8505), .ZN(n8508) );
  AOI22_X1 U10119 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8527), .B1(n8537), .B2(
        n8868), .ZN(n8507) );
  NOR2_X1 U10120 ( .A1(n8508), .A2(n8507), .ZN(n8530) );
  AOI21_X1 U10121 ( .B1(n8508), .B2(n8507), .A(n8530), .ZN(n8529) );
  INV_X1 U10122 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n10282) );
  MUX2_X1 U10123 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8555), .Z(n8532) );
  XNOR2_X1 U10124 ( .A(n8532), .B(n8527), .ZN(n8514) );
  OR2_X1 U10125 ( .A1(n8510), .A2(n8509), .ZN(n8512) );
  NAND2_X1 U10126 ( .A1(n8512), .A2(n8511), .ZN(n8513) );
  NAND2_X1 U10127 ( .A1(n8514), .A2(n8513), .ZN(n8533) );
  OAI21_X1 U10128 ( .B1(n8514), .B2(n8513), .A(n8533), .ZN(n8515) );
  NAND2_X1 U10129 ( .A1(n8515), .A2(n10146), .ZN(n8517) );
  OAI211_X1 U10130 ( .C1(n8565), .C2(n10282), .A(n8517), .B(n8516), .ZN(n8526)
         );
  NOR2_X1 U10131 ( .A1(n8519), .A2(n8518), .ZN(n8521) );
  NOR2_X1 U10132 ( .A1(n8537), .A2(n8787), .ZN(n8522) );
  AOI21_X1 U10133 ( .B1(n8537), .B2(n8787), .A(n8522), .ZN(n8523) );
  AOI21_X1 U10134 ( .B1(n4581), .B2(n8523), .A(n8538), .ZN(n8524) );
  NOR2_X1 U10135 ( .A1(n8524), .A2(n8571), .ZN(n8525) );
  AOI211_X1 U10136 ( .C1(n10155), .C2(n8527), .A(n8526), .B(n8525), .ZN(n8528)
         );
  OAI21_X1 U10137 ( .B1(n8529), .B2(n10152), .A(n8528), .ZN(P2_U3198) );
  XNOR2_X1 U10138 ( .A(n8567), .B(n8548), .ZN(n8531) );
  AOI21_X1 U10139 ( .B1(n8865), .B2(n8531), .A(n8549), .ZN(n8547) );
  MUX2_X1 U10140 ( .A(n8775), .B(n8865), .S(n8555), .Z(n8554) );
  XOR2_X1 U10141 ( .A(n8567), .B(n8554), .Z(n8536) );
  OR2_X1 U10142 ( .A1(n8537), .A2(n8532), .ZN(n8534) );
  NAND2_X1 U10143 ( .A1(n8534), .A2(n8533), .ZN(n8535) );
  NAND2_X1 U10144 ( .A1(n8536), .A2(n8535), .ZN(n8552) );
  OAI21_X1 U10145 ( .B1(n8536), .B2(n8535), .A(n8552), .ZN(n8544) );
  INV_X1 U10146 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n10286) );
  NOR2_X1 U10147 ( .A1(n8565), .A2(n10286), .ZN(n8543) );
  XNOR2_X1 U10148 ( .A(n8567), .B(n8566), .ZN(n8539) );
  AOI21_X1 U10149 ( .B1(n8539), .B2(n8775), .A(n8569), .ZN(n8541) );
  OAI21_X1 U10150 ( .B1(n8571), .B2(n8541), .A(n8540), .ZN(n8542) );
  AOI211_X1 U10151 ( .C1(n10146), .C2(n8544), .A(n8543), .B(n8542), .ZN(n8546)
         );
  NAND2_X1 U10152 ( .A1(n10155), .A2(n8567), .ZN(n8545) );
  OAI211_X1 U10153 ( .C1(n8547), .C2(n10152), .A(n8546), .B(n8545), .ZN(
        P2_U3199) );
  NOR2_X1 U10154 ( .A1(n8567), .A2(n8548), .ZN(n8550) );
  NAND2_X1 U10155 ( .A1(n8586), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8577) );
  OAI21_X1 U10156 ( .B1(n8586), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8577), .ZN(
        n8551) );
  AOI21_X1 U10157 ( .B1(n4580), .B2(n8551), .A(n8578), .ZN(n8576) );
  INV_X1 U10158 ( .A(n8552), .ZN(n8553) );
  MUX2_X1 U10159 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8555), .Z(n8557) );
  AND2_X1 U10160 ( .A1(n8556), .A2(n8557), .ZN(n8587) );
  INV_X1 U10161 ( .A(n8556), .ZN(n8559) );
  INV_X1 U10162 ( .A(n8557), .ZN(n8558) );
  NAND2_X1 U10163 ( .A1(n8559), .A2(n8558), .ZN(n8585) );
  INV_X1 U10164 ( .A(n8585), .ZN(n8560) );
  OAI21_X1 U10165 ( .B1(n8561), .B2(n8562), .A(n8598), .ZN(n8573) );
  INV_X1 U10166 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10309) );
  NAND3_X1 U10167 ( .A1(n8562), .A2(n10146), .A3(n8586), .ZN(n8563) );
  OAI211_X1 U10168 ( .C1(n8565), .C2(n10309), .A(n8564), .B(n8563), .ZN(n8572)
         );
  NOR2_X1 U10169 ( .A1(n8567), .A2(n8566), .ZN(n8568) );
  NAND2_X1 U10170 ( .A1(n8586), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8581) );
  OAI21_X1 U10171 ( .B1(n8586), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8581), .ZN(
        n8570) );
  OAI21_X1 U10172 ( .B1(n8576), .B2(n10152), .A(n8575), .ZN(P2_U3200) );
  XNOR2_X1 U10173 ( .A(n8597), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8590) );
  INV_X1 U10174 ( .A(n8590), .ZN(n8579) );
  XNOR2_X1 U10175 ( .A(n8580), .B(n8579), .ZN(n8603) );
  INV_X1 U10176 ( .A(n8581), .ZN(n8582) );
  XNOR2_X1 U10177 ( .A(n8597), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8589) );
  XNOR2_X1 U10178 ( .A(n8584), .B(n8589), .ZN(n8601) );
  OAI21_X1 U10179 ( .B1(n8587), .B2(n8586), .A(n8585), .ZN(n8592) );
  MUX2_X1 U10180 ( .A(n8590), .B(n8589), .S(n8588), .Z(n8591) );
  XNOR2_X1 U10181 ( .A(n8592), .B(n8591), .ZN(n8594) );
  NOR2_X1 U10182 ( .A1(n8594), .A2(n8593), .ZN(n8600) );
  NAND2_X1 U10183 ( .A1(n10145), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8596) );
  OAI211_X1 U10184 ( .C1(n8598), .C2(n8597), .A(n8596), .B(n8595), .ZN(n8599)
         );
  OAI21_X1 U10185 ( .B1(n8603), .B2(n10152), .A(n8602), .ZN(P2_U3201) );
  INV_X1 U10186 ( .A(n8823), .ZN(n8885) );
  INV_X1 U10187 ( .A(n8604), .ZN(n8605) );
  NAND2_X1 U10188 ( .A1(n8605), .A2(n8800), .ZN(n8612) );
  NAND2_X1 U10189 ( .A1(n8607), .A2(n8606), .ZN(n8883) );
  AOI21_X1 U10190 ( .B1(n8612), .B2(n8883), .A(n8636), .ZN(n8609) );
  AOI21_X1 U10191 ( .B1(n8636), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8609), .ZN(
        n8608) );
  OAI21_X1 U10192 ( .B1(n8885), .B2(n10171), .A(n8608), .ZN(P2_U3202) );
  AOI21_X1 U10193 ( .B1(n8636), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8609), .ZN(
        n8610) );
  OAI21_X1 U10194 ( .B1(n8888), .B2(n10171), .A(n8610), .ZN(P2_U3203) );
  NAND2_X1 U10195 ( .A1(n8611), .A2(n10174), .ZN(n8617) );
  OAI21_X1 U10196 ( .B1(n10174), .B2(n8613), .A(n8612), .ZN(n8614) );
  AOI21_X1 U10197 ( .B1(n8615), .B2(n8801), .A(n8614), .ZN(n8616) );
  OAI211_X1 U10198 ( .C1(n8619), .C2(n8618), .A(n8617), .B(n8616), .ZN(
        P2_U3204) );
  XNOR2_X1 U10199 ( .A(n8620), .B(n8622), .ZN(n8894) );
  MUX2_X1 U10200 ( .A(n8624), .B(n8889), .S(n10174), .Z(n8627) );
  AOI22_X1 U10201 ( .A1(n8891), .A2(n8801), .B1(n8800), .B2(n8625), .ZN(n8626)
         );
  OAI211_X1 U10202 ( .C1(n8894), .C2(n8822), .A(n8627), .B(n8626), .ZN(
        P2_U3205) );
  XNOR2_X1 U10203 ( .A(n8628), .B(n8629), .ZN(n8900) );
  OAI21_X1 U10204 ( .B1(n8630), .B2(n8629), .A(n8813), .ZN(n8632) );
  AOI22_X1 U10205 ( .A1(n8633), .A2(n8810), .B1(n8808), .B2(n8664), .ZN(n8634)
         );
  MUX2_X1 U10206 ( .A(n8896), .B(n8637), .S(n8636), .Z(n8640) );
  AOI22_X1 U10207 ( .A1(n8897), .A2(n8801), .B1(n8800), .B2(n8638), .ZN(n8639)
         );
  OAI211_X1 U10208 ( .C1(n8900), .C2(n8822), .A(n8640), .B(n8639), .ZN(
        P2_U3206) );
  XNOR2_X1 U10209 ( .A(n8642), .B(n8641), .ZN(n8906) );
  XNOR2_X1 U10210 ( .A(n8644), .B(n8643), .ZN(n8646) );
  AOI222_X1 U10211 ( .A1(n8813), .A2(n8646), .B1(n8679), .B2(n8808), .C1(n8645), .C2(n8810), .ZN(n8901) );
  MUX2_X1 U10212 ( .A(n8647), .B(n8901), .S(n8817), .Z(n8650) );
  AOI22_X1 U10213 ( .A1(n8903), .A2(n8801), .B1(n8800), .B2(n8648), .ZN(n8649)
         );
  OAI211_X1 U10214 ( .C1(n8906), .C2(n8822), .A(n8650), .B(n8649), .ZN(
        P2_U3207) );
  NAND2_X1 U10215 ( .A1(n8652), .A2(n8651), .ZN(n8705) );
  NAND2_X1 U10216 ( .A1(n8705), .A2(n8653), .ZN(n8692) );
  NAND2_X1 U10217 ( .A1(n8692), .A2(n8654), .ZN(n8656) );
  NAND2_X1 U10218 ( .A1(n8656), .A2(n8655), .ZN(n8678) );
  AND2_X1 U10219 ( .A1(n8660), .A2(n8658), .ZN(n8663) );
  NAND2_X1 U10220 ( .A1(n8660), .A2(n8659), .ZN(n8661) );
  OAI21_X1 U10221 ( .B1(n8663), .B2(n8662), .A(n8661), .ZN(n8665) );
  AOI222_X1 U10222 ( .A1(n8813), .A2(n8665), .B1(n8693), .B2(n8808), .C1(n8664), .C2(n8810), .ZN(n8907) );
  INV_X1 U10223 ( .A(n8815), .ZN(n8667) );
  AOI22_X1 U10224 ( .A1(n8909), .A2(n8667), .B1(n8800), .B2(n8666), .ZN(n8668)
         );
  AOI21_X1 U10225 ( .B1(n8907), .B2(n8668), .A(n8636), .ZN(n8673) );
  XNOR2_X1 U10226 ( .A(n8670), .B(n8669), .ZN(n8912) );
  OAI22_X1 U10227 ( .A1(n8912), .A2(n8822), .B1(n8671), .B2(n8817), .ZN(n8672)
         );
  OR2_X1 U10228 ( .A1(n8673), .A2(n8672), .ZN(P2_U3208) );
  NAND2_X1 U10229 ( .A1(n8675), .A2(n8674), .ZN(n8676) );
  XNOR2_X1 U10230 ( .A(n8676), .B(n8677), .ZN(n8918) );
  XNOR2_X1 U10231 ( .A(n8678), .B(n8677), .ZN(n8680) );
  AOI222_X1 U10232 ( .A1(n8813), .A2(n8680), .B1(n8679), .B2(n8810), .C1(n8706), .C2(n8808), .ZN(n8913) );
  OAI21_X1 U10233 ( .B1(n8681), .B2(n8815), .A(n8913), .ZN(n8682) );
  NAND2_X1 U10234 ( .A1(n8682), .A2(n10174), .ZN(n8685) );
  AOI22_X1 U10235 ( .A1(n8683), .A2(n8800), .B1(n8636), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n8684) );
  OAI211_X1 U10236 ( .C1(n8918), .C2(n8822), .A(n8685), .B(n8684), .ZN(
        P2_U3209) );
  NAND2_X1 U10237 ( .A1(n8686), .A2(n8687), .ZN(n8689) );
  XNOR2_X1 U10238 ( .A(n8692), .B(n8691), .ZN(n8694) );
  AOI222_X1 U10239 ( .A1(n8813), .A2(n8694), .B1(n8693), .B2(n8810), .C1(n8723), .C2(n8808), .ZN(n8919) );
  MUX2_X1 U10240 ( .A(n8695), .B(n8919), .S(n10174), .Z(n8698) );
  AOI22_X1 U10241 ( .A1(n8921), .A2(n8801), .B1(n8800), .B2(n8696), .ZN(n8697)
         );
  OAI211_X1 U10242 ( .C1(n8924), .C2(n8822), .A(n8698), .B(n8697), .ZN(
        P2_U3210) );
  AND2_X1 U10243 ( .A1(n4574), .A2(n8700), .ZN(n8701) );
  XNOR2_X1 U10244 ( .A(n8701), .B(n8703), .ZN(n8930) );
  NAND3_X1 U10245 ( .A1(n8722), .A2(n8703), .A3(n8702), .ZN(n8704) );
  NAND2_X1 U10246 ( .A1(n8705), .A2(n8704), .ZN(n8708) );
  AOI222_X1 U10247 ( .A1(n8813), .A2(n8708), .B1(n8707), .B2(n8808), .C1(n8706), .C2(n8810), .ZN(n8925) );
  MUX2_X1 U10248 ( .A(n8709), .B(n8925), .S(n10174), .Z(n8712) );
  AOI22_X1 U10249 ( .A1(n8927), .A2(n8801), .B1(n8800), .B2(n8710), .ZN(n8711)
         );
  OAI211_X1 U10250 ( .C1(n8930), .C2(n8822), .A(n8712), .B(n8711), .ZN(
        P2_U3211) );
  NAND2_X1 U10251 ( .A1(n8686), .A2(n8713), .ZN(n8715) );
  NAND2_X1 U10252 ( .A1(n8715), .A2(n8714), .ZN(n8716) );
  XNOR2_X1 U10253 ( .A(n8716), .B(n8718), .ZN(n8936) );
  INV_X1 U10254 ( .A(n8718), .ZN(n8720) );
  NAND3_X1 U10255 ( .A1(n8717), .A2(n8720), .A3(n8719), .ZN(n8721) );
  NAND2_X1 U10256 ( .A1(n8722), .A2(n8721), .ZN(n8724) );
  AOI222_X1 U10257 ( .A1(n8813), .A2(n8724), .B1(n8745), .B2(n8808), .C1(n8723), .C2(n8810), .ZN(n8931) );
  MUX2_X1 U10258 ( .A(n8725), .B(n8931), .S(n10174), .Z(n8728) );
  AOI22_X1 U10259 ( .A1(n8933), .A2(n8801), .B1(n8800), .B2(n8726), .ZN(n8727)
         );
  OAI211_X1 U10260 ( .C1(n8936), .C2(n8822), .A(n8728), .B(n8727), .ZN(
        P2_U3212) );
  XOR2_X1 U10261 ( .A(n8731), .B(n8686), .Z(n8939) );
  INV_X1 U10262 ( .A(n8717), .ZN(n8729) );
  AOI21_X1 U10263 ( .B1(n8731), .B2(n8730), .A(n8729), .ZN(n8732) );
  OAI222_X1 U10264 ( .A1(n8770), .A2(n8733), .B1(n8768), .B2(n8754), .C1(n8765), .C2(n8732), .ZN(n8937) );
  INV_X1 U10265 ( .A(n8937), .ZN(n8734) );
  MUX2_X1 U10266 ( .A(n8735), .B(n8734), .S(n8817), .Z(n8739) );
  AOI22_X1 U10267 ( .A1(n8737), .A2(n8801), .B1(n8800), .B2(n8736), .ZN(n8738)
         );
  OAI211_X1 U10268 ( .C1(n8939), .C2(n8822), .A(n8739), .B(n8738), .ZN(
        P2_U3213) );
  OAI21_X1 U10269 ( .B1(n8741), .B2(n8743), .A(n8740), .ZN(n8947) );
  INV_X1 U10270 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8747) );
  XNOR2_X1 U10271 ( .A(n8742), .B(n8743), .ZN(n8746) );
  AOI222_X1 U10272 ( .A1(n8813), .A2(n8746), .B1(n8745), .B2(n8810), .C1(n8744), .C2(n8808), .ZN(n8942) );
  MUX2_X1 U10273 ( .A(n8747), .B(n8942), .S(n10174), .Z(n8750) );
  AOI22_X1 U10274 ( .A1(n8944), .A2(n8801), .B1(n8800), .B2(n8748), .ZN(n8749)
         );
  OAI211_X1 U10275 ( .C1(n8947), .C2(n8822), .A(n8750), .B(n8749), .ZN(
        P2_U3214) );
  XNOR2_X1 U10276 ( .A(n8751), .B(n8755), .ZN(n8752) );
  OAI222_X1 U10277 ( .A1(n8770), .A2(n8754), .B1(n8768), .B2(n8753), .C1(n8752), .C2(n8765), .ZN(n8859) );
  INV_X1 U10278 ( .A(n8860), .ZN(n8757) );
  AND2_X1 U10279 ( .A1(n8756), .A2(n8755), .ZN(n8858) );
  NOR3_X1 U10280 ( .A1(n8757), .A2(n8858), .A3(n8822), .ZN(n8761) );
  AOI22_X1 U10281 ( .A1(n8636), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8800), .B2(
        n8758), .ZN(n8759) );
  OAI21_X1 U10282 ( .B1(n8952), .B2(n10171), .A(n8759), .ZN(n8760) );
  AOI211_X1 U10283 ( .C1(n8859), .C2(n8817), .A(n8761), .B(n8760), .ZN(n8762)
         );
  INV_X1 U10284 ( .A(n8762), .ZN(P2_U3215) );
  XNOR2_X1 U10285 ( .A(n8763), .B(n8766), .ZN(n8958) );
  INV_X1 U10286 ( .A(n8764), .ZN(n8767) );
  AOI21_X1 U10287 ( .B1(n8767), .B2(n8766), .A(n8765), .ZN(n8774) );
  OAI22_X1 U10288 ( .A1(n8771), .A2(n8770), .B1(n8769), .B2(n8768), .ZN(n8772)
         );
  AOI21_X1 U10289 ( .B1(n8774), .B2(n8773), .A(n8772), .ZN(n8953) );
  MUX2_X1 U10290 ( .A(n8775), .B(n8953), .S(n8817), .Z(n8778) );
  AOI22_X1 U10291 ( .A1(n8955), .A2(n8801), .B1(n8800), .B2(n8776), .ZN(n8777)
         );
  OAI211_X1 U10292 ( .C1(n8958), .C2(n8822), .A(n8778), .B(n8777), .ZN(
        P2_U3216) );
  XNOR2_X1 U10293 ( .A(n8780), .B(n8779), .ZN(n8964) );
  OAI211_X1 U10294 ( .C1(n8783), .C2(n8782), .A(n8781), .B(n8813), .ZN(n8786)
         );
  AOI22_X1 U10295 ( .A1(n8784), .A2(n8810), .B1(n8808), .B2(n8811), .ZN(n8785)
         );
  MUX2_X1 U10296 ( .A(n8960), .B(n8787), .S(n8636), .Z(n8790) );
  AOI22_X1 U10297 ( .A1(n8961), .A2(n8801), .B1(n8800), .B2(n8788), .ZN(n8789)
         );
  OAI211_X1 U10298 ( .C1(n8964), .C2(n8822), .A(n8790), .B(n8789), .ZN(
        P2_U3217) );
  XOR2_X1 U10299 ( .A(n8793), .B(n8791), .Z(n8970) );
  XNOR2_X1 U10300 ( .A(n8792), .B(n8793), .ZN(n8796) );
  AOI222_X1 U10301 ( .A1(n8813), .A2(n8796), .B1(n8795), .B2(n8810), .C1(n8794), .C2(n8808), .ZN(n8965) );
  MUX2_X1 U10302 ( .A(n8797), .B(n8965), .S(n10174), .Z(n8803) );
  INV_X1 U10303 ( .A(n8798), .ZN(n8799) );
  AOI22_X1 U10304 ( .A1(n8967), .A2(n8801), .B1(n8800), .B2(n8799), .ZN(n8802)
         );
  OAI211_X1 U10305 ( .C1(n8970), .C2(n8822), .A(n8803), .B(n8802), .ZN(
        P2_U3218) );
  XNOR2_X1 U10306 ( .A(n8805), .B(n8804), .ZN(n8978) );
  XNOR2_X1 U10307 ( .A(n8807), .B(n8806), .ZN(n8812) );
  AOI222_X1 U10308 ( .A1(n8813), .A2(n8812), .B1(n8811), .B2(n8810), .C1(n8809), .C2(n8808), .ZN(n8971) );
  INV_X1 U10309 ( .A(n8971), .ZN(n8819) );
  INV_X1 U10310 ( .A(n8974), .ZN(n8816) );
  OAI22_X1 U10311 ( .A1(n8816), .A2(n8815), .B1(n8814), .B2(n10169), .ZN(n8818) );
  OAI21_X1 U10312 ( .B1(n8819), .B2(n8818), .A(n8817), .ZN(n8821) );
  NAND2_X1 U10313 ( .A1(n8636), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8820) );
  OAI211_X1 U10314 ( .C1(n8978), .C2(n8822), .A(n8821), .B(n8820), .ZN(
        P2_U3219) );
  NAND2_X1 U10315 ( .A1(n8823), .A2(n8875), .ZN(n8825) );
  INV_X1 U10316 ( .A(n8883), .ZN(n8824) );
  NAND2_X1 U10317 ( .A1(n8824), .A2(n10233), .ZN(n8827) );
  OAI211_X1 U10318 ( .C1(n10233), .C2(n7470), .A(n8825), .B(n8827), .ZN(
        P2_U3490) );
  NAND2_X1 U10319 ( .A1(n8826), .A2(n8875), .ZN(n8828) );
  OAI211_X1 U10320 ( .C1(n10233), .C2(n6447), .A(n8828), .B(n8827), .ZN(
        P2_U3489) );
  INV_X1 U10321 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8829) );
  MUX2_X1 U10322 ( .A(n8829), .B(n8889), .S(n10233), .Z(n8831) );
  NAND2_X1 U10323 ( .A1(n8891), .A2(n8875), .ZN(n8830) );
  OAI211_X1 U10324 ( .C1(n8894), .C2(n8878), .A(n8831), .B(n8830), .ZN(
        P2_U3487) );
  INV_X1 U10325 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8832) );
  MUX2_X1 U10326 ( .A(n8832), .B(n8896), .S(n10233), .Z(n8834) );
  NAND2_X1 U10327 ( .A1(n8897), .A2(n8875), .ZN(n8833) );
  OAI211_X1 U10328 ( .C1(n8900), .C2(n8878), .A(n8834), .B(n8833), .ZN(
        P2_U3486) );
  INV_X1 U10329 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8835) );
  MUX2_X1 U10330 ( .A(n8835), .B(n8901), .S(n10233), .Z(n8837) );
  NAND2_X1 U10331 ( .A1(n8903), .A2(n8875), .ZN(n8836) );
  OAI211_X1 U10332 ( .C1(n8906), .C2(n8878), .A(n8837), .B(n8836), .ZN(
        P2_U3485) );
  INV_X1 U10333 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8838) );
  MUX2_X1 U10334 ( .A(n8838), .B(n8907), .S(n10233), .Z(n8840) );
  NAND2_X1 U10335 ( .A1(n8909), .A2(n8875), .ZN(n8839) );
  OAI211_X1 U10336 ( .C1(n8912), .C2(n8878), .A(n8840), .B(n8839), .ZN(
        P2_U3484) );
  INV_X1 U10337 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8841) );
  MUX2_X1 U10338 ( .A(n8841), .B(n8913), .S(n10233), .Z(n8843) );
  NAND2_X1 U10339 ( .A1(n8915), .A2(n8875), .ZN(n8842) );
  OAI211_X1 U10340 ( .C1(n8878), .C2(n8918), .A(n8843), .B(n8842), .ZN(
        P2_U3483) );
  INV_X1 U10341 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8844) );
  MUX2_X1 U10342 ( .A(n8844), .B(n8919), .S(n10233), .Z(n8846) );
  NAND2_X1 U10343 ( .A1(n8921), .A2(n8875), .ZN(n8845) );
  OAI211_X1 U10344 ( .C1(n8924), .C2(n8878), .A(n8846), .B(n8845), .ZN(
        P2_U3482) );
  INV_X1 U10345 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8847) );
  MUX2_X1 U10346 ( .A(n8847), .B(n8925), .S(n10233), .Z(n8849) );
  NAND2_X1 U10347 ( .A1(n8927), .A2(n8875), .ZN(n8848) );
  OAI211_X1 U10348 ( .C1(n8930), .C2(n8878), .A(n8849), .B(n8848), .ZN(
        P2_U3481) );
  INV_X1 U10349 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8850) );
  MUX2_X1 U10350 ( .A(n8850), .B(n8931), .S(n10233), .Z(n8852) );
  NAND2_X1 U10351 ( .A1(n8933), .A2(n8875), .ZN(n8851) );
  OAI211_X1 U10352 ( .C1(n8878), .C2(n8936), .A(n8852), .B(n8851), .ZN(
        P2_U3480) );
  MUX2_X1 U10353 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8937), .S(n10233), .Z(
        n8854) );
  OAI22_X1 U10354 ( .A1(n8939), .A2(n8878), .B1(n8938), .B2(n8864), .ZN(n8853)
         );
  OR2_X1 U10355 ( .A1(n8854), .A2(n8853), .ZN(P2_U3479) );
  INV_X1 U10356 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8855) );
  MUX2_X1 U10357 ( .A(n8855), .B(n8942), .S(n10233), .Z(n8857) );
  NAND2_X1 U10358 ( .A1(n8944), .A2(n8875), .ZN(n8856) );
  OAI211_X1 U10359 ( .C1(n8878), .C2(n8947), .A(n8857), .B(n8856), .ZN(
        P2_U3478) );
  INV_X1 U10360 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8862) );
  NOR2_X1 U10361 ( .A1(n8858), .A2(n10217), .ZN(n8861) );
  AOI21_X1 U10362 ( .B1(n8861), .B2(n8860), .A(n8859), .ZN(n8948) );
  MUX2_X1 U10363 ( .A(n8862), .B(n8948), .S(n10233), .Z(n8863) );
  OAI21_X1 U10364 ( .B1(n8952), .B2(n8864), .A(n8863), .ZN(P2_U3477) );
  MUX2_X1 U10365 ( .A(n8865), .B(n8953), .S(n10233), .Z(n8867) );
  NAND2_X1 U10366 ( .A1(n8955), .A2(n8875), .ZN(n8866) );
  OAI211_X1 U10367 ( .C1(n8958), .C2(n8878), .A(n8867), .B(n8866), .ZN(
        P2_U3476) );
  MUX2_X1 U10368 ( .A(n8960), .B(n8868), .S(n10231), .Z(n8870) );
  NAND2_X1 U10369 ( .A1(n8961), .A2(n8875), .ZN(n8869) );
  OAI211_X1 U10370 ( .C1(n8964), .C2(n8878), .A(n8870), .B(n8869), .ZN(
        P2_U3475) );
  MUX2_X1 U10371 ( .A(n8871), .B(n8965), .S(n10233), .Z(n8873) );
  NAND2_X1 U10372 ( .A1(n8967), .A2(n8875), .ZN(n8872) );
  OAI211_X1 U10373 ( .C1(n8970), .C2(n8878), .A(n8873), .B(n8872), .ZN(
        P2_U3474) );
  MUX2_X1 U10374 ( .A(n8874), .B(n8971), .S(n10233), .Z(n8877) );
  NAND2_X1 U10375 ( .A1(n8974), .A2(n8875), .ZN(n8876) );
  OAI211_X1 U10376 ( .C1(n8878), .C2(n8978), .A(n8877), .B(n8876), .ZN(
        P2_U3473) );
  OAI22_X1 U10377 ( .A1(n8880), .A2(n10217), .B1(n8879), .B2(n10215), .ZN(
        n8881) );
  OR2_X1 U10378 ( .A1(n8882), .A2(n8881), .ZN(n8979) );
  MUX2_X1 U10379 ( .A(n8979), .B(P2_REG1_REG_12__SCAN_IN), .S(n10231), .Z(
        P2_U3471) );
  NOR2_X1 U10380 ( .A1(n8883), .A2(n10223), .ZN(n8886) );
  AOI21_X1 U10381 ( .B1(n10223), .B2(P2_REG0_REG_31__SCAN_IN), .A(n8886), .ZN(
        n8884) );
  OAI21_X1 U10382 ( .B1(n8885), .B2(n8951), .A(n8884), .ZN(P2_U3458) );
  AOI21_X1 U10383 ( .B1(n10223), .B2(P2_REG0_REG_30__SCAN_IN), .A(n8886), .ZN(
        n8887) );
  OAI21_X1 U10384 ( .B1(n8888), .B2(n8951), .A(n8887), .ZN(P2_U3457) );
  INV_X1 U10385 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8890) );
  MUX2_X1 U10386 ( .A(n8890), .B(n8889), .S(n10221), .Z(n8893) );
  NAND2_X1 U10387 ( .A1(n8891), .A2(n8973), .ZN(n8892) );
  OAI211_X1 U10388 ( .C1(n8894), .C2(n8977), .A(n8893), .B(n8892), .ZN(
        P2_U3455) );
  INV_X1 U10389 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8895) );
  MUX2_X1 U10390 ( .A(n8896), .B(n8895), .S(n10223), .Z(n8899) );
  NAND2_X1 U10391 ( .A1(n8897), .A2(n8973), .ZN(n8898) );
  OAI211_X1 U10392 ( .C1(n8900), .C2(n8977), .A(n8899), .B(n8898), .ZN(
        P2_U3454) );
  INV_X1 U10393 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8902) );
  MUX2_X1 U10394 ( .A(n8902), .B(n8901), .S(n10221), .Z(n8905) );
  NAND2_X1 U10395 ( .A1(n8903), .A2(n8973), .ZN(n8904) );
  OAI211_X1 U10396 ( .C1(n8906), .C2(n8977), .A(n8905), .B(n8904), .ZN(
        P2_U3453) );
  INV_X1 U10397 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8908) );
  MUX2_X1 U10398 ( .A(n8908), .B(n8907), .S(n10221), .Z(n8911) );
  NAND2_X1 U10399 ( .A1(n8909), .A2(n8973), .ZN(n8910) );
  OAI211_X1 U10400 ( .C1(n8912), .C2(n8977), .A(n8911), .B(n8910), .ZN(
        P2_U3452) );
  INV_X1 U10401 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8914) );
  MUX2_X1 U10402 ( .A(n8914), .B(n8913), .S(n10221), .Z(n8917) );
  NAND2_X1 U10403 ( .A1(n8915), .A2(n8973), .ZN(n8916) );
  OAI211_X1 U10404 ( .C1(n8918), .C2(n8977), .A(n8917), .B(n8916), .ZN(
        P2_U3451) );
  INV_X1 U10405 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8920) );
  MUX2_X1 U10406 ( .A(n8920), .B(n8919), .S(n10221), .Z(n8923) );
  NAND2_X1 U10407 ( .A1(n8921), .A2(n8973), .ZN(n8922) );
  OAI211_X1 U10408 ( .C1(n8924), .C2(n8977), .A(n8923), .B(n8922), .ZN(
        P2_U3450) );
  INV_X1 U10409 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8926) );
  MUX2_X1 U10410 ( .A(n8926), .B(n8925), .S(n10221), .Z(n8929) );
  NAND2_X1 U10411 ( .A1(n8927), .A2(n8973), .ZN(n8928) );
  OAI211_X1 U10412 ( .C1(n8930), .C2(n8977), .A(n8929), .B(n8928), .ZN(
        P2_U3449) );
  INV_X1 U10413 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8932) );
  MUX2_X1 U10414 ( .A(n8932), .B(n8931), .S(n10221), .Z(n8935) );
  NAND2_X1 U10415 ( .A1(n8933), .A2(n8973), .ZN(n8934) );
  OAI211_X1 U10416 ( .C1(n8936), .C2(n8977), .A(n8935), .B(n8934), .ZN(
        P2_U3448) );
  MUX2_X1 U10417 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8937), .S(n10221), .Z(
        n8941) );
  OAI22_X1 U10418 ( .A1(n8939), .A2(n8977), .B1(n8938), .B2(n8951), .ZN(n8940)
         );
  OR2_X1 U10419 ( .A1(n8941), .A2(n8940), .ZN(P2_U3447) );
  INV_X1 U10420 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8943) );
  MUX2_X1 U10421 ( .A(n8943), .B(n8942), .S(n10221), .Z(n8946) );
  NAND2_X1 U10422 ( .A1(n8944), .A2(n8973), .ZN(n8945) );
  OAI211_X1 U10423 ( .C1(n8947), .C2(n8977), .A(n8946), .B(n8945), .ZN(
        P2_U3446) );
  INV_X1 U10424 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8949) );
  MUX2_X1 U10425 ( .A(n8949), .B(n8948), .S(n10221), .Z(n8950) );
  OAI21_X1 U10426 ( .B1(n8952), .B2(n8951), .A(n8950), .ZN(P2_U3444) );
  INV_X1 U10427 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8954) );
  MUX2_X1 U10428 ( .A(n8954), .B(n8953), .S(n10221), .Z(n8957) );
  NAND2_X1 U10429 ( .A1(n8955), .A2(n8973), .ZN(n8956) );
  OAI211_X1 U10430 ( .C1(n8958), .C2(n8977), .A(n8957), .B(n8956), .ZN(
        P2_U3441) );
  MUX2_X1 U10431 ( .A(n8960), .B(n8959), .S(n10223), .Z(n8963) );
  NAND2_X1 U10432 ( .A1(n8961), .A2(n8973), .ZN(n8962) );
  OAI211_X1 U10433 ( .C1(n8964), .C2(n8977), .A(n8963), .B(n8962), .ZN(
        P2_U3438) );
  INV_X1 U10434 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8966) );
  MUX2_X1 U10435 ( .A(n8966), .B(n8965), .S(n10221), .Z(n8969) );
  NAND2_X1 U10436 ( .A1(n8967), .A2(n8973), .ZN(n8968) );
  OAI211_X1 U10437 ( .C1(n8970), .C2(n8977), .A(n8969), .B(n8968), .ZN(
        P2_U3435) );
  INV_X1 U10438 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8972) );
  MUX2_X1 U10439 ( .A(n8972), .B(n8971), .S(n10221), .Z(n8976) );
  NAND2_X1 U10440 ( .A1(n8974), .A2(n8973), .ZN(n8975) );
  OAI211_X1 U10441 ( .C1(n8978), .C2(n8977), .A(n8976), .B(n8975), .ZN(
        P2_U3432) );
  MUX2_X1 U10442 ( .A(n8979), .B(P2_REG0_REG_12__SCAN_IN), .S(n10223), .Z(
        P2_U3426) );
  INV_X1 U10443 ( .A(n8980), .ZN(n9904) );
  NOR4_X1 U10444 ( .A1(n8982), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n8981), .ZN(n8983) );
  AOI21_X1 U10445 ( .B1(n8984), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8983), .ZN(
        n8985) );
  OAI21_X1 U10446 ( .B1(n9904), .B2(n8986), .A(n8985), .ZN(P2_U3264) );
  INV_X1 U10447 ( .A(n8987), .ZN(n8988) );
  AOI22_X1 U10448 ( .A1(n9362), .A2(n9103), .B1(n9101), .B2(n9363), .ZN(n9587)
         );
  AOI22_X1 U10449 ( .A1(n9595), .A2(n9105), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n8993) );
  OAI21_X1 U10450 ( .B1(n9587), .B2(n9914), .A(n8993), .ZN(n8994) );
  AOI21_X1 U10451 ( .B1(n9849), .B2(n9924), .A(n8994), .ZN(n8995) );
  NAND2_X1 U10452 ( .A1(n8996), .A2(n8997), .ZN(n8998) );
  XOR2_X1 U10453 ( .A(n8999), .B(n8998), .Z(n9005) );
  OAI22_X1 U10454 ( .A1(n9001), .A2(n9091), .B1(n9000), .B2(n9089), .ZN(n9946)
         );
  AOI22_X1 U10455 ( .A1(n9117), .A2(n9946), .B1(P1_REG3_REG_14__SCAN_IN), .B2(
        P1_U3086), .ZN(n9002) );
  OAI21_X1 U10456 ( .B1(n9948), .B2(n9926), .A(n9002), .ZN(n9003) );
  AOI21_X1 U10457 ( .B1(n9951), .B2(n9924), .A(n9003), .ZN(n9004) );
  OAI21_X1 U10458 ( .B1(n9005), .B2(n9919), .A(n9004), .ZN(P1_U3215) );
  AOI21_X1 U10459 ( .B1(n9007), .B2(n9006), .A(n9061), .ZN(n9013) );
  AND2_X1 U10460 ( .A1(n9367), .A2(n9101), .ZN(n9008) );
  AOI21_X1 U10461 ( .B1(n9365), .B2(n9103), .A(n9008), .ZN(n9788) );
  INV_X1 U10462 ( .A(n9009), .ZN(n9652) );
  AOI22_X1 U10463 ( .A1(n9652), .A2(n9105), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n9010) );
  OAI21_X1 U10464 ( .B1(n9788), .B2(n9914), .A(n9010), .ZN(n9011) );
  AOI21_X1 U10465 ( .B1(n9862), .B2(n9924), .A(n9011), .ZN(n9012) );
  OAI21_X1 U10466 ( .B1(n9013), .B2(n9919), .A(n9012), .ZN(P1_U3216) );
  OAI21_X1 U10467 ( .B1(n9015), .B2(n4523), .A(n9014), .ZN(n9016) );
  NAND2_X1 U10468 ( .A1(n9016), .A2(n9097), .ZN(n9021) );
  AND2_X1 U10469 ( .A1(n9370), .A2(n9101), .ZN(n9017) );
  AOI21_X1 U10470 ( .B1(n9024), .B2(n9103), .A(n9017), .ZN(n9710) );
  OAI22_X1 U10471 ( .A1(n9710), .A2(n9914), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9018), .ZN(n9019) );
  AOI21_X1 U10472 ( .B1(n9713), .B2(n9105), .A(n9019), .ZN(n9020) );
  OAI211_X1 U10473 ( .C1(n9879), .C2(n9070), .A(n9021), .B(n9020), .ZN(
        P1_U3219) );
  XNOR2_X1 U10474 ( .A(n9023), .B(n9022), .ZN(n9029) );
  AOI22_X1 U10475 ( .A1(n9367), .A2(n9103), .B1(n9101), .B2(n9024), .ZN(n9678)
         );
  OAI22_X1 U10476 ( .A1(n9678), .A2(n9914), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9025), .ZN(n9026) );
  AOI21_X1 U10477 ( .B1(n9684), .B2(n9105), .A(n9026), .ZN(n9028) );
  NAND2_X1 U10478 ( .A1(n9683), .A2(n9924), .ZN(n9027) );
  OAI211_X1 U10479 ( .C1(n9029), .C2(n9919), .A(n9028), .B(n9027), .ZN(
        P1_U3223) );
  OAI21_X1 U10480 ( .B1(n9031), .B2(n9030), .A(n9100), .ZN(n9035) );
  AOI22_X1 U10481 ( .A1(n9363), .A2(n9103), .B1(n9101), .B2(n9365), .ZN(n9617)
         );
  NAND2_X1 U10482 ( .A1(n9857), .A2(n9924), .ZN(n9033) );
  AOI22_X1 U10483 ( .A1(n9625), .A2(n9105), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n9032) );
  OAI211_X1 U10484 ( .C1(n9617), .C2(n9914), .A(n9033), .B(n9032), .ZN(n9034)
         );
  AOI21_X1 U10485 ( .B1(n9035), .B2(n9097), .A(n9034), .ZN(n9036) );
  INV_X1 U10486 ( .A(n9036), .ZN(P1_U3225) );
  NAND2_X1 U10487 ( .A1(n4599), .A2(n9040), .ZN(n9039) );
  AOI22_X1 U10488 ( .A1(n4643), .A2(n9040), .B1(n9038), .B2(n9039), .ZN(n9047)
         );
  AOI22_X1 U10489 ( .A1(n9117), .A2(n9041), .B1(P1_REG3_REG_16__SCAN_IN), .B2(
        P1_U3086), .ZN(n9042) );
  OAI21_X1 U10490 ( .B1(n9043), .B2(n9926), .A(n9042), .ZN(n9044) );
  AOI21_X1 U10491 ( .B1(n9045), .B2(n9924), .A(n9044), .ZN(n9046) );
  OAI21_X1 U10492 ( .B1(n9047), .B2(n9919), .A(n9046), .ZN(P1_U3226) );
  OAI21_X1 U10493 ( .B1(n9050), .B2(n9049), .A(n9048), .ZN(n9051) );
  NAND2_X1 U10494 ( .A1(n9051), .A2(n9097), .ZN(n9057) );
  NAND2_X1 U10495 ( .A1(n9370), .A2(n9103), .ZN(n9053) );
  NAND2_X1 U10496 ( .A1(n9372), .A2(n9101), .ZN(n9052) );
  NAND2_X1 U10497 ( .A1(n9053), .A2(n9052), .ZN(n9750) );
  NOR2_X1 U10498 ( .A1(n9926), .A2(n9741), .ZN(n9054) );
  AOI211_X1 U10499 ( .C1(n9117), .C2(n9750), .A(n9055), .B(n9054), .ZN(n9056)
         );
  OAI211_X1 U10500 ( .C1(n9887), .C2(n9070), .A(n9057), .B(n9056), .ZN(
        P1_U3228) );
  INV_X1 U10501 ( .A(n9058), .ZN(n9063) );
  NOR3_X1 U10502 ( .A1(n9061), .A2(n9060), .A3(n9059), .ZN(n9062) );
  OAI21_X1 U10503 ( .B1(n9063), .B2(n9062), .A(n9097), .ZN(n9069) );
  OAI22_X1 U10504 ( .A1(n9064), .A2(n9091), .B1(n9082), .B2(n9089), .ZN(n9634)
         );
  INV_X1 U10505 ( .A(n9640), .ZN(n9066) );
  OAI22_X1 U10506 ( .A1(n9066), .A2(n9926), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9065), .ZN(n9067) );
  AOI21_X1 U10507 ( .B1(n9634), .B2(n9117), .A(n9067), .ZN(n9068) );
  OAI211_X1 U10508 ( .C1(n6604), .C2(n9070), .A(n9069), .B(n9068), .ZN(
        P1_U3229) );
  XNOR2_X1 U10509 ( .A(n9072), .B(n9071), .ZN(n9073) );
  XNOR2_X1 U10510 ( .A(n9074), .B(n9073), .ZN(n9078) );
  OAI22_X1 U10511 ( .A1(n9196), .A2(n9091), .B1(n9092), .B2(n9089), .ZN(n9693)
         );
  AOI22_X1 U10512 ( .A1(n9693), .A2(n9117), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n9075) );
  OAI21_X1 U10513 ( .B1(n9700), .B2(n9926), .A(n9075), .ZN(n9076) );
  AOI21_X1 U10514 ( .B1(n9698), .B2(n9924), .A(n9076), .ZN(n9077) );
  OAI21_X1 U10515 ( .B1(n9078), .B2(n9919), .A(n9077), .ZN(P1_U3233) );
  NAND2_X1 U10516 ( .A1(n4565), .A2(n9079), .ZN(n9081) );
  XNOR2_X1 U10517 ( .A(n9081), .B(n9080), .ZN(n9086) );
  OAI22_X1 U10518 ( .A1(n9082), .A2(n9091), .B1(n9196), .B2(n9089), .ZN(n9664)
         );
  AOI22_X1 U10519 ( .A1(n9664), .A2(n9117), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n9083) );
  OAI21_X1 U10520 ( .B1(n9671), .B2(n9926), .A(n9083), .ZN(n9084) );
  AOI21_X1 U10521 ( .B1(n9669), .B2(n9924), .A(n9084), .ZN(n9085) );
  OAI21_X1 U10522 ( .B1(n9086), .B2(n9919), .A(n9085), .ZN(P1_U3235) );
  AOI21_X1 U10523 ( .B1(n4576), .B2(n4633), .A(n9087), .ZN(n9088) );
  AOI21_X1 U10524 ( .B1(n4523), .B2(n4588), .A(n9088), .ZN(n9096) );
  OAI22_X1 U10525 ( .A1(n9092), .A2(n9091), .B1(n9090), .B2(n9089), .ZN(n9724)
         );
  AOI22_X1 U10526 ( .A1(n9724), .A2(n9117), .B1(P1_REG3_REG_18__SCAN_IN), .B2(
        P1_U3086), .ZN(n9093) );
  OAI21_X1 U10527 ( .B1(n9729), .B2(n9926), .A(n9093), .ZN(n9094) );
  AOI21_X1 U10528 ( .B1(n9816), .B2(n9924), .A(n9094), .ZN(n9095) );
  OAI21_X1 U10529 ( .B1(n9096), .B2(n9919), .A(n9095), .ZN(P1_U3238) );
  NAND2_X1 U10530 ( .A1(n8989), .A2(n9097), .ZN(n9111) );
  AOI21_X1 U10531 ( .B1(n9100), .B2(n9099), .A(n9098), .ZN(n9110) );
  AND2_X1 U10532 ( .A1(n9364), .A2(n9101), .ZN(n9102) );
  AOI21_X1 U10533 ( .B1(n9104), .B2(n9103), .A(n9102), .ZN(n9601) );
  INV_X1 U10534 ( .A(n9610), .ZN(n9106) );
  AOI22_X1 U10535 ( .A1(n9106), .A2(n9105), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n9107) );
  OAI21_X1 U10536 ( .B1(n9601), .B2(n9914), .A(n9107), .ZN(n9108) );
  AOI21_X1 U10537 ( .B1(n9853), .B2(n9924), .A(n9108), .ZN(n9109) );
  OAI21_X1 U10538 ( .B1(n9111), .B2(n9110), .A(n9109), .ZN(P1_U3240) );
  NAND2_X1 U10539 ( .A1(n9113), .A2(n9112), .ZN(n9114) );
  XOR2_X1 U10540 ( .A(n9115), .B(n9114), .Z(n9123) );
  AOI22_X1 U10541 ( .A1(n9117), .A2(n9116), .B1(P1_REG3_REG_15__SCAN_IN), .B2(
        P1_U3086), .ZN(n9118) );
  OAI21_X1 U10542 ( .B1(n9119), .B2(n9926), .A(n9118), .ZN(n9120) );
  AOI21_X1 U10543 ( .B1(n9121), .B2(n9924), .A(n9120), .ZN(n9122) );
  OAI21_X1 U10544 ( .B1(n9123), .B2(n9919), .A(n9122), .ZN(P1_U3241) );
  AND2_X1 U10545 ( .A1(n9583), .A2(n9207), .ZN(n9275) );
  NAND2_X1 U10546 ( .A1(n9632), .A2(n9222), .ZN(n9201) );
  INV_X1 U10547 ( .A(n9184), .ZN(n9332) );
  NOR2_X1 U10548 ( .A1(n9124), .A2(n9332), .ZN(n9186) );
  AND3_X1 U10549 ( .A1(n9128), .A2(n9347), .A3(n9127), .ZN(n9130) );
  NAND3_X1 U10550 ( .A1(n9131), .A2(n9130), .A3(n9129), .ZN(n9144) );
  OAI21_X1 U10551 ( .B1(n9140), .B2(n9382), .A(n10067), .ZN(n9138) );
  NAND2_X1 U10552 ( .A1(n9383), .A2(n9347), .ZN(n9134) );
  OAI21_X1 U10553 ( .B1(n9134), .B2(n9132), .A(n9139), .ZN(n9137) );
  NAND2_X1 U10554 ( .A1(n9382), .A2(n9347), .ZN(n9133) );
  OAI21_X1 U10555 ( .B1(n9134), .B2(n10067), .A(n9133), .ZN(n9136) );
  AOI22_X1 U10556 ( .A1(n9138), .A2(n9137), .B1(n9136), .B2(n9135), .ZN(n9143)
         );
  OAI22_X1 U10557 ( .A1(n9140), .A2(n9139), .B1(n9347), .B2(n9382), .ZN(n9141)
         );
  NAND2_X1 U10558 ( .A1(n9141), .A2(n10072), .ZN(n9142) );
  NAND2_X1 U10559 ( .A1(n9148), .A2(n9147), .ZN(n9149) );
  MUX2_X1 U10560 ( .A(n9150), .B(n9149), .S(n9222), .Z(n9155) );
  MUX2_X1 U10561 ( .A(n9152), .B(n9151), .S(n9222), .Z(n9153) );
  INV_X1 U10562 ( .A(n9153), .ZN(n9154) );
  AOI21_X1 U10563 ( .B1(n9160), .B2(n9162), .A(n9157), .ZN(n9158) );
  NAND2_X1 U10564 ( .A1(n9165), .A2(n9163), .ZN(n9308) );
  NOR2_X1 U10565 ( .A1(n9158), .A2(n9308), .ZN(n9159) );
  NAND2_X1 U10566 ( .A1(n9167), .A2(n9164), .ZN(n9311) );
  OAI21_X1 U10567 ( .B1(n9159), .B2(n9311), .A(n9312), .ZN(n9170) );
  NAND3_X1 U10568 ( .A1(n9166), .A2(n9312), .A3(n9165), .ZN(n9168) );
  NAND2_X1 U10569 ( .A1(n9168), .A2(n9167), .ZN(n9169) );
  AOI211_X1 U10570 ( .C1(n9176), .C2(n9175), .A(n9172), .B(n9171), .ZN(n9174)
         );
  INV_X1 U10571 ( .A(n9175), .ZN(n9315) );
  NAND2_X1 U10572 ( .A1(n9178), .A2(n9177), .ZN(n9318) );
  INV_X1 U10573 ( .A(n9181), .ZN(n9322) );
  NAND2_X1 U10574 ( .A1(n9194), .A2(n9183), .ZN(n9324) );
  OAI211_X1 U10575 ( .C1(n9193), .C2(n9324), .A(n9184), .B(n9192), .ZN(n9185)
         );
  MUX2_X1 U10576 ( .A(n9186), .B(n9185), .S(n9222), .Z(n9190) );
  NOR2_X1 U10577 ( .A1(n9698), .A2(n9187), .ZN(n9198) );
  OAI21_X1 U10578 ( .B1(n9198), .B2(n9327), .A(n9222), .ZN(n9189) );
  NAND2_X1 U10579 ( .A1(n9199), .A2(n9188), .ZN(n9267) );
  AOI22_X1 U10580 ( .A1(n9190), .A2(n9189), .B1(n9222), .B2(n9267), .ZN(n9197)
         );
  NAND2_X1 U10581 ( .A1(n9192), .A2(n9191), .ZN(n9295) );
  NOR2_X1 U10582 ( .A1(n9193), .A2(n9295), .ZN(n9195) );
  INV_X1 U10583 ( .A(n9194), .ZN(n9328) );
  NOR2_X1 U10584 ( .A1(n9683), .A2(n9196), .ZN(n9271) );
  NOR2_X1 U10585 ( .A1(n9271), .A2(n9198), .ZN(n9260) );
  NAND2_X1 U10586 ( .A1(n9203), .A2(n9200), .ZN(n9261) );
  AND2_X1 U10587 ( .A1(n9632), .A2(n9202), .ZN(n9268) );
  INV_X1 U10588 ( .A(n9203), .ZN(n9204) );
  NOR3_X1 U10589 ( .A1(n9268), .A2(n9204), .A3(n9222), .ZN(n9205) );
  MUX2_X1 U10590 ( .A(n9269), .B(n9262), .S(n9222), .Z(n9208) );
  OR2_X1 U10591 ( .A1(n9853), .A2(n9210), .ZN(n9258) );
  INV_X1 U10592 ( .A(n9258), .ZN(n9212) );
  OAI211_X1 U10593 ( .C1(n9212), .C2(n9211), .A(n9347), .B(n9583), .ZN(n9214)
         );
  NAND2_X1 U10594 ( .A1(n9216), .A2(n9215), .ZN(n9281) );
  OAI21_X1 U10595 ( .B1(n9281), .B2(n9259), .A(n9282), .ZN(n9217) );
  AOI22_X1 U10596 ( .A1(n9218), .A2(n9282), .B1(n9347), .B2(n9217), .ZN(n9220)
         );
  MUX2_X1 U10597 ( .A(n9283), .B(n9257), .S(n9222), .Z(n9219) );
  INV_X1 U10598 ( .A(n9223), .ZN(n9221) );
  NAND2_X1 U10599 ( .A1(n9545), .A2(n9360), .ZN(n9227) );
  NAND2_X1 U10600 ( .A1(n9360), .A2(n9286), .ZN(n9287) );
  NAND3_X1 U10601 ( .A1(n9224), .A2(n9355), .A3(n9287), .ZN(n9226) );
  NAND2_X1 U10602 ( .A1(n9545), .A2(n9225), .ZN(n9348) );
  OAI211_X1 U10603 ( .C1(n9228), .C2(n9227), .A(n9226), .B(n9348), .ZN(n9346)
         );
  OAI21_X1 U10604 ( .B1(n9346), .B2(n5284), .A(n9347), .ZN(n9293) );
  INV_X1 U10605 ( .A(n9355), .ZN(n9256) );
  XOR2_X1 U10606 ( .A(n9360), .B(n9554), .Z(n9255) );
  INV_X1 U10607 ( .A(n9620), .ZN(n9615) );
  INV_X1 U10608 ( .A(n9631), .ZN(n9249) );
  NOR4_X1 U10609 ( .A1(n10014), .A2(n10001), .A3(n9229), .A4(n5964), .ZN(n9231) );
  INV_X1 U10610 ( .A(n9982), .ZN(n9973) );
  NAND3_X1 U10611 ( .A1(n9231), .A2(n9973), .A3(n9230), .ZN(n9234) );
  NOR3_X1 U10612 ( .A1(n9234), .A2(n9233), .A3(n9232), .ZN(n9235) );
  NAND4_X1 U10613 ( .A1(n9238), .A2(n9237), .A3(n9236), .A4(n9235), .ZN(n9239)
         );
  NOR4_X1 U10614 ( .A1(n9242), .A2(n9241), .A3(n9240), .A4(n9239), .ZN(n9243)
         );
  NAND4_X1 U10615 ( .A1(n9245), .A2(n9942), .A3(n9244), .A4(n9243), .ZN(n9246)
         );
  NOR4_X1 U10616 ( .A1(n9717), .A2(n9324), .A3(n9295), .A4(n9246), .ZN(n9247)
         );
  NAND4_X1 U10617 ( .A1(n9662), .A2(n9247), .A3(n9691), .A4(n9680), .ZN(n9248)
         );
  NOR4_X1 U10618 ( .A1(n9615), .A2(n9250), .A3(n9249), .A4(n9248), .ZN(n9251)
         );
  NAND4_X1 U10619 ( .A1(n9572), .A2(n9252), .A3(n9251), .A4(n9604), .ZN(n9253)
         );
  INV_X1 U10620 ( .A(n9348), .ZN(n9339) );
  NAND2_X1 U10621 ( .A1(n9259), .A2(n9258), .ZN(n9278) );
  INV_X1 U10622 ( .A(n9260), .ZN(n9266) );
  NAND3_X1 U10623 ( .A1(n9269), .A2(n9632), .A3(n9261), .ZN(n9263) );
  AND2_X1 U10624 ( .A1(n9263), .A2(n9262), .ZN(n9265) );
  NAND2_X1 U10625 ( .A1(n9265), .A2(n9264), .ZN(n9274) );
  NOR3_X1 U10626 ( .A1(n9278), .A2(n9266), .A3(n9274), .ZN(n9284) );
  INV_X1 U10627 ( .A(n9267), .ZN(n9270) );
  OAI211_X1 U10628 ( .C1(n9271), .C2(n9270), .A(n9269), .B(n9268), .ZN(n9272)
         );
  INV_X1 U10629 ( .A(n9272), .ZN(n9273) );
  NOR2_X1 U10630 ( .A1(n9274), .A2(n9273), .ZN(n9277) );
  INV_X1 U10631 ( .A(n9275), .ZN(n9276) );
  NOR2_X1 U10632 ( .A1(n9277), .A2(n9276), .ZN(n9279) );
  NOR2_X1 U10633 ( .A1(n9279), .A2(n9278), .ZN(n9280) );
  OR2_X1 U10634 ( .A1(n9281), .A2(n9280), .ZN(n9333) );
  OAI211_X1 U10635 ( .C1(n9284), .C2(n9333), .A(n9283), .B(n9282), .ZN(n9335)
         );
  NOR2_X1 U10636 ( .A1(n9333), .A2(n9692), .ZN(n9285) );
  OAI22_X1 U10637 ( .A1(n8161), .A2(n9286), .B1(n9335), .B2(n9285), .ZN(n9288)
         );
  OAI22_X1 U10638 ( .A1(n9338), .A2(n9288), .B1(n9554), .B2(n9287), .ZN(n9290)
         );
  NOR2_X1 U10639 ( .A1(n5284), .A2(n9294), .ZN(n9342) );
  INV_X1 U10640 ( .A(n5962), .ZN(n9344) );
  INV_X1 U10641 ( .A(n9295), .ZN(n9330) );
  AND4_X1 U10642 ( .A1(n9299), .A2(n9298), .A3(n9297), .A4(n5964), .ZN(n9303)
         );
  AND4_X1 U10643 ( .A1(n9303), .A2(n9302), .A3(n9301), .A4(n9300), .ZN(n9306)
         );
  OAI211_X1 U10644 ( .C1(n9307), .C2(n9306), .A(n9305), .B(n9304), .ZN(n9310)
         );
  INV_X1 U10645 ( .A(n9308), .ZN(n9309) );
  NAND2_X1 U10646 ( .A1(n9310), .A2(n9309), .ZN(n9314) );
  INV_X1 U10647 ( .A(n9311), .ZN(n9313) );
  AOI21_X1 U10648 ( .B1(n9314), .B2(n9313), .A(n5008), .ZN(n9317) );
  AOI21_X1 U10649 ( .B1(n9317), .B2(n9316), .A(n9315), .ZN(n9320) );
  AOI21_X1 U10650 ( .B1(n9320), .B2(n9319), .A(n9318), .ZN(n9323) );
  NOR3_X1 U10651 ( .A1(n9323), .A2(n9322), .A3(n9321), .ZN(n9326) );
  INV_X1 U10652 ( .A(n9324), .ZN(n9325) );
  OAI21_X1 U10653 ( .B1(n4831), .B2(n9326), .A(n9325), .ZN(n9329) );
  AOI211_X1 U10654 ( .C1(n9330), .C2(n9329), .A(n9328), .B(n9327), .ZN(n9331)
         );
  NOR3_X1 U10655 ( .A1(n9333), .A2(n9332), .A3(n9331), .ZN(n9334) );
  NOR2_X1 U10656 ( .A1(n9335), .A2(n9334), .ZN(n9337) );
  OAI22_X1 U10657 ( .A1(n9338), .A2(n9337), .B1(n9336), .B2(n9554), .ZN(n9340)
         );
  OAI21_X1 U10658 ( .B1(n9340), .B2(n9339), .A(n9355), .ZN(n9341) );
  MUX2_X1 U10659 ( .A(n9342), .B(n9344), .S(n9341), .Z(n9343) );
  NAND3_X1 U10660 ( .A1(n9936), .A2(n9344), .A3(n9402), .ZN(n9345) );
  OAI211_X1 U10661 ( .C1(n9351), .C2(n9358), .A(n9345), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9357) );
  OAI21_X1 U10662 ( .B1(n9348), .B2(n9347), .A(n9346), .ZN(n9354) );
  NOR4_X1 U10663 ( .A1(n9352), .A2(n9351), .A3(n9350), .A4(n9349), .ZN(n9353)
         );
  OAI211_X1 U10664 ( .C1(n9355), .C2(n5284), .A(n9354), .B(n9353), .ZN(n9356)
         );
  OAI211_X1 U10665 ( .C1(n9359), .C2(n9358), .A(n9357), .B(n9356), .ZN(
        P1_U3242) );
  MUX2_X1 U10666 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9360), .S(n9385), .Z(
        P1_U3584) );
  MUX2_X1 U10667 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9361), .S(n9385), .Z(
        P1_U3583) );
  MUX2_X1 U10668 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9362), .S(n9385), .Z(
        P1_U3582) );
  MUX2_X1 U10669 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9363), .S(n9385), .Z(
        P1_U3580) );
  MUX2_X1 U10670 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9364), .S(n9385), .Z(
        P1_U3579) );
  MUX2_X1 U10671 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9365), .S(n9385), .Z(
        P1_U3578) );
  MUX2_X1 U10672 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9366), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10673 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9367), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10674 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9368), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10675 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9369), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10676 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9370), .S(n9385), .Z(
        P1_U3572) );
  MUX2_X1 U10677 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9371), .S(n9385), .Z(
        P1_U3571) );
  MUX2_X1 U10678 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9372), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10679 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9373), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10680 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9374), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10681 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9375), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10682 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9376), .S(n9385), .Z(
        P1_U3566) );
  MUX2_X1 U10683 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9377), .S(n9385), .Z(
        P1_U3565) );
  MUX2_X1 U10684 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9378), .S(n9385), .Z(
        P1_U3564) );
  MUX2_X1 U10685 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9379), .S(n9385), .Z(
        P1_U3563) );
  MUX2_X1 U10686 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9380), .S(n9385), .Z(
        P1_U3562) );
  MUX2_X1 U10687 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9381), .S(n9385), .Z(
        P1_U3561) );
  MUX2_X1 U10688 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9382), .S(n9385), .Z(
        P1_U3560) );
  MUX2_X1 U10689 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9383), .S(n9385), .Z(
        P1_U3559) );
  MUX2_X1 U10690 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9384), .S(n9385), .Z(
        P1_U3557) );
  MUX2_X1 U10691 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n9386), .S(n9385), .Z(
        P1_U3554) );
  OAI211_X1 U10692 ( .C1(n9389), .C2(n9388), .A(n9531), .B(n9387), .ZN(n9396)
         );
  OAI211_X1 U10693 ( .C1(n9391), .C2(n9401), .A(n9507), .B(n9390), .ZN(n9395)
         );
  AOI22_X1 U10694 ( .A1(n9936), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9394) );
  NAND2_X1 U10695 ( .A1(n9530), .A2(n9392), .ZN(n9393) );
  NAND4_X1 U10696 ( .A1(n9396), .A2(n9395), .A3(n9394), .A4(n9393), .ZN(
        P1_U3244) );
  NAND3_X1 U10697 ( .A1(n9398), .A2(n9397), .A3(n4519), .ZN(n9404) );
  NOR2_X1 U10698 ( .A1(n4519), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9400) );
  NOR2_X1 U10699 ( .A1(n9400), .A2(n9399), .ZN(n9931) );
  NOR2_X1 U10700 ( .A1(n9931), .A2(n10534), .ZN(n9928) );
  AOI21_X1 U10701 ( .B1(n9402), .B2(n9401), .A(n9928), .ZN(n9403) );
  NAND3_X1 U10702 ( .A1(n9404), .A2(P1_U3973), .A3(n9403), .ZN(n9445) );
  NOR2_X1 U10703 ( .A1(n9405), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9406) );
  AOI21_X1 U10704 ( .B1(n9936), .B2(P1_ADDR_REG_2__SCAN_IN), .A(n9406), .ZN(
        n9407) );
  OAI21_X1 U10705 ( .B1(n9503), .B2(n9408), .A(n9407), .ZN(n9409) );
  INV_X1 U10706 ( .A(n9409), .ZN(n9417) );
  OAI211_X1 U10707 ( .C1(n9411), .C2(n9410), .A(n9531), .B(n9423), .ZN(n9416)
         );
  OAI211_X1 U10708 ( .C1(n9414), .C2(n9413), .A(n9507), .B(n9412), .ZN(n9415)
         );
  NAND4_X1 U10709 ( .A1(n9445), .A2(n9417), .A3(n9416), .A4(n9415), .ZN(
        P1_U3245) );
  OAI211_X1 U10710 ( .C1(n9420), .C2(n9419), .A(n9507), .B(n9418), .ZN(n9430)
         );
  MUX2_X1 U10711 ( .A(n6797), .B(P1_REG1_REG_3__SCAN_IN), .S(n9426), .Z(n9421)
         );
  NAND3_X1 U10712 ( .A1(n9423), .A2(n9422), .A3(n9421), .ZN(n9424) );
  NAND3_X1 U10713 ( .A1(n9531), .A2(n9440), .A3(n9424), .ZN(n9429) );
  AND2_X1 U10714 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9425) );
  AOI21_X1 U10715 ( .B1(n9936), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n9425), .ZN(
        n9428) );
  NAND2_X1 U10716 ( .A1(n9530), .A2(n9426), .ZN(n9427) );
  NAND4_X1 U10717 ( .A1(n9430), .A2(n9429), .A3(n9428), .A4(n9427), .ZN(
        P1_U3246) );
  AOI21_X1 U10718 ( .B1(n9936), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n9431), .ZN(
        n9432) );
  OAI21_X1 U10719 ( .B1(n9503), .B2(n9437), .A(n9432), .ZN(n9433) );
  INV_X1 U10720 ( .A(n9433), .ZN(n9444) );
  OAI211_X1 U10721 ( .C1(n9436), .C2(n9435), .A(n9507), .B(n9434), .ZN(n9443)
         );
  MUX2_X1 U10722 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6800), .S(n9437), .Z(n9438)
         );
  NAND3_X1 U10723 ( .A1(n9440), .A2(n9439), .A3(n9438), .ZN(n9441) );
  NAND3_X1 U10724 ( .A1(n9531), .A2(n9457), .A3(n9441), .ZN(n9442) );
  NAND4_X1 U10725 ( .A1(n9445), .A2(n9444), .A3(n9443), .A4(n9442), .ZN(
        P1_U3247) );
  NOR2_X1 U10726 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9446), .ZN(n9449) );
  NOR2_X1 U10727 ( .A1(n9503), .A2(n9447), .ZN(n9448) );
  AOI211_X1 U10728 ( .C1(n9936), .C2(P1_ADDR_REG_5__SCAN_IN), .A(n9449), .B(
        n9448), .ZN(n9461) );
  OAI211_X1 U10729 ( .C1(n9452), .C2(n9451), .A(n9507), .B(n9450), .ZN(n9460)
         );
  INV_X1 U10730 ( .A(n9453), .ZN(n9456) );
  MUX2_X1 U10731 ( .A(n6803), .B(P1_REG1_REG_5__SCAN_IN), .S(n9454), .Z(n9455)
         );
  NAND3_X1 U10732 ( .A1(n9457), .A2(n9456), .A3(n9455), .ZN(n9458) );
  NAND3_X1 U10733 ( .A1(n9531), .A2(n9471), .A3(n9458), .ZN(n9459) );
  NAND3_X1 U10734 ( .A1(n9461), .A2(n9460), .A3(n9459), .ZN(P1_U3248) );
  AND2_X1 U10735 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9464) );
  NOR2_X1 U10736 ( .A1(n9503), .A2(n9462), .ZN(n9463) );
  AOI211_X1 U10737 ( .C1(n9936), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n9464), .B(
        n9463), .ZN(n9476) );
  OAI211_X1 U10738 ( .C1(n9467), .C2(n9466), .A(n9507), .B(n9465), .ZN(n9475)
         );
  INV_X1 U10739 ( .A(n9468), .ZN(n9473) );
  NAND3_X1 U10740 ( .A1(n9471), .A2(n9470), .A3(n9469), .ZN(n9472) );
  NAND3_X1 U10741 ( .A1(n9531), .A2(n9473), .A3(n9472), .ZN(n9474) );
  NAND3_X1 U10742 ( .A1(n9476), .A2(n9475), .A3(n9474), .ZN(P1_U3249) );
  NOR2_X1 U10743 ( .A1(n9503), .A2(n9477), .ZN(n9478) );
  AOI211_X1 U10744 ( .C1(n9936), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n9479), .B(
        n9478), .ZN(n9489) );
  OAI211_X1 U10745 ( .C1(n9482), .C2(n9481), .A(n9531), .B(n9480), .ZN(n9488)
         );
  AOI211_X1 U10746 ( .C1(n9485), .C2(n9484), .A(n9483), .B(n9534), .ZN(n9486)
         );
  INV_X1 U10747 ( .A(n9486), .ZN(n9487) );
  NAND3_X1 U10748 ( .A1(n9489), .A2(n9488), .A3(n9487), .ZN(P1_U3254) );
  AOI211_X1 U10749 ( .C1(n9492), .C2(n9491), .A(n9490), .B(n9534), .ZN(n9493)
         );
  INV_X1 U10750 ( .A(n9493), .ZN(n9502) );
  INV_X1 U10751 ( .A(n9494), .ZN(n9495) );
  AOI21_X1 U10752 ( .B1(n9936), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n9495), .ZN(
        n9501) );
  NAND2_X1 U10753 ( .A1(n9530), .A2(n9496), .ZN(n9500) );
  OAI211_X1 U10754 ( .C1(n9498), .C2(n9497), .A(n9531), .B(n9510), .ZN(n9499)
         );
  NAND4_X1 U10755 ( .A1(n9502), .A2(n9501), .A3(n9500), .A4(n9499), .ZN(
        P1_U3256) );
  AND2_X1 U10756 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9505) );
  NOR2_X1 U10757 ( .A1(n9503), .A2(n9514), .ZN(n9504) );
  AOI211_X1 U10758 ( .C1(n9936), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n9505), .B(
        n9504), .ZN(n9519) );
  OAI211_X1 U10759 ( .C1(n9509), .C2(n9508), .A(n9507), .B(n9506), .ZN(n9518)
         );
  INV_X1 U10760 ( .A(n9510), .ZN(n9511) );
  AOI21_X1 U10761 ( .B1(n9514), .B2(P1_REG1_REG_14__SCAN_IN), .A(n9511), .ZN(
        n9512) );
  OAI211_X1 U10762 ( .C1(P1_REG1_REG_14__SCAN_IN), .C2(n9514), .A(n9513), .B(
        n9512), .ZN(n9515) );
  NAND3_X1 U10763 ( .A1(n9531), .A2(n9516), .A3(n9515), .ZN(n9517) );
  NAND3_X1 U10764 ( .A1(n9519), .A2(n9518), .A3(n9517), .ZN(P1_U3257) );
  NAND2_X1 U10765 ( .A1(n9524), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9520) );
  NAND2_X1 U10766 ( .A1(n9521), .A2(n9520), .ZN(n9523) );
  XNOR2_X1 U10767 ( .A(n9523), .B(n9522), .ZN(n9535) );
  INV_X1 U10768 ( .A(n9535), .ZN(n9529) );
  NAND2_X1 U10769 ( .A1(n9524), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9525) );
  NAND2_X1 U10770 ( .A1(n9526), .A2(n9525), .ZN(n9527) );
  XNOR2_X1 U10771 ( .A(n9527), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9532) );
  OAI22_X1 U10772 ( .A1(n9529), .A2(n9534), .B1(n9532), .B2(n9528), .ZN(n9537)
         );
  AOI21_X1 U10773 ( .B1(n9532), .B2(n9531), .A(n9530), .ZN(n9533) );
  OAI21_X1 U10774 ( .B1(n9535), .B2(n9534), .A(n9533), .ZN(n9536) );
  MUX2_X1 U10775 ( .A(n9537), .B(n9536), .S(n5285), .Z(n9538) );
  INV_X1 U10776 ( .A(n9538), .ZN(n9540) );
  NAND2_X1 U10777 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n9539) );
  OAI211_X1 U10778 ( .C1(n9541), .C2(n4987), .A(n9540), .B(n9539), .ZN(
        P1_U3262) );
  INV_X1 U10779 ( .A(n9542), .ZN(n9756) );
  NAND2_X1 U10780 ( .A1(n9734), .A2(n9756), .ZN(n9551) );
  OAI21_X1 U10781 ( .B1(n9734), .B2(n9543), .A(n9551), .ZN(n9544) );
  AOI21_X1 U10782 ( .B1(n9545), .B2(n9950), .A(n9544), .ZN(n9546) );
  OAI21_X1 U10783 ( .B1(n9547), .B2(n9746), .A(n9546), .ZN(P1_U3263) );
  INV_X1 U10784 ( .A(n9548), .ZN(n9549) );
  AOI211_X1 U10785 ( .C1(n9554), .C2(n9550), .A(n10003), .B(n9549), .ZN(n9757)
         );
  INV_X1 U10786 ( .A(n9757), .ZN(n9556) );
  OAI21_X1 U10787 ( .B1(n9734), .B2(n9552), .A(n9551), .ZN(n9553) );
  AOI21_X1 U10788 ( .B1(n9554), .B2(n9950), .A(n9553), .ZN(n9555) );
  OAI21_X1 U10789 ( .B1(n9556), .B2(n9746), .A(n9555), .ZN(P1_U3264) );
  OAI22_X1 U10790 ( .A1(n9558), .A2(n9699), .B1(n9557), .B2(n9734), .ZN(n9559)
         );
  AOI21_X1 U10791 ( .B1(n9560), .B2(n9950), .A(n9559), .ZN(n9561) );
  OAI21_X1 U10792 ( .B1(n9562), .B2(n9746), .A(n9561), .ZN(n9563) );
  AOI21_X1 U10793 ( .B1(n9564), .B2(n10006), .A(n9563), .ZN(n9565) );
  OAI21_X1 U10794 ( .B1(n9566), .B2(n10033), .A(n9565), .ZN(P1_U3356) );
  OAI21_X1 U10795 ( .B1(n9572), .B2(n9568), .A(n9567), .ZN(n9571) );
  INV_X1 U10796 ( .A(n9569), .ZN(n9570) );
  AOI21_X1 U10797 ( .B1(n9571), .B2(n9996), .A(n9570), .ZN(n9762) );
  XNOR2_X1 U10798 ( .A(n9573), .B(n9572), .ZN(n9763) );
  OAI22_X1 U10799 ( .A1(n9575), .A2(n9699), .B1(n9574), .B2(n9734), .ZN(n9576)
         );
  AOI21_X1 U10800 ( .B1(n9760), .B2(n9950), .A(n9576), .ZN(n9580) );
  AOI21_X1 U10801 ( .B1(n9760), .B2(n9593), .A(n10003), .ZN(n9578) );
  NAND2_X1 U10802 ( .A1(n9759), .A2(n10025), .ZN(n9579) );
  OAI211_X1 U10803 ( .C1(n9763), .C2(n9737), .A(n9580), .B(n9579), .ZN(n9581)
         );
  INV_X1 U10804 ( .A(n9581), .ZN(n9582) );
  OAI21_X1 U10805 ( .B1(n10033), .B2(n9762), .A(n9582), .ZN(P1_U3265) );
  NAND3_X1 U10806 ( .A1(n9584), .A2(n9583), .A3(n9591), .ZN(n9585) );
  NAND2_X1 U10807 ( .A1(n9586), .A2(n9585), .ZN(n9589) );
  INV_X1 U10808 ( .A(n9587), .ZN(n9588) );
  AOI21_X1 U10809 ( .B1(n9589), .B2(n9996), .A(n9588), .ZN(n9766) );
  OAI21_X1 U10810 ( .B1(n9592), .B2(n9591), .A(n9590), .ZN(n9764) );
  AOI21_X1 U10811 ( .B1(n9607), .B2(n9849), .A(n10003), .ZN(n9594) );
  NAND2_X1 U10812 ( .A1(n9594), .A2(n9593), .ZN(n9765) );
  AOI22_X1 U10813 ( .A1(n9595), .A2(n10019), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n10033), .ZN(n9597) );
  NAND2_X1 U10814 ( .A1(n9849), .A2(n9950), .ZN(n9596) );
  OAI211_X1 U10815 ( .C1(n9765), .C2(n9746), .A(n9597), .B(n9596), .ZN(n9598)
         );
  AOI21_X1 U10816 ( .B1(n9764), .B2(n10006), .A(n9598), .ZN(n9599) );
  OAI21_X1 U10817 ( .B1(n10033), .B2(n9766), .A(n9599), .ZN(P1_U3266) );
  XNOR2_X1 U10818 ( .A(n9600), .B(n9604), .ZN(n9603) );
  INV_X1 U10819 ( .A(n9601), .ZN(n9602) );
  AOI21_X1 U10820 ( .B1(n9603), .B2(n9996), .A(n9602), .ZN(n9772) );
  INV_X1 U10821 ( .A(n9604), .ZN(n9605) );
  XNOR2_X1 U10822 ( .A(n9606), .B(n9605), .ZN(n9770) );
  OAI211_X1 U10823 ( .C1(n9608), .C2(n9624), .A(n10073), .B(n9607), .ZN(n9771)
         );
  OAI22_X1 U10824 ( .A1(n9610), .A2(n9699), .B1(n9609), .B2(n9734), .ZN(n9611)
         );
  AOI21_X1 U10825 ( .B1(n9853), .B2(n9950), .A(n9611), .ZN(n9612) );
  OAI21_X1 U10826 ( .B1(n9771), .B2(n9746), .A(n9612), .ZN(n9613) );
  AOI21_X1 U10827 ( .B1(n9770), .B2(n10006), .A(n9613), .ZN(n9614) );
  OAI21_X1 U10828 ( .B1(n10033), .B2(n9772), .A(n9614), .ZN(P1_U3267) );
  XNOR2_X1 U10829 ( .A(n9616), .B(n9615), .ZN(n9619) );
  INV_X1 U10830 ( .A(n9617), .ZN(n9618) );
  AOI21_X1 U10831 ( .B1(n9619), .B2(n9996), .A(n9618), .ZN(n9779) );
  XNOR2_X1 U10832 ( .A(n9621), .B(n9620), .ZN(n9776) );
  NAND2_X1 U10833 ( .A1(n9857), .A2(n9638), .ZN(n9622) );
  NAND2_X1 U10834 ( .A1(n9622), .A2(n10073), .ZN(n9623) );
  OR2_X1 U10835 ( .A1(n9624), .A2(n9623), .ZN(n9777) );
  AOI22_X1 U10836 ( .A1(n9625), .A2(n10019), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n10033), .ZN(n9627) );
  NAND2_X1 U10837 ( .A1(n9857), .A2(n9950), .ZN(n9626) );
  OAI211_X1 U10838 ( .C1(n9777), .C2(n9746), .A(n9627), .B(n9626), .ZN(n9628)
         );
  AOI21_X1 U10839 ( .B1(n9776), .B2(n10006), .A(n9628), .ZN(n9629) );
  OAI21_X1 U10840 ( .B1(n9779), .B2(n10033), .A(n9629), .ZN(P1_U3268) );
  XNOR2_X1 U10841 ( .A(n9630), .B(n9631), .ZN(n9786) );
  AOI21_X1 U10842 ( .B1(n9648), .B2(n9632), .A(n9631), .ZN(n9633) );
  NOR3_X1 U10843 ( .A1(n4542), .A2(n9633), .A3(n10016), .ZN(n9635) );
  NOR2_X1 U10844 ( .A1(n9635), .A2(n9634), .ZN(n9785) );
  INV_X1 U10845 ( .A(n9785), .ZN(n9644) );
  NAND2_X1 U10846 ( .A1(n9782), .A2(n9655), .ZN(n9637) );
  AND2_X1 U10847 ( .A1(n9638), .A2(n9637), .ZN(n9783) );
  NAND2_X1 U10848 ( .A1(n9783), .A2(n9639), .ZN(n9642) );
  AOI22_X1 U10849 ( .A1(n9640), .A2(n10019), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n10033), .ZN(n9641) );
  OAI211_X1 U10850 ( .C1(n6604), .C2(n10029), .A(n9642), .B(n9641), .ZN(n9643)
         );
  AOI21_X1 U10851 ( .B1(n9644), .B2(n9734), .A(n9643), .ZN(n9645) );
  OAI21_X1 U10852 ( .B1(n9737), .B2(n9786), .A(n9645), .ZN(P1_U3269) );
  INV_X1 U10853 ( .A(n9788), .ZN(n9651) );
  OR2_X1 U10854 ( .A1(n9646), .A2(n9653), .ZN(n9647) );
  NAND2_X1 U10855 ( .A1(n9648), .A2(n9647), .ZN(n9649) );
  NAND2_X1 U10856 ( .A1(n9649), .A2(n9996), .ZN(n9790) );
  INV_X1 U10857 ( .A(n9790), .ZN(n9650) );
  AOI211_X1 U10858 ( .C1(n10019), .C2(n9652), .A(n9651), .B(n9650), .ZN(n9660)
         );
  XNOR2_X1 U10859 ( .A(n9654), .B(n9653), .ZN(n9787) );
  AOI21_X1 U10860 ( .B1(n9862), .B2(n9667), .A(n10003), .ZN(n9656) );
  NAND2_X1 U10861 ( .A1(n9656), .A2(n9655), .ZN(n9789) );
  AOI22_X1 U10862 ( .A1(n9862), .A2(n9950), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n10033), .ZN(n9657) );
  OAI21_X1 U10863 ( .B1(n9789), .B2(n9746), .A(n9657), .ZN(n9658) );
  AOI21_X1 U10864 ( .B1(n9787), .B2(n10006), .A(n9658), .ZN(n9659) );
  OAI21_X1 U10865 ( .B1(n9660), .B2(n10033), .A(n9659), .ZN(P1_U3270) );
  XOR2_X1 U10866 ( .A(n9661), .B(n9662), .Z(n9797) );
  INV_X1 U10867 ( .A(n9797), .ZN(n9676) );
  XOR2_X1 U10868 ( .A(n9663), .B(n9662), .Z(n9666) );
  INV_X1 U10869 ( .A(n9664), .ZN(n9665) );
  OAI21_X1 U10870 ( .B1(n9666), .B2(n10016), .A(n9665), .ZN(n9795) );
  NAND2_X1 U10871 ( .A1(n9795), .A2(n9734), .ZN(n9675) );
  INV_X1 U10872 ( .A(n9667), .ZN(n9668) );
  AOI211_X1 U10873 ( .C1(n9669), .C2(n4926), .A(n10003), .B(n9668), .ZN(n9796)
         );
  NOR2_X1 U10874 ( .A1(n9867), .A2(n10029), .ZN(n9673) );
  OAI22_X1 U10875 ( .A1(n9671), .A2(n9699), .B1(n9734), .B2(n9670), .ZN(n9672)
         );
  AOI211_X1 U10876 ( .C1(n9796), .C2(n10025), .A(n9673), .B(n9672), .ZN(n9674)
         );
  OAI211_X1 U10877 ( .C1(n9676), .C2(n9737), .A(n9675), .B(n9674), .ZN(
        P1_U3271) );
  XOR2_X1 U10878 ( .A(n9677), .B(n9680), .Z(n9679) );
  OAI21_X1 U10879 ( .B1(n9679), .B2(n10016), .A(n9678), .ZN(n9800) );
  INV_X1 U10880 ( .A(n9800), .ZN(n9689) );
  XNOR2_X1 U10881 ( .A(n9681), .B(n9680), .ZN(n9802) );
  INV_X1 U10882 ( .A(n9683), .ZN(n9871) );
  AOI211_X1 U10883 ( .C1(n9683), .C2(n9696), .A(n10003), .B(n9682), .ZN(n9801)
         );
  NAND2_X1 U10884 ( .A1(n9801), .A2(n10025), .ZN(n9686) );
  AOI22_X1 U10885 ( .A1(P1_REG2_REG_21__SCAN_IN), .A2(n10033), .B1(n9684), 
        .B2(n10019), .ZN(n9685) );
  OAI211_X1 U10886 ( .C1(n9871), .C2(n10029), .A(n9686), .B(n9685), .ZN(n9687)
         );
  AOI21_X1 U10887 ( .B1(n9802), .B2(n10006), .A(n9687), .ZN(n9688) );
  OAI21_X1 U10888 ( .B1(n9689), .B2(n10033), .A(n9688), .ZN(P1_U3272) );
  XOR2_X1 U10889 ( .A(n9691), .B(n9690), .Z(n9807) );
  INV_X1 U10890 ( .A(n9807), .ZN(n9706) );
  XOR2_X1 U10891 ( .A(n9692), .B(n9691), .Z(n9695) );
  INV_X1 U10892 ( .A(n9693), .ZN(n9694) );
  OAI21_X1 U10893 ( .B1(n9695), .B2(n10016), .A(n9694), .ZN(n9805) );
  NAND2_X1 U10894 ( .A1(n9805), .A2(n9734), .ZN(n9705) );
  INV_X1 U10895 ( .A(n9696), .ZN(n9697) );
  AOI211_X1 U10896 ( .C1(n9698), .C2(n9712), .A(n10003), .B(n9697), .ZN(n9806)
         );
  INV_X1 U10897 ( .A(n9698), .ZN(n9875) );
  NOR2_X1 U10898 ( .A1(n9875), .A2(n10029), .ZN(n9703) );
  OAI22_X1 U10899 ( .A1(n9734), .A2(n9701), .B1(n9700), .B2(n9699), .ZN(n9702)
         );
  AOI211_X1 U10900 ( .C1(n9806), .C2(n10025), .A(n9703), .B(n9702), .ZN(n9704)
         );
  OAI211_X1 U10901 ( .C1(n9737), .C2(n9706), .A(n9705), .B(n9704), .ZN(
        P1_U3273) );
  NAND2_X1 U10902 ( .A1(n9707), .A2(n9717), .ZN(n9708) );
  NAND3_X1 U10903 ( .A1(n9709), .A2(n9996), .A3(n9708), .ZN(n9711) );
  OAI211_X1 U10904 ( .C1(n9879), .C2(n9728), .A(n10073), .B(n9712), .ZN(n9811)
         );
  INV_X1 U10905 ( .A(n9811), .ZN(n9716) );
  AOI22_X1 U10906 ( .A1(n10033), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9713), 
        .B2(n10019), .ZN(n9714) );
  OAI21_X1 U10907 ( .B1(n9879), .B2(n10029), .A(n9714), .ZN(n9715) );
  AOI21_X1 U10908 ( .B1(n9716), .B2(n10025), .A(n9715), .ZN(n9720) );
  XNOR2_X1 U10909 ( .A(n9718), .B(n5021), .ZN(n9810) );
  NAND2_X1 U10910 ( .A1(n9810), .A2(n10006), .ZN(n9719) );
  OAI211_X1 U10911 ( .C1(n9813), .C2(n10033), .A(n9720), .B(n9719), .ZN(
        P1_U3274) );
  XNOR2_X1 U10912 ( .A(n9721), .B(n9723), .ZN(n9820) );
  INV_X1 U10913 ( .A(n9820), .ZN(n9736) );
  XOR2_X1 U10914 ( .A(n9723), .B(n9722), .Z(n9726) );
  INV_X1 U10915 ( .A(n9724), .ZN(n9725) );
  OAI21_X1 U10916 ( .B1(n9726), .B2(n10016), .A(n9725), .ZN(n9818) );
  AND2_X1 U10917 ( .A1(n9816), .A2(n9739), .ZN(n9727) );
  OR3_X1 U10918 ( .A1(n9728), .A2(n9727), .A3(n10003), .ZN(n9817) );
  INV_X1 U10919 ( .A(n9729), .ZN(n9730) );
  AOI22_X1 U10920 ( .A1(n10033), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9730), 
        .B2(n10019), .ZN(n9732) );
  NAND2_X1 U10921 ( .A1(n9816), .A2(n9950), .ZN(n9731) );
  OAI211_X1 U10922 ( .C1(n9817), .C2(n9746), .A(n9732), .B(n9731), .ZN(n9733)
         );
  AOI21_X1 U10923 ( .B1(n9818), .B2(n9734), .A(n9733), .ZN(n9735) );
  OAI21_X1 U10924 ( .B1(n9737), .B2(n9736), .A(n9735), .ZN(P1_U3275) );
  XNOR2_X1 U10925 ( .A(n9738), .B(n9748), .ZN(n9823) );
  OAI211_X1 U10926 ( .C1(n9887), .C2(n9740), .A(n10073), .B(n9739), .ZN(n9824)
         );
  INV_X1 U10927 ( .A(n9741), .ZN(n9742) );
  AOI22_X1 U10928 ( .A1(n10033), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9742), 
        .B2(n10019), .ZN(n9745) );
  NAND2_X1 U10929 ( .A1(n9743), .A2(n9950), .ZN(n9744) );
  OAI211_X1 U10930 ( .C1(n9824), .C2(n9746), .A(n9745), .B(n9744), .ZN(n9754)
         );
  OAI211_X1 U10931 ( .C1(n9749), .C2(n9748), .A(n9747), .B(n9996), .ZN(n9752)
         );
  INV_X1 U10932 ( .A(n9750), .ZN(n9751) );
  NOR2_X1 U10933 ( .A1(n9825), .A2(n10033), .ZN(n9753) );
  AOI211_X1 U10934 ( .C1(n9823), .C2(n10006), .A(n9754), .B(n9753), .ZN(n9755)
         );
  INV_X1 U10935 ( .A(n9755), .ZN(P1_U3276) );
  NOR2_X1 U10936 ( .A1(n9757), .A2(n9756), .ZN(n9843) );
  MUX2_X1 U10937 ( .A(n6596), .B(n9843), .S(n10141), .Z(n9758) );
  OAI21_X1 U10938 ( .B1(n8161), .B2(n9837), .A(n9758), .ZN(P1_U3552) );
  INV_X1 U10939 ( .A(n10112), .ZN(n10078) );
  AOI21_X1 U10940 ( .B1(n10095), .B2(n9760), .A(n9759), .ZN(n9761) );
  OAI211_X1 U10941 ( .C1(n9763), .C2(n10078), .A(n9762), .B(n9761), .ZN(n9846)
         );
  MUX2_X1 U10942 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9846), .S(n10141), .Z(
        P1_U3550) );
  NAND2_X1 U10943 ( .A1(n9764), .A2(n10112), .ZN(n9767) );
  NAND3_X1 U10944 ( .A1(n9767), .A2(n9766), .A3(n9765), .ZN(n9847) );
  MUX2_X1 U10945 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9847), .S(n10141), .Z(
        n9768) );
  AOI21_X1 U10946 ( .B1(n6616), .B2(n9849), .A(n9768), .ZN(n9769) );
  INV_X1 U10947 ( .A(n9769), .ZN(P1_U3549) );
  NAND2_X1 U10948 ( .A1(n9770), .A2(n10112), .ZN(n9773) );
  NAND3_X1 U10949 ( .A1(n9773), .A2(n9772), .A3(n9771), .ZN(n9851) );
  MUX2_X1 U10950 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9851), .S(n10141), .Z(
        n9774) );
  AOI21_X1 U10951 ( .B1(n6616), .B2(n9853), .A(n9774), .ZN(n9775) );
  INV_X1 U10952 ( .A(n9775), .ZN(P1_U3548) );
  NAND2_X1 U10953 ( .A1(n9776), .A2(n10112), .ZN(n9778) );
  NAND3_X1 U10954 ( .A1(n9779), .A2(n9778), .A3(n9777), .ZN(n9855) );
  MUX2_X1 U10955 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9855), .S(n10141), .Z(
        n9780) );
  AOI21_X1 U10956 ( .B1(n6616), .B2(n9857), .A(n9780), .ZN(n9781) );
  INV_X1 U10957 ( .A(n9781), .ZN(P1_U3547) );
  AOI22_X1 U10958 ( .A1(n9783), .A2(n10073), .B1(n10095), .B2(n9782), .ZN(
        n9784) );
  OAI211_X1 U10959 ( .C1(n10078), .C2(n9786), .A(n9785), .B(n9784), .ZN(n9859)
         );
  MUX2_X1 U10960 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9859), .S(n10141), .Z(
        P1_U3546) );
  NAND2_X1 U10961 ( .A1(n9787), .A2(n10112), .ZN(n9792) );
  AND2_X1 U10962 ( .A1(n9789), .A2(n9788), .ZN(n9791) );
  NAND3_X1 U10963 ( .A1(n9792), .A2(n9791), .A3(n9790), .ZN(n9860) );
  MUX2_X1 U10964 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9860), .S(n10141), .Z(
        n9793) );
  AOI21_X1 U10965 ( .B1(n6616), .B2(n9862), .A(n9793), .ZN(n9794) );
  INV_X1 U10966 ( .A(n9794), .ZN(P1_U3545) );
  INV_X1 U10967 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9798) );
  AOI211_X1 U10968 ( .C1(n10112), .C2(n9797), .A(n9796), .B(n9795), .ZN(n9864)
         );
  MUX2_X1 U10969 ( .A(n9798), .B(n9864), .S(n10141), .Z(n9799) );
  OAI21_X1 U10970 ( .B1(n9867), .B2(n9837), .A(n9799), .ZN(P1_U3544) );
  INV_X1 U10971 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9803) );
  AOI211_X1 U10972 ( .C1(n10112), .C2(n9802), .A(n9801), .B(n9800), .ZN(n9868)
         );
  MUX2_X1 U10973 ( .A(n9803), .B(n9868), .S(n10141), .Z(n9804) );
  OAI21_X1 U10974 ( .B1(n9871), .B2(n9837), .A(n9804), .ZN(P1_U3543) );
  INV_X1 U10975 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9808) );
  AOI211_X1 U10976 ( .C1(n9807), .C2(n10112), .A(n9806), .B(n9805), .ZN(n9872)
         );
  MUX2_X1 U10977 ( .A(n9808), .B(n9872), .S(n10141), .Z(n9809) );
  OAI21_X1 U10978 ( .B1(n9875), .B2(n9837), .A(n9809), .ZN(P1_U3542) );
  NAND2_X1 U10979 ( .A1(n9810), .A2(n10112), .ZN(n9812) );
  NAND3_X1 U10980 ( .A1(n9813), .A2(n9812), .A3(n9811), .ZN(n9876) );
  MUX2_X1 U10981 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9876), .S(n10141), .Z(
        n9814) );
  INV_X1 U10982 ( .A(n9814), .ZN(n9815) );
  OAI21_X1 U10983 ( .B1(n9879), .B2(n9837), .A(n9815), .ZN(P1_U3541) );
  INV_X1 U10984 ( .A(n9816), .ZN(n9883) );
  INV_X1 U10985 ( .A(n9817), .ZN(n9819) );
  AOI211_X1 U10986 ( .C1(n10112), .C2(n9820), .A(n9819), .B(n9818), .ZN(n9880)
         );
  MUX2_X1 U10987 ( .A(n9821), .B(n9880), .S(n10141), .Z(n9822) );
  OAI21_X1 U10988 ( .B1(n9883), .B2(n9837), .A(n9822), .ZN(P1_U3540) );
  NAND2_X1 U10989 ( .A1(n9823), .A2(n10112), .ZN(n9826) );
  MUX2_X1 U10990 ( .A(n7594), .B(n9885), .S(n10141), .Z(n9827) );
  OAI21_X1 U10991 ( .B1(n9887), .B2(n9837), .A(n9827), .ZN(P1_U3539) );
  AOI211_X1 U10992 ( .C1(n9830), .C2(n10112), .A(n9829), .B(n9828), .ZN(n9888)
         );
  MUX2_X1 U10993 ( .A(n9831), .B(n9888), .S(n10141), .Z(n9832) );
  OAI21_X1 U10994 ( .B1(n9891), .B2(n9837), .A(n9832), .ZN(P1_U3538) );
  AOI211_X1 U10995 ( .C1(n10112), .C2(n9835), .A(n9834), .B(n9833), .ZN(n9892)
         );
  MUX2_X1 U10996 ( .A(n5651), .B(n9892), .S(n10141), .Z(n9836) );
  OAI21_X1 U10997 ( .B1(n9895), .B2(n9837), .A(n9836), .ZN(P1_U3537) );
  MUX2_X1 U10998 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9838), .S(n10141), .Z(
        P1_U3522) );
  INV_X1 U10999 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9839) );
  MUX2_X1 U11000 ( .A(n9840), .B(n9839), .S(n10123), .Z(n9841) );
  OAI21_X1 U11001 ( .B1(n9842), .B2(n9894), .A(n9841), .ZN(P1_U3521) );
  INV_X1 U11002 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9844) );
  MUX2_X1 U11003 ( .A(n9844), .B(n9843), .S(n10125), .Z(n9845) );
  OAI21_X1 U11004 ( .B1(n8161), .B2(n9894), .A(n9845), .ZN(P1_U3520) );
  MUX2_X1 U11005 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9846), .S(n10125), .Z(
        P1_U3518) );
  MUX2_X1 U11006 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9847), .S(n10125), .Z(
        n9848) );
  AOI21_X1 U11007 ( .B1(n6623), .B2(n9849), .A(n9848), .ZN(n9850) );
  INV_X1 U11008 ( .A(n9850), .ZN(P1_U3517) );
  MUX2_X1 U11009 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9851), .S(n10125), .Z(
        n9852) );
  AOI21_X1 U11010 ( .B1(n6623), .B2(n9853), .A(n9852), .ZN(n9854) );
  INV_X1 U11011 ( .A(n9854), .ZN(P1_U3516) );
  MUX2_X1 U11012 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9855), .S(n10125), .Z(
        n9856) );
  AOI21_X1 U11013 ( .B1(n6623), .B2(n9857), .A(n9856), .ZN(n9858) );
  INV_X1 U11014 ( .A(n9858), .ZN(P1_U3515) );
  MUX2_X1 U11015 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9859), .S(n10125), .Z(
        P1_U3514) );
  MUX2_X1 U11016 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9860), .S(n10125), .Z(
        n9861) );
  AOI21_X1 U11017 ( .B1(n6623), .B2(n9862), .A(n9861), .ZN(n9863) );
  INV_X1 U11018 ( .A(n9863), .ZN(P1_U3513) );
  INV_X1 U11019 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9865) );
  MUX2_X1 U11020 ( .A(n9865), .B(n9864), .S(n10125), .Z(n9866) );
  OAI21_X1 U11021 ( .B1(n9867), .B2(n9894), .A(n9866), .ZN(P1_U3512) );
  INV_X1 U11022 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9869) );
  MUX2_X1 U11023 ( .A(n9869), .B(n9868), .S(n10125), .Z(n9870) );
  OAI21_X1 U11024 ( .B1(n9871), .B2(n9894), .A(n9870), .ZN(P1_U3511) );
  INV_X1 U11025 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9873) );
  MUX2_X1 U11026 ( .A(n9873), .B(n9872), .S(n10125), .Z(n9874) );
  OAI21_X1 U11027 ( .B1(n9875), .B2(n9894), .A(n9874), .ZN(P1_U3510) );
  MUX2_X1 U11028 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9876), .S(n10125), .Z(
        n9877) );
  INV_X1 U11029 ( .A(n9877), .ZN(n9878) );
  OAI21_X1 U11030 ( .B1(n9879), .B2(n9894), .A(n9878), .ZN(P1_U3509) );
  INV_X1 U11031 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9881) );
  MUX2_X1 U11032 ( .A(n9881), .B(n9880), .S(n10125), .Z(n9882) );
  OAI21_X1 U11033 ( .B1(n9883), .B2(n9894), .A(n9882), .ZN(P1_U3507) );
  INV_X1 U11034 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9884) );
  MUX2_X1 U11035 ( .A(n9885), .B(n9884), .S(n10123), .Z(n9886) );
  OAI21_X1 U11036 ( .B1(n9887), .B2(n9894), .A(n9886), .ZN(P1_U3504) );
  INV_X1 U11037 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9889) );
  MUX2_X1 U11038 ( .A(n9889), .B(n9888), .S(n10125), .Z(n9890) );
  OAI21_X1 U11039 ( .B1(n9891), .B2(n9894), .A(n9890), .ZN(P1_U3501) );
  MUX2_X1 U11040 ( .A(n5652), .B(n9892), .S(n10125), .Z(n9893) );
  OAI21_X1 U11041 ( .B1(n9895), .B2(n9894), .A(n9893), .ZN(P1_U3498) );
  MUX2_X1 U11042 ( .A(P1_D_REG_1__SCAN_IN), .B(n9898), .S(n10035), .Z(P1_U3440) );
  NOR4_X1 U11043 ( .A1(n9900), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n9899), .ZN(n9901) );
  AOI21_X1 U11044 ( .B1(n9902), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9901), .ZN(
        n9903) );
  OAI21_X1 U11045 ( .B1(n9904), .B2(n9908), .A(n9903), .ZN(P1_U3324) );
  INV_X1 U11046 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10551) );
  OAI222_X1 U11047 ( .A1(n5275), .A2(P1_U3086), .B1(n9908), .B2(n9905), .C1(
        n10551), .C2(n9906), .ZN(P1_U3325) );
  INV_X1 U11048 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10342) );
  OAI222_X1 U11049 ( .A1(P1_U3086), .A2(n9909), .B1(n9908), .B2(n9907), .C1(
        n10342), .C2(n9906), .ZN(P1_U3326) );
  MUX2_X1 U11050 ( .A(n9910), .B(n10534), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3355) );
  INV_X1 U11051 ( .A(n9911), .ZN(n9912) );
  OAI21_X1 U11052 ( .B1(n9914), .B2(n9913), .A(n9912), .ZN(n9923) );
  INV_X1 U11053 ( .A(n9915), .ZN(n9916) );
  NAND3_X1 U11054 ( .A1(n9918), .A2(n9917), .A3(n9916), .ZN(n9920) );
  AOI21_X1 U11055 ( .B1(n9921), .B2(n9920), .A(n9919), .ZN(n9922) );
  AOI211_X1 U11056 ( .C1(n10108), .C2(n9924), .A(n9923), .B(n9922), .ZN(n9925)
         );
  OAI21_X1 U11057 ( .B1(n9927), .B2(n9926), .A(n9925), .ZN(P1_U3224) );
  XNOR2_X1 U11058 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11059 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U11060 ( .A(n9928), .ZN(n9935) );
  NAND2_X1 U11061 ( .A1(n4519), .A2(n9929), .ZN(n9933) );
  NAND2_X1 U11062 ( .A1(n9931), .A2(n9933), .ZN(n9932) );
  MUX2_X1 U11063 ( .A(n9933), .B(n9932), .S(n10534), .Z(n9934) );
  NAND2_X1 U11064 ( .A1(n9935), .A2(n9934), .ZN(n9938) );
  AOI22_X1 U11065 ( .A1(n9936), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9937) );
  OAI21_X1 U11066 ( .B1(n9939), .B2(n9938), .A(n9937), .ZN(P1_U3243) );
  OAI21_X1 U11067 ( .B1(n9942), .B2(n9941), .A(n9940), .ZN(n9947) );
  XNOR2_X1 U11068 ( .A(n9944), .B(n9943), .ZN(n9952) );
  NOR2_X1 U11069 ( .A1(n9952), .A2(n10009), .ZN(n9945) );
  AOI211_X1 U11070 ( .C1(n9996), .C2(n9947), .A(n9946), .B(n9945), .ZN(n10118)
         );
  INV_X1 U11071 ( .A(n9948), .ZN(n9949) );
  AOI222_X1 U11072 ( .A1(n9951), .A2(n9950), .B1(P1_REG2_REG_14__SCAN_IN), 
        .B2(n10033), .C1(n10019), .C2(n9949), .ZN(n9957) );
  INV_X1 U11073 ( .A(n9952), .ZN(n10121) );
  INV_X1 U11074 ( .A(n9953), .ZN(n10026) );
  OAI211_X1 U11075 ( .C1(n10117), .C2(n9954), .A(n10073), .B(n4597), .ZN(
        n10115) );
  INV_X1 U11076 ( .A(n10115), .ZN(n9955) );
  AOI22_X1 U11077 ( .A1(n10121), .A2(n10026), .B1(n10025), .B2(n9955), .ZN(
        n9956) );
  OAI211_X1 U11078 ( .C1(n10033), .C2(n10118), .A(n9957), .B(n9956), .ZN(
        P1_U3279) );
  AOI21_X1 U11079 ( .B1(n9958), .B2(n9968), .A(n10016), .ZN(n9961) );
  AOI21_X1 U11080 ( .B1(n9961), .B2(n9960), .A(n9959), .ZN(n10090) );
  INV_X1 U11081 ( .A(n9963), .ZN(n9964) );
  AOI22_X1 U11082 ( .A1(n10033), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n9964), .B2(
        n10019), .ZN(n9965) );
  OAI21_X1 U11083 ( .B1(n10029), .B2(n4919), .A(n9965), .ZN(n9966) );
  INV_X1 U11084 ( .A(n9966), .ZN(n9972) );
  XNOR2_X1 U11085 ( .A(n9967), .B(n9968), .ZN(n10092) );
  OAI211_X1 U11086 ( .C1(n4920), .C2(n4919), .A(n10073), .B(n9969), .ZN(n10089) );
  INV_X1 U11087 ( .A(n10089), .ZN(n9970) );
  AOI22_X1 U11088 ( .A1(n10092), .A2(n10006), .B1(n10025), .B2(n9970), .ZN(
        n9971) );
  OAI211_X1 U11089 ( .C1(n10033), .C2(n10090), .A(n9972), .B(n9971), .ZN(
        P1_U3285) );
  XNOR2_X1 U11090 ( .A(n9974), .B(n9973), .ZN(n9976) );
  AOI21_X1 U11091 ( .B1(n9976), .B2(n9996), .A(n9975), .ZN(n10062) );
  INV_X1 U11092 ( .A(n9977), .ZN(n9978) );
  AOI22_X1 U11093 ( .A1(n10033), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n9978), .B2(
        n10019), .ZN(n9979) );
  OAI21_X1 U11094 ( .B1(n10029), .B2(n10063), .A(n9979), .ZN(n9980) );
  INV_X1 U11095 ( .A(n9980), .ZN(n9990) );
  XNOR2_X1 U11096 ( .A(n9981), .B(n9982), .ZN(n10065) );
  NAND2_X1 U11097 ( .A1(n9984), .A2(n9983), .ZN(n9985) );
  NAND2_X1 U11098 ( .A1(n9985), .A2(n10073), .ZN(n9986) );
  OR2_X1 U11099 ( .A1(n9987), .A2(n9986), .ZN(n10061) );
  INV_X1 U11100 ( .A(n10061), .ZN(n9988) );
  AOI22_X1 U11101 ( .A1(n10065), .A2(n10006), .B1(n10025), .B2(n9988), .ZN(
        n9989) );
  OAI211_X1 U11102 ( .C1(n10033), .C2(n10062), .A(n9990), .B(n9989), .ZN(
        P1_U3289) );
  OAI21_X1 U11103 ( .B1(n9993), .B2(n9992), .A(n9991), .ZN(n9997) );
  INV_X1 U11104 ( .A(n9994), .ZN(n9995) );
  AOI21_X1 U11105 ( .B1(n9997), .B2(n9996), .A(n9995), .ZN(n10049) );
  AOI22_X1 U11106 ( .A1(n10033), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n10019), .ZN(n9998) );
  OAI21_X1 U11107 ( .B1(n10029), .B2(n10050), .A(n9998), .ZN(n9999) );
  INV_X1 U11108 ( .A(n9999), .ZN(n10008) );
  XNOR2_X1 U11109 ( .A(n10000), .B(n10001), .ZN(n10052) );
  INV_X1 U11110 ( .A(n10024), .ZN(n10004) );
  AOI211_X1 U11111 ( .C1(n10005), .C2(n10004), .A(n10003), .B(n10002), .ZN(
        n10047) );
  AOI22_X1 U11112 ( .A1(n10006), .A2(n10052), .B1(n10025), .B2(n10047), .ZN(
        n10007) );
  OAI211_X1 U11113 ( .C1(n10033), .C2(n10049), .A(n10008), .B(n10007), .ZN(
        P1_U3291) );
  INV_X1 U11114 ( .A(n10009), .ZN(n10088) );
  XNOR2_X1 U11115 ( .A(n10014), .B(n10010), .ZN(n10045) );
  INV_X1 U11116 ( .A(n10011), .ZN(n10012) );
  AOI21_X1 U11117 ( .B1(n10014), .B2(n10013), .A(n10012), .ZN(n10017) );
  OAI21_X1 U11118 ( .B1(n10017), .B2(n10016), .A(n10015), .ZN(n10018) );
  AOI21_X1 U11119 ( .B1(n10088), .B2(n10045), .A(n10018), .ZN(n10042) );
  AOI22_X1 U11120 ( .A1(n10019), .A2(P1_REG3_REG_1__SCAN_IN), .B1(
        P1_REG2_REG_1__SCAN_IN), .B2(n10033), .ZN(n10032) );
  NAND2_X1 U11121 ( .A1(n10021), .A2(n10020), .ZN(n10022) );
  NAND2_X1 U11122 ( .A1(n10073), .A2(n10022), .ZN(n10023) );
  NOR2_X1 U11123 ( .A1(n10024), .A2(n10023), .ZN(n10039) );
  NAND2_X1 U11124 ( .A1(n10025), .A2(n10039), .ZN(n10028) );
  NAND2_X1 U11125 ( .A1(n10026), .A2(n10045), .ZN(n10027) );
  OAI211_X1 U11126 ( .C1(n10041), .C2(n10029), .A(n10028), .B(n10027), .ZN(
        n10030) );
  INV_X1 U11127 ( .A(n10030), .ZN(n10031) );
  OAI211_X1 U11128 ( .C1(n10033), .C2(n10042), .A(n10032), .B(n10031), .ZN(
        P1_U3292) );
  AND2_X1 U11129 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10034), .ZN(P1_U3294) );
  AND2_X1 U11130 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10034), .ZN(P1_U3295) );
  AND2_X1 U11131 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10034), .ZN(P1_U3296) );
  AND2_X1 U11132 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10034), .ZN(P1_U3297) );
  AND2_X1 U11133 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10034), .ZN(P1_U3298) );
  AND2_X1 U11134 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10034), .ZN(P1_U3299) );
  AND2_X1 U11135 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10034), .ZN(P1_U3300) );
  AND2_X1 U11136 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10034), .ZN(P1_U3301) );
  AND2_X1 U11137 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10034), .ZN(P1_U3302) );
  AND2_X1 U11138 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10034), .ZN(P1_U3303) );
  AND2_X1 U11139 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10034), .ZN(P1_U3304) );
  AND2_X1 U11140 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10034), .ZN(P1_U3305) );
  AND2_X1 U11141 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10034), .ZN(P1_U3306) );
  AND2_X1 U11142 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10034), .ZN(P1_U3307) );
  AND2_X1 U11143 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10034), .ZN(P1_U3308) );
  AND2_X1 U11144 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10034), .ZN(P1_U3309) );
  AND2_X1 U11145 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10034), .ZN(P1_U3310) );
  AND2_X1 U11146 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10034), .ZN(P1_U3311) );
  AND2_X1 U11147 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10034), .ZN(P1_U3312) );
  AND2_X1 U11148 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10034), .ZN(P1_U3313) );
  AND2_X1 U11149 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10034), .ZN(P1_U3314) );
  AND2_X1 U11150 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10034), .ZN(P1_U3315) );
  AND2_X1 U11151 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10034), .ZN(P1_U3316) );
  AND2_X1 U11152 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10034), .ZN(P1_U3317) );
  AND2_X1 U11153 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10034), .ZN(P1_U3318) );
  AND2_X1 U11154 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10034), .ZN(P1_U3319) );
  INV_X1 U11155 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10604) );
  NOR2_X1 U11156 ( .A1(n10035), .A2(n10604), .ZN(P1_U3320) );
  INV_X1 U11157 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10562) );
  NOR2_X1 U11158 ( .A1(n10035), .A2(n10562), .ZN(P1_U3321) );
  INV_X1 U11159 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10575) );
  NOR2_X1 U11160 ( .A1(n10035), .A2(n10575), .ZN(P1_U3322) );
  INV_X1 U11161 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10393) );
  NOR2_X1 U11162 ( .A1(n10035), .A2(n10393), .ZN(P1_U3323) );
  INV_X1 U11163 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10037) );
  AOI21_X1 U11164 ( .B1(n10038), .B2(n10037), .A(n10036), .ZN(P1_U3439) );
  INV_X1 U11165 ( .A(n10039), .ZN(n10040) );
  OAI21_X1 U11166 ( .B1(n10041), .B2(n10116), .A(n10040), .ZN(n10044) );
  INV_X1 U11167 ( .A(n10042), .ZN(n10043) );
  AOI211_X1 U11168 ( .C1(n10122), .C2(n10045), .A(n10044), .B(n10043), .ZN(
        n10126) );
  INV_X1 U11169 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10046) );
  AOI22_X1 U11170 ( .A1(n10125), .A2(n10126), .B1(n10046), .B2(n10123), .ZN(
        P1_U3456) );
  INV_X1 U11171 ( .A(n10047), .ZN(n10048) );
  OAI211_X1 U11172 ( .C1(n10050), .C2(n10116), .A(n10049), .B(n10048), .ZN(
        n10051) );
  AOI21_X1 U11173 ( .B1(n10112), .B2(n10052), .A(n10051), .ZN(n10127) );
  INV_X1 U11174 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10053) );
  AOI22_X1 U11175 ( .A1(n10125), .A2(n10127), .B1(n10053), .B2(n10123), .ZN(
        P1_U3459) );
  OAI21_X1 U11176 ( .B1(n10055), .B2(n10116), .A(n10054), .ZN(n10058) );
  INV_X1 U11177 ( .A(n10056), .ZN(n10057) );
  AOI211_X1 U11178 ( .C1(n10059), .C2(n10112), .A(n10058), .B(n10057), .ZN(
        n10128) );
  INV_X1 U11179 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10060) );
  AOI22_X1 U11180 ( .A1(n10125), .A2(n10128), .B1(n10060), .B2(n10123), .ZN(
        P1_U3462) );
  OAI211_X1 U11181 ( .C1(n10063), .C2(n10116), .A(n10062), .B(n10061), .ZN(
        n10064) );
  AOI21_X1 U11182 ( .B1(n10112), .B2(n10065), .A(n10064), .ZN(n10129) );
  AOI22_X1 U11183 ( .A1(n10125), .A2(n10129), .B1(n5381), .B2(n10123), .ZN(
        P1_U3465) );
  AOI21_X1 U11184 ( .B1(n10095), .B2(n10067), .A(n10066), .ZN(n10068) );
  OAI211_X1 U11185 ( .C1(n10078), .C2(n10070), .A(n10069), .B(n10068), .ZN(
        n10071) );
  INV_X1 U11186 ( .A(n10071), .ZN(n10130) );
  AOI22_X1 U11187 ( .A1(n10125), .A2(n10130), .B1(n5408), .B2(n10123), .ZN(
        P1_U3468) );
  AOI22_X1 U11188 ( .A1(n10074), .A2(n10073), .B1(n10095), .B2(n10072), .ZN(
        n10075) );
  OAI211_X1 U11189 ( .C1(n10078), .C2(n10077), .A(n10076), .B(n10075), .ZN(
        n10079) );
  INV_X1 U11190 ( .A(n10079), .ZN(n10132) );
  AOI22_X1 U11191 ( .A1(n10125), .A2(n10132), .B1(n5445), .B2(n10123), .ZN(
        P1_U3471) );
  INV_X1 U11192 ( .A(n10085), .ZN(n10087) );
  AOI21_X1 U11193 ( .B1(n10095), .B2(n10081), .A(n10080), .ZN(n10082) );
  OAI211_X1 U11194 ( .C1(n10085), .C2(n10084), .A(n10083), .B(n10082), .ZN(
        n10086) );
  AOI21_X1 U11195 ( .B1(n10088), .B2(n10087), .A(n10086), .ZN(n10134) );
  AOI22_X1 U11196 ( .A1(n10125), .A2(n10134), .B1(n5429), .B2(n10123), .ZN(
        P1_U3474) );
  OAI211_X1 U11197 ( .C1(n4919), .C2(n10116), .A(n10090), .B(n10089), .ZN(
        n10091) );
  AOI21_X1 U11198 ( .B1(n10112), .B2(n10092), .A(n10091), .ZN(n10135) );
  INV_X1 U11199 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10093) );
  AOI22_X1 U11200 ( .A1(n10125), .A2(n10135), .B1(n10093), .B2(n10123), .ZN(
        P1_U3477) );
  AND2_X1 U11201 ( .A1(n10094), .A2(n10112), .ZN(n10099) );
  AND2_X1 U11202 ( .A1(n10096), .A2(n10095), .ZN(n10098) );
  NOR4_X1 U11203 ( .A1(n10100), .A2(n10099), .A3(n10098), .A4(n10097), .ZN(
        n10136) );
  INV_X1 U11204 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10101) );
  AOI22_X1 U11205 ( .A1(n10125), .A2(n10136), .B1(n10101), .B2(n10123), .ZN(
        P1_U3480) );
  OAI21_X1 U11206 ( .B1(n10103), .B2(n10116), .A(n10102), .ZN(n10105) );
  AOI211_X1 U11207 ( .C1(n10112), .C2(n10106), .A(n10105), .B(n10104), .ZN(
        n10137) );
  INV_X1 U11208 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10107) );
  AOI22_X1 U11209 ( .A1(n10125), .A2(n10137), .B1(n10107), .B2(n10123), .ZN(
        P1_U3483) );
  OAI211_X1 U11210 ( .C1(n4932), .C2(n10116), .A(n10110), .B(n10109), .ZN(
        n10111) );
  AOI21_X1 U11211 ( .B1(n10113), .B2(n10112), .A(n10111), .ZN(n10138) );
  INV_X1 U11212 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10114) );
  AOI22_X1 U11213 ( .A1(n10125), .A2(n10138), .B1(n10114), .B2(n10123), .ZN(
        P1_U3489) );
  OAI21_X1 U11214 ( .B1(n10117), .B2(n10116), .A(n10115), .ZN(n10120) );
  INV_X1 U11215 ( .A(n10118), .ZN(n10119) );
  AOI211_X1 U11216 ( .C1(n10122), .C2(n10121), .A(n10120), .B(n10119), .ZN(
        n10140) );
  INV_X1 U11217 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10124) );
  AOI22_X1 U11218 ( .A1(n10125), .A2(n10140), .B1(n10124), .B2(n10123), .ZN(
        P1_U3495) );
  AOI22_X1 U11219 ( .A1(n10141), .A2(n10126), .B1(n6794), .B2(n10139), .ZN(
        P1_U3523) );
  AOI22_X1 U11220 ( .A1(n10141), .A2(n10127), .B1(n6793), .B2(n10139), .ZN(
        P1_U3524) );
  AOI22_X1 U11221 ( .A1(n10141), .A2(n10128), .B1(n6797), .B2(n10139), .ZN(
        P1_U3525) );
  AOI22_X1 U11222 ( .A1(n10141), .A2(n10129), .B1(n6800), .B2(n10139), .ZN(
        P1_U3526) );
  AOI22_X1 U11223 ( .A1(n10141), .A2(n10130), .B1(n6803), .B2(n10139), .ZN(
        P1_U3527) );
  AOI22_X1 U11224 ( .A1(n10141), .A2(n10132), .B1(n10131), .B2(n10139), .ZN(
        P1_U3528) );
  AOI22_X1 U11225 ( .A1(n10141), .A2(n10134), .B1(n10133), .B2(n10139), .ZN(
        P1_U3529) );
  AOI22_X1 U11226 ( .A1(n10141), .A2(n10135), .B1(n6792), .B2(n10139), .ZN(
        P1_U3530) );
  AOI22_X1 U11227 ( .A1(n10141), .A2(n10136), .B1(n5500), .B2(n10139), .ZN(
        P1_U3531) );
  AOI22_X1 U11228 ( .A1(n10141), .A2(n10137), .B1(n6879), .B2(n10139), .ZN(
        P1_U3532) );
  AOI22_X1 U11229 ( .A1(n10141), .A2(n10138), .B1(n7077), .B2(n10139), .ZN(
        P1_U3534) );
  AOI22_X1 U11230 ( .A1(n10141), .A2(n10140), .B1(n5631), .B2(n10139), .ZN(
        P1_U3536) );
  INV_X1 U11231 ( .A(n10142), .ZN(n10143) );
  AOI21_X1 U11232 ( .B1(n6660), .B2(n10144), .A(n10143), .ZN(n10153) );
  NAND2_X1 U11233 ( .A1(n10145), .A2(P2_ADDR_REG_1__SCAN_IN), .ZN(n10151) );
  OAI211_X1 U11234 ( .C1(n10149), .C2(n10148), .A(n10147), .B(n10146), .ZN(
        n10150) );
  OAI211_X1 U11235 ( .C1(n10153), .C2(n10152), .A(n10151), .B(n10150), .ZN(
        n10154) );
  AOI21_X1 U11236 ( .B1(n10156), .B2(n10155), .A(n10154), .ZN(n10163) );
  INV_X1 U11237 ( .A(n10157), .ZN(n10159) );
  OAI21_X1 U11238 ( .B1(n10159), .B2(P2_REG2_REG_1__SCAN_IN), .A(n10158), .ZN(
        n10160) );
  NAND2_X1 U11239 ( .A1(n10161), .A2(n10160), .ZN(n10162) );
  OAI211_X1 U11240 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n7319), .A(n10163), .B(
        n10162), .ZN(P2_U3183) );
  AOI21_X1 U11241 ( .B1(n10166), .B2(n10165), .A(n10164), .ZN(n10167) );
  OAI222_X1 U11242 ( .A1(n10171), .A2(n10170), .B1(n10169), .B2(n10168), .C1(
        n8636), .C2(n10167), .ZN(n10172) );
  INV_X1 U11243 ( .A(n10172), .ZN(n10173) );
  OAI21_X1 U11244 ( .B1(n10174), .B2(n6074), .A(n10173), .ZN(P2_U3229) );
  INV_X1 U11245 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10178) );
  OAI22_X1 U11246 ( .A1(n10175), .A2(n10208), .B1(n7318), .B2(n10215), .ZN(
        n10176) );
  NOR2_X1 U11247 ( .A1(n10177), .A2(n10176), .ZN(n10224) );
  AOI22_X1 U11248 ( .A1(n10223), .A2(n10178), .B1(n10224), .B2(n10221), .ZN(
        P2_U3393) );
  INV_X1 U11249 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10185) );
  INV_X1 U11250 ( .A(n10179), .ZN(n10183) );
  INV_X1 U11251 ( .A(n10180), .ZN(n10182) );
  AOI211_X1 U11252 ( .C1(n10184), .C2(n10183), .A(n10182), .B(n10181), .ZN(
        n10225) );
  AOI22_X1 U11253 ( .A1(n10223), .A2(n10185), .B1(n10225), .B2(n10221), .ZN(
        P2_U3396) );
  INV_X1 U11254 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10190) );
  OAI22_X1 U11255 ( .A1(n10187), .A2(n10217), .B1(n10186), .B2(n10215), .ZN(
        n10188) );
  NOR2_X1 U11256 ( .A1(n10189), .A2(n10188), .ZN(n10226) );
  AOI22_X1 U11257 ( .A1(n10223), .A2(n10190), .B1(n10226), .B2(n10221), .ZN(
        P2_U3399) );
  INV_X1 U11258 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10197) );
  INV_X1 U11259 ( .A(n10191), .ZN(n10195) );
  OAI21_X1 U11260 ( .B1(n10193), .B2(n10215), .A(n10192), .ZN(n10194) );
  AOI21_X1 U11261 ( .B1(n10196), .B2(n10195), .A(n10194), .ZN(n10227) );
  AOI22_X1 U11262 ( .A1(n10223), .A2(n10197), .B1(n10227), .B2(n10221), .ZN(
        P2_U3405) );
  INV_X1 U11263 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10202) );
  NOR2_X1 U11264 ( .A1(n10198), .A2(n10208), .ZN(n10200) );
  AOI211_X1 U11265 ( .C1(n10213), .C2(n10201), .A(n10200), .B(n10199), .ZN(
        n10228) );
  AOI22_X1 U11266 ( .A1(n10223), .A2(n10202), .B1(n10228), .B2(n10221), .ZN(
        P2_U3411) );
  INV_X1 U11267 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10207) );
  OAI22_X1 U11268 ( .A1(n10204), .A2(n10217), .B1(n10203), .B2(n10215), .ZN(
        n10205) );
  NOR2_X1 U11269 ( .A1(n10206), .A2(n10205), .ZN(n10229) );
  AOI22_X1 U11270 ( .A1(n10223), .A2(n10207), .B1(n10229), .B2(n10221), .ZN(
        P2_U3414) );
  INV_X1 U11271 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10214) );
  NOR2_X1 U11272 ( .A1(n10209), .A2(n10208), .ZN(n10211) );
  AOI211_X1 U11273 ( .C1(n10213), .C2(n10212), .A(n10211), .B(n10210), .ZN(
        n10230) );
  AOI22_X1 U11274 ( .A1(n10223), .A2(n10214), .B1(n10230), .B2(n10221), .ZN(
        P2_U3420) );
  INV_X1 U11275 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10222) );
  OAI22_X1 U11276 ( .A1(n10218), .A2(n10217), .B1(n10216), .B2(n10215), .ZN(
        n10219) );
  NOR2_X1 U11277 ( .A1(n10220), .A2(n10219), .ZN(n10232) );
  AOI22_X1 U11278 ( .A1(n10223), .A2(n10222), .B1(n10232), .B2(n10221), .ZN(
        P2_U3423) );
  AOI22_X1 U11279 ( .A1(n10233), .A2(n10224), .B1(n6660), .B2(n10231), .ZN(
        P2_U3460) );
  AOI22_X1 U11280 ( .A1(n10233), .A2(n10225), .B1(n6021), .B2(n10231), .ZN(
        P2_U3461) );
  AOI22_X1 U11281 ( .A1(n10233), .A2(n10226), .B1(n6057), .B2(n10231), .ZN(
        P2_U3462) );
  AOI22_X1 U11282 ( .A1(n10233), .A2(n10227), .B1(n6659), .B2(n10231), .ZN(
        P2_U3464) );
  AOI22_X1 U11283 ( .A1(n10233), .A2(n10228), .B1(n6675), .B2(n10231), .ZN(
        P2_U3466) );
  AOI22_X1 U11284 ( .A1(n10233), .A2(n10229), .B1(n6134), .B2(n10231), .ZN(
        P2_U3467) );
  AOI22_X1 U11285 ( .A1(n10233), .A2(n10230), .B1(n6167), .B2(n10231), .ZN(
        P2_U3469) );
  AOI22_X1 U11286 ( .A1(n10233), .A2(n10232), .B1(n6176), .B2(n10231), .ZN(
        P2_U3470) );
  AOI21_X1 U11287 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10239) );
  INV_X1 U11288 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10235) );
  NAND2_X1 U11289 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n10234) );
  NOR2_X1 U11290 ( .A1(n10235), .A2(n10234), .ZN(n10237) );
  NOR2_X1 U11291 ( .A1(n10239), .A2(n10237), .ZN(n10236) );
  XOR2_X1 U11292 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10236), .Z(ADD_1068_U5) );
  XOR2_X1 U11293 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  NOR2_X1 U11294 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10288) );
  NOR2_X1 U11295 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10285) );
  NOR2_X1 U11296 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10281) );
  NOR2_X1 U11297 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10277) );
  NOR2_X1 U11298 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10273) );
  NOR2_X1 U11299 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10269) );
  NOR2_X1 U11300 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10265) );
  NOR2_X1 U11301 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10261) );
  NOR2_X1 U11302 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n10257) );
  NOR2_X1 U11303 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10253) );
  NOR2_X1 U11304 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10251) );
  NOR2_X1 U11305 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n10249) );
  NOR2_X1 U11306 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10247) );
  NOR2_X1 U11307 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10245) );
  NAND2_X1 U11308 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n10243) );
  XOR2_X1 U11309 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10701) );
  NAND2_X1 U11310 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n10241) );
  NOR2_X1 U11311 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n10237), .ZN(n10238) );
  NOR2_X1 U11312 ( .A1(n10239), .A2(n10238), .ZN(n10691) );
  XOR2_X1 U11313 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10690) );
  NAND2_X1 U11314 ( .A1(n10691), .A2(n10690), .ZN(n10240) );
  NAND2_X1 U11315 ( .A1(n10241), .A2(n10240), .ZN(n10700) );
  NAND2_X1 U11316 ( .A1(n10701), .A2(n10700), .ZN(n10242) );
  NAND2_X1 U11317 ( .A1(n10243), .A2(n10242), .ZN(n10703) );
  XNOR2_X1 U11318 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10702) );
  NOR2_X1 U11319 ( .A1(n10703), .A2(n10702), .ZN(n10244) );
  NOR2_X1 U11320 ( .A1(n10245), .A2(n10244), .ZN(n10693) );
  XNOR2_X1 U11321 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10692) );
  NOR2_X1 U11322 ( .A1(n10693), .A2(n10692), .ZN(n10246) );
  NOR2_X1 U11323 ( .A1(n10247), .A2(n10246), .ZN(n10699) );
  XNOR2_X1 U11324 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n10698) );
  NOR2_X1 U11325 ( .A1(n10699), .A2(n10698), .ZN(n10248) );
  NOR2_X1 U11326 ( .A1(n10249), .A2(n10248), .ZN(n10695) );
  XNOR2_X1 U11327 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10694) );
  NOR2_X1 U11328 ( .A1(n10695), .A2(n10694), .ZN(n10250) );
  NOR2_X1 U11329 ( .A1(n10251), .A2(n10250), .ZN(n10697) );
  XNOR2_X1 U11330 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10696) );
  NOR2_X1 U11331 ( .A1(n10697), .A2(n10696), .ZN(n10252) );
  NOR2_X1 U11332 ( .A1(n10253), .A2(n10252), .ZN(n10689) );
  INV_X1 U11333 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10255) );
  AOI22_X1 U11334 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10255), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n10254), .ZN(n10688) );
  NOR2_X1 U11335 ( .A1(n10689), .A2(n10688), .ZN(n10256) );
  NOR2_X1 U11336 ( .A1(n10257), .A2(n10256), .ZN(n10305) );
  INV_X1 U11337 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10259) );
  AOI22_X1 U11338 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n10259), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n10258), .ZN(n10304) );
  NOR2_X1 U11339 ( .A1(n10305), .A2(n10304), .ZN(n10260) );
  NOR2_X1 U11340 ( .A1(n10261), .A2(n10260), .ZN(n10303) );
  INV_X1 U11341 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10263) );
  AOI22_X1 U11342 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n10263), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n10262), .ZN(n10302) );
  NOR2_X1 U11343 ( .A1(n10303), .A2(n10302), .ZN(n10264) );
  NOR2_X1 U11344 ( .A1(n10265), .A2(n10264), .ZN(n10301) );
  INV_X1 U11345 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10267) );
  INV_X1 U11346 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n10266) );
  AOI22_X1 U11347 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n10267), .B1(
        P1_ADDR_REG_12__SCAN_IN), .B2(n10266), .ZN(n10300) );
  NOR2_X1 U11348 ( .A1(n10301), .A2(n10300), .ZN(n10268) );
  NOR2_X1 U11349 ( .A1(n10269), .A2(n10268), .ZN(n10299) );
  INV_X1 U11350 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10271) );
  AOI22_X1 U11351 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(n10271), .B1(
        P1_ADDR_REG_13__SCAN_IN), .B2(n10270), .ZN(n10298) );
  NOR2_X1 U11352 ( .A1(n10299), .A2(n10298), .ZN(n10272) );
  NOR2_X1 U11353 ( .A1(n10273), .A2(n10272), .ZN(n10297) );
  INV_X1 U11354 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10275) );
  AOI22_X1 U11355 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n10275), .B1(
        P1_ADDR_REG_14__SCAN_IN), .B2(n10274), .ZN(n10296) );
  NOR2_X1 U11356 ( .A1(n10297), .A2(n10296), .ZN(n10276) );
  NOR2_X1 U11357 ( .A1(n10277), .A2(n10276), .ZN(n10295) );
  INV_X1 U11358 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10279) );
  AOI22_X1 U11359 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n10279), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n10278), .ZN(n10294) );
  NOR2_X1 U11360 ( .A1(n10295), .A2(n10294), .ZN(n10280) );
  NOR2_X1 U11361 ( .A1(n10281), .A2(n10280), .ZN(n10293) );
  INV_X1 U11362 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10283) );
  AOI22_X1 U11363 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n10283), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n10282), .ZN(n10292) );
  NOR2_X1 U11364 ( .A1(n10293), .A2(n10292), .ZN(n10284) );
  NOR2_X1 U11365 ( .A1(n10285), .A2(n10284), .ZN(n10291) );
  AOI22_X1 U11366 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n7592), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(n10286), .ZN(n10290) );
  NOR2_X1 U11367 ( .A1(n10291), .A2(n10290), .ZN(n10287) );
  NOR2_X1 U11368 ( .A1(n10288), .A2(n10287), .ZN(n10306) );
  NAND2_X1 U11369 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10306), .ZN(n10307) );
  OAI21_X1 U11370 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n10306), .A(n10307), 
        .ZN(n10289) );
  XNOR2_X1 U11371 ( .A(n10289), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1068_U55)
         );
  XNOR2_X1 U11372 ( .A(n10291), .B(n10290), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11373 ( .A(n10293), .B(n10292), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11374 ( .A(n10295), .B(n10294), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11375 ( .A(n10297), .B(n10296), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11376 ( .A(n10299), .B(n10298), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11377 ( .A(n10301), .B(n10300), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11378 ( .A(n10303), .B(n10302), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11379 ( .A(n10305), .B(n10304), .ZN(ADD_1068_U63) );
  XOR2_X1 U11380 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .Z(n10687) );
  NOR2_X1 U11381 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10306), .ZN(n10308) );
  OAI21_X1 U11382 ( .B1(n10309), .B2(n10308), .A(n10307), .ZN(n10685) );
  OAI22_X1 U11383 ( .A1(SI_10_), .A2(keyinput_g22), .B1(P1_IR_REG_9__SCAN_IN), 
        .B2(keyinput_g99), .ZN(n10310) );
  AOI221_X1 U11384 ( .B1(SI_10_), .B2(keyinput_g22), .C1(keyinput_g99), .C2(
        P1_IR_REG_9__SCAN_IN), .A(n10310), .ZN(n10317) );
  OAI22_X1 U11385 ( .A1(SI_29_), .A2(keyinput_g3), .B1(SI_13_), .B2(
        keyinput_g19), .ZN(n10311) );
  AOI221_X1 U11386 ( .B1(SI_29_), .B2(keyinput_g3), .C1(keyinput_g19), .C2(
        SI_13_), .A(n10311), .ZN(n10316) );
  OAI22_X1 U11387 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_g49), .B1(
        keyinput_g80), .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n10312) );
  AOI221_X1 U11388 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_g49), .C1(
        P2_DATAO_REG_16__SCAN_IN), .C2(keyinput_g80), .A(n10312), .ZN(n10315)
         );
  OAI22_X1 U11389 ( .A1(SI_26_), .A2(keyinput_g6), .B1(P1_IR_REG_24__SCAN_IN), 
        .B2(keyinput_g114), .ZN(n10313) );
  AOI221_X1 U11390 ( .B1(SI_26_), .B2(keyinput_g6), .C1(keyinput_g114), .C2(
        P1_IR_REG_24__SCAN_IN), .A(n10313), .ZN(n10314) );
  NAND4_X1 U11391 ( .A1(n10317), .A2(n10316), .A3(n10315), .A4(n10314), .ZN(
        n10350) );
  OAI22_X1 U11392 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(keyinput_g112), .B1(
        P1_IR_REG_25__SCAN_IN), .B2(keyinput_g115), .ZN(n10318) );
  AOI221_X1 U11393 ( .B1(P1_IR_REG_22__SCAN_IN), .B2(keyinput_g112), .C1(
        keyinput_g115), .C2(P1_IR_REG_25__SCAN_IN), .A(n10318), .ZN(n10325) );
  OAI22_X1 U11394 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(keyinput_g55), .B1(
        keyinput_g23), .B2(SI_9_), .ZN(n10319) );
  AOI221_X1 U11395 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_g55), .C1(
        SI_9_), .C2(keyinput_g23), .A(n10319), .ZN(n10324) );
  OAI22_X1 U11396 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(keyinput_g45), .B1(
        P1_IR_REG_31__SCAN_IN), .B2(keyinput_g121), .ZN(n10320) );
  AOI221_X1 U11397 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_g45), .C1(
        keyinput_g121), .C2(P1_IR_REG_31__SCAN_IN), .A(n10320), .ZN(n10323) );
  OAI22_X1 U11398 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(keyinput_g35), .B1(
        keyinput_g40), .B2(P2_REG3_REG_3__SCAN_IN), .ZN(n10321) );
  AOI221_X1 U11399 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput_g35), .C1(
        P2_REG3_REG_3__SCAN_IN), .C2(keyinput_g40), .A(n10321), .ZN(n10322) );
  NAND4_X1 U11400 ( .A1(n10325), .A2(n10324), .A3(n10323), .A4(n10322), .ZN(
        n10349) );
  OAI22_X1 U11401 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(keyinput_g58), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(keyinput_g83), .ZN(n10326) );
  AOI221_X1 U11402 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput_g58), .C1(
        keyinput_g83), .C2(P2_DATAO_REG_13__SCAN_IN), .A(n10326), .ZN(n10333)
         );
  OAI22_X1 U11403 ( .A1(SI_25_), .A2(keyinput_g7), .B1(keyinput_g109), .B2(
        P1_IR_REG_19__SCAN_IN), .ZN(n10327) );
  AOI221_X1 U11404 ( .B1(SI_25_), .B2(keyinput_g7), .C1(P1_IR_REG_19__SCAN_IN), 
        .C2(keyinput_g109), .A(n10327), .ZN(n10332) );
  OAI22_X1 U11405 ( .A1(P2_RD_REG_SCAN_IN), .A2(keyinput_g33), .B1(
        keyinput_g29), .B2(SI_3_), .ZN(n10328) );
  AOI221_X1 U11406 ( .B1(P2_RD_REG_SCAN_IN), .B2(keyinput_g33), .C1(SI_3_), 
        .C2(keyinput_g29), .A(n10328), .ZN(n10331) );
  OAI22_X1 U11407 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_g43), .B1(
        P1_IR_REG_14__SCAN_IN), .B2(keyinput_g104), .ZN(n10329) );
  AOI221_X1 U11408 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_g43), .C1(
        keyinput_g104), .C2(P1_IR_REG_14__SCAN_IN), .A(n10329), .ZN(n10330) );
  NAND4_X1 U11409 ( .A1(n10333), .A2(n10332), .A3(n10331), .A4(n10330), .ZN(
        n10348) );
  INV_X1 U11410 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10334) );
  XNOR2_X1 U11411 ( .A(n10334), .B(keyinput_g123), .ZN(n10339) );
  XOR2_X1 U11412 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_g54), .Z(n10338) );
  XNOR2_X1 U11413 ( .A(n10335), .B(keyinput_g111), .ZN(n10337) );
  XNOR2_X1 U11414 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_g74), .ZN(n10336) );
  NOR4_X1 U11415 ( .A1(n10339), .A2(n10338), .A3(n10337), .A4(n10336), .ZN(
        n10346) );
  INV_X1 U11416 ( .A(n10534), .ZN(n10341) );
  OAI22_X1 U11417 ( .A1(n10342), .A2(keyinput_g67), .B1(n10341), .B2(
        keyinput_g90), .ZN(n10340) );
  AOI221_X1 U11418 ( .B1(n10342), .B2(keyinput_g67), .C1(keyinput_g90), .C2(
        n10341), .A(n10340), .ZN(n10345) );
  OAI22_X1 U11419 ( .A1(SI_17_), .A2(keyinput_g15), .B1(P1_D_REG_4__SCAN_IN), 
        .B2(keyinput_g126), .ZN(n10343) );
  AOI221_X1 U11420 ( .B1(SI_17_), .B2(keyinput_g15), .C1(keyinput_g126), .C2(
        P1_D_REG_4__SCAN_IN), .A(n10343), .ZN(n10344) );
  NAND3_X1 U11421 ( .A1(n10346), .A2(n10345), .A3(n10344), .ZN(n10347) );
  NOR4_X1 U11422 ( .A1(n10350), .A2(n10349), .A3(n10348), .A4(n10347), .ZN(
        n10683) );
  OAI22_X1 U11423 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(keyinput_g69), .B1(
        keyinput_g2), .B2(SI_30_), .ZN(n10351) );
  AOI221_X1 U11424 ( .B1(P2_DATAO_REG_27__SCAN_IN), .B2(keyinput_g69), .C1(
        SI_30_), .C2(keyinput_g2), .A(n10351), .ZN(n10358) );
  OAI22_X1 U11425 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_g60), .B1(
        P1_IR_REG_15__SCAN_IN), .B2(keyinput_g105), .ZN(n10352) );
  AOI221_X1 U11426 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .C1(
        keyinput_g105), .C2(P1_IR_REG_15__SCAN_IN), .A(n10352), .ZN(n10357) );
  OAI22_X1 U11427 ( .A1(SI_19_), .A2(keyinput_g13), .B1(keyinput_g122), .B2(
        P1_D_REG_0__SCAN_IN), .ZN(n10353) );
  AOI221_X1 U11428 ( .B1(SI_19_), .B2(keyinput_g13), .C1(P1_D_REG_0__SCAN_IN), 
        .C2(keyinput_g122), .A(n10353), .ZN(n10356) );
  OAI22_X1 U11429 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(keyinput_g71), .B1(
        P1_IR_REG_26__SCAN_IN), .B2(keyinput_g116), .ZN(n10354) );
  AOI221_X1 U11430 ( .B1(P2_DATAO_REG_25__SCAN_IN), .B2(keyinput_g71), .C1(
        keyinput_g116), .C2(P1_IR_REG_26__SCAN_IN), .A(n10354), .ZN(n10355) );
  NAND4_X1 U11431 ( .A1(n10358), .A2(n10357), .A3(n10356), .A4(n10355), .ZN(
        n10486) );
  OAI22_X1 U11432 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(keyinput_g87), .B1(
        P1_IR_REG_18__SCAN_IN), .B2(keyinput_g108), .ZN(n10359) );
  AOI221_X1 U11433 ( .B1(P2_DATAO_REG_9__SCAN_IN), .B2(keyinput_g87), .C1(
        keyinput_g108), .C2(P1_IR_REG_18__SCAN_IN), .A(n10359), .ZN(n10384) );
  OAI22_X1 U11434 ( .A1(SI_15_), .A2(keyinput_g17), .B1(keyinput_g110), .B2(
        P1_IR_REG_20__SCAN_IN), .ZN(n10360) );
  AOI221_X1 U11435 ( .B1(SI_15_), .B2(keyinput_g17), .C1(P1_IR_REG_20__SCAN_IN), .C2(keyinput_g110), .A(n10360), .ZN(n10363) );
  OAI22_X1 U11436 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput_g42), .B1(
        keyinput_g68), .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n10361) );
  AOI221_X1 U11437 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput_g42), .C1(
        P2_DATAO_REG_28__SCAN_IN), .C2(keyinput_g68), .A(n10361), .ZN(n10362)
         );
  OAI211_X1 U11438 ( .C1(n10645), .C2(keyinput_g84), .A(n10363), .B(n10362), 
        .ZN(n10364) );
  AOI21_X1 U11439 ( .B1(n10645), .B2(keyinput_g84), .A(n10364), .ZN(n10383) );
  AOI22_X1 U11440 ( .A1(SI_21_), .A2(keyinput_g11), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(keyinput_g50), .ZN(n10365) );
  OAI221_X1 U11441 ( .B1(SI_21_), .B2(keyinput_g11), .C1(
        P2_REG3_REG_17__SCAN_IN), .C2(keyinput_g50), .A(n10365), .ZN(n10372)
         );
  AOI22_X1 U11442 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(keyinput_g100), .B1(SI_22_), .B2(keyinput_g10), .ZN(n10366) );
  OAI221_X1 U11443 ( .B1(P1_IR_REG_10__SCAN_IN), .B2(keyinput_g100), .C1(
        SI_22_), .C2(keyinput_g10), .A(n10366), .ZN(n10371) );
  AOI22_X1 U11444 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(keyinput_g94), .B1(
        P2_REG3_REG_10__SCAN_IN), .B2(keyinput_g39), .ZN(n10367) );
  OAI221_X1 U11445 ( .B1(P1_IR_REG_4__SCAN_IN), .B2(keyinput_g94), .C1(
        P2_REG3_REG_10__SCAN_IN), .C2(keyinput_g39), .A(n10367), .ZN(n10370)
         );
  AOI22_X1 U11446 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_g59), .B1(SI_6_), 
        .B2(keyinput_g26), .ZN(n10368) );
  OAI221_X1 U11447 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .C1(SI_6_), .C2(keyinput_g26), .A(n10368), .ZN(n10369) );
  NOR4_X1 U11448 ( .A1(n10372), .A2(n10371), .A3(n10370), .A4(n10369), .ZN(
        n10382) );
  AOI22_X1 U11449 ( .A1(SI_31_), .A2(keyinput_g1), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(keyinput_g85), .ZN(n10373) );
  OAI221_X1 U11450 ( .B1(SI_31_), .B2(keyinput_g1), .C1(
        P2_DATAO_REG_11__SCAN_IN), .C2(keyinput_g85), .A(n10373), .ZN(n10380)
         );
  AOI22_X1 U11451 ( .A1(P1_D_REG_5__SCAN_IN), .A2(keyinput_g127), .B1(SI_4_), 
        .B2(keyinput_g28), .ZN(n10374) );
  OAI221_X1 U11452 ( .B1(P1_D_REG_5__SCAN_IN), .B2(keyinput_g127), .C1(SI_4_), 
        .C2(keyinput_g28), .A(n10374), .ZN(n10379) );
  AOI22_X1 U11453 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(keyinput_g103), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(keyinput_g44), .ZN(n10375) );
  OAI221_X1 U11454 ( .B1(P1_IR_REG_13__SCAN_IN), .B2(keyinput_g103), .C1(
        P2_REG3_REG_1__SCAN_IN), .C2(keyinput_g44), .A(n10375), .ZN(n10378) );
  AOI22_X1 U11455 ( .A1(P1_D_REG_3__SCAN_IN), .A2(keyinput_g125), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(keyinput_g75), .ZN(n10376) );
  OAI221_X1 U11456 ( .B1(P1_D_REG_3__SCAN_IN), .B2(keyinput_g125), .C1(
        P2_DATAO_REG_21__SCAN_IN), .C2(keyinput_g75), .A(n10376), .ZN(n10377)
         );
  NOR4_X1 U11457 ( .A1(n10380), .A2(n10379), .A3(n10378), .A4(n10377), .ZN(
        n10381) );
  NAND4_X1 U11458 ( .A1(n10384), .A2(n10383), .A3(n10382), .A4(n10381), .ZN(
        n10485) );
  AOI22_X1 U11459 ( .A1(n6199), .A2(keyinput_g56), .B1(keyinput_g5), .B2(
        n10657), .ZN(n10385) );
  OAI221_X1 U11460 ( .B1(n6199), .B2(keyinput_g56), .C1(n10657), .C2(
        keyinput_g5), .A(n10385), .ZN(n10391) );
  INV_X1 U11461 ( .A(SI_16_), .ZN(n10387) );
  AOI22_X1 U11462 ( .A1(n10388), .A2(keyinput_g63), .B1(keyinput_g16), .B2(
        n10387), .ZN(n10386) );
  OAI221_X1 U11463 ( .B1(n10388), .B2(keyinput_g63), .C1(n10387), .C2(
        keyinput_g16), .A(n10386), .ZN(n10390) );
  XOR2_X1 U11464 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_g97), .Z(n10389) );
  OR3_X1 U11465 ( .A1(n10391), .A2(n10390), .A3(n10389), .ZN(n10396) );
  AOI22_X1 U11466 ( .A1(n5252), .A2(keyinput_g107), .B1(n10568), .B2(
        keyinput_g76), .ZN(n10392) );
  OAI221_X1 U11467 ( .B1(n5252), .B2(keyinput_g107), .C1(n10568), .C2(
        keyinput_g76), .A(n10392), .ZN(n10395) );
  XNOR2_X1 U11468 ( .A(n10393), .B(keyinput_g124), .ZN(n10394) );
  NOR3_X1 U11469 ( .A1(n10396), .A2(n10395), .A3(n10394), .ZN(n10433) );
  AOI22_X1 U11470 ( .A1(n10398), .A2(keyinput_g61), .B1(keyinput_g86), .B2(
        n10635), .ZN(n10397) );
  OAI221_X1 U11471 ( .B1(n10398), .B2(keyinput_g61), .C1(n10635), .C2(
        keyinput_g86), .A(n10397), .ZN(n10407) );
  AOI22_X1 U11472 ( .A1(n5269), .A2(keyinput_g120), .B1(n5214), .B2(
        keyinput_g95), .ZN(n10399) );
  OAI221_X1 U11473 ( .B1(n5269), .B2(keyinput_g120), .C1(n5214), .C2(
        keyinput_g95), .A(n10399), .ZN(n10406) );
  INV_X1 U11474 ( .A(SI_7_), .ZN(n10401) );
  AOI22_X1 U11475 ( .A1(n10607), .A2(keyinput_g36), .B1(keyinput_g25), .B2(
        n10401), .ZN(n10400) );
  OAI221_X1 U11476 ( .B1(n10607), .B2(keyinput_g36), .C1(n10401), .C2(
        keyinput_g25), .A(n10400), .ZN(n10405) );
  XNOR2_X1 U11477 ( .A(P2_REG3_REG_22__SCAN_IN), .B(keyinput_g57), .ZN(n10403)
         );
  XNOR2_X1 U11478 ( .A(SI_1_), .B(keyinput_g31), .ZN(n10402) );
  NAND2_X1 U11479 ( .A1(n10403), .A2(n10402), .ZN(n10404) );
  NOR4_X1 U11480 ( .A1(n10407), .A2(n10406), .A3(n10405), .A4(n10404), .ZN(
        n10432) );
  INV_X1 U11481 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n10662) );
  AOI22_X1 U11482 ( .A1(n10662), .A2(keyinput_g38), .B1(keyinput_g89), .B2(
        n10409), .ZN(n10408) );
  OAI221_X1 U11483 ( .B1(n10662), .B2(keyinput_g38), .C1(n10409), .C2(
        keyinput_g89), .A(n10408), .ZN(n10417) );
  AOI22_X1 U11484 ( .A1(n10622), .A2(keyinput_g47), .B1(keyinput_g20), .B2(
        n5175), .ZN(n10410) );
  OAI221_X1 U11485 ( .B1(n10622), .B2(keyinput_g47), .C1(n5175), .C2(
        keyinput_g20), .A(n10410), .ZN(n10416) );
  INV_X1 U11486 ( .A(P2_WR_REG_SCAN_IN), .ZN(n10632) );
  AOI22_X1 U11487 ( .A1(n10632), .A2(keyinput_g0), .B1(n10638), .B2(
        keyinput_g82), .ZN(n10411) );
  OAI221_X1 U11488 ( .B1(n10632), .B2(keyinput_g0), .C1(n10638), .C2(
        keyinput_g82), .A(n10411), .ZN(n10415) );
  AOI22_X1 U11489 ( .A1(n10661), .A2(keyinput_g77), .B1(n10413), .B2(
        keyinput_g51), .ZN(n10412) );
  OAI221_X1 U11490 ( .B1(n10661), .B2(keyinput_g77), .C1(n10413), .C2(
        keyinput_g51), .A(n10412), .ZN(n10414) );
  NOR4_X1 U11491 ( .A1(n10417), .A2(n10416), .A3(n10415), .A4(n10414), .ZN(
        n10431) );
  AOI22_X1 U11492 ( .A1(n10419), .A2(keyinput_g12), .B1(keyinput_g102), .B2(
        n5604), .ZN(n10418) );
  OAI221_X1 U11493 ( .B1(n10419), .B2(keyinput_g12), .C1(n5604), .C2(
        keyinput_g102), .A(n10418), .ZN(n10429) );
  AOI22_X1 U11494 ( .A1(n10421), .A2(keyinput_g27), .B1(n10567), .B2(
        keyinput_g73), .ZN(n10420) );
  OAI221_X1 U11495 ( .B1(n10421), .B2(keyinput_g27), .C1(n10567), .C2(
        keyinput_g73), .A(n10420), .ZN(n10428) );
  AOI22_X1 U11496 ( .A1(n10561), .A2(keyinput_g79), .B1(n10423), .B2(
        keyinput_g14), .ZN(n10422) );
  OAI221_X1 U11497 ( .B1(n10561), .B2(keyinput_g79), .C1(n10423), .C2(
        keyinput_g14), .A(n10422), .ZN(n10427) );
  XNOR2_X1 U11498 ( .A(P2_B_REG_SCAN_IN), .B(keyinput_g64), .ZN(n10425) );
  XNOR2_X1 U11499 ( .A(SI_8_), .B(keyinput_g24), .ZN(n10424) );
  NAND2_X1 U11500 ( .A1(n10425), .A2(n10424), .ZN(n10426) );
  NOR4_X1 U11501 ( .A1(n10429), .A2(n10428), .A3(n10427), .A4(n10426), .ZN(
        n10430) );
  NAND4_X1 U11502 ( .A1(n10433), .A2(n10432), .A3(n10431), .A4(n10430), .ZN(
        n10484) );
  AOI22_X1 U11503 ( .A1(n5250), .A2(keyinput_g106), .B1(n10435), .B2(
        keyinput_g4), .ZN(n10434) );
  OAI221_X1 U11504 ( .B1(n5250), .B2(keyinput_g106), .C1(n10435), .C2(
        keyinput_g4), .A(n10434), .ZN(n10446) );
  AOI22_X1 U11505 ( .A1(n10437), .A2(keyinput_g65), .B1(n10588), .B2(
        keyinput_g72), .ZN(n10436) );
  OAI221_X1 U11506 ( .B1(n10437), .B2(keyinput_g65), .C1(n10588), .C2(
        keyinput_g72), .A(n10436), .ZN(n10445) );
  AOI22_X1 U11507 ( .A1(n10440), .A2(keyinput_g52), .B1(keyinput_g70), .B2(
        n10439), .ZN(n10438) );
  OAI221_X1 U11508 ( .B1(n10440), .B2(keyinput_g52), .C1(n10439), .C2(
        keyinput_g70), .A(n10438), .ZN(n10444) );
  XOR2_X1 U11509 ( .A(n6150), .B(keyinput_g53), .Z(n10442) );
  XNOR2_X1 U11510 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput_g113), .ZN(n10441)
         );
  NAND2_X1 U11511 ( .A1(n10442), .A2(n10441), .ZN(n10443) );
  NOR4_X1 U11512 ( .A1(n10446), .A2(n10445), .A3(n10444), .A4(n10443), .ZN(
        n10482) );
  INV_X1 U11513 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10654) );
  AOI22_X1 U11514 ( .A1(n10448), .A2(keyinput_g62), .B1(keyinput_g48), .B2(
        n10654), .ZN(n10447) );
  OAI221_X1 U11515 ( .B1(n10448), .B2(keyinput_g62), .C1(n10654), .C2(
        keyinput_g48), .A(n10447), .ZN(n10456) );
  XOR2_X1 U11516 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_g93), .Z(n10455) );
  XOR2_X1 U11517 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(keyinput_g66), .Z(n10454)
         );
  XNOR2_X1 U11518 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_g96), .ZN(n10452) );
  XNOR2_X1 U11519 ( .A(SI_2_), .B(keyinput_g30), .ZN(n10451) );
  XNOR2_X1 U11520 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_g117), .ZN(n10450)
         );
  XNOR2_X1 U11521 ( .A(SI_23_), .B(keyinput_g9), .ZN(n10449) );
  NAND4_X1 U11522 ( .A1(n10452), .A2(n10451), .A3(n10450), .A4(n10449), .ZN(
        n10453) );
  NOR4_X1 U11523 ( .A1(n10456), .A2(n10455), .A3(n10454), .A4(n10453), .ZN(
        n10481) );
  INV_X1 U11524 ( .A(SI_14_), .ZN(n10458) );
  AOI22_X1 U11525 ( .A1(n10459), .A2(keyinput_g46), .B1(keyinput_g18), .B2(
        n10458), .ZN(n10457) );
  OAI221_X1 U11526 ( .B1(n10459), .B2(keyinput_g46), .C1(n10458), .C2(
        keyinput_g18), .A(n10457), .ZN(n10469) );
  AOI22_X1 U11527 ( .A1(n10461), .A2(keyinput_g21), .B1(n10606), .B2(
        keyinput_g78), .ZN(n10460) );
  OAI221_X1 U11528 ( .B1(n10461), .B2(keyinput_g21), .C1(n10606), .C2(
        keyinput_g78), .A(n10460), .ZN(n10468) );
  INV_X1 U11529 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10600) );
  AOI22_X1 U11530 ( .A1(n10463), .A2(keyinput_g81), .B1(n10600), .B2(
        keyinput_g37), .ZN(n10462) );
  OAI221_X1 U11531 ( .B1(n10463), .B2(keyinput_g81), .C1(n10600), .C2(
        keyinput_g37), .A(n10462), .ZN(n10467) );
  XOR2_X1 U11532 ( .A(n5535), .B(keyinput_g98), .Z(n10465) );
  XNOR2_X1 U11533 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_g101), .ZN(n10464)
         );
  NAND2_X1 U11534 ( .A1(n10465), .A2(n10464), .ZN(n10466) );
  NOR4_X1 U11535 ( .A1(n10469), .A2(n10468), .A3(n10467), .A4(n10466), .ZN(
        n10480) );
  INV_X1 U11536 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n10593) );
  AOI22_X1 U11537 ( .A1(n5272), .A2(keyinput_g119), .B1(n10593), .B2(
        keyinput_g91), .ZN(n10470) );
  OAI221_X1 U11538 ( .B1(n5272), .B2(keyinput_g119), .C1(n10593), .C2(
        keyinput_g91), .A(n10470), .ZN(n10478) );
  AOI22_X1 U11539 ( .A1(n10565), .A2(keyinput_g41), .B1(keyinput_g8), .B2(
        n10577), .ZN(n10471) );
  OAI221_X1 U11540 ( .B1(n10565), .B2(keyinput_g41), .C1(n10577), .C2(
        keyinput_g8), .A(n10471), .ZN(n10477) );
  XNOR2_X1 U11541 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput_g88), .ZN(n10475)
         );
  XNOR2_X1 U11542 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_g118), .ZN(n10474)
         );
  XNOR2_X1 U11543 ( .A(P2_STATE_REG_SCAN_IN), .B(keyinput_g34), .ZN(n10473) );
  XNOR2_X1 U11544 ( .A(SI_0_), .B(keyinput_g32), .ZN(n10472) );
  NAND4_X1 U11545 ( .A1(n10475), .A2(n10474), .A3(n10473), .A4(n10472), .ZN(
        n10476) );
  NOR3_X1 U11546 ( .A1(n10478), .A2(n10477), .A3(n10476), .ZN(n10479) );
  NAND4_X1 U11547 ( .A1(n10482), .A2(n10481), .A3(n10480), .A4(n10479), .ZN(
        n10483) );
  NOR4_X1 U11548 ( .A1(n10486), .A2(n10485), .A3(n10484), .A4(n10483), .ZN(
        n10682) );
  XOR2_X1 U11549 ( .A(SI_18_), .B(keyinput_f14), .Z(n10493) );
  AOI22_X1 U11550 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(keyinput_f96), .B1(
        P2_REG3_REG_10__SCAN_IN), .B2(keyinput_f39), .ZN(n10487) );
  OAI221_X1 U11551 ( .B1(P1_IR_REG_6__SCAN_IN), .B2(keyinput_f96), .C1(
        P2_REG3_REG_10__SCAN_IN), .C2(keyinput_f39), .A(n10487), .ZN(n10492)
         );
  AOI22_X1 U11552 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(keyinput_f116), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(keyinput_f59), .ZN(n10488) );
  OAI221_X1 U11553 ( .B1(P1_IR_REG_26__SCAN_IN), .B2(keyinput_f116), .C1(
        P2_REG3_REG_2__SCAN_IN), .C2(keyinput_f59), .A(n10488), .ZN(n10491) );
  AOI22_X1 U11554 ( .A1(SI_5_), .A2(keyinput_f27), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(keyinput_f52), .ZN(n10489) );
  OAI221_X1 U11555 ( .B1(SI_5_), .B2(keyinput_f27), .C1(P2_REG3_REG_4__SCAN_IN), .C2(keyinput_f52), .A(n10489), .ZN(n10490) );
  NOR4_X1 U11556 ( .A1(n10493), .A2(n10492), .A3(n10491), .A4(n10490), .ZN(
        n10521) );
  AOI22_X1 U11557 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(keyinput_f65), .B1(
        P2_REG3_REG_9__SCAN_IN), .B2(keyinput_f53), .ZN(n10494) );
  OAI221_X1 U11558 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(keyinput_f65), .C1(
        P2_REG3_REG_9__SCAN_IN), .C2(keyinput_f53), .A(n10494), .ZN(n10501) );
  AOI22_X1 U11559 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(keyinput_f104), .B1(
        P2_REG3_REG_6__SCAN_IN), .B2(keyinput_f61), .ZN(n10495) );
  OAI221_X1 U11560 ( .B1(P1_IR_REG_14__SCAN_IN), .B2(keyinput_f104), .C1(
        P2_REG3_REG_6__SCAN_IN), .C2(keyinput_f61), .A(n10495), .ZN(n10500) );
  AOI22_X1 U11561 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(keyinput_f67), .B1(
        P2_REG3_REG_11__SCAN_IN), .B2(keyinput_f58), .ZN(n10496) );
  OAI221_X1 U11562 ( .B1(P2_DATAO_REG_29__SCAN_IN), .B2(keyinput_f67), .C1(
        P2_REG3_REG_11__SCAN_IN), .C2(keyinput_f58), .A(n10496), .ZN(n10499)
         );
  AOI22_X1 U11563 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(keyinput_f101), .B1(
        P2_STATE_REG_SCAN_IN), .B2(keyinput_f34), .ZN(n10497) );
  OAI221_X1 U11564 ( .B1(P1_IR_REG_11__SCAN_IN), .B2(keyinput_f101), .C1(
        P2_STATE_REG_SCAN_IN), .C2(keyinput_f34), .A(n10497), .ZN(n10498) );
  NOR4_X1 U11565 ( .A1(n10501), .A2(n10500), .A3(n10499), .A4(n10498), .ZN(
        n10520) );
  AOI22_X1 U11566 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_f54), .B1(SI_3_), 
        .B2(keyinput_f29), .ZN(n10502) );
  OAI221_X1 U11567 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_f54), .C1(SI_3_), .C2(keyinput_f29), .A(n10502), .ZN(n10509) );
  AOI22_X1 U11568 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(keyinput_f111), .B1(SI_11_), .B2(keyinput_f21), .ZN(n10503) );
  OAI221_X1 U11569 ( .B1(P1_IR_REG_21__SCAN_IN), .B2(keyinput_f111), .C1(
        SI_11_), .C2(keyinput_f21), .A(n10503), .ZN(n10508) );
  AOI22_X1 U11570 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(keyinput_f108), .B1(
        P2_REG3_REG_26__SCAN_IN), .B2(keyinput_f62), .ZN(n10504) );
  OAI221_X1 U11571 ( .B1(P1_IR_REG_18__SCAN_IN), .B2(keyinput_f108), .C1(
        P2_REG3_REG_26__SCAN_IN), .C2(keyinput_f62), .A(n10504), .ZN(n10507)
         );
  AOI22_X1 U11572 ( .A1(SI_14_), .A2(keyinput_f18), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(keyinput_f70), .ZN(n10505) );
  OAI221_X1 U11573 ( .B1(SI_14_), .B2(keyinput_f18), .C1(
        P2_DATAO_REG_26__SCAN_IN), .C2(keyinput_f70), .A(n10505), .ZN(n10506)
         );
  NOR4_X1 U11574 ( .A1(n10509), .A2(n10508), .A3(n10507), .A4(n10506), .ZN(
        n10519) );
  AOI22_X1 U11575 ( .A1(SI_0_), .A2(keyinput_f32), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(keyinput_f71), .ZN(n10510) );
  OAI221_X1 U11576 ( .B1(SI_0_), .B2(keyinput_f32), .C1(
        P2_DATAO_REG_25__SCAN_IN), .C2(keyinput_f71), .A(n10510), .ZN(n10517)
         );
  AOI22_X1 U11577 ( .A1(SI_22_), .A2(keyinput_f10), .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_f43), .ZN(n10511) );
  OAI221_X1 U11578 ( .B1(SI_22_), .B2(keyinput_f10), .C1(
        P2_REG3_REG_8__SCAN_IN), .C2(keyinput_f43), .A(n10511), .ZN(n10516) );
  AOI22_X1 U11579 ( .A1(P1_D_REG_0__SCAN_IN), .A2(keyinput_f122), .B1(SI_17_), 
        .B2(keyinput_f15), .ZN(n10512) );
  OAI221_X1 U11580 ( .B1(P1_D_REG_0__SCAN_IN), .B2(keyinput_f122), .C1(SI_17_), 
        .C2(keyinput_f15), .A(n10512), .ZN(n10515) );
  AOI22_X1 U11581 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(keyinput_f109), .B1(
        P2_B_REG_SCAN_IN), .B2(keyinput_f64), .ZN(n10513) );
  OAI221_X1 U11582 ( .B1(P1_IR_REG_19__SCAN_IN), .B2(keyinput_f109), .C1(
        P2_B_REG_SCAN_IN), .C2(keyinput_f64), .A(n10513), .ZN(n10514) );
  NOR4_X1 U11583 ( .A1(n10517), .A2(n10516), .A3(n10515), .A4(n10514), .ZN(
        n10518) );
  NAND4_X1 U11584 ( .A1(n10521), .A2(n10520), .A3(n10519), .A4(n10518), .ZN(
        n10676) );
  AOI22_X1 U11585 ( .A1(SI_13_), .A2(keyinput_f19), .B1(P2_RD_REG_SCAN_IN), 
        .B2(keyinput_f33), .ZN(n10522) );
  OAI221_X1 U11586 ( .B1(SI_13_), .B2(keyinput_f19), .C1(P2_RD_REG_SCAN_IN), 
        .C2(keyinput_f33), .A(n10522), .ZN(n10529) );
  AOI22_X1 U11587 ( .A1(SI_25_), .A2(keyinput_f7), .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput_f56), .ZN(n10523) );
  OAI221_X1 U11588 ( .B1(SI_25_), .B2(keyinput_f7), .C1(
        P2_REG3_REG_13__SCAN_IN), .C2(keyinput_f56), .A(n10523), .ZN(n10528)
         );
  AOI22_X1 U11589 ( .A1(SI_2_), .A2(keyinput_f30), .B1(P2_DATAO_REG_7__SCAN_IN), .B2(keyinput_f89), .ZN(n10524) );
  OAI221_X1 U11590 ( .B1(SI_2_), .B2(keyinput_f30), .C1(
        P2_DATAO_REG_7__SCAN_IN), .C2(keyinput_f89), .A(n10524), .ZN(n10527)
         );
  AOI22_X1 U11591 ( .A1(SI_23_), .A2(keyinput_f9), .B1(P2_REG3_REG_7__SCAN_IN), 
        .B2(keyinput_f35), .ZN(n10525) );
  OAI221_X1 U11592 ( .B1(SI_23_), .B2(keyinput_f9), .C1(P2_REG3_REG_7__SCAN_IN), .C2(keyinput_f35), .A(n10525), .ZN(n10526) );
  NOR4_X1 U11593 ( .A1(n10529), .A2(n10528), .A3(n10527), .A4(n10526), .ZN(
        n10559) );
  AOI22_X1 U11594 ( .A1(P1_D_REG_2__SCAN_IN), .A2(keyinput_f124), .B1(
        P2_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .ZN(n10530) );
  OAI221_X1 U11595 ( .B1(P1_D_REG_2__SCAN_IN), .B2(keyinput_f124), .C1(
        P2_REG3_REG_24__SCAN_IN), .C2(keyinput_f51), .A(n10530), .ZN(n10538)
         );
  AOI22_X1 U11596 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(keyinput_f114), .B1(SI_16_), .B2(keyinput_f16), .ZN(n10531) );
  OAI221_X1 U11597 ( .B1(P1_IR_REG_24__SCAN_IN), .B2(keyinput_f114), .C1(
        SI_16_), .C2(keyinput_f16), .A(n10531), .ZN(n10537) );
  AOI22_X1 U11598 ( .A1(SI_31_), .A2(keyinput_f1), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(keyinput_f81), .ZN(n10532) );
  OAI221_X1 U11599 ( .B1(SI_31_), .B2(keyinput_f1), .C1(
        P2_DATAO_REG_15__SCAN_IN), .C2(keyinput_f81), .A(n10532), .ZN(n10536)
         );
  AOI22_X1 U11600 ( .A1(n10534), .A2(keyinput_f90), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(keyinput_f75), .ZN(n10533) );
  OAI221_X1 U11601 ( .B1(n10534), .B2(keyinput_f90), .C1(
        P2_DATAO_REG_21__SCAN_IN), .C2(keyinput_f75), .A(n10533), .ZN(n10535)
         );
  NOR4_X1 U11602 ( .A1(n10538), .A2(n10537), .A3(n10536), .A4(n10535), .ZN(
        n10558) );
  AOI22_X1 U11603 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(keyinput_f120), .B1(SI_6_), 
        .B2(keyinput_f26), .ZN(n10539) );
  OAI221_X1 U11604 ( .B1(P1_IR_REG_30__SCAN_IN), .B2(keyinput_f120), .C1(SI_6_), .C2(keyinput_f26), .A(n10539), .ZN(n10546) );
  AOI22_X1 U11605 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(keyinput_f103), .B1(SI_12_), .B2(keyinput_f20), .ZN(n10540) );
  OAI221_X1 U11606 ( .B1(P1_IR_REG_13__SCAN_IN), .B2(keyinput_f103), .C1(
        SI_12_), .C2(keyinput_f20), .A(n10540), .ZN(n10545) );
  AOI22_X1 U11607 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(keyinput_f110), .B1(
        P2_REG3_REG_21__SCAN_IN), .B2(keyinput_f45), .ZN(n10541) );
  OAI221_X1 U11608 ( .B1(P1_IR_REG_20__SCAN_IN), .B2(keyinput_f110), .C1(
        P2_REG3_REG_21__SCAN_IN), .C2(keyinput_f45), .A(n10541), .ZN(n10544)
         );
  AOI22_X1 U11609 ( .A1(P1_D_REG_1__SCAN_IN), .A2(keyinput_f123), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(keyinput_f83), .ZN(n10542) );
  OAI221_X1 U11610 ( .B1(P1_D_REG_1__SCAN_IN), .B2(keyinput_f123), .C1(
        P2_DATAO_REG_13__SCAN_IN), .C2(keyinput_f83), .A(n10542), .ZN(n10543)
         );
  NOR4_X1 U11611 ( .A1(n10546), .A2(n10545), .A3(n10544), .A4(n10543), .ZN(
        n10557) );
  AOI22_X1 U11612 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(keyinput_f95), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(keyinput_f74), .ZN(n10547) );
  OAI221_X1 U11613 ( .B1(P1_IR_REG_5__SCAN_IN), .B2(keyinput_f95), .C1(
        P2_DATAO_REG_22__SCAN_IN), .C2(keyinput_f74), .A(n10547), .ZN(n10555)
         );
  AOI22_X1 U11614 ( .A1(SI_9_), .A2(keyinput_f23), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(keyinput_f85), .ZN(n10548) );
  OAI221_X1 U11615 ( .B1(SI_9_), .B2(keyinput_f23), .C1(
        P2_DATAO_REG_11__SCAN_IN), .C2(keyinput_f85), .A(n10548), .ZN(n10554)
         );
  AOI22_X1 U11616 ( .A1(SI_19_), .A2(keyinput_f13), .B1(SI_29_), .B2(
        keyinput_f3), .ZN(n10549) );
  OAI221_X1 U11617 ( .B1(SI_19_), .B2(keyinput_f13), .C1(SI_29_), .C2(
        keyinput_f3), .A(n10549), .ZN(n10553) );
  AOI22_X1 U11618 ( .A1(SI_20_), .A2(keyinput_f12), .B1(n10551), .B2(
        keyinput_f66), .ZN(n10550) );
  OAI221_X1 U11619 ( .B1(SI_20_), .B2(keyinput_f12), .C1(n10551), .C2(
        keyinput_f66), .A(n10550), .ZN(n10552) );
  NOR4_X1 U11620 ( .A1(n10555), .A2(n10554), .A3(n10553), .A4(n10552), .ZN(
        n10556) );
  NAND4_X1 U11621 ( .A1(n10559), .A2(n10558), .A3(n10557), .A4(n10556), .ZN(
        n10675) );
  AOI22_X1 U11622 ( .A1(n10562), .A2(keyinput_f126), .B1(n10561), .B2(
        keyinput_f79), .ZN(n10560) );
  OAI221_X1 U11623 ( .B1(n10562), .B2(keyinput_f126), .C1(n10561), .C2(
        keyinput_f79), .A(n10560), .ZN(n10573) );
  AOI22_X1 U11624 ( .A1(n10565), .A2(keyinput_f41), .B1(keyinput_f17), .B2(
        n10564), .ZN(n10563) );
  OAI221_X1 U11625 ( .B1(n10565), .B2(keyinput_f41), .C1(n10564), .C2(
        keyinput_f17), .A(n10563), .ZN(n10572) );
  AOI22_X1 U11626 ( .A1(n10568), .A2(keyinput_f76), .B1(n10567), .B2(
        keyinput_f73), .ZN(n10566) );
  OAI221_X1 U11627 ( .B1(n10568), .B2(keyinput_f76), .C1(n10567), .C2(
        keyinput_f73), .A(n10566), .ZN(n10571) );
  AOI22_X1 U11628 ( .A1(n5252), .A2(keyinput_f107), .B1(n5534), .B2(
        keyinput_f99), .ZN(n10569) );
  OAI221_X1 U11629 ( .B1(n5252), .B2(keyinput_f107), .C1(n5534), .C2(
        keyinput_f99), .A(n10569), .ZN(n10570) );
  NOR4_X1 U11630 ( .A1(n10573), .A2(n10572), .A3(n10571), .A4(n10570), .ZN(
        n10615) );
  AOI22_X1 U11631 ( .A1(n5272), .A2(keyinput_f119), .B1(n10575), .B2(
        keyinput_f125), .ZN(n10574) );
  OAI221_X1 U11632 ( .B1(n5272), .B2(keyinput_f119), .C1(n10575), .C2(
        keyinput_f125), .A(n10574), .ZN(n10585) );
  AOI22_X1 U11633 ( .A1(n10578), .A2(keyinput_f6), .B1(keyinput_f8), .B2(
        n10577), .ZN(n10576) );
  OAI221_X1 U11634 ( .B1(n10578), .B2(keyinput_f6), .C1(n10577), .C2(
        keyinput_f8), .A(n10576), .ZN(n10584) );
  XNOR2_X1 U11635 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput_f87), .ZN(n10582)
         );
  XNOR2_X1 U11636 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_f118), .ZN(n10581)
         );
  XNOR2_X1 U11637 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_f117), .ZN(n10580)
         );
  XNOR2_X1 U11638 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput_f46), .ZN(n10579)
         );
  NAND4_X1 U11639 ( .A1(n10582), .A2(n10581), .A3(n10580), .A4(n10579), .ZN(
        n10583) );
  NOR3_X1 U11640 ( .A1(n10585), .A2(n10584), .A3(n10583), .ZN(n10614) );
  AOI22_X1 U11641 ( .A1(n10588), .A2(keyinput_f72), .B1(keyinput_f28), .B2(
        n10587), .ZN(n10586) );
  OAI221_X1 U11642 ( .B1(n10588), .B2(keyinput_f72), .C1(n10587), .C2(
        keyinput_f28), .A(n10586), .ZN(n10597) );
  XOR2_X1 U11643 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_f100), .Z(n10596) );
  XNOR2_X1 U11644 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(keyinput_f80), .ZN(n10592) );
  XNOR2_X1 U11645 ( .A(SI_1_), .B(keyinput_f31), .ZN(n10591) );
  XNOR2_X1 U11646 ( .A(SI_7_), .B(keyinput_f25), .ZN(n10590) );
  XNOR2_X1 U11647 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput_f113), .ZN(n10589)
         );
  NAND4_X1 U11648 ( .A1(n10592), .A2(n10591), .A3(n10590), .A4(n10589), .ZN(
        n10595) );
  XNOR2_X1 U11649 ( .A(keyinput_f91), .B(n10593), .ZN(n10594) );
  NOR4_X1 U11650 ( .A1(n10597), .A2(n10596), .A3(n10595), .A4(n10594), .ZN(
        n10613) );
  INV_X1 U11651 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n10599) );
  AOI22_X1 U11652 ( .A1(n10600), .A2(keyinput_f37), .B1(n10599), .B2(
        keyinput_f42), .ZN(n10598) );
  OAI221_X1 U11653 ( .B1(n10600), .B2(keyinput_f37), .C1(n10599), .C2(
        keyinput_f42), .A(n10598), .ZN(n10611) );
  AOI22_X1 U11654 ( .A1(n10602), .A2(keyinput_f11), .B1(n5912), .B2(
        keyinput_f68), .ZN(n10601) );
  OAI221_X1 U11655 ( .B1(n10602), .B2(keyinput_f11), .C1(n5912), .C2(
        keyinput_f68), .A(n10601), .ZN(n10610) );
  AOI22_X1 U11656 ( .A1(n10604), .A2(keyinput_f127), .B1(n7319), .B2(
        keyinput_f44), .ZN(n10603) );
  OAI221_X1 U11657 ( .B1(n10604), .B2(keyinput_f127), .C1(n7319), .C2(
        keyinput_f44), .A(n10603), .ZN(n10609) );
  AOI22_X1 U11658 ( .A1(n10607), .A2(keyinput_f36), .B1(keyinput_f78), .B2(
        n10606), .ZN(n10605) );
  OAI221_X1 U11659 ( .B1(n10607), .B2(keyinput_f36), .C1(n10606), .C2(
        keyinput_f78), .A(n10605), .ZN(n10608) );
  NOR4_X1 U11660 ( .A1(n10611), .A2(n10610), .A3(n10609), .A4(n10608), .ZN(
        n10612) );
  NAND4_X1 U11661 ( .A1(n10615), .A2(n10614), .A3(n10613), .A4(n10612), .ZN(
        n10674) );
  AOI22_X1 U11662 ( .A1(n5604), .A2(keyinput_f102), .B1(n10617), .B2(
        keyinput_f24), .ZN(n10616) );
  OAI221_X1 U11663 ( .B1(n5604), .B2(keyinput_f102), .C1(n10617), .C2(
        keyinput_f24), .A(n10616), .ZN(n10628) );
  AOI22_X1 U11664 ( .A1(n5224), .A2(keyinput_f115), .B1(n10619), .B2(
        keyinput_f22), .ZN(n10618) );
  OAI221_X1 U11665 ( .B1(n5224), .B2(keyinput_f115), .C1(n10619), .C2(
        keyinput_f22), .A(n10618), .ZN(n10627) );
  INV_X1 U11666 ( .A(SI_30_), .ZN(n10621) );
  AOI22_X1 U11667 ( .A1(n10622), .A2(keyinput_f47), .B1(keyinput_f2), .B2(
        n10621), .ZN(n10620) );
  OAI221_X1 U11668 ( .B1(n10622), .B2(keyinput_f47), .C1(n10621), .C2(
        keyinput_f2), .A(n10620), .ZN(n10626) );
  XNOR2_X1 U11669 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_f121), .ZN(n10624)
         );
  XNOR2_X1 U11670 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_f105), .ZN(n10623)
         );
  NAND2_X1 U11671 ( .A1(n10624), .A2(n10623), .ZN(n10625) );
  NOR4_X1 U11672 ( .A1(n10628), .A2(n10627), .A3(n10626), .A4(n10625), .ZN(
        n10672) );
  INV_X1 U11673 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10630) );
  AOI22_X1 U11674 ( .A1(n10630), .A2(keyinput_f57), .B1(keyinput_f106), .B2(
        n5250), .ZN(n10629) );
  OAI221_X1 U11675 ( .B1(n10630), .B2(keyinput_f57), .C1(n5250), .C2(
        keyinput_f106), .A(n10629), .ZN(n10642) );
  AOI22_X1 U11676 ( .A1(n10632), .A2(keyinput_f0), .B1(n5535), .B2(
        keyinput_f98), .ZN(n10631) );
  OAI221_X1 U11677 ( .B1(n10632), .B2(keyinput_f0), .C1(n5535), .C2(
        keyinput_f98), .A(n10631), .ZN(n10641) );
  AOI22_X1 U11678 ( .A1(n10635), .A2(keyinput_f86), .B1(n10634), .B2(
        keyinput_f40), .ZN(n10633) );
  OAI221_X1 U11679 ( .B1(n10635), .B2(keyinput_f86), .C1(n10634), .C2(
        keyinput_f40), .A(n10633), .ZN(n10640) );
  INV_X1 U11680 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10637) );
  AOI22_X1 U11681 ( .A1(n10638), .A2(keyinput_f82), .B1(n10637), .B2(
        keyinput_f60), .ZN(n10636) );
  OAI221_X1 U11682 ( .B1(n10638), .B2(keyinput_f82), .C1(n10637), .C2(
        keyinput_f60), .A(n10636), .ZN(n10639) );
  NOR4_X1 U11683 ( .A1(n10642), .A2(n10641), .A3(n10640), .A4(n10639), .ZN(
        n10671) );
  AOI22_X1 U11684 ( .A1(n5402), .A2(keyinput_f94), .B1(n6086), .B2(
        keyinput_f49), .ZN(n10643) );
  OAI221_X1 U11685 ( .B1(n5402), .B2(keyinput_f94), .C1(n6086), .C2(
        keyinput_f49), .A(n10643), .ZN(n10652) );
  AOI22_X1 U11686 ( .A1(n5880), .A2(keyinput_f69), .B1(keyinput_f84), .B2(
        n10645), .ZN(n10644) );
  OAI221_X1 U11687 ( .B1(n5880), .B2(keyinput_f69), .C1(n10645), .C2(
        keyinput_f84), .A(n10644), .ZN(n10651) );
  XNOR2_X1 U11688 ( .A(SI_28_), .B(keyinput_f4), .ZN(n10649) );
  XNOR2_X1 U11689 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_f97), .ZN(n10648) );
  XNOR2_X1 U11690 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_f112), .ZN(n10647)
         );
  XNOR2_X1 U11691 ( .A(P2_REG3_REG_15__SCAN_IN), .B(keyinput_f63), .ZN(n10646)
         );
  NAND4_X1 U11692 ( .A1(n10649), .A2(n10648), .A3(n10647), .A4(n10646), .ZN(
        n10650) );
  NOR3_X1 U11693 ( .A1(n10652), .A2(n10651), .A3(n10650), .ZN(n10670) );
  AOI22_X1 U11694 ( .A1(n10655), .A2(keyinput_f88), .B1(n10654), .B2(
        keyinput_f48), .ZN(n10653) );
  OAI221_X1 U11695 ( .B1(n10655), .B2(keyinput_f88), .C1(n10654), .C2(
        keyinput_f48), .A(n10653), .ZN(n10668) );
  AOI22_X1 U11696 ( .A1(n10658), .A2(keyinput_f55), .B1(keyinput_f5), .B2(
        n10657), .ZN(n10656) );
  OAI221_X1 U11697 ( .B1(n10658), .B2(keyinput_f55), .C1(n10657), .C2(
        keyinput_f5), .A(n10656), .ZN(n10667) );
  AOI22_X1 U11698 ( .A1(n10661), .A2(keyinput_f77), .B1(n10660), .B2(
        keyinput_f50), .ZN(n10659) );
  OAI221_X1 U11699 ( .B1(n10661), .B2(keyinput_f77), .C1(n10660), .C2(
        keyinput_f50), .A(n10659), .ZN(n10666) );
  XOR2_X1 U11700 ( .A(n10662), .B(keyinput_f38), .Z(n10664) );
  XNOR2_X1 U11701 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_f93), .ZN(n10663) );
  NAND2_X1 U11702 ( .A1(n10664), .A2(n10663), .ZN(n10665) );
  NOR4_X1 U11703 ( .A1(n10668), .A2(n10667), .A3(n10666), .A4(n10665), .ZN(
        n10669) );
  NAND4_X1 U11704 ( .A1(n10672), .A2(n10671), .A3(n10670), .A4(n10669), .ZN(
        n10673) );
  OR4_X1 U11705 ( .A1(n10676), .A2(n10675), .A3(n10674), .A4(n10673), .ZN(
        n10678) );
  AOI21_X1 U11706 ( .B1(keyinput_f92), .B2(n10678), .A(keyinput_g92), .ZN(
        n10680) );
  INV_X1 U11707 ( .A(keyinput_f92), .ZN(n10677) );
  AOI21_X1 U11708 ( .B1(n10678), .B2(n10677), .A(n5340), .ZN(n10679) );
  AOI22_X1 U11709 ( .A1(n5340), .A2(n10680), .B1(keyinput_g92), .B2(n10679), 
        .ZN(n10681) );
  AOI21_X1 U11710 ( .B1(n10683), .B2(n10682), .A(n10681), .ZN(n10684) );
  XNOR2_X1 U11711 ( .A(n10685), .B(n10684), .ZN(n10686) );
  XNOR2_X1 U11712 ( .A(n10687), .B(n10686), .ZN(ADD_1068_U4) );
  XNOR2_X1 U11713 ( .A(n10689), .B(n10688), .ZN(ADD_1068_U47) );
  XOR2_X1 U11714 ( .A(n10691), .B(n10690), .Z(ADD_1068_U54) );
  XNOR2_X1 U11715 ( .A(n10693), .B(n10692), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11716 ( .A(n10695), .B(n10694), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11717 ( .A(n10697), .B(n10696), .ZN(ADD_1068_U48) );
  XNOR2_X1 U11718 ( .A(n10699), .B(n10698), .ZN(ADD_1068_U50) );
  XOR2_X1 U11719 ( .A(n10701), .B(n10700), .Z(ADD_1068_U53) );
  XNOR2_X1 U11720 ( .A(n10703), .B(n10702), .ZN(ADD_1068_U52) );
  BUF_X4 U5027 ( .A(n6445), .Z(n8555) );
  CLKBUF_X1 U5037 ( .A(n5380), .Z(n5792) );
  CLKBUF_X2 U5044 ( .A(n6022), .Z(n4505) );
endmodule

