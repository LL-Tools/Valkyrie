

module b22_C_gen_AntiSAT_k_128_9 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, 
        SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, 
        SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, 
        SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, 
        SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, 
        P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, 
        P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, 
        P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, 
        P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, 
        P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, 
        P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, 
        P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, 
        P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, 
        P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, 
        P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, 
        P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, 
        P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, 
        P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, 
        P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, 
        P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, 
        P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, 
        P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, 
        P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, 
        P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, 
        P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, 
        P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, 
        P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, 
        P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, 
        P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, 
        P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, 
        P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, 
        P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, 
        P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, 
        P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, 
        P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, 
        P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, 
        P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, 
        P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, 
        P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, 
        P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, 
        P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, 
        P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, 
        P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, 
        P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, 
        P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, 
        P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, 
        P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, 
        P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, 
        P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, 
        P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, 
        P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, 
        P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, 
        P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0,
         keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5,
         keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10,
         keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15,
         keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20,
         keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25,
         keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30,
         keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35,
         keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40,
         keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45,
         keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50,
         keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55,
         keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60,
         keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1,
         keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6,
         keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11,
         keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16,
         keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21,
         keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26,
         keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31,
         keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36,
         keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41,
         keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46,
         keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51,
         keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56,
         keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61,
         keyinput_g62, keyinput_g63;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6467, n6468, n6469, n6470, n6471, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148;

  INV_X4 U7215 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  AND2_X1 U7216 ( .A1(n12262), .A2(n12133), .ZN(n13680) );
  NAND2_X2 U7217 ( .A1(n9009), .A2(n9008), .ZN(n14212) );
  NOR2_X1 U7218 ( .A1(n14602), .A2(n14601), .ZN(n14600) );
  INV_X2 U7219 ( .A(n12027), .ZN(n12265) );
  NAND2_X1 U7220 ( .A1(n8293), .A2(n8292), .ZN(n14789) );
  INV_X1 U7222 ( .A(n8759), .ZN(n8958) );
  XNOR2_X1 U7223 ( .A(n8956), .B(P1_IR_REG_19__SCAN_IN), .ZN(n9168) );
  CLKBUF_X1 U7224 ( .A(n8685), .Z(n10447) );
  CLKBUF_X2 U7225 ( .A(n7523), .Z(n10346) );
  NAND2_X1 U7226 ( .A1(n8603), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8605) );
  AND3_X1 U7227 ( .A1(n6729), .A2(n6731), .A3(n8703), .ZN(n6707) );
  NAND3_X1 U7228 ( .A1(n8134), .A2(n8214), .A3(n8133), .ZN(n8381) );
  CLKBUF_X1 U7229 ( .A(n14980), .Z(n6467) );
  NOR2_X1 U7230 ( .A1(n10355), .A2(n12820), .ZN(n14980) );
  CLKBUF_X1 U7231 ( .A(n13683), .Z(n6468) );
  OAI21_X1 U7232 ( .B1(n10113), .B2(n10713), .A(n14477), .ZN(n13683) );
  CLKBUF_X1 U7233 ( .A(n11711), .Z(n6469) );
  NAND2_X2 U7234 ( .A1(n7123), .A2(n7122), .ZN(n11324) );
  AOI21_X1 U7235 ( .B1(n6784), .B2(n14725), .A(n8614), .ZN(n13484) );
  INV_X1 U7236 ( .A(n9496), .ZN(n9567) );
  AND2_X1 U7237 ( .A1(n8682), .A2(n8681), .ZN(n8685) );
  INV_X1 U7238 ( .A(n12282), .ZN(n12090) );
  NAND2_X1 U7239 ( .A1(n12371), .A2(n12377), .ZN(n12507) );
  AND3_X1 U7240 ( .A1(n7555), .A2(n7554), .A3(n7553), .ZN(n10493) );
  AND2_X1 U7241 ( .A1(n7968), .A2(n6565), .ZN(n7473) );
  INV_X1 U7242 ( .A(n9457), .ZN(n8233) );
  NAND2_X1 U7243 ( .A1(n14700), .A2(n8331), .ZN(n7123) );
  INV_X1 U7244 ( .A(n12284), .ZN(n12125) );
  NAND2_X1 U7245 ( .A1(n6474), .A2(n14244), .ZN(n9109) );
  INV_X1 U7246 ( .A(n7542), .ZN(n9435) );
  NOR2_X1 U7247 ( .A1(n11605), .A2(n7381), .ZN(n11606) );
  INV_X1 U7248 ( .A(n12820), .ZN(n12776) );
  INV_X1 U7249 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n7460) );
  OR2_X1 U7250 ( .A1(n7715), .A2(n7912), .ZN(n7918) );
  INV_X1 U7251 ( .A(n8739), .ZN(n8957) );
  INV_X2 U7252 ( .A(n8991), .ZN(n9334) );
  OAI21_X1 U7253 ( .B1(n8739), .B2(n14256), .A(n8751), .ZN(n11188) );
  AND2_X2 U7254 ( .A1(n6707), .A2(n6730), .ZN(n9070) );
  AOI21_X1 U7255 ( .B1(P3_ADDR_REG_6__SCAN_IN), .B2(n9695), .A(n9694), .ZN(
        n9696) );
  MUX2_X1 U7256 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7962), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n7965) );
  INV_X1 U7257 ( .A(n8043), .ZN(n8050) );
  INV_X1 U7258 ( .A(n13382), .ZN(n13502) );
  NAND2_X1 U7259 ( .A1(n9018), .A2(n9017), .ZN(n14208) );
  INV_X1 U7260 ( .A(n15018), .ZN(n12698) );
  INV_X1 U7261 ( .A(n12820), .ZN(n6473) );
  AND2_X1 U7262 ( .A1(n8863), .A2(n8862), .ZN(n13652) );
  NAND2_X1 U7263 ( .A1(n14254), .A2(n8739), .ZN(n14218) );
  XOR2_X1 U7265 ( .A(n8683), .B(n9660), .Z(n6470) );
  XNOR2_X1 U7266 ( .A(n8720), .B(n8719), .ZN(n9114) );
  NOR2_X2 U7267 ( .A1(n14309), .A2(n14308), .ZN(n14307) );
  OAI21_X2 U7268 ( .B1(n7884), .B2(n6509), .A(n7886), .ZN(n7899) );
  XNOR2_X2 U7269 ( .A(n9746), .B(n6876), .ZN(n14274) );
  AOI21_X2 U7270 ( .B1(n12576), .B2(n7018), .A(n7014), .ZN(n7013) );
  AND2_X2 U7271 ( .A1(n6574), .A2(n7094), .ZN(n13333) );
  OAI21_X2 U7272 ( .B1(n10347), .B2(n10356), .A(n11666), .ZN(n11667) );
  OR2_X2 U7273 ( .A1(n13124), .A2(n12534), .ZN(n9960) );
  XNOR2_X2 U7274 ( .A(n12188), .B(n12186), .ZN(n13152) );
  INV_X2 U7275 ( .A(n7935), .ZN(n15044) );
  NAND2_X2 U7276 ( .A1(n15135), .A2(n9743), .ZN(n9746) );
  INV_X1 U7277 ( .A(n12314), .ZN(n6471) );
  AND2_X2 U7278 ( .A1(n12352), .A2(n12350), .ZN(n12509) );
  OAI21_X2 U7279 ( .B1(n11541), .B2(n11540), .A(n11539), .ZN(n11599) );
  OAI21_X2 U7280 ( .B1(n11599), .B2(n7041), .A(n7039), .ZN(n11837) );
  NOR2_X2 U7281 ( .A1(n9688), .A2(n9689), .ZN(n9690) );
  NOR2_X2 U7282 ( .A1(n14451), .A2(n14450), .ZN(n14449) );
  NAND2_X2 U7283 ( .A1(n14445), .A2(n6872), .ZN(n14450) );
  OAI21_X2 U7284 ( .B1(n9732), .B2(n9733), .A(n6888), .ZN(n9681) );
  XNOR2_X2 U7285 ( .A(n6753), .B(P1_ADDR_REG_1__SCAN_IN), .ZN(n9732) );
  XNOR2_X2 U7286 ( .A(n6995), .B(n10981), .ZN(n10971) );
  NAND3_X2 U7287 ( .A1(n6994), .A2(n8204), .A3(n8202), .ZN(n6995) );
  NAND4_X4 U7288 ( .A1(n8194), .A2(n8193), .A3(n8192), .A4(n8191), .ZN(n13308)
         );
  INV_X2 U7289 ( .A(n12092), .ZN(n12285) );
  INV_X4 U7290 ( .A(n11076), .ZN(n12092) );
  OAI22_X2 U7291 ( .A1(n8223), .A2(n8224), .B1(n10128), .B2(n8053), .ZN(n8242)
         );
  XNOR2_X2 U7292 ( .A(n9758), .B(n9757), .ZN(n14280) );
  NAND2_X2 U7293 ( .A1(n14276), .A2(n9756), .ZN(n9758) );
  XNOR2_X2 U7294 ( .A(n7461), .B(n7469), .ZN(n7930) );
  XNOR2_X2 U7295 ( .A(n8605), .B(n8604), .ZN(n8681) );
  XNOR2_X1 U7296 ( .A(n11606), .B(n11668), .ZN(n14855) );
  INV_X2 U7298 ( .A(n7931), .ZN(n12820) );
  NAND2_X1 U7299 ( .A1(n13520), .A2(n8675), .ZN(n13402) );
  NAND2_X1 U7300 ( .A1(n12671), .A2(n6535), .ZN(n12614) );
  OAI21_X1 U7301 ( .B1(n11124), .B2(n8653), .A(n8654), .ZN(n10827) );
  NAND2_X1 U7302 ( .A1(n15024), .A2(n12361), .ZN(n15011) );
  NAND2_X1 U7303 ( .A1(n10970), .A2(n10971), .ZN(n10863) );
  AND2_X1 U7304 ( .A1(n10718), .A2(n12066), .ZN(n7389) );
  INV_X1 U7305 ( .A(n14766), .ZN(n10869) );
  INV_X1 U7306 ( .A(n13770), .ZN(n11078) );
  INV_X2 U7307 ( .A(n12092), .ZN(n12275) );
  AND2_X1 U7308 ( .A1(n10077), .A2(n10075), .ZN(n11076) );
  INV_X1 U7309 ( .A(n14721), .ZN(n14746) );
  NAND2_X1 U7310 ( .A1(n14745), .A2(n8681), .ZN(n12193) );
  CLKBUF_X2 U7311 ( .A(n8768), .Z(n9107) );
  INV_X4 U7312 ( .A(n10196), .ZN(n8477) );
  NOR2_X1 U7313 ( .A1(n9666), .A2(n11533), .ZN(n14745) );
  CLKBUF_X2 U7314 ( .A(n7550), .Z(n9431) );
  CLKBUF_X2 U7315 ( .A(n7529), .Z(n7926) );
  AND2_X1 U7316 ( .A1(n8717), .A2(n14244), .ZN(n8767) );
  NAND2_X4 U7317 ( .A1(n7930), .A2(n7931), .ZN(n10341) );
  INV_X1 U7318 ( .A(n8712), .ZN(n6474) );
  INV_X1 U7319 ( .A(n8158), .ZN(n13579) );
  BUF_X1 U7321 ( .A(n14272), .Z(n6476) );
  INV_X4 U7322 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  AOI21_X1 U7323 ( .B1(n9642), .B2(n9641), .A(n9640), .ZN(n9673) );
  MUX2_X1 U7324 ( .A(n13078), .B(n13077), .S(n15120), .Z(n13079) );
  OAI211_X1 U7325 ( .C1(n13480), .C2(n14817), .A(n13483), .B(n13484), .ZN(
        n13563) );
  NOR2_X1 U7326 ( .A1(n8694), .A2(n8693), .ZN(n8695) );
  NAND2_X1 U7327 ( .A1(n12203), .A2(n12202), .ZN(n13251) );
  MUX2_X1 U7328 ( .A(n14194), .B(n14193), .S(n14549), .Z(n14195) );
  AND2_X1 U7329 ( .A1(n7049), .A2(n12260), .ZN(n13722) );
  MUX2_X1 U7330 ( .A(n14096), .B(n14193), .S(n14560), .Z(n14097) );
  AOI211_X1 U7331 ( .C1(n14212), .C2(n6468), .A(n13682), .B(n13681), .ZN(
        n13684) );
  INV_X1 U7332 ( .A(n6997), .ZN(n13369) );
  AOI21_X2 U7333 ( .B1(n13389), .B2(n13398), .A(n6648), .ZN(n13375) );
  NAND2_X1 U7334 ( .A1(n6999), .A2(n6998), .ZN(n6997) );
  AOI21_X1 U7335 ( .B1(n13152), .B2(n13153), .A(n12189), .ZN(n13217) );
  CLKBUF_X1 U7336 ( .A(n13612), .Z(n13705) );
  NAND2_X1 U7337 ( .A1(n7862), .A2(n7861), .ZN(n12592) );
  NAND2_X1 U7338 ( .A1(n9049), .A2(n9048), .ZN(n13926) );
  NAND2_X1 U7339 ( .A1(n14285), .A2(n6746), .ZN(n14260) );
  XNOR2_X1 U7340 ( .A(n13502), .B(n13255), .ZN(n13374) );
  NAND2_X1 U7341 ( .A1(n6986), .A2(n6985), .ZN(n7397) );
  NOR2_X1 U7342 ( .A1(n13265), .A2(n13268), .ZN(n13266) );
  XNOR2_X1 U7343 ( .A(n8534), .B(n6806), .ZN(n11939) );
  NAND2_X1 U7344 ( .A1(n12614), .A2(n10001), .ZN(n12617) );
  XNOR2_X1 U7345 ( .A(n6631), .B(n8482), .ZN(n12251) );
  NAND2_X1 U7346 ( .A1(n11512), .A2(n11511), .ZN(n11722) );
  NAND2_X1 U7347 ( .A1(n13316), .A2(n12248), .ZN(n6631) );
  XNOR2_X1 U7348 ( .A(n12781), .B(n12795), .ZN(n12753) );
  NAND3_X1 U7349 ( .A1(n6946), .A2(n6945), .A3(n6944), .ZN(n7803) );
  OAI21_X1 U7350 ( .B1(n14442), .B2(n14443), .A(n6875), .ZN(n6874) );
  NAND2_X1 U7351 ( .A1(n8377), .A2(n8376), .ZN(n11449) );
  OAI21_X1 U7352 ( .B1(n11503), .B2(n11502), .A(n11501), .ZN(n11512) );
  OAI21_X1 U7353 ( .B1(n11306), .B2(n6975), .A(n6972), .ZN(n11455) );
  NAND2_X1 U7354 ( .A1(n7492), .A2(n7491), .ZN(n7494) );
  NAND2_X1 U7355 ( .A1(n11331), .A2(n8659), .ZN(n11306) );
  AND2_X1 U7356 ( .A1(n6641), .A2(n6640), .ZN(n14437) );
  NAND2_X1 U7357 ( .A1(n14976), .A2(n11680), .ZN(n11802) );
  AND2_X1 U7358 ( .A1(n15012), .A2(n7605), .ZN(n11255) );
  NAND4_X1 U7359 ( .A1(n6939), .A2(P1_DATAO_REG_13__SCAN_IN), .A3(n6941), .A4(
        n6938), .ZN(n7712) );
  XNOR2_X1 U7360 ( .A(n9754), .B(n6871), .ZN(n14278) );
  NAND2_X1 U7361 ( .A1(n15139), .A2(n9751), .ZN(n9754) );
  AOI21_X1 U7362 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n9703), .A(n9702), .ZN(
        n9704) );
  NOR2_X1 U7363 ( .A1(n10882), .A2(n14789), .ZN(n11152) );
  INV_X2 U7364 ( .A(n14733), .ZN(n14736) );
  NAND2_X1 U7365 ( .A1(n7702), .A2(n7701), .ZN(n7704) );
  NAND2_X1 U7366 ( .A1(n6626), .A2(n6816), .ZN(n11197) );
  NAND2_X1 U7367 ( .A1(n8338), .A2(n8337), .ZN(n14813) );
  OR2_X1 U7368 ( .A1(n14924), .A2(n6897), .ZN(n6895) );
  NOR2_X1 U7369 ( .A1(n14274), .A2(n14275), .ZN(n14273) );
  AND2_X1 U7370 ( .A1(n13310), .A2(n14746), .ZN(n11176) );
  NOR2_X1 U7371 ( .A1(n10721), .A2(n7389), .ZN(n10692) );
  NAND2_X2 U7372 ( .A1(n10665), .A2(n15009), .ZN(n15080) );
  OR2_X1 U7373 ( .A1(n10866), .A2(n11457), .ZN(n10459) );
  AND2_X1 U7374 ( .A1(n10616), .A2(n14746), .ZN(n11173) );
  INV_X1 U7375 ( .A(n10616), .ZN(n13310) );
  NAND4_X1 U7376 ( .A1(n8241), .A2(n8240), .A3(n8239), .A4(n8238), .ZN(n13306)
         );
  NAND2_X2 U7377 ( .A1(n6996), .A2(n8218), .ZN(n10981) );
  NAND2_X1 U7378 ( .A1(n8763), .A2(n6655), .ZN(n10714) );
  AND2_X1 U7379 ( .A1(n8216), .A2(n8217), .ZN(n6996) );
  CLKBUF_X1 U7380 ( .A(n8233), .Z(n6481) );
  BUF_X4 U7381 ( .A(n8233), .Z(n6482) );
  NAND3_X1 U7382 ( .A1(n7535), .A2(n7534), .A3(n7533), .ZN(n10404) );
  INV_X4 U7383 ( .A(n9472), .ZN(n9635) );
  NAND4_X1 U7384 ( .A1(n8758), .A2(n8757), .A3(n8756), .A4(n8755), .ZN(n13772)
         );
  INV_X4 U7385 ( .A(n8469), .ZN(n8576) );
  NAND2_X1 U7386 ( .A1(n7377), .A2(n8718), .ZN(n13773) );
  INV_X2 U7387 ( .A(n8465), .ZN(n8575) );
  NAND4_X2 U7388 ( .A1(n8746), .A2(n8745), .A3(n8744), .A4(n8743), .ZN(n13776)
         );
  NAND2_X1 U7389 ( .A1(n8742), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n8745) );
  INV_X1 U7390 ( .A(n10087), .ZN(n10085) );
  AOI21_X1 U7391 ( .B1(n6794), .B2(n6791), .A(n6790), .ZN(n6789) );
  NAND2_X1 U7392 ( .A1(n8607), .A2(n8606), .ZN(n14725) );
  CLKBUF_X3 U7393 ( .A(n7540), .Z(n12315) );
  AND2_X1 U7394 ( .A1(n7475), .A2(n7480), .ZN(n7540) );
  NAND2_X2 U7395 ( .A1(n10341), .A2(n8050), .ZN(n7804) );
  OAI21_X1 U7396 ( .B1(n9131), .B2(n7374), .A(n9130), .ZN(n11941) );
  INV_X1 U7397 ( .A(n7480), .ZN(n13133) );
  XNOR2_X1 U7398 ( .A(n7914), .B(P3_IR_REG_22__SCAN_IN), .ZN(n12543) );
  CLKBUF_X1 U7399 ( .A(n9168), .Z(n14023) );
  AND2_X1 U7400 ( .A1(n8717), .A2(n8716), .ZN(n8983) );
  INV_X1 U7401 ( .A(n7481), .ZN(n7475) );
  MUX2_X1 U7402 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8142), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n8143) );
  AND2_X2 U7403 ( .A1(n7474), .A2(n13128), .ZN(n7480) );
  INV_X1 U7404 ( .A(n11251), .ZN(n9343) );
  INV_X1 U7405 ( .A(n9153), .ZN(n9131) );
  XNOR2_X1 U7406 ( .A(n7920), .B(n7919), .ZN(n10898) );
  MUX2_X1 U7407 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7472), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n7474) );
  NAND2_X1 U7408 ( .A1(n9069), .A2(n9068), .ZN(n11251) );
  XNOR2_X1 U7409 ( .A(n8146), .B(n8145), .ZN(n13588) );
  INV_X1 U7410 ( .A(n8716), .ZN(n14244) );
  OR2_X1 U7411 ( .A1(n9151), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n9153) );
  MUX2_X1 U7412 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8723), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n8725) );
  OR2_X1 U7413 ( .A1(n8144), .A2(n8151), .ZN(n8146) );
  OAI21_X1 U7414 ( .B1(n8603), .B2(P2_IR_REG_20__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8602) );
  OR2_X1 U7415 ( .A1(n7473), .A2(n7460), .ZN(n6867) );
  NAND2_X1 U7416 ( .A1(n8724), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8720) );
  NAND2_X2 U7417 ( .A1(n6706), .A2(P3_U3151), .ZN(n12303) );
  INV_X4 U7418 ( .A(n8726), .ZN(n6706) );
  NAND2_X2 U7419 ( .A1(n8050), .A2(P3_U3151), .ZN(n13138) );
  INV_X2 U7420 ( .A(n8050), .ZN(n6475) );
  AND2_X1 U7421 ( .A1(n7383), .A2(n6523), .ZN(n7127) );
  AND2_X1 U7422 ( .A1(n7383), .A2(n7124), .ZN(n7126) );
  AND2_X1 U7423 ( .A1(n6523), .A2(n7125), .ZN(n7124) );
  AND2_X1 U7424 ( .A1(n8600), .A2(n8138), .ZN(n7383) );
  AND3_X1 U7425 ( .A1(n8137), .A2(n8136), .A3(n8135), .ZN(n8600) );
  AND4_X1 U7426 ( .A1(n8702), .A2(n8701), .A3(n8929), .A4(n8915), .ZN(n8703)
         );
  NOR2_X1 U7427 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(n8149), .ZN(n7125) );
  AND2_X1 U7428 ( .A1(n8196), .A2(n8132), .ZN(n8214) );
  INV_X1 U7429 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n7496) );
  XOR2_X1 U7430 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), .Z(
        n9730) );
  NOR2_X1 U7431 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n8196) );
  INV_X1 U7432 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7466) );
  BUF_X1 U7433 ( .A(P3_IR_REG_0__SCAN_IN), .Z(n13142) );
  INV_X1 U7434 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n6753) );
  INV_X1 U7435 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n7746) );
  NOR2_X1 U7436 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n8129) );
  NOR3_X1 U7437 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .A3(
        P2_IR_REG_4__SCAN_IN), .ZN(n8133) );
  NOR2_X1 U7438 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), .ZN(
        n7454) );
  NOR2_X1 U7439 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .ZN(
        n7453) );
  NOR2_X1 U7440 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n6814) );
  INV_X4 U7441 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X2 U7442 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n8727) );
  NOR2_X1 U7443 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n7448) );
  NOR2_X1 U7444 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_5__SCAN_IN), .ZN(
        n7449) );
  NOR2_X1 U7445 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), .ZN(
        n7450) );
  OAI21_X2 U7446 ( .B1(n14289), .B2(n13057), .A(n14295), .ZN(n12799) );
  OAI21_X1 U7447 ( .B1(n11435), .B2(n11443), .A(n8375), .ZN(n8377) );
  AOI21_X2 U7449 ( .B1(n12867), .B2(n7897), .A(n6519), .ZN(n8029) );
  NOR2_X2 U7450 ( .A1(n10298), .A2(n10297), .ZN(n10296) );
  INV_X4 U7451 ( .A(n9109), .ZN(n8742) );
  XNOR2_X1 U7452 ( .A(n7552), .B(n7551), .ZN(n14272) );
  NOR2_X2 U7453 ( .A1(n12963), .A2(n12964), .ZN(n12962) );
  OAI22_X2 U7454 ( .A1(n12976), .A2(n12980), .B1(n12989), .B2(n13113), .ZN(
        n12963) );
  NOR2_X2 U7455 ( .A1(n10747), .A2(n10714), .ZN(n10799) );
  AOI21_X2 U7456 ( .B1(n12801), .B2(n14310), .A(n12800), .ZN(n12813) );
  NAND2_X1 U7457 ( .A1(n14745), .A2(n8681), .ZN(n6477) );
  INV_X2 U7458 ( .A(n11440), .ZN(n11505) );
  NAND2_X1 U7459 ( .A1(n8608), .A2(n13588), .ZN(n6478) );
  NAND2_X1 U7460 ( .A1(n8608), .A2(n13588), .ZN(n6479) );
  NAND2_X1 U7461 ( .A1(n8608), .A2(n13588), .ZN(n10196) );
  NAND2_X1 U7462 ( .A1(n10449), .A2(n10448), .ZN(n6480) );
  OAI21_X2 U7463 ( .B1(n11674), .B2(n11637), .A(n14916), .ZN(n11675) );
  AOI211_X2 U7464 ( .C1(n14109), .C2(n14526), .A(n14108), .B(n14107), .ZN(
        n14110) );
  AOI21_X2 U7465 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(n9768), .A(n14449), .ZN(
        n14455) );
  OAI22_X2 U7466 ( .A1(n11449), .A2(n7108), .B1(n11504), .B2(n7107), .ZN(
        n11756) );
  NOR2_X2 U7467 ( .A1(n14455), .A2(n14454), .ZN(n14453) );
  OAI22_X2 U7468 ( .A1(n13404), .A2(n8532), .B1(n13411), .B2(n13287), .ZN(
        n13389) );
  OR2_X4 U7469 ( .A1(n6870), .A2(n6869), .ZN(n11180) );
  OR2_X1 U7470 ( .A1(n13033), .A2(n12940), .ZN(n12446) );
  INV_X1 U7471 ( .A(n7246), .ZN(n7242) );
  NOR2_X1 U7472 ( .A1(n7596), .A2(n6826), .ZN(n6824) );
  NAND2_X1 U7473 ( .A1(n7452), .A2(n6827), .ZN(n6826) );
  INV_X1 U7474 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n6827) );
  INV_X1 U7475 ( .A(n8767), .ZN(n8991) );
  AND2_X1 U7476 ( .A1(n11856), .A2(n9251), .ZN(n7354) );
  NAND2_X1 U7477 ( .A1(n8060), .A2(n8059), .ZN(n8271) );
  AOI21_X1 U7478 ( .B1(n6833), .B2(n6838), .A(n6832), .ZN(n6831) );
  INV_X1 U7479 ( .A(n8766), .ZN(n9338) );
  NAND2_X1 U7480 ( .A1(n9198), .A2(n9199), .ZN(n7339) );
  INV_X1 U7481 ( .A(n7309), .ZN(n7308) );
  OR4_X1 U7482 ( .A1(n8899), .A2(n9172), .A3(n9171), .A4(n9233), .ZN(n9250) );
  AND2_X1 U7483 ( .A1(n7210), .A2(n9538), .ZN(n7209) );
  NAND2_X1 U7484 ( .A1(n9592), .A2(n9591), .ZN(n9593) );
  INV_X1 U7485 ( .A(n9589), .ZN(n9592) );
  AOI21_X1 U7486 ( .B1(n7191), .B2(n7188), .A(n7187), .ZN(n7186) );
  INV_X1 U7487 ( .A(n9598), .ZN(n7187) );
  NOR2_X1 U7488 ( .A1(n7196), .A2(n7188), .ZN(n7190) );
  NOR2_X1 U7489 ( .A1(n6982), .A2(n9650), .ZN(n6981) );
  NOR2_X1 U7490 ( .A1(n6515), .A2(n6983), .ZN(n6982) );
  AOI21_X1 U7491 ( .B1(n6789), .B2(n6792), .A(n6545), .ZN(n6788) );
  AND2_X1 U7492 ( .A1(n6795), .A2(n7376), .ZN(n6794) );
  NAND2_X1 U7493 ( .A1(n8346), .A2(n8079), .ZN(n6795) );
  OR2_X1 U7494 ( .A1(n9445), .A2(n11029), .ZN(n12491) );
  OR2_X1 U7495 ( .A1(n7997), .A2(n12560), .ZN(n12481) );
  INV_X1 U7496 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n7913) );
  XNOR2_X1 U7497 ( .A(n9634), .B(n9636), .ZN(n9658) );
  AND2_X1 U7498 ( .A1(n7116), .A2(n7114), .ZN(n7113) );
  INV_X1 U7499 ( .A(n13443), .ZN(n7114) );
  INV_X1 U7500 ( .A(n8661), .ZN(n6976) );
  AND2_X1 U7501 ( .A1(n8683), .A2(n9669), .ZN(n9475) );
  NAND2_X1 U7502 ( .A1(n7299), .A2(n7298), .ZN(n9348) );
  NAND2_X1 U7503 ( .A1(n9320), .A2(n9319), .ZN(n7298) );
  OAI21_X1 U7504 ( .B1(n9317), .B2(n7301), .A(n6643), .ZN(n7299) );
  NOR2_X1 U7505 ( .A1(n7300), .A2(n9316), .ZN(n7301) );
  NOR2_X1 U7506 ( .A1(n14030), .A2(n6695), .ZN(n6694) );
  INV_X1 U7507 ( .A(n8977), .ZN(n6695) );
  OR2_X1 U7508 ( .A1(n14419), .A2(n12029), .ZN(n9245) );
  INV_X1 U7509 ( .A(n13773), .ZN(n10693) );
  INV_X1 U7510 ( .A(n9087), .ZN(n7348) );
  AOI21_X1 U7511 ( .B1(n7323), .B2(n9322), .A(n6608), .ZN(n7322) );
  INV_X1 U7512 ( .A(n6799), .ZN(n6811) );
  NAND2_X1 U7513 ( .A1(n8524), .A2(n8118), .ZN(n6799) );
  INV_X1 U7514 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7271) );
  INV_X1 U7515 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9064) );
  INV_X1 U7516 ( .A(n8500), .ZN(n8107) );
  NAND2_X1 U7517 ( .A1(n8444), .A2(n8445), .ZN(n6717) );
  XNOR2_X1 U7518 ( .A(n8096), .B(SI_17_), .ZN(n8445) );
  NAND2_X1 U7519 ( .A1(n8075), .A2(n8074), .ZN(n8347) );
  NAND2_X1 U7520 ( .A1(n13066), .A2(n12835), .ZN(n12502) );
  AND4_X1 U7521 ( .A1(n7882), .A2(n7881), .A3(n7880), .A4(n7879), .ZN(n7948)
         );
  OR2_X1 U7522 ( .A1(n14940), .A2(n11642), .ZN(n6897) );
  NAND2_X1 U7523 ( .A1(n11614), .A2(n6898), .ZN(n6896) );
  INV_X1 U7524 ( .A(n14940), .ZN(n6898) );
  AND4_X1 U7525 ( .A1(n7870), .A2(n7869), .A3(n7868), .A4(n7867), .ZN(n12885)
         );
  AOI21_X1 U7526 ( .B1(n6837), .B2(n6835), .A(n6834), .ZN(n6833) );
  INV_X1 U7527 ( .A(n12442), .ZN(n6835) );
  INV_X1 U7528 ( .A(n12446), .ZN(n6834) );
  OR2_X1 U7529 ( .A1(n12943), .A2(n12955), .ZN(n12442) );
  AOI21_X1 U7530 ( .B1(n7241), .B2(n7654), .A(n6495), .ZN(n7239) );
  NAND2_X1 U7531 ( .A1(n7921), .A2(n12336), .ZN(n15060) );
  NAND2_X1 U7532 ( .A1(n7639), .A2(n7638), .ZN(n11353) );
  AOI21_X1 U7533 ( .B1(n11252), .B2(n6855), .A(n6854), .ZN(n6853) );
  INV_X1 U7534 ( .A(n12369), .ZN(n6855) );
  INV_X1 U7535 ( .A(n12371), .ZN(n6854) );
  AND2_X1 U7536 ( .A1(n7957), .A2(n7958), .ZN(n11829) );
  INV_X1 U7537 ( .A(n7804), .ZN(n12322) );
  INV_X1 U7538 ( .A(n15060), .ZN(n15045) );
  INV_X1 U7539 ( .A(n14339), .ZN(n15063) );
  OAI21_X1 U7540 ( .B1(n10168), .B2(P3_D_REG_1__SCAN_IN), .A(n7975), .ZN(
        n10659) );
  OR2_X1 U7541 ( .A1(n7470), .A2(n7460), .ZN(n7461) );
  NAND2_X1 U7542 ( .A1(n7843), .A2(n7842), .ZN(n7846) );
  INV_X1 U7543 ( .A(n6929), .ZN(n6928) );
  OAI21_X1 U7544 ( .B1(n7680), .B2(n6930), .A(n7501), .ZN(n6929) );
  NOR2_X1 U7545 ( .A1(n13144), .A2(n7157), .ZN(n7156) );
  INV_X1 U7546 ( .A(n12204), .ZN(n7157) );
  NAND2_X1 U7547 ( .A1(n12211), .A2(n7154), .ZN(n7153) );
  INV_X1 U7548 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n7134) );
  AND2_X1 U7549 ( .A1(n6774), .A2(n6578), .ZN(n7096) );
  INV_X1 U7550 ( .A(n7100), .ZN(n7097) );
  XNOR2_X1 U7551 ( .A(n13492), .B(n6785), .ZN(n13355) );
  NAND2_X1 U7552 ( .A1(n8385), .A2(n8384), .ZN(n11504) );
  NAND2_X1 U7553 ( .A1(n10827), .A2(n10833), .ZN(n8656) );
  OAI22_X1 U7554 ( .A1(n9474), .A2(n11176), .B1(n13308), .B2(n11180), .ZN(
        n10969) );
  OAI21_X1 U7555 ( .B1(n9168), .B2(n9167), .A(n10076), .ZN(n12066) );
  XNOR2_X1 U7556 ( .A(n11074), .B(n11075), .ZN(n11116) );
  NAND3_X1 U7557 ( .A1(n11876), .A2(n11843), .A3(n11841), .ZN(n11877) );
  AND4_X1 U7558 ( .A1(n8927), .A2(n8926), .A3(n8925), .A4(n8924), .ZN(n12048)
         );
  NOR2_X1 U7559 ( .A1(n13907), .A2(n14198), .ZN(n13895) );
  NAND2_X1 U7560 ( .A1(n13908), .A2(n14106), .ZN(n13907) );
  NAND2_X1 U7561 ( .A1(n9057), .A2(n13899), .ZN(n9393) );
  AOI21_X1 U7562 ( .B1(n6489), .B2(n6693), .A(n6533), .ZN(n6689) );
  OR2_X1 U7563 ( .A1(n14155), .A2(n13754), .ZN(n6696) );
  NAND2_X1 U7564 ( .A1(n6698), .A2(n6697), .ZN(n8955) );
  AOI21_X1 U7565 ( .B1(n6699), .B2(n6507), .A(n6590), .ZN(n6697) );
  NAND2_X1 U7566 ( .A1(n6660), .A2(n6661), .ZN(n14086) );
  INV_X1 U7567 ( .A(n6662), .ZN(n6661) );
  OAI21_X1 U7568 ( .B1(n7352), .B2(n6663), .A(n9092), .ZN(n6662) );
  NAND2_X1 U7569 ( .A1(n6683), .A2(n7062), .ZN(n11247) );
  AOI21_X1 U7570 ( .B1(n7063), .B2(n7065), .A(n6540), .ZN(n7062) );
  NAND2_X1 U7571 ( .A1(n10964), .A2(n7063), .ZN(n6683) );
  NAND2_X1 U7572 ( .A1(n6669), .A2(n6668), .ZN(n11239) );
  AOI21_X1 U7573 ( .B1(n6671), .B2(n6672), .A(n6529), .ZN(n6668) );
  NAND2_X1 U7574 ( .A1(n11201), .A2(n6675), .ZN(n6670) );
  NAND2_X1 U7575 ( .A1(n6667), .A2(n6671), .ZN(n11046) );
  OR2_X1 U7576 ( .A1(n6672), .A2(n11201), .ZN(n6667) );
  OR2_X1 U7577 ( .A1(n11201), .A2(n9083), .ZN(n6677) );
  NAND2_X1 U7578 ( .A1(n8765), .A2(n7081), .ZN(n7080) );
  NOR2_X1 U7579 ( .A1(n8778), .A2(n7082), .ZN(n7081) );
  INV_X1 U7580 ( .A(n8764), .ZN(n7082) );
  OR2_X1 U7581 ( .A1(n9328), .A2(n9327), .ZN(n9353) );
  AND2_X1 U7582 ( .A1(n8560), .A2(n8559), .ZN(n13592) );
  NAND2_X1 U7583 ( .A1(n7288), .A2(n8063), .ZN(n8286) );
  NAND2_X1 U7584 ( .A1(n8271), .A2(n8270), .ZN(n7288) );
  AOI21_X1 U7585 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n9711), .A(n9710), .ZN(
        n9723) );
  NOR2_X1 U7586 ( .A1(n9764), .A2(n9763), .ZN(n9710) );
  OR2_X1 U7587 ( .A1(n7932), .A2(n12488), .ZN(n14341) );
  INV_X1 U7588 ( .A(n7948), .ZN(n12870) );
  AND2_X1 U7589 ( .A1(n8025), .A2(n8024), .ZN(n12853) );
  OR2_X1 U7590 ( .A1(n8023), .A2(n12526), .ZN(n8024) );
  INV_X1 U7591 ( .A(n8613), .ZN(n8614) );
  XNOR2_X1 U7592 ( .A(n8680), .B(n8679), .ZN(n13480) );
  INV_X1 U7593 ( .A(n9657), .ZN(n8679) );
  NOR2_X1 U7594 ( .A1(n9198), .A2(n9199), .ZN(n7338) );
  NAND2_X1 U7595 ( .A1(n7217), .A2(n9498), .ZN(n7215) );
  INV_X1 U7596 ( .A(n9497), .ZN(n7217) );
  NAND2_X1 U7597 ( .A1(n7331), .A2(n9213), .ZN(n7330) );
  NAND2_X1 U7598 ( .A1(n7316), .A2(n9223), .ZN(n7315) );
  NAND2_X1 U7599 ( .A1(n9255), .A2(n9256), .ZN(n7309) );
  NOR2_X1 U7600 ( .A1(n7306), .A2(n7305), .ZN(n7304) );
  AOI22_X1 U7601 ( .A1(n7306), .A2(n7310), .B1(n9258), .B2(n7303), .ZN(n7302)
         );
  OR2_X1 U7602 ( .A1(n9539), .A2(n9538), .ZN(n9540) );
  NOR2_X1 U7603 ( .A1(n7328), .A2(n9270), .ZN(n7325) );
  AOI21_X1 U7604 ( .B1(n9270), .B2(n7328), .A(n7327), .ZN(n7326) );
  NAND2_X1 U7605 ( .A1(n9564), .A2(n9566), .ZN(n7219) );
  AND2_X1 U7606 ( .A1(n7196), .A2(n7192), .ZN(n7191) );
  NAND2_X1 U7607 ( .A1(n7195), .A2(n7193), .ZN(n7192) );
  INV_X1 U7608 ( .A(n13178), .ZN(n7176) );
  INV_X1 U7609 ( .A(n7191), .ZN(n7189) );
  NOR2_X1 U7610 ( .A1(n7194), .A2(n9597), .ZN(n7195) );
  NAND2_X1 U7611 ( .A1(n7185), .A2(n7184), .ZN(n7183) );
  INV_X1 U7612 ( .A(n7190), .ZN(n7184) );
  AND2_X1 U7613 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(n8536), .ZN(n8539) );
  INV_X1 U7614 ( .A(n8666), .ZN(n6983) );
  INV_X1 U7615 ( .A(n8119), .ZN(n6808) );
  AND2_X1 U7616 ( .A1(n6801), .A2(n6805), .ZN(n6800) );
  INV_X1 U7617 ( .A(n8553), .ZN(n6805) );
  NAND2_X1 U7618 ( .A1(n6806), .A2(SI_24_), .ZN(n6801) );
  NOR2_X1 U7619 ( .A1(n6806), .A2(SI_24_), .ZN(n6802) );
  AND2_X1 U7620 ( .A1(n7289), .A2(n6789), .ZN(n6725) );
  INV_X1 U7621 ( .A(n15072), .ZN(n7539) );
  AND2_X1 U7622 ( .A1(n12635), .A2(n7019), .ZN(n7018) );
  NAND2_X1 U7623 ( .A1(n7022), .A2(n7021), .ZN(n7019) );
  AOI21_X1 U7624 ( .B1(n12497), .B2(n12496), .A(n12495), .ZN(n12498) );
  OAI21_X1 U7625 ( .B1(n6476), .B2(n10356), .A(n6625), .ZN(n10360) );
  NAND2_X1 U7626 ( .A1(n6476), .A2(n10356), .ZN(n6625) );
  AND2_X1 U7627 ( .A1(n12868), .A2(n7261), .ZN(n7260) );
  NAND2_X1 U7628 ( .A1(n12457), .A2(n7857), .ZN(n7261) );
  INV_X1 U7629 ( .A(n7857), .ZN(n7262) );
  AND2_X1 U7630 ( .A1(n12457), .A2(n12881), .ZN(n12463) );
  INV_X1 U7631 ( .A(n7231), .ZN(n7230) );
  INV_X1 U7632 ( .A(n7234), .ZN(n7228) );
  INV_X1 U7633 ( .A(n7809), .ZN(n7478) );
  NAND2_X1 U7634 ( .A1(n12951), .A2(n7232), .ZN(n7231) );
  INV_X1 U7635 ( .A(n7371), .ZN(n7232) );
  NOR2_X1 U7636 ( .A1(n7941), .A2(n6864), .ZN(n6863) );
  INV_X1 U7637 ( .A(n12406), .ZN(n6864) );
  NAND2_X1 U7638 ( .A1(n15068), .A2(n15059), .ZN(n15058) );
  AND2_X1 U7639 ( .A1(n7459), .A2(n7267), .ZN(n7266) );
  NOR2_X1 U7640 ( .A1(P3_IR_REG_28__SCAN_IN), .A2(P3_IR_REG_27__SCAN_IN), .ZN(
        n7267) );
  AND2_X1 U7641 ( .A1(n7457), .A2(n7964), .ZN(n7969) );
  INV_X1 U7642 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7457) );
  INV_X1 U7643 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n7964) );
  NOR2_X1 U7644 ( .A1(n7918), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n7915) );
  INV_X1 U7645 ( .A(n7417), .ZN(n6960) );
  INV_X1 U7646 ( .A(n12182), .ZN(n7173) );
  AND2_X1 U7647 ( .A1(n7177), .A2(n7176), .ZN(n7175) );
  INV_X1 U7648 ( .A(n11163), .ZN(n7142) );
  INV_X1 U7649 ( .A(n12209), .ZN(n12199) );
  NAND2_X1 U7650 ( .A1(n6481), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7088) );
  AND2_X1 U7651 ( .A1(n8563), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8163) );
  NAND2_X1 U7652 ( .A1(n13436), .A2(n6992), .ZN(n6991) );
  NAND2_X1 U7653 ( .A1(n8673), .A2(n8672), .ZN(n6992) );
  NOR2_X1 U7654 ( .A1(n13537), .A2(n12171), .ZN(n6884) );
  INV_X1 U7655 ( .A(n6516), .ZN(n6968) );
  INV_X1 U7656 ( .A(n8285), .ZN(n7091) );
  NOR2_X1 U7657 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n6993) );
  NOR2_X1 U7658 ( .A1(n8597), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n8623) );
  INV_X1 U7659 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8637) );
  OAI21_X1 U7660 ( .B1(n12083), .B2(n6732), .A(n6503), .ZN(n13612) );
  NAND2_X1 U7661 ( .A1(n7053), .A2(n11427), .ZN(n7052) );
  INV_X1 U7662 ( .A(n11425), .ZN(n7053) );
  NOR2_X1 U7663 ( .A1(n11425), .A2(n11426), .ZN(n7054) );
  NAND2_X1 U7664 ( .A1(n9402), .A2(n9399), .ZN(n9400) );
  NOR2_X1 U7665 ( .A1(n9398), .A2(n9397), .ZN(n9399) );
  INV_X1 U7667 ( .A(n14106), .ZN(n9368) );
  NOR2_X1 U7668 ( .A1(n7070), .A2(n7069), .ZN(n7068) );
  INV_X1 U7669 ( .A(n9007), .ZN(n7069) );
  INV_X1 U7670 ( .A(n9096), .ZN(n7357) );
  AND2_X1 U7671 ( .A1(n9390), .A2(n9095), .ZN(n7358) );
  INV_X1 U7672 ( .A(n6823), .ZN(n6822) );
  NAND2_X1 U7673 ( .A1(n14233), .A2(n12049), .ZN(n6823) );
  AND2_X1 U7674 ( .A1(n9245), .A2(n9241), .ZN(n9384) );
  AOI21_X1 U7675 ( .B1(n6673), .B2(n6676), .A(n11059), .ZN(n6671) );
  AND2_X1 U7676 ( .A1(n9343), .A2(n11150), .ZN(n10075) );
  NOR2_X1 U7677 ( .A1(n9123), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n7061) );
  AND2_X1 U7678 ( .A1(n8087), .A2(n8090), .ZN(n8088) );
  NAND2_X1 U7679 ( .A1(n6726), .A2(n6788), .ZN(n8086) );
  NAND2_X1 U7680 ( .A1(n8347), .A2(n6789), .ZN(n6726) );
  NAND2_X1 U7681 ( .A1(n8071), .A2(n8070), .ZN(n6715) );
  AOI21_X1 U7682 ( .B1(n7286), .B2(n8287), .A(n6550), .ZN(n7285) );
  INV_X1 U7683 ( .A(n8063), .ZN(n7286) );
  NOR2_X1 U7684 ( .A1(n7287), .A2(n7284), .ZN(n7283) );
  INV_X1 U7685 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n9691) );
  XNOR2_X1 U7686 ( .A(n9690), .B(n9691), .ZN(n9740) );
  NOR2_X1 U7687 ( .A1(n9699), .A2(n9698), .ZN(n9753) );
  AND2_X1 U7688 ( .A1(n6630), .A2(n6629), .ZN(n9764) );
  NAND2_X1 U7689 ( .A1(n9708), .A2(P3_ADDR_REG_11__SCAN_IN), .ZN(n6629) );
  OR2_X1 U7690 ( .A1(n9762), .A2(n9761), .ZN(n6630) );
  OAI21_X1 U7691 ( .B1(P3_ADDR_REG_16__SCAN_IN), .B2(n9717), .A(n9716), .ZN(
        n9772) );
  OR2_X1 U7692 ( .A1(n7891), .A2(n7890), .ZN(n7905) );
  INV_X1 U7693 ( .A(n7030), .ZN(n7029) );
  OAI21_X1 U7694 ( .B1(n10061), .B2(n6581), .A(n10062), .ZN(n7030) );
  NOR2_X1 U7695 ( .A1(n11387), .A2(n7034), .ZN(n7033) );
  INV_X1 U7696 ( .A(n7037), .ZN(n7034) );
  OAI21_X1 U7697 ( .B1(n12597), .B2(n7012), .A(n7010), .ZN(n12556) );
  AOI21_X1 U7698 ( .B1(n12661), .B2(n7011), .A(n10027), .ZN(n7010) );
  INV_X1 U7699 ( .A(n12661), .ZN(n7012) );
  INV_X1 U7700 ( .A(n10025), .ZN(n7011) );
  NAND2_X1 U7701 ( .A1(n9986), .A2(n7387), .ZN(n11904) );
  AND2_X1 U7702 ( .A1(n10025), .A2(n10023), .ZN(n12595) );
  OAI21_X1 U7703 ( .B1(n12565), .B2(n10020), .A(n10019), .ZN(n12593) );
  OR2_X1 U7704 ( .A1(n11904), .A2(n9987), .ZN(n7028) );
  OR2_X1 U7705 ( .A1(n10016), .A2(n10015), .ZN(n7023) );
  AND2_X1 U7706 ( .A1(n9958), .A2(n9957), .ZN(n9959) );
  NAND2_X1 U7707 ( .A1(n10404), .A2(n10668), .ZN(n15059) );
  XNOR2_X1 U7708 ( .A(n11678), .B(n11615), .ZN(n14971) );
  AND3_X2 U7709 ( .A1(n6895), .A2(n6896), .A3(n6584), .ZN(n11616) );
  NOR2_X1 U7710 ( .A1(n14990), .A2(n14989), .ZN(n14988) );
  OR2_X1 U7711 ( .A1(n14988), .A2(n6891), .ZN(n6890) );
  AND2_X1 U7712 ( .A1(n11665), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n6891) );
  NOR2_X1 U7713 ( .A1(n12703), .A2(n6889), .ZN(n12722) );
  NOR2_X1 U7714 ( .A1(n12706), .A2(n7696), .ZN(n6889) );
  NAND2_X1 U7715 ( .A1(n12752), .A2(n12758), .ZN(n12781) );
  OR2_X2 U7716 ( .A1(n12753), .A2(n6910), .ZN(n6909) );
  OR2_X1 U7717 ( .A1(n14301), .A2(n12754), .ZN(n6910) );
  NAND2_X1 U7718 ( .A1(n12782), .A2(n6908), .ZN(n6907) );
  INV_X1 U7719 ( .A(n14301), .ZN(n6908) );
  OR2_X1 U7720 ( .A1(n12753), .A2(n12754), .ZN(n6912) );
  INV_X1 U7721 ( .A(n6915), .ZN(n6913) );
  OAI21_X1 U7722 ( .B1(n9444), .B2(n9443), .A(n12481), .ZN(n12305) );
  AND2_X1 U7723 ( .A1(n12451), .A2(n12452), .ZN(n12912) );
  NAND2_X1 U7724 ( .A1(n12937), .A2(n12442), .ZN(n6839) );
  NAND2_X1 U7725 ( .A1(n7800), .A2(n12687), .ZN(n7234) );
  AND4_X1 U7726 ( .A1(n7485), .A2(n7484), .A3(n7483), .A4(n7482), .ZN(n12940)
         );
  OR2_X1 U7727 ( .A1(n12962), .A2(n7231), .ZN(n12950) );
  AND2_X1 U7728 ( .A1(n12428), .A2(n12433), .ZN(n12964) );
  NAND2_X1 U7729 ( .A1(n7943), .A2(n6865), .ZN(n12967) );
  NOR2_X1 U7730 ( .A1(n12970), .A2(n6866), .ZN(n6865) );
  AOI21_X1 U7731 ( .B1(n14326), .B2(n7249), .A(n7248), .ZN(n12976) );
  AND2_X1 U7732 ( .A1(n7252), .A2(n12986), .ZN(n7249) );
  OAI21_X1 U7733 ( .B1(n7250), .B2(n12990), .A(n6551), .ZN(n7248) );
  AND2_X1 U7734 ( .A1(n12430), .A2(n12427), .ZN(n12980) );
  AND4_X1 U7735 ( .A1(n7784), .A2(n7783), .A3(n7782), .A4(n7781), .ZN(n12989)
         );
  NOR2_X1 U7736 ( .A1(n13003), .A2(n12518), .ZN(n7252) );
  INV_X1 U7737 ( .A(n7251), .ZN(n7250) );
  OAI21_X1 U7738 ( .B1(n13003), .B2(n7256), .A(n7254), .ZN(n7251) );
  NAND2_X1 U7739 ( .A1(n9993), .A2(n7255), .ZN(n7254) );
  AND4_X1 U7740 ( .A1(n7770), .A2(n7769), .A3(n7768), .A4(n7767), .ZN(n13001)
         );
  AND2_X1 U7741 ( .A1(n12417), .A2(n12422), .ZN(n13003) );
  AOI21_X1 U7742 ( .B1(n6863), .B2(n12514), .A(n6861), .ZN(n6860) );
  INV_X1 U7743 ( .A(n12407), .ZN(n6861) );
  INV_X1 U7744 ( .A(n6863), .ZN(n6862) );
  NAND2_X1 U7745 ( .A1(n11828), .A2(n11827), .ZN(n11826) );
  NAND2_X1 U7746 ( .A1(n6841), .A2(n6840), .ZN(n11586) );
  AOI22_X1 U7747 ( .A1(n6843), .A2(n6850), .B1(n6846), .B2(n6848), .ZN(n6840)
         );
  OR2_X1 U7748 ( .A1(n6846), .A2(n6843), .ZN(n6842) );
  NAND2_X1 U7749 ( .A1(n11353), .A2(n7241), .ZN(n7235) );
  OAI21_X1 U7750 ( .B1(n11353), .B2(n7238), .A(n7236), .ZN(n11587) );
  INV_X1 U7751 ( .A(n7239), .ZN(n7238) );
  AOI21_X1 U7752 ( .B1(n7239), .B2(n7240), .A(n7237), .ZN(n7236) );
  NAND2_X1 U7753 ( .A1(n11350), .A2(n12503), .ZN(n11352) );
  AND2_X1 U7754 ( .A1(n12382), .A2(n12383), .ZN(n12503) );
  NAND2_X1 U7755 ( .A1(n6853), .A2(n12507), .ZN(n6852) );
  NAND2_X1 U7756 ( .A1(n12381), .A2(n7637), .ZN(n11226) );
  AND4_X1 U7757 ( .A1(n7612), .A2(n7611), .A3(n7610), .A4(n7609), .ZN(n15018)
         );
  AND2_X1 U7758 ( .A1(n7603), .A2(n7584), .ZN(n7263) );
  INV_X1 U7759 ( .A(n15015), .ZN(n7603) );
  AND2_X1 U7760 ( .A1(n12369), .A2(n12364), .ZN(n15015) );
  AND4_X1 U7761 ( .A1(n7593), .A2(n7592), .A3(n7591), .A4(n7590), .ZN(n15029)
         );
  NAND2_X1 U7762 ( .A1(n10915), .A2(n7572), .ZN(n15028) );
  INV_X1 U7763 ( .A(n12700), .ZN(n15017) );
  INV_X1 U7764 ( .A(n9431), .ZN(n12312) );
  NAND2_X1 U7765 ( .A1(n7877), .A2(n7876), .ZN(n7949) );
  OR2_X1 U7766 ( .A1(n9431), .A2(n11691), .ZN(n7861) );
  NAND2_X1 U7767 ( .A1(n7974), .A2(n7983), .ZN(n10168) );
  OAI22_X1 U7768 ( .A1(n12300), .A2(n12299), .B1(P2_DATAO_REG_29__SCAN_IN), 
        .B2(n13582), .ZN(n12309) );
  NAND2_X1 U7769 ( .A1(n6963), .A2(n6962), .ZN(n9427) );
  AOI21_X1 U7770 ( .B1(n6509), .B2(n6964), .A(n6609), .ZN(n6962) );
  NAND2_X1 U7771 ( .A1(n7846), .A2(n6607), .ZN(n7859) );
  NAND2_X1 U7772 ( .A1(n6616), .A2(n6528), .ZN(n7456) );
  INV_X1 U7773 ( .A(n7912), .ZN(n6616) );
  OAI21_X1 U7774 ( .B1(n7831), .B2(n7830), .A(n7829), .ZN(n7843) );
  NAND2_X1 U7775 ( .A1(n7816), .A2(n7815), .ZN(n7831) );
  NAND2_X1 U7776 ( .A1(n7803), .A2(n7442), .ZN(n7445) );
  NAND2_X1 U7777 ( .A1(n6947), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7442) );
  NAND2_X1 U7778 ( .A1(n7494), .A2(n7441), .ZN(n6947) );
  NAND2_X1 U7779 ( .A1(n7445), .A2(n7444), .ZN(n7816) );
  NAND2_X1 U7780 ( .A1(n6949), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6948) );
  INV_X1 U7781 ( .A(n7441), .ZN(n6949) );
  INV_X1 U7782 ( .A(n7494), .ZN(n6943) );
  NAND2_X1 U7783 ( .A1(n7494), .A2(n6599), .ZN(n6945) );
  NAND2_X1 U7784 ( .A1(n7788), .A2(n7439), .ZN(n7492) );
  NAND2_X1 U7785 ( .A1(n7744), .A2(n7432), .ZN(n7758) );
  NAND2_X1 U7786 ( .A1(n7758), .A2(n7757), .ZN(n7760) );
  NAND2_X1 U7787 ( .A1(n7730), .A2(n7430), .ZN(n7742) );
  NAND2_X1 U7788 ( .A1(n7712), .A2(n7428), .ZN(n7728) );
  NAND2_X1 U7789 ( .A1(n6940), .A2(n10401), .ZN(n7428) );
  NAND2_X1 U7790 ( .A1(n7704), .A2(n7427), .ZN(n6940) );
  NAND2_X1 U7791 ( .A1(n6937), .A2(n10401), .ZN(n6939) );
  AND2_X1 U7792 ( .A1(n7425), .A2(n7424), .ZN(n7501) );
  INV_X1 U7793 ( .A(n7423), .ZN(n6930) );
  AND2_X1 U7794 ( .A1(n7423), .A2(n7422), .ZN(n7680) );
  NAND2_X1 U7795 ( .A1(n7681), .A2(n7680), .ZN(n7683) );
  OR2_X1 U7796 ( .A1(n7646), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n7666) );
  OR2_X1 U7797 ( .A1(n7666), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n7685) );
  INV_X1 U7798 ( .A(n7648), .ZN(n6956) );
  OAI21_X1 U7799 ( .B1(n7628), .B2(n7416), .A(n7417), .ZN(n7649) );
  NAND2_X1 U7800 ( .A1(n7628), .A2(n7417), .ZN(n6957) );
  AND2_X1 U7801 ( .A1(n7404), .A2(n7403), .ZN(n7563) );
  NOR2_X2 U7802 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n7523) );
  NAND2_X1 U7803 ( .A1(n8514), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8527) );
  INV_X1 U7804 ( .A(n13171), .ZN(n13254) );
  AOI21_X1 U7805 ( .B1(n7179), .B2(n7370), .A(n6598), .ZN(n7177) );
  INV_X1 U7806 ( .A(n7179), .ZN(n7178) );
  NAND2_X1 U7807 ( .A1(n7167), .A2(n7169), .ZN(n7166) );
  INV_X1 U7808 ( .A(n13204), .ZN(n7167) );
  NAND2_X1 U7809 ( .A1(n7139), .A2(n7137), .ZN(n11395) );
  AND2_X1 U7810 ( .A1(n7140), .A2(n7138), .ZN(n7137) );
  INV_X1 U7811 ( .A(n11374), .ZN(n7138) );
  AND2_X1 U7812 ( .A1(n9666), .A2(n11533), .ZN(n10473) );
  NAND2_X1 U7813 ( .A1(n9618), .A2(n9617), .ZN(n9627) );
  NOR4_X1 U7814 ( .A1(n13355), .A2(n13338), .A3(n13374), .A4(n9655), .ZN(n9659) );
  AND2_X1 U7815 ( .A1(n8158), .A2(n13583), .ZN(n8278) );
  AND2_X1 U7816 ( .A1(n8678), .A2(n8585), .ZN(n13338) );
  NAND2_X1 U7817 ( .A1(n13341), .A2(n13146), .ZN(n8585) );
  NAND2_X1 U7818 ( .A1(n13382), .A2(n13255), .ZN(n6998) );
  NAND2_X1 U7819 ( .A1(n7104), .A2(n7106), .ZN(n7103) );
  NAND2_X1 U7820 ( .A1(n13370), .A2(n6796), .ZN(n7104) );
  NAND2_X1 U7821 ( .A1(n13374), .A2(n7105), .ZN(n6796) );
  NOR2_X1 U7822 ( .A1(n7102), .A2(n7101), .ZN(n7100) );
  INV_X1 U7823 ( .A(n7106), .ZN(n7102) );
  INV_X1 U7824 ( .A(n7105), .ZN(n7101) );
  AND2_X1 U7825 ( .A1(n13507), .A2(n13187), .ZN(n6648) );
  NAND2_X1 U7826 ( .A1(n13526), .A2(n13235), .ZN(n6650) );
  NOR2_X1 U7827 ( .A1(n13526), .A2(n13235), .ZN(n6649) );
  INV_X1 U7828 ( .A(n13435), .ZN(n6651) );
  NAND2_X1 U7829 ( .A1(n6505), .A2(n8487), .ZN(n7116) );
  NAND2_X1 U7830 ( .A1(n7118), .A2(n8487), .ZN(n7117) );
  INV_X1 U7831 ( .A(n8470), .ZN(n7118) );
  NAND2_X1 U7832 ( .A1(n13543), .A2(n13292), .ZN(n7120) );
  NAND2_X1 U7833 ( .A1(n7397), .A2(n8670), .ZN(n13458) );
  NAND2_X1 U7834 ( .A1(n11971), .A2(n8669), .ZN(n11952) );
  OR2_X1 U7835 ( .A1(n13547), .A2(n8454), .ZN(n6621) );
  NAND2_X1 U7836 ( .A1(n8417), .A2(n8416), .ZN(n12161) );
  INV_X1 U7837 ( .A(n8664), .ZN(n6984) );
  AND2_X1 U7838 ( .A1(n9522), .A2(n8332), .ZN(n7122) );
  INV_X1 U7839 ( .A(n11157), .ZN(n6969) );
  NAND2_X1 U7840 ( .A1(n8283), .A2(n10826), .ZN(n10835) );
  NAND2_X1 U7841 ( .A1(n10981), .A2(n10866), .ZN(n10864) );
  NAND2_X1 U7842 ( .A1(n8434), .A2(n8433), .ZN(n13553) );
  XNOR2_X1 U7843 ( .A(n8152), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8158) );
  NAND2_X1 U7844 ( .A1(n7128), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8152) );
  OR2_X1 U7845 ( .A1(n8625), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n8630) );
  NAND2_X1 U7846 ( .A1(n7129), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8476) );
  AND2_X1 U7847 ( .A1(n7132), .A2(n7131), .ZN(n7130) );
  AND2_X1 U7848 ( .A1(n6496), .A2(n7133), .ZN(n7132) );
  INV_X1 U7849 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n7133) );
  OR2_X1 U7850 ( .A1(n8893), .A2(n8892), .ZN(n8906) );
  NAND2_X1 U7851 ( .A1(n8960), .A2(n8959), .ZN(n12069) );
  NAND2_X1 U7852 ( .A1(n11547), .A2(n11548), .ZN(n7043) );
  AND2_X1 U7853 ( .A1(n11557), .A2(n7043), .ZN(n7042) );
  NAND2_X1 U7854 ( .A1(n13686), .A2(n13685), .ZN(n12083) );
  INV_X1 U7855 ( .A(n11837), .ZN(n11840) );
  AOI21_X1 U7856 ( .B1(n7055), .B2(n6736), .A(n6544), .ZN(n6735) );
  INV_X1 U7857 ( .A(n7058), .ZN(n6736) );
  INV_X1 U7858 ( .A(n7055), .ZN(n6737) );
  NOR2_X1 U7859 ( .A1(n13715), .A2(n7056), .ZN(n7055) );
  INV_X1 U7860 ( .A(n12062), .ZN(n7056) );
  NAND2_X1 U7861 ( .A1(n9363), .A2(n9362), .ZN(n9404) );
  AND3_X1 U7862 ( .A1(n8953), .A2(n8952), .A3(n8951), .ZN(n13625) );
  AND4_X1 U7863 ( .A1(n8773), .A2(n8772), .A3(n8771), .A4(n8770), .ZN(n11071)
         );
  NAND2_X1 U7864 ( .A1(n8766), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n8734) );
  OR2_X1 U7865 ( .A1(n7074), .A2(n6488), .ZN(n7072) );
  NOR2_X1 U7866 ( .A1(n6488), .A2(n13948), .ZN(n7073) );
  INV_X1 U7867 ( .A(n13979), .ZN(n7070) );
  NAND2_X1 U7868 ( .A1(n13994), .A2(n7068), .ZN(n13984) );
  NAND2_X1 U7869 ( .A1(n6818), .A2(n6817), .ZN(n13985) );
  INV_X1 U7870 ( .A(n14212), .ZN(n6817) );
  OR2_X1 U7871 ( .A1(n13996), .A2(n13997), .ZN(n13994) );
  NAND2_X1 U7872 ( .A1(n14028), .A2(n7358), .ZN(n14021) );
  NAND2_X1 U7873 ( .A1(n6692), .A2(n6696), .ZN(n6691) );
  INV_X1 U7874 ( .A(n6694), .ZN(n6692) );
  INV_X1 U7875 ( .A(n6696), .ZN(n6693) );
  NAND2_X1 U7876 ( .A1(n14052), .A2(n6694), .ZN(n6690) );
  NAND2_X1 U7877 ( .A1(n14046), .A2(n9094), .ZN(n14029) );
  NAND2_X1 U7878 ( .A1(n14029), .A2(n14030), .ZN(n14028) );
  NAND2_X1 U7879 ( .A1(n14063), .A2(n7359), .ZN(n14046) );
  NOR2_X1 U7880 ( .A1(n14043), .A2(n7360), .ZN(n7359) );
  INV_X1 U7881 ( .A(n9266), .ZN(n7360) );
  NAND2_X1 U7882 ( .A1(n7084), .A2(n7083), .ZN(n14052) );
  AND2_X1 U7883 ( .A1(n14043), .A2(n8967), .ZN(n7083) );
  NAND2_X1 U7884 ( .A1(n8955), .A2(n7085), .ZN(n7084) );
  NOR2_X1 U7885 ( .A1(n14064), .A2(n7086), .ZN(n7085) );
  INV_X1 U7886 ( .A(n8954), .ZN(n7086) );
  NAND2_X1 U7887 ( .A1(n14087), .A2(n7361), .ZN(n14063) );
  AND2_X1 U7888 ( .A1(n14064), .A2(n9260), .ZN(n7361) );
  OR2_X1 U7889 ( .A1(n14086), .A2(n9387), .ZN(n14087) );
  NOR2_X1 U7890 ( .A1(n7353), .A2(n6666), .ZN(n6665) );
  INV_X1 U7891 ( .A(n9245), .ZN(n6666) );
  INV_X1 U7892 ( .A(n7354), .ZN(n7353) );
  AOI21_X1 U7893 ( .B1(n7354), .B2(n9386), .A(n6542), .ZN(n7352) );
  OR2_X1 U7894 ( .A1(n12041), .A2(n11523), .ZN(n9251) );
  NOR2_X1 U7895 ( .A1(n8912), .A2(n7078), .ZN(n7077) );
  NAND2_X1 U7896 ( .A1(n11863), .A2(n11862), .ZN(n11861) );
  AOI21_X1 U7897 ( .B1(n6494), .B2(n6536), .A(n6484), .ZN(n6658) );
  NAND2_X1 U7898 ( .A1(n11289), .A2(n9380), .ZN(n9086) );
  OAI22_X1 U7899 ( .A1(n11239), .A2(n11246), .B1(n11049), .B2(n11883), .ZN(
        n11289) );
  NAND2_X1 U7900 ( .A1(n6674), .A2(n6511), .ZN(n6673) );
  NAND2_X1 U7901 ( .A1(n10953), .A2(n6678), .ZN(n6674) );
  NAND2_X1 U7902 ( .A1(n9083), .A2(n9084), .ZN(n6678) );
  INV_X1 U7903 ( .A(n7064), .ZN(n7063) );
  OAI21_X1 U7904 ( .B1(n10963), .B2(n7065), .A(n11059), .ZN(n7064) );
  INV_X1 U7905 ( .A(n8826), .ZN(n7065) );
  NAND2_X1 U7906 ( .A1(n11194), .A2(n8812), .ZN(n10964) );
  NAND2_X1 U7907 ( .A1(n10964), .A2(n10963), .ZN(n10962) );
  NAND2_X1 U7908 ( .A1(n9082), .A2(n9081), .ZN(n11201) );
  AND2_X1 U7909 ( .A1(n9372), .A2(n11981), .ZN(n7079) );
  NAND2_X1 U7910 ( .A1(n10799), .A2(n14520), .ZN(n11991) );
  INV_X1 U7911 ( .A(n7067), .ZN(n7351) );
  NAND2_X1 U7912 ( .A1(n6684), .A2(n6687), .ZN(n10745) );
  OR2_X1 U7913 ( .A1(n10085), .A2(n13774), .ZN(n6687) );
  NAND2_X1 U7914 ( .A1(n6686), .A2(n6685), .ZN(n6684) );
  INV_X1 U7915 ( .A(n10728), .ZN(n6686) );
  AND2_X1 U7916 ( .A1(n8740), .A2(n6530), .ZN(n10087) );
  OAI22_X1 U7917 ( .A1(n10144), .A2(n6706), .B1(n10134), .B2(n8726), .ZN(n6705) );
  NAND2_X1 U7918 ( .A1(n8980), .A2(n8979), .ZN(n14155) );
  INV_X1 U7919 ( .A(n14526), .ZN(n14534) );
  XNOR2_X1 U7920 ( .A(n8708), .B(P1_IR_REG_30__SCAN_IN), .ZN(n8712) );
  OR2_X1 U7921 ( .A1(n14235), .A2(n14236), .ZN(n8708) );
  AND2_X1 U7922 ( .A1(n9353), .A2(n9329), .ZN(n12257) );
  XNOR2_X1 U7923 ( .A(n8710), .B(P1_IR_REG_29__SCAN_IN), .ZN(n8716) );
  NAND2_X1 U7924 ( .A1(n7321), .A2(n7320), .ZN(n9323) );
  INV_X1 U7925 ( .A(n7323), .ZN(n7320) );
  INV_X1 U7926 ( .A(n8721), .ZN(n8722) );
  NAND2_X1 U7927 ( .A1(n9070), .A2(n7059), .ZN(n9133) );
  AND2_X1 U7928 ( .A1(n7061), .A2(n7060), .ZN(n7059) );
  INV_X1 U7929 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n7060) );
  NOR2_X1 U7930 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n9128) );
  INV_X1 U7931 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9127) );
  NAND2_X1 U7932 ( .A1(n6799), .A2(SI_24_), .ZN(n6807) );
  NAND2_X1 U7933 ( .A1(n6811), .A2(n6810), .ZN(n6809) );
  NAND2_X1 U7934 ( .A1(n8116), .A2(n8115), .ZN(n8118) );
  NAND2_X1 U7935 ( .A1(n6775), .A2(n8114), .ZN(n8117) );
  NAND2_X1 U7936 ( .A1(n9066), .A2(n9151), .ZN(n9167) );
  MUX2_X1 U7937 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9063), .S(
        P1_IR_REG_22__SCAN_IN), .Z(n9066) );
  NAND2_X1 U7938 ( .A1(n9070), .A2(n9062), .ZN(n6728) );
  AND2_X1 U7939 ( .A1(n8503), .A2(n8502), .ZN(n11148) );
  NAND2_X1 U7940 ( .A1(n7333), .A2(n8108), .ZN(n8501) );
  NAND2_X1 U7941 ( .A1(n6717), .A2(n8097), .ZN(n6716) );
  AND2_X1 U7942 ( .A1(n8097), .A2(SI_18_), .ZN(n7296) );
  OR2_X1 U7943 ( .A1(n8347), .A2(n6792), .ZN(n6787) );
  XNOR2_X1 U7944 ( .A(n8052), .B(SI_3_), .ZN(n8223) );
  XNOR2_X1 U7945 ( .A(n9732), .B(n6752), .ZN(n9735) );
  INV_X1 U7946 ( .A(n9733), .ZN(n6752) );
  NAND2_X1 U7947 ( .A1(n9677), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n6888) );
  XNOR2_X1 U7948 ( .A(n9740), .B(n6642), .ZN(n9742) );
  INV_X1 U7949 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6642) );
  NAND2_X1 U7950 ( .A1(n6749), .A2(n14435), .ZN(n9765) );
  OAI21_X1 U7951 ( .B1(n14437), .B2(n14436), .A(n6750), .ZN(n6749) );
  INV_X1 U7952 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n6750) );
  NOR2_X1 U7953 ( .A1(n9721), .A2(n9720), .ZN(n9713) );
  OAI21_X1 U7954 ( .B1(n14287), .B2(n14286), .A(n6747), .ZN(n6746) );
  INV_X1 U7955 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n6747) );
  NOR2_X1 U7956 ( .A1(n12556), .A2(n12555), .ZN(n12557) );
  AND4_X1 U7957 ( .A1(n7814), .A2(n7813), .A3(n7812), .A4(n7811), .ZN(n12955)
         );
  AND2_X1 U7958 ( .A1(n12556), .A2(n12555), .ZN(n12558) );
  AND4_X1 U7959 ( .A1(n7626), .A2(n7625), .A3(n7624), .A4(n7623), .ZN(n11354)
         );
  AND3_X1 U7960 ( .A1(n7602), .A2(n7601), .A3(n7600), .ZN(n15020) );
  NAND2_X1 U7961 ( .A1(n7806), .A2(n7805), .ZN(n12943) );
  AND4_X1 U7962 ( .A1(n7700), .A2(n7699), .A3(n7698), .A4(n7697), .ZN(n14340)
         );
  AND2_X1 U7963 ( .A1(n10030), .A2(n10029), .ZN(n12670) );
  AOI21_X1 U7964 ( .B1(n12333), .B2(n7390), .A(n12332), .ZN(n12335) );
  NAND4_X1 U7965 ( .A1(n7516), .A2(n7515), .A3(n7514), .A4(n7513), .ZN(n12693)
         );
  XNOR2_X1 U7966 ( .A(n6890), .B(n11803), .ZN(n11619) );
  NOR2_X1 U7967 ( .A1(n11619), .A2(n7512), .ZN(n11799) );
  NOR2_X1 U7968 ( .A1(n11801), .A2(n11800), .ZN(n12703) );
  XNOR2_X1 U7969 ( .A(n12722), .B(n12736), .ZN(n12704) );
  AOI21_X1 U7970 ( .B1(n9442), .B2(n15060), .A(n9441), .ZN(n12554) );
  OAI21_X1 U7971 ( .B1(n12853), .B2(n11829), .A(n8032), .ZN(n8033) );
  OR2_X1 U7972 ( .A1(n9431), .A2(n11887), .ZN(n7888) );
  OAI21_X1 U7973 ( .B1(n8006), .B2(n15045), .A(n8005), .ZN(n12859) );
  INV_X1 U7974 ( .A(n7949), .ZN(n12862) );
  NAND2_X1 U7975 ( .A1(n13587), .A2(n9460), .ZN(n6786) );
  NAND2_X1 U7976 ( .A1(n8526), .A2(n8525), .ZN(n13514) );
  NOR2_X1 U7977 ( .A1(n7146), .A2(n13267), .ZN(n7144) );
  NOR2_X1 U7978 ( .A1(n7151), .A2(n7148), .ZN(n7146) );
  NOR2_X1 U7979 ( .A1(n12211), .A2(n7149), .ZN(n7148) );
  INV_X1 U7980 ( .A(n7156), .ZN(n7149) );
  NAND2_X1 U7981 ( .A1(n7150), .A2(n7153), .ZN(n7147) );
  NAND2_X1 U7982 ( .A1(n8312), .A2(n8311), .ZN(n11154) );
  NAND2_X1 U7983 ( .A1(n8367), .A2(n8366), .ZN(n11443) );
  XNOR2_X1 U7984 ( .A(n12185), .B(n12183), .ZN(n13233) );
  INV_X1 U7985 ( .A(n12184), .ZN(n12183) );
  NAND2_X1 U7986 ( .A1(n8351), .A2(n8350), .ZN(n11382) );
  NAND2_X1 U7987 ( .A1(n8273), .A2(n8272), .ZN(n10911) );
  NAND2_X1 U7988 ( .A1(n8562), .A2(n8561), .ZN(n13497) );
  NAND2_X1 U7989 ( .A1(n10477), .A2(n14724), .ZN(n13262) );
  NAND2_X1 U7990 ( .A1(n14679), .A2(n14678), .ZN(n14677) );
  NAND2_X1 U7991 ( .A1(n9459), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n7275) );
  NAND2_X1 U7992 ( .A1(n12219), .A2(n9460), .ZN(n7276) );
  OAI22_X1 U7993 ( .A1(n8225), .A2(n10145), .B1(n10196), .B2(n10217), .ZN(
        n6870) );
  NOR2_X1 U7994 ( .A1(n8206), .A2(n10144), .ZN(n6869) );
  OR2_X1 U7995 ( .A1(n14743), .A2(n10844), .ZN(n14724) );
  NAND2_X2 U7996 ( .A1(n8891), .A2(n8890), .ZN(n14419) );
  NAND2_X1 U7997 ( .A1(n14407), .A2(n12014), .ZN(n13642) );
  NAND2_X1 U7998 ( .A1(n6743), .A2(n12137), .ZN(n6742) );
  NAND2_X1 U7999 ( .A1(n13680), .A2(n6537), .ZN(n6743) );
  NAND2_X1 U8000 ( .A1(n13643), .A2(n12020), .ZN(n13693) );
  OAI21_X1 U8001 ( .B1(n13881), .B2(n13880), .A(n6770), .ZN(n6769) );
  AOI21_X1 U8002 ( .B1(n13882), .B2(n13883), .A(n14465), .ZN(n6770) );
  XNOR2_X1 U8003 ( .A(n13895), .B(n6815), .ZN(n13887) );
  NAND2_X2 U8004 ( .A1(n10181), .A2(n10112), .ZN(n14477) );
  NAND2_X1 U8005 ( .A1(n9039), .A2(n9038), .ZN(n14203) );
  INV_X1 U8006 ( .A(n14560), .ZN(n14558) );
  NAND2_X1 U8007 ( .A1(n12296), .A2(n8774), .ZN(n9049) );
  NAND2_X1 U8008 ( .A1(n14203), .A2(n9158), .ZN(n6681) );
  NAND2_X1 U8009 ( .A1(n14115), .A2(n6682), .ZN(n14202) );
  AND2_X1 U8010 ( .A1(n14114), .A2(n14113), .ZN(n6682) );
  XNOR2_X1 U8011 ( .A(n9735), .B(n10200), .ZN(n15147) );
  XNOR2_X1 U8012 ( .A(n6748), .B(n9765), .ZN(n14440) );
  INV_X1 U8013 ( .A(n9766), .ZN(n6748) );
  NAND2_X1 U8014 ( .A1(n14440), .A2(n14648), .ZN(n14439) );
  OAI21_X1 U8015 ( .B1(n14446), .B2(n14447), .A(n6873), .ZN(n6872) );
  INV_X1 U8016 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n6873) );
  NAND2_X1 U8017 ( .A1(n14260), .A2(n14259), .ZN(n14258) );
  INV_X1 U8018 ( .A(n7338), .ZN(n7334) );
  NAND2_X1 U8019 ( .A1(n7337), .A2(n7335), .ZN(n9201) );
  NOR2_X1 U8020 ( .A1(n7338), .A2(n7336), .ZN(n7335) );
  NAND2_X1 U8021 ( .A1(n9497), .A2(n9499), .ZN(n7216) );
  OR2_X1 U8022 ( .A1(n7222), .A2(n9509), .ZN(n7221) );
  INV_X1 U8023 ( .A(n9508), .ZN(n7222) );
  NAND2_X1 U8024 ( .A1(n9224), .A2(n7314), .ZN(n7313) );
  INV_X1 U8025 ( .A(n9223), .ZN(n7314) );
  OR2_X1 U8026 ( .A1(n7225), .A2(n9520), .ZN(n7224) );
  INV_X1 U8027 ( .A(n9519), .ZN(n7225) );
  AOI21_X1 U8028 ( .B1(n7310), .B2(n7309), .A(n6547), .ZN(n7307) );
  NOR2_X1 U8029 ( .A1(n7308), .A2(n9369), .ZN(n7306) );
  NOR2_X1 U8030 ( .A1(n7308), .A2(n9259), .ZN(n7305) );
  NOR2_X1 U8031 ( .A1(n9533), .A2(n7212), .ZN(n7213) );
  NAND2_X1 U8032 ( .A1(n7212), .A2(n9533), .ZN(n7211) );
  NAND2_X1 U8033 ( .A1(n7213), .A2(n7211), .ZN(n7210) );
  INV_X1 U8034 ( .A(n9267), .ZN(n7327) );
  NAND2_X1 U8035 ( .A1(n7198), .A2(n7197), .ZN(n9547) );
  NAND2_X1 U8036 ( .A1(n9542), .A2(n9544), .ZN(n7197) );
  NAND2_X1 U8037 ( .A1(n9553), .A2(n9555), .ZN(n7200) );
  OR2_X1 U8038 ( .A1(n9280), .A2(n9281), .ZN(n7341) );
  NAND2_X1 U8039 ( .A1(n9576), .A2(n9578), .ZN(n7202) );
  NAND2_X1 U8040 ( .A1(n7281), .A2(n9307), .ZN(n7280) );
  INV_X1 U8041 ( .A(n9306), .ZN(n7281) );
  NAND2_X1 U8042 ( .A1(n7203), .A2(n7206), .ZN(n9589) );
  NAND2_X1 U8043 ( .A1(n7207), .A2(n9585), .ZN(n7206) );
  INV_X1 U8044 ( .A(n7186), .ZN(n7185) );
  MUX2_X1 U8045 ( .A(n14203), .B(n13748), .S(n9176), .Z(n9311) );
  INV_X1 U8046 ( .A(n8085), .ZN(n7290) );
  INV_X1 U8047 ( .A(n8092), .ZN(n7295) );
  NAND2_X1 U8048 ( .A1(n15064), .A2(n15051), .ZN(n12351) );
  OR2_X1 U8049 ( .A1(n12696), .A2(n11360), .ZN(n7246) );
  NAND2_X1 U8050 ( .A1(n7245), .A2(n7244), .ZN(n7243) );
  INV_X1 U8051 ( .A(n11353), .ZN(n7245) );
  INV_X1 U8052 ( .A(n13906), .ZN(n9396) );
  XNOR2_X1 U8053 ( .A(n9168), .B(n9167), .ZN(n9341) );
  NOR2_X1 U8054 ( .A1(n6500), .A2(n6543), .ZN(n6643) );
  NOR2_X1 U8055 ( .A1(n8906), .A2(n8905), .ZN(n8919) );
  AND2_X1 U8056 ( .A1(n8705), .A2(n8704), .ZN(n9122) );
  INV_X1 U8057 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7269) );
  INV_X1 U8058 ( .A(n8428), .ZN(n7293) );
  INV_X1 U8059 ( .A(n8088), .ZN(n7294) );
  INV_X1 U8060 ( .A(n6558), .ZN(n6778) );
  NOR2_X1 U8061 ( .A1(n7778), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n7779) );
  NAND2_X1 U8062 ( .A1(n14881), .A2(n6532), .ZN(n11671) );
  NAND2_X1 U8063 ( .A1(n12757), .A2(n12755), .ZN(n12794) );
  NAND2_X1 U8064 ( .A1(n12788), .A2(n12810), .ZN(n6921) );
  OR2_X1 U8065 ( .A1(n7949), .A2(n7948), .ZN(n12467) );
  INV_X1 U8066 ( .A(n12452), .ZN(n6832) );
  OR2_X1 U8067 ( .A1(n7807), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n7809) );
  INV_X1 U8068 ( .A(n12382), .ZN(n6848) );
  AOI21_X1 U8069 ( .B1(n6845), .B2(n6849), .A(n6844), .ZN(n6843) );
  INV_X1 U8070 ( .A(n12503), .ZN(n6845) );
  INV_X1 U8071 ( .A(n6847), .ZN(n6846) );
  OAI21_X1 U8072 ( .B1(n12503), .B2(n6848), .A(n12387), .ZN(n6847) );
  NAND2_X1 U8073 ( .A1(n12351), .A2(n12346), .ZN(n7935) );
  NAND2_X1 U8074 ( .A1(n7243), .A2(n7241), .ZN(n11567) );
  NOR2_X1 U8075 ( .A1(n10168), .A2(n7994), .ZN(n8013) );
  NOR2_X1 U8076 ( .A1(n7898), .A2(n6965), .ZN(n6964) );
  INV_X1 U8077 ( .A(n7886), .ZN(n6965) );
  AND2_X1 U8078 ( .A1(n7459), .A2(n7463), .ZN(n7265) );
  NOR2_X1 U8079 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), .ZN(
        n7455) );
  INV_X1 U8080 ( .A(n6935), .ZN(n6934) );
  OAI21_X1 U8081 ( .B1(n7757), .B2(n6936), .A(n7436), .ZN(n6935) );
  INV_X1 U8082 ( .A(n7434), .ZN(n6936) );
  NOR2_X2 U8084 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n7577) );
  INV_X1 U8085 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7447) );
  AOI21_X1 U8086 ( .B1(n13170), .B2(n7180), .A(n13224), .ZN(n7179) );
  AOI22_X1 U8087 ( .A1(n7186), .A2(n7189), .B1(n7190), .B2(n7195), .ZN(n7182)
         );
  AND2_X1 U8088 ( .A1(n9616), .A2(n9615), .ZN(n9617) );
  AND2_X1 U8089 ( .A1(n8166), .A2(n8165), .ZN(n12212) );
  INV_X1 U8090 ( .A(n13355), .ZN(n7098) );
  NOR2_X1 U8091 ( .A1(n8463), .A2(n13314), .ZN(n8462) );
  NAND2_X1 U8092 ( .A1(n6887), .A2(n6886), .ZN(n11715) );
  AND2_X1 U8093 ( .A1(n8339), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8352) );
  NOR2_X1 U8094 ( .A1(n8340), .A2(n11167), .ZN(n8339) );
  AOI21_X1 U8095 ( .B1(n6981), .B2(n6983), .A(n6539), .ZN(n6978) );
  INV_X1 U8096 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7131) );
  OR2_X1 U8097 ( .A1(n8335), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n8348) );
  OR2_X1 U8098 ( .A1(n8364), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n8307) );
  AOI21_X1 U8099 ( .B1(n7042), .B2(n7040), .A(n11835), .ZN(n7039) );
  INV_X1 U8100 ( .A(n7042), .ZN(n7041) );
  INV_X1 U8101 ( .A(n11600), .ZN(n7040) );
  AND2_X1 U8102 ( .A1(n12055), .A2(n6582), .ZN(n7058) );
  INV_X1 U8103 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8905) );
  NAND2_X1 U8104 ( .A1(n11694), .A2(n6766), .ZN(n11696) );
  OR2_X1 U8105 ( .A1(n11695), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6766) );
  AND2_X1 U8106 ( .A1(n6665), .A2(n9090), .ZN(n6659) );
  INV_X1 U8107 ( .A(n8900), .ZN(n7078) );
  NAND2_X1 U8108 ( .A1(n7347), .A2(n9087), .ZN(n7346) );
  INV_X1 U8109 ( .A(n9085), .ZN(n7344) );
  INV_X1 U8110 ( .A(n6673), .ZN(n6672) );
  NOR2_X1 U8111 ( .A1(n8587), .A2(n7319), .ZN(n7318) );
  INV_X1 U8112 ( .A(n8126), .ZN(n7319) );
  NOR2_X1 U8113 ( .A1(n8586), .A2(SI_28_), .ZN(n7323) );
  AOI21_X1 U8114 ( .B1(n6800), .B2(n6802), .A(n6603), .ZN(n6798) );
  NAND2_X1 U8115 ( .A1(n8109), .A2(SI_21_), .ZN(n8111) );
  INV_X1 U8116 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n8696) );
  INV_X1 U8117 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n8701) );
  INV_X1 U8118 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8915) );
  XNOR2_X1 U8119 ( .A(n8393), .B(SI_14_), .ZN(n8410) );
  INV_X1 U8120 ( .A(n6794), .ZN(n6792) );
  INV_X1 U8121 ( .A(n8083), .ZN(n6790) );
  INV_X1 U8122 ( .A(n8079), .ZN(n6791) );
  OR2_X1 U8123 ( .A1(n8848), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n8861) );
  INV_X1 U8124 ( .A(n7285), .ZN(n6776) );
  CLKBUF_X1 U8125 ( .A(n8813), .Z(n8814) );
  OAI21_X1 U8126 ( .B1(n6475), .B2(n10129), .A(n8051), .ZN(n8052) );
  OAI21_X1 U8127 ( .B1(n8043), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n8040), .ZN(
        n8041) );
  INV_X1 U8128 ( .A(n9730), .ZN(n9680) );
  INV_X1 U8129 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n9683) );
  XNOR2_X1 U8130 ( .A(n9686), .B(n9687), .ZN(n9728) );
  INV_X1 U8131 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n9697) );
  AOI21_X1 U8132 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n9701), .A(n9700), .ZN(
        n9727) );
  NOR2_X1 U8133 ( .A1(n7620), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7640) );
  NAND2_X1 U8134 ( .A1(n9979), .A2(n12387), .ZN(n7035) );
  NAND2_X1 U8135 ( .A1(n7015), .A2(n10011), .ZN(n7014) );
  NAND2_X1 U8136 ( .A1(n7018), .A2(n7020), .ZN(n7015) );
  INV_X1 U8137 ( .A(n12607), .ZN(n9997) );
  OR2_X1 U8138 ( .A1(n7765), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n7778) );
  NAND2_X1 U8139 ( .A1(n7038), .A2(n12696), .ZN(n7037) );
  NOR2_X1 U8140 ( .A1(n12574), .A2(n12687), .ZN(n7022) );
  INV_X1 U8141 ( .A(n7021), .ZN(n7020) );
  NOR2_X1 U8142 ( .A1(n7693), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7720) );
  NAND2_X1 U8143 ( .A1(n15067), .A2(n12345), .ZN(n10522) );
  AOI21_X1 U8144 ( .B1(n7009), .B2(n7008), .A(n7006), .ZN(n7005) );
  INV_X1 U8145 ( .A(n10988), .ZN(n7006) );
  INV_X1 U8146 ( .A(n7008), .ZN(n7007) );
  NAND2_X1 U8147 ( .A1(n7863), .A2(n9925), .ZN(n7891) );
  INV_X1 U8148 ( .A(n7864), .ZN(n7863) );
  NAND2_X1 U8149 ( .A1(n7751), .A2(n7750), .ZN(n7765) );
  INV_X1 U8150 ( .A(n12502), .ZN(n12528) );
  AOI21_X1 U8151 ( .B1(n10509), .B2(n10358), .A(n10357), .ZN(n10501) );
  AOI21_X1 U8152 ( .B1(n14858), .B2(n14857), .A(n14856), .ZN(n14874) );
  XNOR2_X1 U8153 ( .A(n11671), .B(n11672), .ZN(n14899) );
  AOI21_X1 U8154 ( .B1(n14892), .B2(n14891), .A(n14890), .ZN(n14909) );
  OR2_X1 U8155 ( .A1(n14905), .A2(n11632), .ZN(n6904) );
  OR2_X1 U8156 ( .A1(n14889), .A2(n11632), .ZN(n6906) );
  NOR2_X1 U8157 ( .A1(n14904), .A2(n11611), .ZN(n11613) );
  AOI21_X1 U8158 ( .B1(n14927), .B2(n14926), .A(n14925), .ZN(n14943) );
  INV_X1 U8159 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n11273) );
  OR2_X1 U8160 ( .A1(n14924), .A2(n11642), .ZN(n6900) );
  NAND2_X1 U8161 ( .A1(n14950), .A2(n6585), .ZN(n11678) );
  AOI21_X1 U8162 ( .B1(n14961), .B2(n14960), .A(n14959), .ZN(n14984) );
  NOR2_X1 U8163 ( .A1(n11617), .A2(n14957), .ZN(n14990) );
  NAND2_X1 U8164 ( .A1(n11806), .A2(n11807), .ZN(n12705) );
  NAND2_X1 U8165 ( .A1(n12705), .A2(n6624), .ZN(n12726) );
  NAND2_X1 U8166 ( .A1(n12708), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n6624) );
  NOR2_X1 U8167 ( .A1(n12762), .A2(n12761), .ZN(n12773) );
  NOR2_X1 U8168 ( .A1(n7745), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n7761) );
  AND3_X1 U8169 ( .A1(n6909), .A2(n6907), .A3(n6614), .ZN(n12785) );
  NAND2_X1 U8170 ( .A1(n12821), .A2(n6916), .ZN(n6915) );
  INV_X1 U8171 ( .A(n6921), .ZN(n6916) );
  AOI21_X1 U8172 ( .B1(n12778), .B2(n12798), .A(n14316), .ZN(n12825) );
  NAND2_X1 U8173 ( .A1(n6921), .A2(n12819), .ZN(n6920) );
  NAND2_X1 U8174 ( .A1(n9433), .A2(n9432), .ZN(n9445) );
  AOI21_X1 U8175 ( .B1(n7260), .B2(n7262), .A(n7259), .ZN(n7258) );
  INV_X1 U8176 ( .A(n8002), .ZN(n7259) );
  AND2_X1 U8177 ( .A1(n12467), .A2(n12475), .ZN(n12525) );
  INV_X1 U8178 ( .A(n12868), .ZN(n12873) );
  NAND2_X1 U8179 ( .A1(n7834), .A2(n9893), .ZN(n7849) );
  OR2_X1 U8180 ( .A1(n7849), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n7864) );
  INV_X1 U8181 ( .A(n7226), .ZN(n12925) );
  AOI21_X1 U8182 ( .B1(n12937), .B2(n7228), .A(n7233), .ZN(n7227) );
  NAND2_X1 U8183 ( .A1(n12937), .A2(n7230), .ZN(n7229) );
  NAND2_X1 U8184 ( .A1(n6858), .A2(n6856), .ZN(n13004) );
  AOI21_X1 U8185 ( .B1(n6493), .B2(n6862), .A(n6857), .ZN(n6856) );
  INV_X1 U8186 ( .A(n12412), .ZN(n6857) );
  NAND2_X1 U8187 ( .A1(n7692), .A2(n7691), .ZN(n11823) );
  OR2_X1 U8188 ( .A1(n7672), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7674) );
  OR2_X1 U8189 ( .A1(n7674), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7693) );
  AND2_X1 U8190 ( .A1(n12397), .A2(n12402), .ZN(n14337) );
  AND2_X1 U8191 ( .A1(n7640), .A2(n11273), .ZN(n7656) );
  NAND2_X1 U8192 ( .A1(n7656), .A2(n7655), .ZN(n7672) );
  OR2_X1 U8193 ( .A1(n7606), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7620) );
  INV_X1 U8194 ( .A(n12509), .ZN(n7570) );
  AND2_X1 U8195 ( .A1(n7528), .A2(n6553), .ZN(n6644) );
  OR2_X1 U8196 ( .A1(n7804), .A2(n10150), .ZN(n7527) );
  INV_X1 U8197 ( .A(n11829), .ZN(n15070) );
  NOR2_X1 U8198 ( .A1(n12541), .A2(n15115), .ZN(n10664) );
  OAI211_X1 U8199 ( .C1(n13123), .C2(n10663), .A(n10662), .B(n10661), .ZN(
        n10665) );
  INV_X1 U8200 ( .A(n12818), .ZN(n12334) );
  OR2_X1 U8201 ( .A1(n15073), .A2(n12543), .ZN(n15116) );
  NAND2_X1 U8202 ( .A1(n11352), .A2(n12382), .ZN(n11566) );
  NAND2_X1 U8203 ( .A1(n7960), .A2(n12342), .ZN(n15115) );
  INV_X1 U8204 ( .A(n15115), .ZN(n15071) );
  INV_X1 U8205 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7264) );
  NAND2_X1 U8206 ( .A1(n9430), .A2(n9429), .ZN(n12300) );
  OR2_X1 U8207 ( .A1(n9427), .A2(n9426), .ZN(n9430) );
  NAND2_X1 U8208 ( .A1(n7874), .A2(n7873), .ZN(n7884) );
  XNOR2_X1 U8209 ( .A(n7973), .B(P3_IR_REG_26__SCAN_IN), .ZN(n7983) );
  NAND2_X1 U8210 ( .A1(n7859), .A2(n6617), .ZN(n7872) );
  OAI21_X1 U8211 ( .B1(n7846), .B2(P1_DATAO_REG_24__SCAN_IN), .A(n6952), .ZN(
        n6617) );
  INV_X1 U8212 ( .A(n6953), .ZN(n6952) );
  OAI21_X1 U8213 ( .B1(n7845), .B2(P1_DATAO_REG_24__SCAN_IN), .A(n11940), .ZN(
        n6953) );
  INV_X1 U8214 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n7979) );
  OAI21_X1 U8215 ( .B1(n7978), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7980) );
  NAND2_X1 U8216 ( .A1(n7915), .A2(n7913), .ZN(n7978) );
  AND2_X1 U8217 ( .A1(n7815), .A2(n7443), .ZN(n7444) );
  INV_X1 U8218 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n7919) );
  AND2_X1 U8219 ( .A1(n6948), .A2(n11149), .ZN(n6944) );
  AND2_X1 U8220 ( .A1(n7441), .A2(n7440), .ZN(n7491) );
  INV_X1 U8221 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n7497) );
  NAND2_X1 U8222 ( .A1(n6933), .A2(n6931), .ZN(n7786) );
  AOI21_X1 U8223 ( .B1(n6934), .B2(n6936), .A(n6932), .ZN(n6931) );
  NAND2_X1 U8224 ( .A1(n7758), .A2(n6934), .ZN(n6933) );
  INV_X1 U8225 ( .A(n7437), .ZN(n6932) );
  AND2_X1 U8226 ( .A1(n7439), .A2(n7438), .ZN(n7785) );
  NAND2_X1 U8227 ( .A1(n7786), .A2(n7785), .ZN(n7788) );
  NAND2_X1 U8228 ( .A1(n6635), .A2(n6634), .ZN(n7745) );
  INV_X1 U8229 ( .A(n7715), .ZN(n6635) );
  AND2_X1 U8230 ( .A1(n7432), .A2(n7431), .ZN(n7741) );
  NAND2_X1 U8231 ( .A1(n7742), .A2(n7741), .ZN(n7744) );
  AND2_X1 U8232 ( .A1(n7430), .A2(n7429), .ZN(n7727) );
  NAND2_X1 U8233 ( .A1(n7728), .A2(n7727), .ZN(n7730) );
  NAND2_X1 U8234 ( .A1(n7704), .A2(n6588), .ZN(n6938) );
  NAND2_X1 U8235 ( .A1(n6942), .A2(n10401), .ZN(n6941) );
  INV_X1 U8236 ( .A(n7427), .ZN(n6942) );
  NOR2_X1 U8237 ( .A1(n6645), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n6825) );
  NAND2_X1 U8238 ( .A1(n6927), .A2(n6925), .ZN(n7702) );
  AOI21_X1 U8239 ( .B1(n6928), .B2(n6930), .A(n6926), .ZN(n6925) );
  INV_X1 U8240 ( .A(n7425), .ZN(n6926) );
  AOI21_X1 U8241 ( .B1(n7648), .B2(n6960), .A(n6959), .ZN(n6958) );
  NAND2_X1 U8242 ( .A1(n7627), .A2(n7648), .ZN(n6961) );
  INV_X1 U8243 ( .A(n7419), .ZN(n6959) );
  AND2_X1 U8244 ( .A1(n7421), .A2(n7420), .ZN(n7662) );
  NOR2_X1 U8245 ( .A1(n6645), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n7630) );
  INV_X1 U8246 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n7629) );
  AND2_X1 U8247 ( .A1(n7410), .A2(n7409), .ZN(n7594) );
  AND2_X1 U8248 ( .A1(n7407), .A2(n7406), .ZN(n7580) );
  NAND2_X1 U8249 ( .A1(n7155), .A2(n7158), .ZN(n7152) );
  NAND2_X1 U8250 ( .A1(n13195), .A2(n13194), .ZN(n13206) );
  NAND2_X1 U8251 ( .A1(n11103), .A2(n11102), .ZN(n11164) );
  INV_X1 U8252 ( .A(n11105), .ZN(n11103) );
  OR2_X1 U8253 ( .A1(n8387), .A2(n8386), .ZN(n8399) );
  AND2_X1 U8254 ( .A1(n7174), .A2(n7172), .ZN(n7171) );
  NAND2_X1 U8255 ( .A1(n12181), .A2(n7173), .ZN(n7172) );
  AOI21_X1 U8256 ( .B1(n11106), .B2(n7141), .A(n6502), .ZN(n7140) );
  AND2_X1 U8257 ( .A1(n7166), .A2(n6594), .ZN(n7164) );
  AND2_X1 U8258 ( .A1(n13194), .A2(n7169), .ZN(n7168) );
  OR2_X1 U8259 ( .A1(n10907), .A2(n10908), .ZN(n10905) );
  OR2_X1 U8260 ( .A1(n8399), .A2(n11039), .ZN(n8419) );
  AND4_X1 U8261 ( .A1(n8544), .A2(n8543), .A3(n8542), .A4(n8541), .ZN(n13187)
         );
  NAND2_X1 U8262 ( .A1(n8576), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n7087) );
  AOI21_X1 U8263 ( .B1(n14570), .B2(n10313), .A(n10312), .ZN(n10311) );
  OR2_X1 U8264 ( .A1(n8318), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n8335) );
  NOR2_X1 U8265 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n8130) );
  AND2_X1 U8266 ( .A1(n14636), .A2(n14635), .ZN(n14633) );
  AOI21_X1 U8267 ( .B1(n14388), .B2(n11035), .A(n14633), .ZN(n14651) );
  OAI21_X1 U8268 ( .B1(n12239), .B2(n12238), .A(n12237), .ZN(n12240) );
  AND2_X1 U8269 ( .A1(n8163), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8688) );
  AND2_X1 U8270 ( .A1(n8590), .A2(n8589), .ZN(n9458) );
  AND2_X1 U8271 ( .A1(n10473), .A2(n8609), .ZN(n13171) );
  NAND2_X1 U8272 ( .A1(n6718), .A2(n6719), .ZN(n13339) );
  AOI21_X1 U8273 ( .B1(n6721), .B2(n6720), .A(n6541), .ZN(n6719) );
  INV_X1 U8274 ( .A(n6517), .ZN(n6720) );
  NOR2_X1 U8275 ( .A1(n13487), .A2(n6881), .ZN(n6879) );
  INV_X1 U8276 ( .A(n13338), .ZN(n7093) );
  AND2_X1 U8277 ( .A1(n8572), .A2(n8566), .ZN(n13366) );
  NAND2_X1 U8278 ( .A1(n13392), .A2(n6518), .ZN(n13363) );
  NAND2_X1 U8279 ( .A1(n13502), .A2(n13255), .ZN(n7105) );
  AND2_X1 U8280 ( .A1(n13392), .A2(n13382), .ZN(n13378) );
  AND2_X1 U8281 ( .A1(n8540), .A2(n8547), .ZN(n13394) );
  INV_X1 U8282 ( .A(n6990), .ZN(n6989) );
  OAI21_X1 U8283 ( .B1(n6991), .B2(n8672), .A(n8674), .ZN(n6990) );
  INV_X1 U8284 ( .A(n9653), .ZN(n13424) );
  AOI21_X1 U8285 ( .B1(n7113), .B2(n7117), .A(n6504), .ZN(n7111) );
  AND2_X1 U8286 ( .A1(n8687), .A2(n6485), .ZN(n6883) );
  NAND2_X1 U8287 ( .A1(n11964), .A2(n6884), .ZN(n13467) );
  AND2_X1 U8288 ( .A1(n11964), .A2(n13543), .ZN(n13465) );
  NOR2_X1 U8289 ( .A1(n14377), .A2(n13297), .ZN(n7108) );
  INV_X1 U8290 ( .A(n6887), .ZN(n11760) );
  AOI21_X1 U8291 ( .B1(n6974), .B2(n6973), .A(n6548), .ZN(n6972) );
  INV_X1 U8292 ( .A(n8660), .ZN(n6973) );
  AND2_X1 U8293 ( .A1(n11327), .A2(n14823), .ZN(n11441) );
  NAND2_X1 U8294 ( .A1(n8360), .A2(n11305), .ZN(n11310) );
  NOR2_X1 U8295 ( .A1(n14712), .A2(n14813), .ZN(n11327) );
  NAND2_X1 U8296 ( .A1(n6878), .A2(n14805), .ZN(n14712) );
  INV_X1 U8297 ( .A(n14711), .ZN(n6878) );
  NAND2_X1 U8298 ( .A1(n6967), .A2(n6966), .ZN(n14709) );
  AOI21_X1 U8299 ( .B1(n6968), .B2(n6487), .A(n6520), .ZN(n6966) );
  OAI21_X1 U8300 ( .B1(n8283), .B2(n7091), .A(n7089), .ZN(n7092) );
  INV_X1 U8301 ( .A(n7090), .ZN(n7089) );
  NAND2_X1 U8302 ( .A1(n11152), .A2(n14797), .ZN(n14711) );
  NAND2_X1 U8303 ( .A1(n8652), .A2(n8651), .ZN(n11124) );
  NAND2_X1 U8304 ( .A1(n8232), .A2(n10861), .ZN(n10999) );
  INV_X1 U8305 ( .A(n9458), .ZN(n13482) );
  NAND2_X1 U8306 ( .A1(n8449), .A2(n8448), .ZN(n13547) );
  AND2_X1 U8307 ( .A1(n10472), .A2(n14745), .ZN(n14814) );
  INV_X1 U8308 ( .A(n14814), .ZN(n14822) );
  INV_X1 U8309 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8140) );
  NAND2_X1 U8310 ( .A1(n8157), .A2(n8156), .ZN(n8159) );
  NAND2_X1 U8311 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n8155), .ZN(n8156) );
  INV_X1 U8312 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8155) );
  XNOR2_X1 U8313 ( .A(n8628), .B(P2_IR_REG_25__SCAN_IN), .ZN(n8639) );
  OR2_X1 U8314 ( .A1(n8112), .A2(SI_22_), .ZN(n7332) );
  NAND2_X1 U8315 ( .A1(n8112), .A2(SI_22_), .ZN(n8113) );
  NAND2_X1 U8316 ( .A1(n8599), .A2(n8636), .ZN(n9669) );
  OR2_X1 U8317 ( .A1(n8227), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n8260) );
  INV_X1 U8318 ( .A(n7048), .ZN(n7047) );
  AOI21_X1 U8319 ( .B1(n7046), .B2(n7048), .A(n12271), .ZN(n7045) );
  INV_X1 U8320 ( .A(n12261), .ZN(n7046) );
  INV_X1 U8321 ( .A(n9001), .ZN(n9002) );
  INV_X1 U8322 ( .A(n10106), .ZN(n10102) );
  NAND2_X1 U8323 ( .A1(n13599), .A2(n13601), .ZN(n13600) );
  NOR2_X1 U8324 ( .A1(n13632), .A2(n7051), .ZN(n7050) );
  INV_X1 U8325 ( .A(n12082), .ZN(n7051) );
  NAND2_X1 U8326 ( .A1(n6738), .A2(n11073), .ZN(n11114) );
  INV_X1 U8327 ( .A(n11116), .ZN(n6738) );
  OR2_X1 U8328 ( .A1(n8962), .A2(n8961), .ZN(n8970) );
  NOR2_X1 U8329 ( .A1(n8866), .A2(n8865), .ZN(n8879) );
  AND2_X1 U8330 ( .A1(n13615), .A2(n12099), .ZN(n13704) );
  INV_X1 U8331 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n8852) );
  OR3_X1 U8332 ( .A1(n8854), .A2(n8853), .A3(n8852), .ZN(n8866) );
  NAND2_X1 U8333 ( .A1(n8934), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8949) );
  NAND2_X1 U8334 ( .A1(n12056), .A2(n7058), .ZN(n7057) );
  NAND2_X1 U8335 ( .A1(n6739), .A2(n7052), .ZN(n6632) );
  AND2_X1 U8336 ( .A1(n13724), .A2(n12260), .ZN(n7048) );
  AND4_X1 U8337 ( .A1(n8911), .A2(n8910), .A3(n8909), .A4(n8908), .ZN(n11523)
         );
  AND4_X1 U8338 ( .A1(n8898), .A2(n8897), .A3(n8896), .A4(n8895), .ZN(n12029)
         );
  AND4_X1 U8339 ( .A1(n8872), .A2(n8871), .A3(n8870), .A4(n8869), .ZN(n12016)
         );
  AND4_X1 U8340 ( .A1(n8859), .A2(n8858), .A3(n8857), .A4(n8856), .ZN(n12007)
         );
  INV_X1 U8341 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9678) );
  NAND2_X1 U8342 ( .A1(n6765), .A2(n6764), .ZN(n6763) );
  NAND2_X1 U8343 ( .A1(n10371), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6764) );
  NOR2_X1 U8344 ( .A1(n12144), .A2(n6761), .ZN(n10533) );
  AND2_X1 U8345 ( .A1(n10382), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6761) );
  NOR2_X1 U8346 ( .A1(n10428), .A2(n6759), .ZN(n10432) );
  AND2_X1 U8347 ( .A1(n10429), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6759) );
  NAND2_X1 U8348 ( .A1(n10432), .A2(n10431), .ZN(n10548) );
  NOR2_X1 U8349 ( .A1(n10676), .A2(n6757), .ZN(n10680) );
  AND2_X1 U8350 ( .A1(n10677), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6757) );
  NAND2_X1 U8351 ( .A1(n10680), .A2(n10679), .ZN(n10816) );
  NAND2_X1 U8352 ( .A1(n10816), .A2(n6756), .ZN(n10818) );
  OR2_X1 U8353 ( .A1(n10817), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6756) );
  NAND2_X1 U8354 ( .A1(n10818), .A2(n10819), .ZN(n11015) );
  XNOR2_X1 U8355 ( .A(n11696), .B(n14464), .ZN(n14461) );
  XOR2_X1 U8356 ( .A(n13747), .B(n9368), .Z(n13906) );
  NOR2_X1 U8357 ( .A1(n13936), .A2(n7075), .ZN(n7074) );
  INV_X1 U8358 ( .A(n9037), .ZN(n7075) );
  NAND2_X1 U8359 ( .A1(n6654), .A2(n9100), .ZN(n13947) );
  NAND2_X1 U8360 ( .A1(n13959), .A2(n13960), .ZN(n6654) );
  OAI21_X1 U8361 ( .B1(n13994), .B2(n6704), .A(n6701), .ZN(n13946) );
  AOI21_X1 U8362 ( .B1(n6702), .B2(n6703), .A(n6526), .ZN(n6701) );
  INV_X1 U8363 ( .A(n7068), .ZN(n6702) );
  AOI21_X1 U8364 ( .B1(n14028), .B2(n6512), .A(n7355), .ZN(n13978) );
  INV_X1 U8365 ( .A(n6818), .ZN(n13999) );
  NOR2_X1 U8366 ( .A1(n6821), .A2(n14083), .ZN(n6820) );
  NAND2_X1 U8367 ( .A1(n14167), .A2(n6822), .ZN(n6821) );
  NOR3_X1 U8368 ( .A1(n11854), .A2(n6823), .A3(n14083), .ZN(n14075) );
  AND2_X1 U8369 ( .A1(n9260), .A2(n9261), .ZN(n14088) );
  INV_X1 U8370 ( .A(n6700), .ZN(n6699) );
  OAI21_X1 U8371 ( .B1(n11862), .B2(n6507), .A(n6547), .ZN(n6700) );
  NOR2_X1 U8372 ( .A1(n11854), .A2(n6823), .ZN(n14077) );
  NAND2_X1 U8373 ( .A1(n11734), .A2(n7354), .ZN(n11855) );
  NOR2_X1 U8374 ( .A1(n11854), .A2(n14189), .ZN(n11924) );
  NAND2_X1 U8375 ( .A1(n9089), .A2(n9245), .ZN(n11735) );
  NAND2_X1 U8376 ( .A1(n11735), .A2(n8912), .ZN(n11734) );
  NAND2_X1 U8377 ( .A1(n11247), .A2(n11246), .ZN(n11245) );
  INV_X1 U8378 ( .A(n9379), .ZN(n11246) );
  OR2_X1 U8379 ( .A1(n6653), .A2(n6652), .ZN(n11982) );
  NOR3_X1 U8380 ( .A1(n7350), .A2(n10751), .A3(n6522), .ZN(n6652) );
  AND2_X1 U8381 ( .A1(n8733), .A2(n7067), .ZN(n10752) );
  AND2_X1 U8382 ( .A1(n9185), .A2(n9174), .ZN(n10753) );
  NAND2_X1 U8383 ( .A1(n10752), .A2(n10753), .ZN(n10751) );
  INV_X1 U8384 ( .A(n13624), .ZN(n13913) );
  OR2_X1 U8385 ( .A1(n13776), .A2(n11188), .ZN(n9371) );
  OAI21_X1 U8386 ( .B1(n10182), .B2(P1_D_REG_0__SCAN_IN), .A(n10186), .ZN(
        n10097) );
  NAND2_X1 U8387 ( .A1(n14028), .A2(n9095), .ZN(n14019) );
  INV_X1 U8388 ( .A(n7345), .ZN(n11475) );
  AOI21_X1 U8389 ( .B1(n11410), .B2(n11411), .A(n7348), .ZN(n7345) );
  AND2_X1 U8390 ( .A1(n8851), .A2(n8850), .ZN(n14426) );
  INV_X1 U8391 ( .A(n14521), .ZN(n14430) );
  NAND2_X1 U8392 ( .A1(n9118), .A2(n9157), .ZN(n14528) );
  INV_X1 U8393 ( .A(n14119), .ZN(n14493) );
  AND2_X1 U8394 ( .A1(n9167), .A2(n11251), .ZN(n9118) );
  AND2_X1 U8395 ( .A1(n10726), .A2(n14541), .ZN(n14521) );
  INV_X1 U8396 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8719) );
  XNOR2_X1 U8397 ( .A(n8588), .B(n8587), .ZN(n12296) );
  NAND2_X1 U8398 ( .A1(n8707), .A2(n9070), .ZN(n8724) );
  XNOR2_X1 U8399 ( .A(n8581), .B(n8583), .ZN(n13587) );
  OAI21_X1 U8400 ( .B1(n6811), .B2(n6804), .A(n6803), .ZN(n8554) );
  NAND2_X1 U8401 ( .A1(n6806), .A2(SI_24_), .ZN(n6803) );
  NOR2_X1 U8402 ( .A1(n6806), .A2(SI_24_), .ZN(n6804) );
  AND2_X1 U8403 ( .A1(n7332), .A2(n8113), .ZN(n8506) );
  AND2_X1 U8404 ( .A1(n9062), .A2(n7343), .ZN(n7342) );
  INV_X1 U8405 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n7343) );
  INV_X1 U8406 ( .A(n8457), .ZN(n8098) );
  NAND2_X1 U8407 ( .A1(n7291), .A2(n8092), .ZN(n8427) );
  NAND2_X1 U8408 ( .A1(n8393), .A2(n8088), .ZN(n7291) );
  OR2_X1 U8409 ( .A1(n8347), .A2(n8346), .ZN(n6793) );
  NAND2_X1 U8410 ( .A1(n7282), .A2(n7285), .ZN(n8304) );
  XNOR2_X1 U8411 ( .A(n8041), .B(SI_1_), .ZN(n8199) );
  INV_X1 U8412 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9734) );
  XNOR2_X1 U8413 ( .A(n9728), .B(n6877), .ZN(n9738) );
  INV_X1 U8414 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n6877) );
  NOR2_X1 U8415 ( .A1(n9693), .A2(n9692), .ZN(n9745) );
  NOR2_X1 U8416 ( .A1(n9706), .A2(n9705), .ZN(n9762) );
  OAI22_X1 U8417 ( .A1(n9723), .A2(n9712), .B1(P1_ADDR_REG_13__SCAN_IN), .B2(
        n9722), .ZN(n9720) );
  AOI22_X1 U8418 ( .A1(n9718), .A2(n9715), .B1(P3_ADDR_REG_15__SCAN_IN), .B2(
        n14474), .ZN(n9769) );
  AND3_X1 U8419 ( .A1(n7636), .A2(n7635), .A3(n7634), .ZN(n11233) );
  NAND2_X1 U8420 ( .A1(n7027), .A2(n7025), .ZN(n11931) );
  AND2_X1 U8421 ( .A1(n11932), .A2(n7026), .ZN(n7025) );
  NAND2_X1 U8422 ( .A1(n7029), .A2(n6583), .ZN(n7026) );
  NAND2_X1 U8423 ( .A1(n7024), .A2(n7029), .ZN(n11933) );
  OR2_X1 U8424 ( .A1(n11904), .A2(n6583), .ZN(n7024) );
  INV_X1 U8425 ( .A(n12693), .ZN(n11825) );
  NAND2_X1 U8426 ( .A1(n7036), .A2(n7032), .ZN(n11493) );
  AND2_X1 U8427 ( .A1(n11494), .A2(n7035), .ZN(n7032) );
  AND2_X1 U8428 ( .A1(n7031), .A2(n7035), .ZN(n11495) );
  AND3_X1 U8429 ( .A1(n7569), .A2(n7568), .A3(n7567), .ZN(n10795) );
  OR2_X1 U8430 ( .A1(n11141), .A2(n11354), .ZN(n9977) );
  NAND2_X1 U8431 ( .A1(n12671), .A2(n9996), .ZN(n12606) );
  NAND2_X1 U8432 ( .A1(n7764), .A2(n7763), .ZN(n12992) );
  AND4_X1 U8433 ( .A1(n7799), .A2(n7798), .A3(n7797), .A4(n7796), .ZN(n12978)
         );
  NAND2_X1 U8434 ( .A1(n11270), .A2(n7037), .ZN(n11386) );
  INV_X1 U8435 ( .A(n7016), .ZN(n12636) );
  AOI21_X1 U8436 ( .B1(n12576), .B2(n7017), .A(n7020), .ZN(n7016) );
  INV_X1 U8437 ( .A(n7022), .ZN(n7017) );
  AND2_X1 U8438 ( .A1(n7028), .A2(n6581), .ZN(n10065) );
  AND4_X1 U8439 ( .A1(n7840), .A2(n7839), .A3(n7838), .A4(n7837), .ZN(n12915)
         );
  NAND2_X1 U8440 ( .A1(n10017), .A2(n7023), .ZN(n12644) );
  NAND2_X1 U8441 ( .A1(n7819), .A2(n7818), .ZN(n12918) );
  INV_X1 U8442 ( .A(n12681), .ZN(n12648) );
  INV_X1 U8443 ( .A(n7003), .ZN(n10989) );
  AOI21_X1 U8444 ( .B1(n10888), .B2(n7004), .A(n7007), .ZN(n7003) );
  INV_X1 U8445 ( .A(n7009), .ZN(n7004) );
  AND4_X1 U8446 ( .A1(n7896), .A2(n7895), .A3(n7894), .A4(n7893), .ZN(n12666)
         );
  NAND2_X1 U8447 ( .A1(n12660), .A2(n12661), .ZN(n12659) );
  BUF_X1 U8448 ( .A(n9958), .Z(n12542) );
  AND4_X1 U8449 ( .A1(n12321), .A2(n9439), .A3(n9438), .A4(n9437), .ZN(n12494)
         );
  AND4_X1 U8450 ( .A1(n12321), .A2(n7929), .A3(n7928), .A4(n7927), .ZN(n11029)
         );
  INV_X1 U8451 ( .A(n12666), .ZN(n12683) );
  INV_X1 U8452 ( .A(n12915), .ZN(n12685) );
  INV_X1 U8453 ( .A(n12955), .ZN(n12926) );
  INV_X1 U8454 ( .A(n15041), .ZN(n12701) );
  INV_X1 U8455 ( .A(n10914), .ZN(n15064) );
  OR2_X1 U8456 ( .A1(n12314), .A2(n7532), .ZN(n7534) );
  AND2_X1 U8457 ( .A1(n7531), .A2(n7530), .ZN(n7535) );
  NOR2_X1 U8458 ( .A1(n10499), .A2(n10614), .ZN(n10498) );
  NOR2_X1 U8459 ( .A1(n14855), .A2(n11621), .ZN(n14854) );
  OAI21_X1 U8460 ( .B1(n14855), .B2(n6893), .A(n6892), .ZN(n14870) );
  NAND2_X1 U8461 ( .A1(n6894), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n6893) );
  INV_X1 U8462 ( .A(n14871), .ZN(n6894) );
  INV_X1 U8463 ( .A(n6906), .ZN(n14888) );
  NAND2_X1 U8464 ( .A1(n6903), .A2(n6901), .ZN(n14904) );
  NAND2_X1 U8465 ( .A1(n11609), .A2(n6902), .ZN(n6901) );
  OR2_X1 U8466 ( .A1(n14889), .A2(n6904), .ZN(n6903) );
  INV_X1 U8467 ( .A(n14905), .ZN(n6902) );
  AND2_X1 U8468 ( .A1(n6906), .A2(n6905), .ZN(n14906) );
  NAND2_X1 U8469 ( .A1(n6896), .A2(n6895), .ZN(n14939) );
  XNOR2_X1 U8470 ( .A(n11616), .B(n11615), .ZN(n14958) );
  NAND2_X1 U8471 ( .A1(n14977), .A2(n14978), .ZN(n14976) );
  NOR2_X1 U8472 ( .A1(n11799), .A2(n11798), .ZN(n11801) );
  INV_X1 U8473 ( .A(n6890), .ZN(n11797) );
  NOR2_X1 U8474 ( .A1(n6521), .A2(n12723), .ZN(n12725) );
  NOR2_X1 U8475 ( .A1(n12725), .A2(n12738), .ZN(n12751) );
  NAND2_X1 U8476 ( .A1(n6909), .A2(n6907), .ZN(n14302) );
  INV_X1 U8477 ( .A(n12782), .ZN(n6911) );
  AOI21_X1 U8478 ( .B1(n6923), .B2(n6914), .A(n6913), .ZN(n6919) );
  INV_X1 U8479 ( .A(n6920), .ZN(n6914) );
  XNOR2_X1 U8480 ( .A(n12305), .B(n12485), .ZN(n12551) );
  NAND2_X1 U8481 ( .A1(n7902), .A2(n7901), .ZN(n7997) );
  NAND2_X1 U8482 ( .A1(n12886), .A2(n7857), .ZN(n12869) );
  NAND2_X1 U8483 ( .A1(n7833), .A2(n7832), .ZN(n13024) );
  NAND2_X1 U8484 ( .A1(n6830), .A2(n6833), .ZN(n12917) );
  OR2_X1 U8485 ( .A1(n12942), .A2(n6838), .ZN(n6830) );
  NAND2_X1 U8486 ( .A1(n6836), .A2(n12442), .ZN(n12934) );
  OR2_X1 U8487 ( .A1(n12942), .A2(n12937), .ZN(n6836) );
  NAND2_X1 U8488 ( .A1(n7468), .A2(n7467), .ZN(n13033) );
  NAND2_X1 U8489 ( .A1(n12950), .A2(n7234), .ZN(n12938) );
  NAND2_X1 U8490 ( .A1(n7943), .A2(n12427), .ZN(n12969) );
  NAND2_X1 U8491 ( .A1(n7247), .A2(n7250), .ZN(n12987) );
  NAND2_X1 U8492 ( .A1(n14326), .A2(n7252), .ZN(n7247) );
  AOI21_X1 U8493 ( .B1(n14326), .B2(n14325), .A(n7253), .ZN(n12998) );
  NAND2_X1 U8494 ( .A1(n6859), .A2(n6860), .ZN(n14324) );
  OR2_X1 U8495 ( .A1(n11828), .A2(n6862), .ZN(n6859) );
  NAND2_X1 U8496 ( .A1(n11826), .A2(n12406), .ZN(n11910) );
  NAND2_X1 U8497 ( .A1(n15036), .A2(n15071), .ZN(n13007) );
  AND3_X1 U8498 ( .A1(n7689), .A2(n7688), .A3(n7687), .ZN(n11593) );
  NAND2_X1 U8499 ( .A1(n7235), .A2(n7239), .ZN(n11588) );
  OAI21_X1 U8500 ( .B1(n7937), .B2(n12507), .A(n6853), .ZN(n11229) );
  NAND2_X1 U8501 ( .A1(n7937), .A2(n12369), .ZN(n11253) );
  NAND2_X1 U8502 ( .A1(n7585), .A2(n7584), .ZN(n15014) );
  INV_X1 U8503 ( .A(n15073), .ZN(n15053) );
  INV_X1 U8504 ( .A(n13007), .ZN(n15004) );
  AOI22_X1 U8505 ( .A1(n13127), .A2(n12322), .B1(n12312), .B2(SI_31_), .ZN(
        n13066) );
  NAND2_X1 U8506 ( .A1(n12326), .A2(n12325), .ZN(n13068) );
  NAND2_X1 U8507 ( .A1(n12554), .A2(n6622), .ZN(n9449) );
  NAND2_X1 U8508 ( .A1(n6623), .A2(n15100), .ZN(n6622) );
  INV_X1 U8509 ( .A(n12551), .ZN(n6623) );
  INV_X1 U8510 ( .A(n12592), .ZN(n13084) );
  INV_X1 U8511 ( .A(n10005), .ZN(n13109) );
  INV_X1 U8512 ( .A(n9998), .ZN(n13113) );
  AND2_X1 U8513 ( .A1(n10339), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13125) );
  XNOR2_X1 U8514 ( .A(n12300), .B(n12298), .ZN(n13132) );
  CLKBUF_X1 U8515 ( .A(n7930), .Z(n13139) );
  NAND2_X1 U8516 ( .A1(n7970), .A2(n7972), .ZN(n11693) );
  NAND2_X1 U8517 ( .A1(n6951), .A2(n11943), .ZN(n6954) );
  INV_X1 U8518 ( .A(n12337), .ZN(n12342) );
  INV_X1 U8519 ( .A(SI_20_), .ZN(n10899) );
  INV_X1 U8520 ( .A(SI_19_), .ZN(n10689) );
  NAND2_X1 U8522 ( .A1(n7760), .A2(n7434), .ZN(n7772) );
  INV_X1 U8523 ( .A(SI_17_), .ZN(n10440) );
  INV_X1 U8524 ( .A(SI_16_), .ZN(n10369) );
  INV_X1 U8525 ( .A(SI_15_), .ZN(n10320) );
  INV_X1 U8526 ( .A(SI_12_), .ZN(n10167) );
  OAI21_X1 U8527 ( .B1(n7681), .B2(n6930), .A(n6928), .ZN(n7504) );
  NAND2_X1 U8528 ( .A1(n7683), .A2(n7423), .ZN(n7502) );
  INV_X1 U8529 ( .A(SI_11_), .ZN(n10163) );
  INV_X1 U8530 ( .A(SI_10_), .ZN(n10148) );
  XNOR2_X1 U8531 ( .A(n7684), .B(n7686), .ZN(n11665) );
  NAND2_X1 U8532 ( .A1(n6957), .A2(n6955), .ZN(n7651) );
  AOI21_X1 U8533 ( .B1(n7416), .B2(n7417), .A(n6956), .ZN(n6955) );
  OR2_X1 U8534 ( .A1(n7523), .A2(n7460), .ZN(n7552) );
  NAND2_X1 U8535 ( .A1(n7524), .A2(n7525), .ZN(n10345) );
  NAND2_X1 U8536 ( .A1(n10908), .A2(n10779), .ZN(n7135) );
  NAND2_X1 U8537 ( .A1(n10905), .A2(n10779), .ZN(n10781) );
  NAND2_X1 U8538 ( .A1(n11722), .A2(n11721), .ZN(n11725) );
  NAND2_X1 U8539 ( .A1(n11164), .A2(n11163), .ZN(n11367) );
  NOR2_X1 U8540 ( .A1(n13169), .A2(n13170), .ZN(n13168) );
  INV_X1 U8541 ( .A(n11180), .ZN(n14755) );
  OAI21_X1 U8542 ( .B1(n13169), .B2(n7178), .A(n7177), .ZN(n13179) );
  NAND2_X1 U8543 ( .A1(n7165), .A2(n7166), .ZN(n13208) );
  NAND2_X1 U8544 ( .A1(n6727), .A2(n8535), .ZN(n13507) );
  NAND2_X1 U8545 ( .A1(n11939), .A2(n9460), .ZN(n6727) );
  NOR2_X1 U8546 ( .A1(n13168), .A2(n7370), .ZN(n13226) );
  NAND2_X1 U8547 ( .A1(n8513), .A2(n8512), .ZN(n13518) );
  NAND2_X1 U8548 ( .A1(n7139), .A2(n7140), .ZN(n11375) );
  NAND2_X1 U8549 ( .A1(n7165), .A2(n7163), .ZN(n13242) );
  AND2_X1 U8550 ( .A1(n13243), .A2(n7164), .ZN(n7163) );
  AND2_X1 U8551 ( .A1(n7165), .A2(n7164), .ZN(n13244) );
  OR2_X1 U8552 ( .A1(n9639), .A2(n9638), .ZN(n9640) );
  NOR2_X1 U8553 ( .A1(n6470), .A2(n9661), .ZN(n9662) );
  INV_X1 U8554 ( .A(n13146), .ZN(n13282) );
  NAND4_X2 U8555 ( .A1(n8222), .A2(n8221), .A3(n8220), .A4(n8219), .ZN(n13307)
         );
  OR2_X1 U8556 ( .A1(n8469), .A2(n8190), .ZN(n8191) );
  AOI21_X1 U8557 ( .B1(n14593), .B2(n14592), .A(n14591), .ZN(n14596) );
  AOI21_X1 U8558 ( .B1(n10266), .B2(n10265), .A(n10264), .ZN(n10584) );
  AOI21_X1 U8559 ( .B1(n14847), .B2(n10586), .A(n14606), .ZN(n14625) );
  AND2_X1 U8560 ( .A1(n10579), .A2(n10578), .ZN(n14639) );
  OR2_X1 U8561 ( .A1(n14654), .A2(n14653), .ZN(n14655) );
  NAND2_X1 U8562 ( .A1(n14677), .A2(n6600), .ZN(n14689) );
  INV_X1 U8563 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n12256) );
  AOI22_X1 U8564 ( .A1(n12257), .A2(n9460), .B1(n9459), .B2(
        P1_DATAO_REG_30__SCAN_IN), .ZN(n13479) );
  NAND2_X1 U8565 ( .A1(n13481), .A2(n13473), .ZN(n8692) );
  NAND2_X1 U8566 ( .A1(n6722), .A2(n6721), .ZN(n13354) );
  NAND2_X1 U8567 ( .A1(n6997), .A2(n6517), .ZN(n6722) );
  NAND2_X1 U8568 ( .A1(n7099), .A2(n7103), .ZN(n13349) );
  NAND2_X1 U8569 ( .A1(n13375), .A2(n7100), .ZN(n7099) );
  INV_X1 U8570 ( .A(n6999), .ZN(n13383) );
  INV_X1 U8571 ( .A(n13507), .ZN(n13396) );
  OAI21_X1 U8572 ( .B1(n13442), .B2(n8673), .A(n8672), .ZN(n13429) );
  NAND2_X1 U8573 ( .A1(n7115), .A2(n7116), .ZN(n13444) );
  OR2_X1 U8574 ( .A1(n8471), .A2(n7117), .ZN(n7115) );
  NAND2_X1 U8575 ( .A1(n7121), .A2(n7120), .ZN(n13460) );
  OR2_X1 U8576 ( .A1(n8471), .A2(n8470), .ZN(n7121) );
  NAND2_X1 U8577 ( .A1(n7110), .A2(n8426), .ZN(n11890) );
  NAND2_X1 U8578 ( .A1(n6980), .A2(n8666), .ZN(n11714) );
  NAND2_X1 U8579 ( .A1(n8665), .A2(n6515), .ZN(n6980) );
  NAND2_X1 U8580 ( .A1(n8665), .A2(n8664), .ZN(n11764) );
  NAND2_X1 U8581 ( .A1(n6977), .A2(n8661), .ZN(n11439) );
  NAND2_X1 U8582 ( .A1(n11306), .A2(n8660), .ZN(n6977) );
  NAND2_X1 U8583 ( .A1(n7123), .A2(n8332), .ZN(n11322) );
  NAND2_X1 U8584 ( .A1(n6970), .A2(n8657), .ZN(n11151) );
  NAND2_X1 U8585 ( .A1(n6971), .A2(n6516), .ZN(n6970) );
  NAND2_X1 U8586 ( .A1(n10835), .A2(n8285), .ZN(n10879) );
  INV_X1 U8587 ( .A(n13473), .ZN(n14714) );
  INV_X1 U8588 ( .A(n13453), .ZN(n14706) );
  NAND2_X1 U8589 ( .A1(n8644), .A2(n14724), .ZN(n14733) );
  AND2_X1 U8590 ( .A1(n10444), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14741) );
  NAND2_X1 U8591 ( .A1(n8159), .A2(n7128), .ZN(n13583) );
  XNOR2_X1 U8592 ( .A(n8631), .B(P2_IR_REG_26__SCAN_IN), .ZN(n13594) );
  OAI21_X1 U8593 ( .B1(n8630), .B2(P2_IR_REG_25__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8631) );
  AND2_X1 U8594 ( .A1(n8626), .A2(n8630), .ZN(n11942) );
  INV_X1 U8595 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8604) );
  INV_X1 U8596 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10874) );
  NAND2_X1 U8597 ( .A1(n8431), .A2(n7132), .ZN(n8475) );
  INV_X1 U8598 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10672) );
  INV_X1 U8599 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10570) );
  INV_X1 U8600 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10656) );
  INV_X1 U8601 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10599) );
  INV_X1 U8602 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10322) );
  INV_X1 U8603 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10236) );
  INV_X1 U8604 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10223) );
  INV_X1 U8605 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10191) );
  INV_X1 U8606 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10174) );
  INV_X1 U8607 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10176) );
  INV_X1 U8608 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10180) );
  INV_X1 U8609 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10141) );
  INV_X1 U8610 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10139) );
  INV_X1 U8611 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10142) );
  INV_X1 U8612 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10178) );
  NAND2_X1 U8613 ( .A1(n8197), .A2(n8212), .ZN(n10217) );
  OAI21_X1 U8614 ( .B1(n12056), .B2(n6737), .A(n6735), .ZN(n13622) );
  NAND2_X1 U8615 ( .A1(n7044), .A2(n7042), .ZN(n11836) );
  NAND2_X1 U8616 ( .A1(n11599), .A2(n11600), .ZN(n7044) );
  NAND2_X1 U8617 ( .A1(n8933), .A2(n8932), .ZN(n13670) );
  NAND2_X1 U8618 ( .A1(n6733), .A2(n6734), .ZN(n13686) );
  AOI21_X1 U8619 ( .B1(n6735), .B2(n6737), .A(n6592), .ZN(n6734) );
  INV_X1 U8620 ( .A(n14426), .ZN(n14413) );
  NAND2_X1 U8621 ( .A1(n14403), .A2(n12011), .ZN(n14407) );
  INV_X1 U8622 ( .A(n13739), .ZN(n14411) );
  NAND2_X1 U8623 ( .A1(n7057), .A2(n12062), .ZN(n13714) );
  NAND2_X1 U8624 ( .A1(n9028), .A2(n9027), .ZN(n14117) );
  NAND2_X1 U8625 ( .A1(n9404), .A2(n9367), .ZN(n9412) );
  INV_X1 U8626 ( .A(n12016), .ZN(n13763) );
  INV_X1 U8627 ( .A(n12007), .ZN(n13764) );
  NAND2_X1 U8628 ( .A1(n6474), .A2(n6534), .ZN(n8735) );
  NAND2_X1 U8629 ( .A1(n13782), .A2(n13781), .ZN(n13780) );
  AND2_X1 U8630 ( .A1(n6763), .A2(n6762), .ZN(n12144) );
  INV_X1 U8631 ( .A(n12145), .ZN(n6762) );
  INV_X1 U8632 ( .A(n6763), .ZN(n12146) );
  NOR2_X1 U8633 ( .A1(n10412), .A2(n6760), .ZN(n10376) );
  AND2_X1 U8634 ( .A1(n10385), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6760) );
  NOR2_X1 U8635 ( .A1(n10376), .A2(n10375), .ZN(n10428) );
  NOR2_X1 U8636 ( .A1(n11211), .A2(n6767), .ZN(n11213) );
  AND2_X1 U8637 ( .A1(n11212), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6767) );
  NAND2_X1 U8638 ( .A1(n11213), .A2(n11214), .ZN(n11694) );
  AND2_X1 U8639 ( .A1(n10391), .A2(n6483), .ZN(n14465) );
  OAI21_X1 U8640 ( .B1(n7466), .B2(n14473), .A(n13885), .ZN(n6772) );
  AND2_X1 U8641 ( .A1(n9166), .A2(n9165), .ZN(n14106) );
  AOI21_X1 U8642 ( .B1(n9117), .B2(n14526), .A(n9116), .ZN(n13921) );
  NAND2_X1 U8643 ( .A1(n13984), .A2(n6703), .ZN(n13962) );
  AND2_X1 U8644 ( .A1(n13984), .A2(n9016), .ZN(n13964) );
  NAND2_X1 U8645 ( .A1(n13994), .A2(n9007), .ZN(n13982) );
  NAND2_X1 U8646 ( .A1(n14021), .A2(n9096), .ZN(n13993) );
  OAI21_X1 U8647 ( .B1(n14052), .B2(n6693), .A(n6489), .ZN(n14010) );
  NAND2_X1 U8648 ( .A1(n6690), .A2(n6696), .ZN(n14008) );
  NAND2_X1 U8649 ( .A1(n14052), .A2(n8977), .ZN(n14031) );
  NAND2_X1 U8650 ( .A1(n14063), .A2(n9266), .ZN(n14044) );
  NAND2_X1 U8651 ( .A1(n7084), .A2(n8967), .ZN(n14050) );
  AND2_X1 U8652 ( .A1(n14087), .A2(n9260), .ZN(n7396) );
  NAND2_X1 U8653 ( .A1(n8955), .A2(n8954), .ZN(n14062) );
  NAND2_X1 U8654 ( .A1(n6664), .A2(n7352), .ZN(n11920) );
  NAND2_X1 U8655 ( .A1(n9089), .A2(n6665), .ZN(n6664) );
  NAND2_X1 U8656 ( .A1(n11861), .A2(n8928), .ZN(n11921) );
  NAND2_X1 U8657 ( .A1(n8904), .A2(n8903), .ZN(n12041) );
  NAND2_X1 U8658 ( .A1(n11518), .A2(n8900), .ZN(n11736) );
  NAND2_X1 U8659 ( .A1(n8842), .A2(n8841), .ZN(n11883) );
  NAND2_X1 U8660 ( .A1(n6670), .A2(n6673), .ZN(n11048) );
  OAI21_X1 U8661 ( .B1(n10964), .B2(n7065), .A(n7063), .ZN(n11058) );
  NAND2_X1 U8662 ( .A1(n10962), .A2(n8826), .ZN(n11060) );
  NAND2_X1 U8663 ( .A1(n6677), .A2(n9084), .ZN(n10954) );
  NAND2_X1 U8664 ( .A1(n7080), .A2(n9372), .ZN(n11984) );
  AND2_X1 U8665 ( .A1(n10729), .A2(n11860), .ZN(n14485) );
  INV_X1 U8666 ( .A(n6656), .ZN(n6655) );
  OAI22_X1 U8667 ( .A1(n8978), .A2(n10143), .B1(n10129), .B2(n8759), .ZN(n6656) );
  INV_X1 U8668 ( .A(n14485), .ZN(n14085) );
  INV_X1 U8669 ( .A(n14482), .ZN(n14082) );
  AND2_X1 U8670 ( .A1(n11414), .A2(n10727), .ZN(n14073) );
  INV_X1 U8671 ( .A(n14073), .ZN(n14092) );
  INV_X1 U8672 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n6710) );
  NAND2_X1 U8673 ( .A1(n8878), .A2(n8877), .ZN(n12024) );
  INV_X1 U8674 ( .A(n14186), .ZN(n14163) );
  NAND2_X1 U8675 ( .A1(n9331), .A2(n9330), .ZN(n14198) );
  NAND2_X1 U8676 ( .A1(n11939), .A2(n8774), .ZN(n9009) );
  NAND2_X1 U8677 ( .A1(n8969), .A2(n8968), .ZN(n14222) );
  NAND2_X1 U8678 ( .A1(n8833), .A2(n8832), .ZN(n11851) );
  NAND2_X1 U8679 ( .A1(n8806), .A2(n8805), .ZN(n14475) );
  XNOR2_X1 U8680 ( .A(n7277), .B(n9355), .ZN(n12219) );
  NAND2_X1 U8681 ( .A1(n9353), .A2(n9352), .ZN(n7277) );
  MUX2_X1 U8682 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9134), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n9135) );
  OR2_X1 U8683 ( .A1(n9127), .A2(n14236), .ZN(n7374) );
  AND2_X1 U8684 ( .A1(n8524), .A2(n8523), .ZN(n11752) );
  INV_X1 U8685 ( .A(n9167), .ZN(n14253) );
  INV_X1 U8686 ( .A(n9070), .ZN(n9071) );
  INV_X1 U8687 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10876) );
  INV_X1 U8688 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10673) );
  INV_X1 U8689 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10571) );
  INV_X1 U8690 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10597) );
  INV_X1 U8691 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10323) );
  INV_X1 U8692 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10237) );
  INV_X1 U8693 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10221) );
  INV_X1 U8694 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10192) );
  INV_X1 U8695 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10171) );
  INV_X1 U8696 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10165) );
  INV_X1 U8697 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10152) );
  INV_X1 U8698 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10136) );
  INV_X1 U8699 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10133) );
  XNOR2_X1 U8700 ( .A(n6758), .B(n8738), .ZN(n10379) );
  NAND2_X1 U8701 ( .A1(n14256), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6758) );
  CLKBUF_X1 U8702 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n14256) );
  INV_X1 U8703 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7465) );
  NOR2_X1 U8704 ( .A1(n15146), .A2(n9736), .ZN(n14263) );
  INV_X1 U8705 ( .A(n9681), .ZN(n9731) );
  NAND2_X1 U8706 ( .A1(n14262), .A2(n6754), .ZN(n15143) );
  OAI21_X1 U8707 ( .B1(n14263), .B2(n14264), .A(n6755), .ZN(n6754) );
  INV_X1 U8708 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n6755) );
  NOR2_X1 U8709 ( .A1(n15143), .A2(n15144), .ZN(n15142) );
  XNOR2_X1 U8710 ( .A(n9738), .B(n14589), .ZN(n15133) );
  XNOR2_X1 U8711 ( .A(n6751), .B(n9741), .ZN(n15137) );
  INV_X1 U8712 ( .A(n9742), .ZN(n6751) );
  INV_X1 U8713 ( .A(n9755), .ZN(n6871) );
  NAND2_X1 U8714 ( .A1(n14278), .A2(n14277), .ZN(n14276) );
  NAND2_X1 U8715 ( .A1(n9760), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n6640) );
  NAND2_X1 U8716 ( .A1(n14439), .A2(n9767), .ZN(n14442) );
  OAI21_X1 U8717 ( .B1(n14260), .B2(n14259), .A(n6745), .ZN(n6744) );
  INV_X1 U8718 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n6745) );
  OAI21_X1 U8719 ( .B1(n12558), .B2(n12557), .A(n12670), .ZN(n12564) );
  NAND2_X1 U8720 ( .A1(n8000), .A2(n7380), .ZN(P3_U3487) );
  AND2_X1 U8721 ( .A1(n7363), .A2(n7999), .ZN(n7380) );
  AOI21_X1 U8722 ( .B1(n13076), .B2(n15131), .A(n8036), .ZN(n8037) );
  OAI22_X1 U8723 ( .A1(n13080), .A2(n13063), .B1(n15131), .B2(n8035), .ZN(
        n8036) );
  MUX2_X1 U8724 ( .A(n8021), .B(n8020), .S(n15131), .Z(n8022) );
  MUX2_X1 U8725 ( .A(n8018), .B(n8020), .S(n15120), .Z(n8019) );
  NAND2_X1 U8726 ( .A1(n7147), .A2(n13241), .ZN(n7145) );
  NAND2_X1 U8727 ( .A1(n14850), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6987) );
  NAND2_X1 U8728 ( .A1(n13563), .A2(n14853), .ZN(n6988) );
  NAND2_X1 U8729 ( .A1(n14829), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6782) );
  NAND2_X1 U8730 ( .A1(n13563), .A2(n14831), .ZN(n6783) );
  NAND2_X1 U8731 ( .A1(n6741), .A2(n6740), .ZN(P1_U3225) );
  AOI21_X1 U8732 ( .B1(n14208), .B2(n6468), .A(n12138), .ZN(n6740) );
  NAND2_X1 U8733 ( .A1(n6742), .A2(n14409), .ZN(n6741) );
  OAI211_X1 U8734 ( .C1(n13884), .C2(n14023), .A(n6771), .B(n6768), .ZN(
        P1_U3262) );
  INV_X1 U8735 ( .A(n6772), .ZN(n6771) );
  NAND2_X1 U8736 ( .A1(n6769), .A2(n14023), .ZN(n6768) );
  OAI21_X1 U8737 ( .B1(n9163), .B2(n14558), .A(n6618), .ZN(n9164) );
  NAND2_X1 U8738 ( .A1(n14558), .A2(n6619), .ZN(n6618) );
  INV_X1 U8739 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6619) );
  NAND2_X1 U8740 ( .A1(n6711), .A2(n6708), .ZN(P1_U3555) );
  AOI21_X1 U8741 ( .B1(n14203), .B2(n14163), .A(n6709), .ZN(n6708) );
  NAND2_X1 U8742 ( .A1(n14202), .A2(n14560), .ZN(n6711) );
  NOR2_X1 U8743 ( .A1(n14560), .A2(n6710), .ZN(n6709) );
  MUX2_X1 U8744 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9163), .S(n14549), .Z(n9155) );
  AOI21_X1 U8745 ( .B1(n14202), .B2(n14549), .A(n6679), .ZN(n14204) );
  NAND2_X1 U8746 ( .A1(n6681), .A2(n6680), .ZN(n6679) );
  NAND2_X1 U8747 ( .A1(n14547), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6680) );
  INV_X1 U8748 ( .A(n14259), .ZN(n6638) );
  INV_X4 U8749 ( .A(n9169), .ZN(n9176) );
  NAND2_X1 U8750 ( .A1(n7066), .A2(n10693), .ZN(n7067) );
  NOR2_X1 U8751 ( .A1(n12024), .A2(n12022), .ZN(n6484) );
  AND2_X1 U8752 ( .A1(n6884), .A2(n13454), .ZN(n6485) );
  AND4_X1 U8753 ( .A1(n12502), .A2(n12479), .A3(n12485), .A4(n6501), .ZN(n6486) );
  AND2_X2 U8754 ( .A1(n9475), .A2(n10447), .ZN(n9472) );
  AND2_X1 U8755 ( .A1(n6969), .A2(n8657), .ZN(n6487) );
  NOR2_X1 U8756 ( .A1(n14203), .A2(n13748), .ZN(n6488) );
  AND2_X1 U8757 ( .A1(n14018), .A2(n6691), .ZN(n6489) );
  INV_X1 U8758 ( .A(n8270), .ZN(n7284) );
  AND2_X1 U8759 ( .A1(n12083), .A2(n7050), .ZN(n6490) );
  OR2_X1 U8760 ( .A1(n11715), .A2(n12161), .ZN(n6491) );
  INV_X1 U8761 ( .A(n13492), .ZN(n6882) );
  XNOR2_X1 U8762 ( .A(n13772), .B(n10714), .ZN(n10706) );
  AND2_X1 U8763 ( .A1(n13392), .A2(n6880), .ZN(n6492) );
  AND2_X1 U8764 ( .A1(n6860), .A2(n12413), .ZN(n6493) );
  AND2_X1 U8765 ( .A1(n9088), .A2(n7346), .ZN(n6494) );
  NAND2_X1 U8766 ( .A1(n8461), .A2(n8460), .ZN(n12171) );
  AND2_X1 U8767 ( .A1(n12695), .A2(n15003), .ZN(n6495) );
  NAND2_X1 U8768 ( .A1(n8792), .A2(n8791), .ZN(n11990) );
  INV_X1 U8769 ( .A(n11990), .ZN(n6627) );
  NAND2_X1 U8770 ( .A1(n6717), .A2(n7296), .ZN(n8472) );
  AND2_X1 U8771 ( .A1(n8430), .A2(n7134), .ZN(n6496) );
  INV_X1 U8772 ( .A(n9202), .ZN(n7336) );
  AND3_X1 U8773 ( .A1(n7519), .A2(n7517), .A3(n7520), .ZN(n6497) );
  INV_X1 U8774 ( .A(n12049), .ZN(n14189) );
  AND2_X1 U8775 ( .A1(n8918), .A2(n8917), .ZN(n12049) );
  AND2_X1 U8776 ( .A1(n8148), .A2(n8147), .ZN(n13341) );
  INV_X1 U8777 ( .A(n13341), .ZN(n13487) );
  INV_X1 U8778 ( .A(n7370), .ZN(n7180) );
  AND2_X1 U8779 ( .A1(n8067), .A2(SI_8_), .ZN(n6498) );
  OR2_X1 U8780 ( .A1(n7050), .A2(n6732), .ZN(n6499) );
  AND2_X1 U8781 ( .A1(n9321), .A2(n7297), .ZN(n6500) );
  INV_X1 U8782 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8145) );
  AND4_X1 U8783 ( .A1(n12526), .A2(n12525), .A3(n12524), .A4(n12873), .ZN(
        n6501) );
  NOR2_X1 U8784 ( .A1(n11365), .A2(n11364), .ZN(n6502) );
  INV_X1 U8785 ( .A(n9993), .ZN(n13122) );
  AND2_X1 U8786 ( .A1(n13704), .A2(n6499), .ZN(n6503) );
  AND2_X1 U8787 ( .A1(n13531), .A2(n7119), .ZN(n6504) );
  AND2_X1 U8788 ( .A1(n8556), .A2(n8555), .ZN(n13382) );
  NAND2_X1 U8789 ( .A1(n6556), .A2(n7120), .ZN(n6505) );
  NAND2_X1 U8790 ( .A1(n8177), .A2(n8176), .ZN(n13526) );
  NAND2_X1 U8791 ( .A1(n11426), .A2(n11425), .ZN(n6506) );
  NAND2_X1 U8792 ( .A1(n8928), .A2(n9369), .ZN(n6507) );
  AND2_X1 U8793 ( .A1(n8507), .A2(SI_22_), .ZN(n6508) );
  INV_X1 U8794 ( .A(n8533), .ZN(n6806) );
  NAND2_X1 U8795 ( .A1(n13162), .A2(n7162), .ZN(n10636) );
  AND2_X1 U8796 ( .A1(n14249), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6509) );
  NAND2_X1 U8797 ( .A1(n10468), .A2(n10467), .ZN(n13162) );
  NAND2_X1 U8798 ( .A1(n13579), .A2(n13583), .ZN(n8469) );
  INV_X1 U8799 ( .A(n12066), .ZN(n12027) );
  NAND2_X1 U8800 ( .A1(n13653), .A2(n13654), .ZN(n12056) );
  INV_X2 U8801 ( .A(n8983), .ZN(n8768) );
  OR2_X2 U8802 ( .A1(n7773), .A2(P3_IR_REG_17__SCAN_IN), .ZN(n6510) );
  NAND2_X1 U8803 ( .A1(n8945), .A2(n8944), .ZN(n14083) );
  OR2_X1 U8804 ( .A1(n11552), .A2(n11050), .ZN(n6511) );
  AND2_X1 U8805 ( .A1(n7276), .A2(n7275), .ZN(n9634) );
  INV_X1 U8806 ( .A(n11411), .ZN(n7347) );
  INV_X1 U8807 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n14236) );
  AND2_X1 U8808 ( .A1(n13997), .A2(n7358), .ZN(n6512) );
  INV_X1 U8809 ( .A(n8287), .ZN(n7287) );
  OR2_X1 U8810 ( .A1(n14065), .A2(n14222), .ZN(n6513) );
  AND2_X1 U8811 ( .A1(n7057), .A2(n7055), .ZN(n6514) );
  NOR2_X1 U8812 ( .A1(n8667), .A2(n6984), .ZN(n6515) );
  NAND2_X1 U8813 ( .A1(n14789), .A2(n13303), .ZN(n6516) );
  NAND2_X1 U8814 ( .A1(n13497), .A2(n13284), .ZN(n6517) );
  INV_X1 U8815 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n7469) );
  AND2_X1 U8816 ( .A1(n13368), .A2(n13382), .ZN(n6518) );
  NOR2_X1 U8817 ( .A1(n12526), .A2(n8027), .ZN(n6519) );
  NAND2_X1 U8818 ( .A1(n8727), .A2(n8728), .ZN(n8760) );
  AND2_X1 U8819 ( .A1(n11154), .A2(n13302), .ZN(n6520) );
  NAND2_X1 U8820 ( .A1(n9358), .A2(n9357), .ZN(n13886) );
  INV_X1 U8821 ( .A(n6838), .ZN(n6837) );
  NAND2_X1 U8822 ( .A1(n6839), .A2(n12447), .ZN(n6838) );
  NOR2_X1 U8823 ( .A1(n12704), .A2(n7722), .ZN(n6521) );
  AND2_X1 U8824 ( .A1(n13771), .A2(n14520), .ZN(n6522) );
  NAND2_X1 U8825 ( .A1(n6793), .A2(n8079), .ZN(n8362) );
  NAND2_X1 U8826 ( .A1(n6787), .A2(n6789), .ZN(n8378) );
  NAND2_X1 U8827 ( .A1(n8321), .A2(n8320), .ZN(n14710) );
  AND4_X1 U8828 ( .A1(n8141), .A2(n8140), .A3(n8637), .A4(n8139), .ZN(n6523)
         );
  INV_X1 U8829 ( .A(n12427), .ZN(n6866) );
  INV_X1 U8830 ( .A(n12505), .ZN(n7237) );
  INV_X1 U8831 ( .A(n6995), .ZN(n10866) );
  AND2_X1 U8832 ( .A1(n12491), .A2(n12487), .ZN(n12485) );
  INV_X1 U8833 ( .A(n12695), .ZN(n12387) );
  NAND2_X1 U8834 ( .A1(n8505), .A2(n8504), .ZN(n13531) );
  INV_X1 U8835 ( .A(n12314), .ZN(n9436) );
  NAND2_X1 U8836 ( .A1(n12083), .A2(n12082), .ZN(n13631) );
  OR3_X1 U8837 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        n13142), .ZN(n6525) );
  NAND2_X1 U8838 ( .A1(n7049), .A2(n7048), .ZN(n13723) );
  AND2_X1 U8839 ( .A1(n14208), .A2(n13750), .ZN(n6526) );
  NAND2_X1 U8840 ( .A1(n13368), .A2(n13188), .ZN(n6527) );
  INV_X1 U8841 ( .A(n9596), .ZN(n7194) );
  INV_X1 U8842 ( .A(n11150), .ZN(n10111) );
  OAI21_X1 U8843 ( .B1(n12262), .B2(n7047), .A(n7045), .ZN(n13599) );
  NAND2_X1 U8844 ( .A1(n8479), .A2(n8478), .ZN(n13537) );
  AND3_X1 U8845 ( .A1(n7455), .A2(n7919), .A3(n7913), .ZN(n6528) );
  AND2_X1 U8846 ( .A1(n11851), .A2(n10955), .ZN(n6529) );
  NAND2_X1 U8847 ( .A1(n8739), .A2(n6705), .ZN(n6530) );
  OR2_X1 U8848 ( .A1(n13553), .A2(n8441), .ZN(n6531) );
  OR2_X1 U8849 ( .A1(n11670), .A2(n11626), .ZN(n6532) );
  NOR2_X1 U8850 ( .A1(n9255), .A2(n9256), .ZN(n7310) );
  NAND2_X1 U8851 ( .A1(n9597), .A2(n7194), .ZN(n7193) );
  INV_X1 U8852 ( .A(n7193), .ZN(n7188) );
  AND2_X1 U8853 ( .A1(n14218), .A2(n13634), .ZN(n6533) );
  INV_X2 U8854 ( .A(n8043), .ZN(n8726) );
  INV_X1 U8855 ( .A(n7654), .ZN(n7244) );
  NOR2_X1 U8856 ( .A1(n11366), .A2(n7142), .ZN(n7141) );
  INV_X1 U8857 ( .A(n9318), .ZN(n7300) );
  INV_X1 U8858 ( .A(n6850), .ZN(n6849) );
  NAND2_X1 U8859 ( .A1(n12382), .A2(n12695), .ZN(n6850) );
  INV_X1 U8860 ( .A(n9535), .ZN(n7212) );
  AND2_X1 U8861 ( .A1(n14244), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6534) );
  INV_X1 U8862 ( .A(n6676), .ZN(n6675) );
  NAND2_X1 U8863 ( .A1(n6511), .A2(n9084), .ZN(n6676) );
  AND2_X1 U8864 ( .A1(n9997), .A2(n9996), .ZN(n6535) );
  OR2_X1 U8865 ( .A1(n7348), .A2(n7344), .ZN(n6536) );
  INV_X1 U8866 ( .A(n7151), .ZN(n7150) );
  OAI21_X1 U8867 ( .B1(n7156), .B2(n7153), .A(n7152), .ZN(n7151) );
  AND2_X1 U8868 ( .A1(n12135), .A2(n12136), .ZN(n6537) );
  INV_X1 U8869 ( .A(n13670), .ZN(n14233) );
  AND2_X1 U8870 ( .A1(n7103), .A2(n7098), .ZN(n6538) );
  NOR2_X1 U8871 ( .A1(n12161), .A2(n13295), .ZN(n6539) );
  NOR2_X1 U8872 ( .A1(n11851), .A2(n13766), .ZN(n6540) );
  NOR2_X1 U8873 ( .A1(n6882), .A2(n6785), .ZN(n6541) );
  NOR2_X1 U8874 ( .A1(n12049), .A2(n13759), .ZN(n6542) );
  AND2_X1 U8875 ( .A1(n7300), .A2(n9316), .ZN(n6543) );
  NAND2_X1 U8876 ( .A1(n6786), .A2(n8584), .ZN(n13492) );
  OR2_X1 U8877 ( .A1(n13620), .A2(n13621), .ZN(n6544) );
  INV_X1 U8878 ( .A(n9214), .ZN(n7331) );
  AND2_X1 U8879 ( .A1(n8379), .A2(SI_13_), .ZN(n6545) );
  INV_X1 U8880 ( .A(n12457), .ZN(n12887) );
  XNOR2_X1 U8881 ( .A(n13020), .B(n6647), .ZN(n12457) );
  OR2_X1 U8882 ( .A1(n13396), .A2(n13187), .ZN(n6546) );
  INV_X1 U8883 ( .A(n9224), .ZN(n7316) );
  NAND2_X1 U8884 ( .A1(n8186), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7537) );
  NAND2_X1 U8885 ( .A1(n13670), .A2(n13758), .ZN(n6547) );
  NOR2_X1 U8886 ( .A1(n11443), .A2(n13298), .ZN(n6548) );
  NAND2_X1 U8887 ( .A1(n7337), .A2(n7334), .ZN(n6549) );
  INV_X1 U8888 ( .A(n7256), .ZN(n7253) );
  NAND2_X1 U8889 ( .A1(n9989), .A2(n12690), .ZN(n7256) );
  INV_X1 U8890 ( .A(n6881), .ZN(n6880) );
  NAND2_X1 U8891 ( .A1(n6518), .A2(n6882), .ZN(n6881) );
  AND2_X1 U8892 ( .A1(n7417), .A2(n7415), .ZN(n7627) );
  INV_X1 U8893 ( .A(n6704), .ZN(n6703) );
  NAND2_X1 U8894 ( .A1(n13963), .A2(n9016), .ZN(n6704) );
  INV_X1 U8895 ( .A(n14503), .ZN(n7066) );
  AND2_X1 U8896 ( .A1(n8065), .A2(SI_7_), .ZN(n6550) );
  NAND2_X1 U8897 ( .A1(n12992), .A2(n12689), .ZN(n6551) );
  INV_X1 U8898 ( .A(n11609), .ZN(n6905) );
  INV_X1 U8899 ( .A(n6975), .ZN(n6974) );
  OR2_X1 U8900 ( .A1(n8662), .A2(n6976), .ZN(n6975) );
  INV_X1 U8901 ( .A(n6923), .ZN(n6922) );
  NAND2_X1 U8902 ( .A1(n12789), .A2(n12810), .ZN(n6923) );
  INV_X1 U8903 ( .A(n7155), .ZN(n7154) );
  NOR2_X1 U8904 ( .A1(n12207), .A2(n12206), .ZN(n7155) );
  AND2_X1 U8905 ( .A1(n14117), .A2(n9101), .ZN(n6552) );
  INV_X1 U8906 ( .A(n9599), .ZN(n7196) );
  INV_X1 U8907 ( .A(n9390), .ZN(n14018) );
  OR2_X1 U8908 ( .A1(n10341), .A2(n10345), .ZN(n6553) );
  AND2_X1 U8909 ( .A1(n11876), .A2(n12006), .ZN(n6554) );
  AND2_X1 U8910 ( .A1(n8899), .A2(n8885), .ZN(n6555) );
  OR2_X1 U8911 ( .A1(n13537), .A2(n8486), .ZN(n6556) );
  AND2_X1 U8912 ( .A1(n13341), .A2(n13282), .ZN(n6557) );
  XOR2_X1 U8913 ( .A(n8068), .B(SI_9_), .Z(n6558) );
  AND2_X1 U8914 ( .A1(n9193), .A2(n10714), .ZN(n6559) );
  AND2_X1 U8915 ( .A1(n7135), .A2(n10780), .ZN(n6560) );
  NOR2_X1 U8916 ( .A1(n12962), .A2(n7371), .ZN(n6561) );
  AND2_X1 U8917 ( .A1(n8426), .A2(n6531), .ZN(n6562) );
  AND2_X1 U8918 ( .A1(n8118), .A2(n6800), .ZN(n6563) );
  AND2_X1 U8919 ( .A1(n11723), .A2(n11721), .ZN(n6564) );
  INV_X1 U8920 ( .A(n14064), .ZN(n14061) );
  AND2_X1 U8921 ( .A1(n9265), .A2(n9266), .ZN(n14064) );
  AND2_X1 U8922 ( .A1(n7266), .A2(n7264), .ZN(n6565) );
  AND2_X1 U8923 ( .A1(n12481), .A2(n12469), .ZN(n12479) );
  OR2_X1 U8924 ( .A1(n9544), .A2(n9542), .ZN(n6566) );
  NOR2_X1 U8925 ( .A1(n7295), .A2(n7290), .ZN(n7289) );
  AND2_X1 U8926 ( .A1(n12017), .A2(n12014), .ZN(n6567) );
  AOI21_X1 U8927 ( .B1(n7294), .B2(n8092), .A(n7293), .ZN(n7292) );
  OR2_X1 U8928 ( .A1(n9510), .A2(n9508), .ZN(n6568) );
  OR2_X1 U8929 ( .A1(n9521), .A2(n9519), .ZN(n6569) );
  AND2_X1 U8930 ( .A1(n6852), .A2(n12504), .ZN(n6570) );
  OR2_X1 U8931 ( .A1(n7331), .A2(n9213), .ZN(n6571) );
  OR2_X1 U8932 ( .A1(n9555), .A2(n9553), .ZN(n6572) );
  NAND2_X1 U8933 ( .A1(n14142), .A2(n12103), .ZN(n6573) );
  INV_X1 U8934 ( .A(n9090), .ZN(n6663) );
  AND2_X1 U8935 ( .A1(n7096), .A2(n7093), .ZN(n6574) );
  NAND2_X1 U8936 ( .A1(n9281), .A2(n9280), .ZN(n6575) );
  AND2_X1 U8937 ( .A1(n13355), .A2(n6527), .ZN(n6721) );
  AND2_X1 U8938 ( .A1(n6912), .A2(n6911), .ZN(n6576) );
  INV_X1 U8939 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7463) );
  NAND2_X1 U8940 ( .A1(n6922), .A2(n12821), .ZN(n6577) );
  NAND2_X1 U8941 ( .A1(n13492), .A2(n6785), .ZN(n6578) );
  OR2_X1 U8942 ( .A1(n7054), .A2(n11117), .ZN(n6579) );
  NAND2_X1 U8943 ( .A1(n12161), .A2(n8425), .ZN(n6580) );
  AND4_X1 U8944 ( .A1(n7856), .A2(n7855), .A3(n7854), .A4(n7853), .ZN(n12601)
         );
  INV_X1 U8945 ( .A(n12601), .ZN(n6647) );
  INV_X1 U8946 ( .A(n13886), .ZN(n6815) );
  AND3_X1 U8947 ( .A1(n7671), .A2(n7670), .A3(n7669), .ZN(n15003) );
  INV_X1 U8948 ( .A(n15003), .ZN(n6844) );
  NAND2_X1 U8949 ( .A1(n11902), .A2(n12692), .ZN(n6581) );
  INV_X1 U8950 ( .A(n13283), .ZN(n6785) );
  NAND2_X1 U8951 ( .A1(n13195), .A2(n7168), .ZN(n7165) );
  INV_X1 U8952 ( .A(n11951), .ZN(n6985) );
  OR2_X1 U8953 ( .A1(n13663), .A2(n13662), .ZN(n6582) );
  NOR2_X1 U8954 ( .A1(n8381), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n8601) );
  OR2_X1 U8955 ( .A1(n10061), .A2(n9987), .ZN(n6583) );
  NAND2_X1 U8956 ( .A1(n9086), .A2(n9085), .ZN(n11410) );
  OR2_X1 U8957 ( .A1(n11677), .A2(n11648), .ZN(n6584) );
  OR2_X1 U8958 ( .A1(n11677), .A2(n11647), .ZN(n6585) );
  INV_X1 U8959 ( .A(n13703), .ZN(n6732) );
  OR2_X1 U8960 ( .A1(n12549), .A2(n13063), .ZN(n6586) );
  OR2_X1 U8961 ( .A1(n12549), .A2(n13121), .ZN(n6587) );
  AND4_X1 U8962 ( .A1(n7490), .A2(n7489), .A3(n7488), .A4(n7487), .ZN(n12966)
         );
  AND4_X1 U8963 ( .A1(n7756), .A2(n7755), .A3(n7754), .A4(n7753), .ZN(n14329)
         );
  INV_X1 U8964 ( .A(n14329), .ZN(n7255) );
  AND2_X1 U8965 ( .A1(n7427), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n6588) );
  NAND2_X1 U8966 ( .A1(n6828), .A2(n6825), .ZN(n7713) );
  NAND2_X1 U8967 ( .A1(n8431), .A2(n8430), .ZN(n8446) );
  AND4_X1 U8968 ( .A1(n7679), .A2(n7678), .A3(n7677), .A4(n7676), .ZN(n14342)
         );
  INV_X1 U8969 ( .A(n14342), .ZN(n12694) );
  INV_X1 U8970 ( .A(n13255), .ZN(n13285) );
  AND4_X1 U8971 ( .A1(n8552), .A2(n8551), .A3(n8550), .A4(n8549), .ZN(n13255)
         );
  AND2_X1 U8972 ( .A1(n11734), .A2(n9251), .ZN(n6589) );
  INV_X1 U8973 ( .A(n9586), .ZN(n7207) );
  INV_X1 U8974 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10401) );
  NOR2_X1 U8975 ( .A1(n14083), .A2(n13757), .ZN(n6590) );
  NAND2_X1 U8976 ( .A1(n8431), .A2(n6496), .ZN(n6591) );
  NAND2_X1 U8977 ( .A1(n11964), .A2(n6485), .ZN(n6885) );
  AND2_X1 U8978 ( .A1(n12075), .A2(n12074), .ZN(n6592) );
  AND2_X1 U8979 ( .A1(n11468), .A2(n8885), .ZN(n6593) );
  NAND2_X1 U8980 ( .A1(n12170), .A2(n12169), .ZN(n6594) );
  OR2_X1 U8981 ( .A1(n7207), .A2(n9585), .ZN(n6595) );
  OR2_X1 U8982 ( .A1(n9566), .A2(n9564), .ZN(n6596) );
  OR2_X1 U8983 ( .A1(n9578), .A2(n9576), .ZN(n6597) );
  INV_X1 U8984 ( .A(n13290), .ZN(n7119) );
  INV_X1 U8985 ( .A(n12706), .ZN(n12708) );
  NAND2_X1 U8986 ( .A1(n8398), .A2(n8397), .ZN(n13557) );
  INV_X1 U8987 ( .A(n13557), .ZN(n6886) );
  INV_X1 U8988 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n6634) );
  AND2_X1 U8989 ( .A1(n12180), .A2(n12179), .ZN(n6598) );
  NAND2_X1 U8990 ( .A1(n11841), .A2(n11876), .ZN(n11842) );
  AND2_X1 U8991 ( .A1(n7441), .A2(n6950), .ZN(n6599) );
  INV_X1 U8992 ( .A(n7241), .ZN(n7240) );
  NOR2_X1 U8993 ( .A1(n7242), .A2(n12511), .ZN(n7241) );
  OR2_X1 U8994 ( .A1(n14671), .A2(n12243), .ZN(n6600) );
  INV_X1 U8995 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6876) );
  AND2_X1 U8996 ( .A1(n6970), .A2(n6487), .ZN(n6601) );
  AND2_X1 U8997 ( .A1(n7243), .A2(n7246), .ZN(n6602) );
  AND2_X1 U8998 ( .A1(n6808), .A2(n11691), .ZN(n6603) );
  AND2_X1 U8999 ( .A1(n7318), .A2(n9322), .ZN(n6604) );
  AND2_X1 U9000 ( .A1(n7385), .A2(n11114), .ZN(n6605) );
  AND2_X1 U9001 ( .A1(n7044), .A2(n7043), .ZN(n6606) );
  INV_X1 U9002 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6950) );
  AND2_X1 U9003 ( .A1(n13912), .A2(n14477), .ZN(n14491) );
  AND2_X2 U9004 ( .A1(n9162), .A2(n10700), .ZN(n14549) );
  INV_X1 U9005 ( .A(n13297), .ZN(n7107) );
  NOR2_X1 U9006 ( .A1(n10355), .A2(n10343), .ZN(n14300) );
  NAND2_X1 U9007 ( .A1(n10101), .A2(n10100), .ZN(n13731) );
  INV_X1 U9008 ( .A(n13731), .ZN(n14409) );
  AND2_X2 U9009 ( .A1(n10857), .A2(n10856), .ZN(n14853) );
  OR3_X1 U9010 ( .A1(n10476), .A2(n10473), .A3(n14814), .ZN(n13267) );
  INV_X1 U9011 ( .A(n6685), .ZN(n10734) );
  NAND2_X1 U9012 ( .A1(n9076), .A2(n9174), .ZN(n6685) );
  AND2_X1 U9013 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n7845), .ZN(n6607) );
  INV_X1 U9014 ( .A(SI_24_), .ZN(n6810) );
  AND2_X1 U9015 ( .A1(n9325), .A2(n13135), .ZN(n6608) );
  AND2_X1 U9016 ( .A1(n14246), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6609) );
  AND2_X1 U9017 ( .A1(n13162), .A2(n10469), .ZN(n6610) );
  AND2_X1 U9018 ( .A1(n6920), .A2(n6915), .ZN(n6611) );
  AND2_X1 U9019 ( .A1(n6900), .A2(n6899), .ZN(n6612) );
  OR2_X1 U9020 ( .A1(n7350), .A2(n10751), .ZN(n6613) );
  OR2_X1 U9021 ( .A1(n14289), .A2(n12784), .ZN(n6614) );
  NOR2_X1 U9022 ( .A1(n8709), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n14235) );
  NOR2_X1 U9023 ( .A1(n14854), .A2(n11607), .ZN(n6615) );
  NAND2_X1 U9024 ( .A1(n13809), .A2(n13810), .ZN(n6765) );
  INV_X1 U9025 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9677) );
  AND2_X1 U9026 ( .A1(n10077), .A2(n10188), .ZN(n10181) );
  OAI211_X1 U9027 ( .C1(n11116), .C2(n6579), .A(n6632), .B(n6506), .ZN(n11538)
         );
  AOI211_X2 U9028 ( .C1(n6467), .C2(n12831), .A(n12830), .B(n12829), .ZN(
        n12832) );
  NAND4_X1 U9029 ( .A1(n7454), .A2(n7453), .A3(n7746), .A4(n7496), .ZN(n7912)
         );
  AOI21_X2 U9030 ( .B1(n12486), .B2(n12485), .A(n12530), .ZN(n12492) );
  NAND2_X1 U9031 ( .A1(n7414), .A2(n7413), .ZN(n7628) );
  NAND2_X1 U9032 ( .A1(n7547), .A2(n7402), .ZN(n7564) );
  AOI21_X2 U9033 ( .B1(n12500), .B2(n12501), .A(n12528), .ZN(n12536) );
  NAND2_X1 U9034 ( .A1(n7663), .A2(n7662), .ZN(n7665) );
  NAND2_X1 U9035 ( .A1(n7665), .A2(n7421), .ZN(n7681) );
  NAND2_X1 U9036 ( .A1(n6620), .A2(n7289), .ZN(n6723) );
  INV_X1 U9037 ( .A(n6788), .ZN(n6620) );
  NAND2_X1 U9038 ( .A1(n6716), .A2(n10546), .ZN(n6773) );
  NAND2_X1 U9039 ( .A1(n6807), .A2(n6809), .ZN(n8534) );
  OAI21_X1 U9040 ( .B1(n13933), .B2(n13932), .A(n9103), .ZN(n13904) );
  INV_X1 U9041 ( .A(n6775), .ZN(n8116) );
  NAND3_X1 U9042 ( .A1(n8117), .A2(SI_23_), .A3(n8118), .ZN(n8524) );
  NAND2_X1 U9043 ( .A1(n7112), .A2(n7111), .ZN(n13435) );
  NAND2_X1 U9044 ( .A1(n10997), .A2(n8231), .ZN(n8647) );
  NOR2_X1 U9045 ( .A1(n13333), .A2(n6557), .ZN(n8596) );
  INV_X1 U9046 ( .A(n11947), .ZN(n8471) );
  OAI21_X2 U9047 ( .B1(n11959), .B2(n11968), .A(n6621), .ZN(n11947) );
  INV_X1 U9048 ( .A(n11756), .ZN(n8405) );
  NAND2_X1 U9049 ( .A1(n6988), .A2(n6987), .ZN(P2_U3528) );
  OAI22_X2 U9050 ( .A1(n13415), .A2(n9653), .B1(n13180), .B2(n13518), .ZN(
        n13404) );
  INV_X2 U9051 ( .A(n10406), .ZN(n15042) );
  NAND2_X2 U9052 ( .A1(n7518), .A2(n6497), .ZN(n10406) );
  NAND2_X2 U9053 ( .A1(n12900), .A2(n7841), .ZN(n12888) );
  OAI21_X1 U9054 ( .B1(n13033), .B2(n12686), .A(n12924), .ZN(n12913) );
  NAND2_X1 U9055 ( .A1(n14933), .A2(n11676), .ZN(n14952) );
  XOR2_X1 U9056 ( .A(n12795), .B(n12794), .Z(n12756) );
  NOR2_X1 U9057 ( .A1(n14282), .A2(n14283), .ZN(n14281) );
  NOR2_X2 U9058 ( .A1(n14279), .A2(n9759), .ZN(n14282) );
  INV_X1 U9059 ( .A(n14260), .ZN(n6639) );
  OAI21_X2 U9060 ( .B1(n14453), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n9771), .ZN(
        n14287) );
  OR2_X2 U9062 ( .A1(n11052), .A2(n11851), .ZN(n11241) );
  NOR2_X2 U9063 ( .A1(n14155), .A2(n6513), .ZN(n14032) );
  INV_X1 U9064 ( .A(n11992), .ZN(n6626) );
  NAND2_X1 U9065 ( .A1(n6628), .A2(n6627), .ZN(n11992) );
  INV_X1 U9066 ( .A(n11991), .ZN(n6628) );
  NAND2_X1 U9067 ( .A1(n6639), .A2(n6638), .ZN(n6637) );
  AND2_X2 U9068 ( .A1(n11298), .A2(n14426), .ZN(n11415) );
  NAND2_X1 U9069 ( .A1(n14441), .A2(n6874), .ZN(n14446) );
  NAND2_X1 U9070 ( .A1(n13952), .A2(n13967), .ZN(n13949) );
  NOR2_X1 U9071 ( .A1(n9725), .A2(n14999), .ZN(n9705) );
  NOR2_X1 U9072 ( .A1(n9727), .A2(n9726), .ZN(n9702) );
  NAND2_X1 U9073 ( .A1(n6744), .A2(n14258), .ZN(n9956) );
  NAND2_X1 U9074 ( .A1(n6812), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8723) );
  NOR2_X1 U9075 ( .A1(n9745), .A2(n9744), .ZN(n9694) );
  NOR2_X1 U9076 ( .A1(n9753), .A2(n9752), .ZN(n9700) );
  NOR2_X1 U9077 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9750), .ZN(n9698) );
  NAND2_X1 U9078 ( .A1(n11877), .A2(n6554), .ZN(n14403) );
  NAND2_X1 U9079 ( .A1(n11070), .A2(n7379), .ZN(n11074) );
  NAND2_X1 U9080 ( .A1(n13612), .A2(n13615), .ZN(n13611) );
  NAND2_X1 U9081 ( .A1(n6731), .A2(n6729), .ZN(n8813) );
  NAND2_X1 U9082 ( .A1(n14709), .A2(n14708), .ZN(n14707) );
  NAND2_X1 U9083 ( .A1(n11969), .A2(n11968), .ZN(n11971) );
  NAND2_X1 U9084 ( .A1(n6979), .A2(n6978), .ZN(n11893) );
  INV_X1 U9085 ( .A(n11952), .ZN(n6986) );
  NAND2_X1 U9086 ( .A1(n10877), .A2(n6487), .ZN(n6967) );
  OAI211_X1 U9087 ( .C1(n8242), .C2(n7274), .A(n6633), .B(n8258), .ZN(n8060)
         );
  NAND2_X1 U9088 ( .A1(n7273), .A2(n8056), .ZN(n6633) );
  NAND2_X1 U9089 ( .A1(n7136), .A2(n6560), .ZN(n10932) );
  NAND2_X1 U9090 ( .A1(n11105), .A2(n7141), .ZN(n7139) );
  NAND2_X1 U9091 ( .A1(n11101), .A2(n11100), .ZN(n11105) );
  INV_X2 U9092 ( .A(n10521), .ZN(n10519) );
  NAND2_X4 U9093 ( .A1(n9959), .A2(n9960), .ZN(n10521) );
  NAND2_X2 U9094 ( .A1(n11272), .A2(n11271), .ZN(n11270) );
  NAND3_X1 U9095 ( .A1(n7523), .A2(n7577), .A3(n7447), .ZN(n7596) );
  AOI21_X1 U9096 ( .B1(n9964), .B2(n10028), .A(n9963), .ZN(n10491) );
  NOR2_X1 U9097 ( .A1(n10791), .A2(n10792), .ZN(n10790) );
  XNOR2_X1 U9098 ( .A(n9749), .B(P2_ADDR_REG_7__SCAN_IN), .ZN(n15141) );
  NOR2_X2 U9099 ( .A1(n14273), .A2(n9747), .ZN(n9749) );
  NAND2_X1 U9100 ( .A1(n15137), .A2(n15136), .ZN(n15135) );
  XNOR2_X1 U9101 ( .A(n6636), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  NAND2_X1 U9102 ( .A1(n14258), .A2(n6637), .ZN(n6636) );
  NAND2_X1 U9103 ( .A1(n14437), .A2(n14436), .ZN(n14435) );
  INV_X1 U9104 ( .A(n14281), .ZN(n6641) );
  NAND2_X1 U9105 ( .A1(n9293), .A2(n9292), .ZN(n9291) );
  NAND2_X1 U9106 ( .A1(n9289), .A2(n9288), .ZN(n9293) );
  INV_X1 U9107 ( .A(n7307), .ZN(n7303) );
  NAND3_X1 U9108 ( .A1(n9305), .A2(n9304), .A3(n7280), .ZN(n7279) );
  NAND2_X1 U9109 ( .A1(n11587), .A2(n7690), .ZN(n14338) );
  AOI21_X2 U9110 ( .B1(n11823), .B2(n12514), .A(n7709), .ZN(n11911) );
  NAND2_X2 U9111 ( .A1(n6644), .A2(n7527), .ZN(n15072) );
  OAI21_X2 U9112 ( .B1(n12888), .B2(n7262), .A(n7260), .ZN(n12867) );
  NAND2_X1 U9113 ( .A1(n6943), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6946) );
  NAND2_X1 U9114 ( .A1(n6646), .A2(n7526), .ZN(n7400) );
  INV_X1 U9115 ( .A(n7537), .ZN(n6646) );
  NAND2_X1 U9116 ( .A1(n6954), .A2(n7859), .ZN(n7858) );
  NAND2_X1 U9117 ( .A1(n12499), .A2(n12498), .ZN(n12500) );
  NAND2_X1 U9118 ( .A1(n6783), .A2(n6782), .ZN(P2_U3496) );
  AOI21_X2 U9119 ( .B1(n6651), .B2(n6650), .A(n6649), .ZN(n13415) );
  XNOR2_X1 U9120 ( .A(n8596), .B(n9657), .ZN(n6784) );
  OAI21_X1 U9121 ( .B1(n7349), .B2(n6522), .A(n9077), .ZN(n6653) );
  NAND2_X1 U9122 ( .A1(n11982), .A2(n11983), .ZN(n9079) );
  NAND2_X1 U9123 ( .A1(n6613), .A2(n7349), .ZN(n10807) );
  AOI21_X2 U9124 ( .B1(n13947), .B2(n13948), .A(n6552), .ZN(n13933) );
  NAND2_X2 U9125 ( .A1(n8739), .A2(n6706), .ZN(n8759) );
  NAND3_X1 U9126 ( .A1(n11289), .A2(n9380), .A3(n6494), .ZN(n6657) );
  NAND2_X1 U9127 ( .A1(n6658), .A2(n6657), .ZN(n11530) );
  NAND2_X1 U9128 ( .A1(n9089), .A2(n6659), .ZN(n6660) );
  NAND2_X1 U9129 ( .A1(n11201), .A2(n6671), .ZN(n6669) );
  NAND2_X1 U9130 ( .A1(n8752), .A2(n10745), .ZN(n8754) );
  NAND2_X1 U9131 ( .A1(n10085), .A2(n8741), .ZN(n9076) );
  NAND2_X1 U9132 ( .A1(n14052), .A2(n6489), .ZN(n6688) );
  NAND2_X1 U9133 ( .A1(n6688), .A2(n6689), .ZN(n13996) );
  OAI21_X1 U9134 ( .B1(n11863), .B2(n6507), .A(n6699), .ZN(n14074) );
  NAND2_X1 U9135 ( .A1(n11863), .A2(n6699), .ZN(n6698) );
  NAND2_X2 U9136 ( .A1(n8739), .A2(n8726), .ZN(n8978) );
  NAND2_X2 U9137 ( .A1(n14248), .A2(n9114), .ZN(n8739) );
  NAND2_X1 U9138 ( .A1(n9070), .A2(n8722), .ZN(n6812) );
  NAND2_X1 U9139 ( .A1(n6713), .A2(n6712), .ZN(n14112) );
  NAND2_X1 U9140 ( .A1(n7076), .A2(n7074), .ZN(n6712) );
  NAND2_X1 U9141 ( .A1(n6714), .A2(n13936), .ZN(n6713) );
  NAND2_X1 U9142 ( .A1(n7076), .A2(n9037), .ZN(n6714) );
  NAND2_X1 U9143 ( .A1(n6715), .A2(n8072), .ZN(n8075) );
  XNOR2_X1 U9144 ( .A(n6715), .B(n8334), .ZN(n10220) );
  NAND3_X1 U9145 ( .A1(n6773), .A2(n8098), .A3(n8472), .ZN(n8455) );
  NAND2_X1 U9146 ( .A1(n13369), .A2(n6721), .ZN(n6718) );
  AND2_X1 U9147 ( .A1(n6722), .A2(n6527), .ZN(n13356) );
  NAND3_X1 U9148 ( .A1(n6724), .A2(n6723), .A3(n7292), .ZN(n8095) );
  NAND2_X1 U9149 ( .A1(n6725), .A2(n8347), .ZN(n6724) );
  NAND2_X1 U9150 ( .A1(n6728), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9067) );
  NAND2_X1 U9151 ( .A1(n9073), .A2(n6728), .ZN(n11150) );
  NAND4_X1 U9152 ( .A1(n8697), .A2(n8699), .A3(n8698), .A4(n8696), .ZN(n8700)
         );
  AND2_X2 U9153 ( .A1(n6814), .A2(n8727), .ZN(n6729) );
  AND4_X2 U9154 ( .A1(n8788), .A2(n8728), .A3(n6813), .A4(n8761), .ZN(n6731)
         );
  INV_X1 U9155 ( .A(n8700), .ZN(n6730) );
  NAND2_X1 U9156 ( .A1(n12056), .A2(n6735), .ZN(n6733) );
  NAND2_X1 U9157 ( .A1(n11538), .A2(n11537), .ZN(n11539) );
  INV_X1 U9158 ( .A(n7385), .ZN(n6739) );
  NOR2_X2 U9159 ( .A1(n14280), .A2(n14618), .ZN(n14279) );
  NOR2_X1 U9160 ( .A1(n15132), .A2(n9739), .ZN(n9741) );
  MUX2_X1 U9161 ( .A(n10370), .B(P1_REG1_REG_1__SCAN_IN), .S(n10379), .Z(
        n13782) );
  NAND2_X1 U9162 ( .A1(n6773), .A2(n8472), .ZN(n8456) );
  NAND3_X1 U9163 ( .A1(n7103), .A2(n7098), .A3(n7097), .ZN(n6774) );
  OAI22_X1 U9164 ( .A1(n8112), .A2(n6508), .B1(n8507), .B2(SI_22_), .ZN(n6775)
         );
  NAND3_X1 U9165 ( .A1(n7332), .A2(n8507), .A3(n8113), .ZN(n8511) );
  AOI21_X1 U9166 ( .B1(n8305), .B2(n6776), .A(n6498), .ZN(n6781) );
  INV_X1 U9167 ( .A(n6777), .ZN(n6779) );
  OAI21_X1 U9168 ( .B1(n8305), .B2(n6498), .A(n6778), .ZN(n6777) );
  OAI21_X1 U9169 ( .B1(n7282), .B2(n8306), .A(n6781), .ZN(n8317) );
  NAND2_X1 U9170 ( .A1(n6780), .A2(n6779), .ZN(n8071) );
  NAND2_X1 U9171 ( .A1(n7282), .A2(n6781), .ZN(n6780) );
  NAND2_X1 U9172 ( .A1(n8524), .A2(n6563), .ZN(n6797) );
  NAND2_X1 U9173 ( .A1(n6797), .A2(n6798), .ZN(n8558) );
  NAND2_X1 U9174 ( .A1(n9135), .A2(n6812), .ZN(n14252) );
  INV_X1 U9175 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n8788) );
  INV_X1 U9176 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6813) );
  NOR2_X2 U9177 ( .A1(n13938), .A2(n13926), .ZN(n13908) );
  INV_X1 U9178 ( .A(n14537), .ZN(n6816) );
  NOR2_X2 U9179 ( .A1(n13985), .A2(n14208), .ZN(n13967) );
  NOR2_X2 U9180 ( .A1(n14015), .A2(n14142), .ZN(n6818) );
  INV_X1 U9181 ( .A(n11854), .ZN(n6819) );
  NAND2_X1 U9182 ( .A1(n6819), .A2(n6820), .ZN(n14065) );
  NAND2_X1 U9183 ( .A1(n6828), .A2(n6824), .ZN(n7495) );
  NOR2_X1 U9184 ( .A1(n7451), .A2(n6645), .ZN(n7705) );
  INV_X1 U9185 ( .A(n7451), .ZN(n6828) );
  NAND2_X1 U9186 ( .A1(n6829), .A2(n6831), .ZN(n7946) );
  NAND2_X1 U9187 ( .A1(n12942), .A2(n6833), .ZN(n6829) );
  NAND2_X1 U9188 ( .A1(n11350), .A2(n6842), .ZN(n6841) );
  NAND2_X1 U9189 ( .A1(n7937), .A2(n6853), .ZN(n6851) );
  NAND2_X1 U9190 ( .A1(n6570), .A2(n6851), .ZN(n11228) );
  NAND2_X1 U9191 ( .A1(n11828), .A2(n6493), .ZN(n6858) );
  NAND2_X1 U9192 ( .A1(n12967), .A2(n12428), .ZN(n12949) );
  INV_X1 U9193 ( .A(n12949), .ZN(n7944) );
  XNOR2_X2 U9194 ( .A(n6867), .B(P3_IR_REG_30__SCAN_IN), .ZN(n7481) );
  NAND2_X1 U9195 ( .A1(n6868), .A2(n7383), .ZN(n8597) );
  NAND2_X1 U9196 ( .A1(n7126), .A2(n6868), .ZN(n7128) );
  AND2_X2 U9197 ( .A1(n7127), .A2(n6868), .ZN(n8144) );
  INV_X2 U9198 ( .A(n8381), .ZN(n6868) );
  NAND2_X2 U9199 ( .A1(n6478), .A2(n6706), .ZN(n8206) );
  NAND2_X2 U9200 ( .A1(n6479), .A2(n8726), .ZN(n8225) );
  INV_X1 U9201 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n6875) );
  NOR2_X2 U9202 ( .A1(n9684), .A2(n9685), .ZN(n9686) );
  NAND2_X1 U9203 ( .A1(n13392), .A2(n6879), .ZN(n13340) );
  NAND2_X1 U9204 ( .A1(n11964), .A2(n6883), .ZN(n13431) );
  INV_X1 U9205 ( .A(n6885), .ZN(n13449) );
  NOR2_X2 U9206 ( .A1(n6491), .A2(n13553), .ZN(n11963) );
  NOR2_X2 U9207 ( .A1(n11456), .A2(n11504), .ZN(n6887) );
  NAND2_X1 U9208 ( .A1(n11607), .A2(n6894), .ZN(n6892) );
  INV_X1 U9209 ( .A(n6900), .ZN(n14923) );
  INV_X1 U9210 ( .A(n11614), .ZN(n6899) );
  XNOR2_X1 U9211 ( .A(n11608), .B(n11672), .ZN(n14889) );
  INV_X1 U9212 ( .A(n6912), .ZN(n12783) );
  NAND2_X1 U9213 ( .A1(n14307), .A2(n6611), .ZN(n6918) );
  AOI21_X1 U9214 ( .B1(n12790), .B2(n12789), .A(n12788), .ZN(n12811) );
  NAND3_X1 U9215 ( .A1(n6918), .A2(n14300), .A3(n6917), .ZN(n6924) );
  NAND3_X1 U9216 ( .A1(n6919), .A2(n6577), .A3(n12790), .ZN(n6917) );
  NAND2_X1 U9217 ( .A1(n6924), .A2(n12832), .ZN(P3_U3201) );
  INV_X1 U9218 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8186) );
  NAND3_X1 U9219 ( .A1(n12331), .A2(n12531), .A3(n6486), .ZN(n12532) );
  NAND2_X1 U9220 ( .A1(n7681), .A2(n6928), .ZN(n6927) );
  INV_X1 U9221 ( .A(n7704), .ZN(n6937) );
  NAND3_X1 U9222 ( .A1(n6939), .A2(n6941), .A3(n6938), .ZN(n7710) );
  NAND3_X1 U9223 ( .A1(n6946), .A2(n6948), .A3(n6945), .ZN(n7801) );
  NAND2_X1 U9224 ( .A1(n7846), .A2(n7845), .ZN(n6951) );
  OAI21_X1 U9225 ( .B1(n7628), .B2(n6961), .A(n6958), .ZN(n7663) );
  NAND2_X1 U9226 ( .A1(n7884), .A2(n6964), .ZN(n6963) );
  NAND2_X2 U9227 ( .A1(n8160), .A2(n8158), .ZN(n8465) );
  AND2_X2 U9228 ( .A1(n8159), .A2(n7128), .ZN(n8160) );
  INV_X1 U9229 ( .A(n10877), .ZN(n6971) );
  INV_X1 U9230 ( .A(n11455), .ZN(n8663) );
  NAND2_X1 U9231 ( .A1(n8665), .A2(n6981), .ZN(n6979) );
  OAI21_X2 U9232 ( .B1(n13442), .B2(n6991), .A(n6989), .ZN(n13425) );
  OR2_X2 U9233 ( .A1(n13425), .A2(n13424), .ZN(n13520) );
  NAND2_X1 U9234 ( .A1(n8144), .A2(n6993), .ZN(n8153) );
  NAND2_X1 U9235 ( .A1(n8144), .A2(n8145), .ZN(n8150) );
  NAND2_X1 U9236 ( .A1(n8153), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8154) );
  AND2_X1 U9237 ( .A1(n8203), .A2(n8205), .ZN(n6994) );
  INV_X1 U9238 ( .A(n10981), .ZN(n14759) );
  OR2_X2 U9239 ( .A1(n13384), .A2(n13385), .ZN(n6999) );
  OAI21_X2 U9240 ( .B1(n13397), .B2(n13398), .A(n6546), .ZN(n13384) );
  AOI21_X2 U9241 ( .B1(n13402), .B2(n8677), .A(n8676), .ZN(n13397) );
  OAI21_X2 U9242 ( .B1(n11893), .B2(n11892), .A(n8668), .ZN(n11969) );
  OAI22_X2 U9243 ( .A1(n13458), .A2(n8671), .B1(n13464), .B2(n8486), .ZN(
        n13442) );
  NAND2_X1 U9244 ( .A1(n14707), .A2(n8658), .ZN(n11333) );
  NAND2_X1 U9245 ( .A1(n13337), .A2(n8678), .ZN(n8680) );
  NAND2_X1 U9246 ( .A1(n11333), .A2(n11332), .ZN(n11331) );
  NAND2_X1 U9247 ( .A1(n7947), .A2(n12459), .ZN(n8001) );
  NAND2_X1 U9248 ( .A1(n7939), .A2(n12395), .ZN(n14336) );
  NAND2_X1 U9249 ( .A1(n15039), .A2(n12346), .ZN(n10913) );
  XNOR2_X2 U9250 ( .A(n7464), .B(n7463), .ZN(n7931) );
  NOR2_X4 U9251 ( .A1(n7495), .A2(n7456), .ZN(n7968) );
  AOI21_X1 U9252 ( .B1(n7375), .B2(n12540), .A(n12539), .ZN(n12547) );
  XNOR2_X1 U9253 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n7526) );
  NAND2_X1 U9254 ( .A1(n8656), .A2(n8655), .ZN(n10877) );
  NAND2_X1 U9255 ( .A1(n8143), .A2(n8153), .ZN(n8608) );
  INV_X4 U9256 ( .A(n8206), .ZN(n9460) );
  NAND2_X1 U9257 ( .A1(n9970), .A2(n9972), .ZN(n7009) );
  OAI21_X1 U9258 ( .B1(n10888), .B2(n7007), .A(n7005), .ZN(n10987) );
  INV_X1 U9259 ( .A(n7000), .ZN(n11142) );
  AOI21_X1 U9260 ( .B1(n10888), .B2(n7005), .A(n7001), .ZN(n7000) );
  NAND2_X1 U9261 ( .A1(n7002), .A2(n9976), .ZN(n7001) );
  NAND2_X1 U9262 ( .A1(n7005), .A2(n7007), .ZN(n7002) );
  NAND2_X1 U9263 ( .A1(n10888), .A2(n9970), .ZN(n10943) );
  OR2_X1 U9264 ( .A1(n9973), .A2(n10944), .ZN(n7008) );
  INV_X1 U9265 ( .A(n7968), .ZN(n7963) );
  NAND2_X1 U9266 ( .A1(n7966), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7967) );
  NAND2_X1 U9267 ( .A1(n7968), .A2(n7964), .ZN(n7966) );
  NAND2_X1 U9268 ( .A1(n12597), .A2(n10025), .ZN(n12660) );
  INV_X1 U9269 ( .A(n7013), .ZN(n12584) );
  NAND2_X1 U9270 ( .A1(n12574), .A2(n12687), .ZN(n7021) );
  NAND3_X1 U9271 ( .A1(n7023), .A2(n10017), .A3(n12588), .ZN(n12642) );
  NAND2_X1 U9272 ( .A1(n10016), .A2(n10015), .ZN(n10017) );
  NAND2_X2 U9273 ( .A1(n12673), .A2(n12672), .ZN(n12671) );
  NAND2_X1 U9274 ( .A1(n11904), .A2(n7029), .ZN(n7027) );
  NAND2_X1 U9275 ( .A1(n11270), .A2(n7033), .ZN(n7036) );
  CLKBUF_X1 U9276 ( .A(n7036), .Z(n7031) );
  INV_X1 U9277 ( .A(n7031), .ZN(n11385) );
  INV_X1 U9278 ( .A(n9978), .ZN(n7038) );
  NAND2_X1 U9279 ( .A1(n12262), .A2(n12261), .ZN(n7049) );
  NAND2_X1 U9280 ( .A1(n14407), .A2(n6567), .ZN(n13643) );
  NAND2_X1 U9281 ( .A1(n12056), .A2(n12055), .ZN(n13665) );
  NAND2_X1 U9282 ( .A1(n11877), .A2(n11876), .ZN(n12004) );
  AND2_X1 U9283 ( .A1(n9070), .A2(n7061), .ZN(n9129) );
  NAND2_X1 U9284 ( .A1(n9133), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9134) );
  INV_X4 U9285 ( .A(n8978), .ZN(n8774) );
  NAND2_X2 U9286 ( .A1(n8725), .A2(n8724), .ZN(n14248) );
  OAI21_X1 U9287 ( .B1(n9169), .B2(n7067), .A(n9182), .ZN(n9183) );
  NAND2_X1 U9288 ( .A1(n10751), .A2(n7067), .ZN(n10707) );
  NAND2_X1 U9289 ( .A1(n13946), .A2(n7073), .ZN(n7071) );
  NAND2_X1 U9290 ( .A1(n7071), .A2(n7072), .ZN(n9059) );
  NAND2_X1 U9291 ( .A1(n13946), .A2(n13945), .ZN(n7076) );
  NAND2_X1 U9292 ( .A1(n11468), .A2(n6555), .ZN(n11518) );
  NAND2_X1 U9293 ( .A1(n11518), .A2(n7077), .ZN(n8914) );
  NAND2_X1 U9294 ( .A1(n7080), .A2(n7079), .ZN(n11986) );
  NAND2_X1 U9295 ( .A1(n8765), .A2(n8764), .ZN(n10798) );
  AND4_X2 U9296 ( .A1(n8185), .A2(n7088), .A3(n8184), .A4(n7087), .ZN(n10616)
         );
  OAI21_X1 U9297 ( .B1(n7091), .B2(n10826), .A(n8301), .ZN(n7090) );
  NAND2_X1 U9298 ( .A1(n7092), .A2(n8303), .ZN(n11156) );
  NAND2_X1 U9299 ( .A1(n7094), .A2(n7096), .ZN(n13334) );
  NAND2_X1 U9300 ( .A1(n7095), .A2(n6538), .ZN(n7094) );
  INV_X1 U9301 ( .A(n13375), .ZN(n7095) );
  OAI21_X1 U9302 ( .B1(n13375), .B2(n13374), .A(n7105), .ZN(n13360) );
  NAND2_X1 U9303 ( .A1(n13497), .A2(n13188), .ZN(n7106) );
  INV_X1 U9304 ( .A(n11711), .ZN(n7109) );
  NAND2_X1 U9305 ( .A1(n7109), .A2(n6580), .ZN(n7110) );
  NAND2_X1 U9306 ( .A1(n7110), .A2(n6562), .ZN(n8443) );
  NAND2_X1 U9307 ( .A1(n8471), .A2(n7113), .ZN(n7112) );
  NAND2_X1 U9308 ( .A1(n8431), .A2(n7130), .ZN(n7129) );
  NAND2_X1 U9309 ( .A1(n10907), .A2(n10779), .ZN(n7136) );
  NAND2_X1 U9310 ( .A1(n11722), .A2(n6564), .ZN(n12160) );
  NAND2_X1 U9311 ( .A1(n13251), .A2(n7144), .ZN(n7143) );
  OAI211_X1 U9312 ( .C1(n13251), .C2(n7145), .A(n7143), .B(n12217), .ZN(
        P2_U3192) );
  NAND2_X1 U9313 ( .A1(n13251), .A2(n12204), .ZN(n13145) );
  INV_X1 U9314 ( .A(n12211), .ZN(n7158) );
  OAI21_X1 U9315 ( .B1(n7161), .B2(n10468), .A(n7159), .ZN(n10638) );
  AND2_X1 U9316 ( .A1(n7160), .A2(n10635), .ZN(n7159) );
  NAND3_X1 U9317 ( .A1(n10470), .A2(n10469), .A3(n13161), .ZN(n7160) );
  INV_X1 U9318 ( .A(n7162), .ZN(n7161) );
  AND2_X1 U9319 ( .A1(n10470), .A2(n10469), .ZN(n7162) );
  INV_X1 U9320 ( .A(n13205), .ZN(n7169) );
  NAND2_X1 U9321 ( .A1(n13169), .A2(n7175), .ZN(n7170) );
  NAND2_X1 U9322 ( .A1(n7170), .A2(n7171), .ZN(n12185) );
  NAND3_X1 U9323 ( .A1(n7177), .A2(n7178), .A3(n7176), .ZN(n7174) );
  NAND2_X1 U9324 ( .A1(n9595), .A2(n7183), .ZN(n7181) );
  NAND2_X1 U9325 ( .A1(n7181), .A2(n7182), .ZN(n9604) );
  NAND3_X1 U9326 ( .A1(n9540), .A2(n9541), .A3(n6566), .ZN(n7198) );
  NAND2_X1 U9327 ( .A1(n7199), .A2(n7200), .ZN(n9558) );
  NAND3_X1 U9328 ( .A1(n9552), .A2(n6572), .A3(n9551), .ZN(n7199) );
  NAND2_X1 U9329 ( .A1(n7201), .A2(n7202), .ZN(n9581) );
  NAND3_X1 U9330 ( .A1(n9575), .A2(n6597), .A3(n9574), .ZN(n7201) );
  NAND2_X1 U9331 ( .A1(n9584), .A2(n9583), .ZN(n7204) );
  NAND2_X1 U9332 ( .A1(n9580), .A2(n9579), .ZN(n7205) );
  NAND3_X1 U9333 ( .A1(n7205), .A2(n7204), .A3(n6595), .ZN(n7203) );
  NAND2_X1 U9334 ( .A1(n9534), .A2(n7211), .ZN(n7208) );
  OAI21_X1 U9335 ( .B1(n9534), .B2(n7213), .A(n7211), .ZN(n9539) );
  NAND2_X1 U9336 ( .A1(n7208), .A2(n7209), .ZN(n9537) );
  NAND2_X1 U9337 ( .A1(n7214), .A2(n7216), .ZN(n9502) );
  NAND3_X1 U9338 ( .A1(n9495), .A2(n7215), .A3(n9494), .ZN(n7214) );
  NAND3_X1 U9339 ( .A1(n9563), .A2(n9562), .A3(n6596), .ZN(n7218) );
  NAND2_X1 U9340 ( .A1(n7218), .A2(n7219), .ZN(n9570) );
  NAND2_X1 U9341 ( .A1(n7220), .A2(n7221), .ZN(n9513) );
  NAND3_X1 U9342 ( .A1(n9507), .A2(n6568), .A3(n9506), .ZN(n7220) );
  NAND3_X1 U9343 ( .A1(n9518), .A2(n6569), .A3(n9517), .ZN(n7223) );
  NAND2_X1 U9344 ( .A1(n7223), .A2(n7224), .ZN(n9526) );
  NAND2_X2 U9345 ( .A1(n12345), .A2(n12348), .ZN(n15068) );
  NAND2_X2 U9346 ( .A1(n15042), .A2(n15072), .ZN(n12348) );
  NAND2_X1 U9347 ( .A1(n10406), .A2(n7539), .ZN(n12345) );
  OAI21_X1 U9348 ( .B1(n12962), .B2(n7229), .A(n7227), .ZN(n7226) );
  AND2_X1 U9349 ( .A1(n12943), .A2(n12926), .ZN(n7233) );
  OAI22_X2 U9350 ( .A1(n11911), .A2(n12517), .B1(n14353), .B2(n14328), .ZN(
        n14326) );
  NAND2_X1 U9351 ( .A1(n7257), .A2(n7258), .ZN(n8003) );
  NAND2_X1 U9352 ( .A1(n12888), .A2(n7260), .ZN(n7257) );
  NAND2_X1 U9353 ( .A1(n12888), .A2(n12887), .ZN(n12886) );
  NAND2_X1 U9354 ( .A1(n7585), .A2(n7263), .ZN(n15012) );
  AND2_X1 U9355 ( .A1(n7968), .A2(n7265), .ZN(n7470) );
  NAND2_X1 U9356 ( .A1(n7968), .A2(n7459), .ZN(n7462) );
  NAND2_X1 U9357 ( .A1(n7968), .A2(n7266), .ZN(n7471) );
  AND2_X2 U9358 ( .A1(n7270), .A2(n7268), .ZN(n8043) );
  NAND4_X1 U9359 ( .A1(n7466), .A2(n12256), .A3(P3_ADDR_REG_19__SCAN_IN), .A4(
        n7269), .ZN(n7268) );
  NAND4_X1 U9360 ( .A1(n7465), .A2(n7271), .A3(P1_ADDR_REG_19__SCAN_IN), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n7270) );
  NAND2_X1 U9361 ( .A1(n7272), .A2(n8056), .ZN(n8257) );
  NAND2_X1 U9362 ( .A1(n8242), .A2(n8243), .ZN(n7272) );
  INV_X1 U9363 ( .A(n8243), .ZN(n7273) );
  INV_X1 U9364 ( .A(n8056), .ZN(n7274) );
  NAND2_X1 U9365 ( .A1(n7279), .A2(n7278), .ZN(n9310) );
  NAND2_X1 U9366 ( .A1(n6524), .A2(n9306), .ZN(n7278) );
  NAND2_X1 U9367 ( .A1(n9310), .A2(n9311), .ZN(n9309) );
  NAND2_X1 U9368 ( .A1(n8271), .A2(n7283), .ZN(n7282) );
  NAND2_X1 U9369 ( .A1(n8086), .A2(n8085), .ZN(n8393) );
  NOR2_X2 U9370 ( .A1(n8813), .A2(n8700), .ZN(n8901) );
  NAND4_X1 U9371 ( .A1(n8707), .A2(n8901), .A3(n8703), .A4(n8719), .ZN(n8709)
         );
  INV_X1 U9372 ( .A(n9319), .ZN(n7297) );
  OAI21_X1 U9373 ( .B1(n9257), .B2(n7304), .A(n7302), .ZN(n7311) );
  NAND2_X1 U9374 ( .A1(n7311), .A2(n14088), .ZN(n9263) );
  NAND2_X1 U9375 ( .A1(n7312), .A2(n7315), .ZN(n9227) );
  NAND3_X1 U9376 ( .A1(n9222), .A2(n7313), .A3(n9221), .ZN(n7312) );
  NAND2_X1 U9377 ( .A1(n8127), .A2(n6604), .ZN(n7317) );
  NAND2_X1 U9378 ( .A1(n8127), .A2(n7318), .ZN(n7321) );
  NAND2_X1 U9379 ( .A1(n8127), .A2(n8126), .ZN(n8588) );
  NAND2_X1 U9380 ( .A1(n7317), .A2(n7322), .ZN(n9328) );
  INV_X1 U9381 ( .A(n7324), .ZN(n9273) );
  AOI21_X1 U9382 ( .B1(n9268), .B2(n7326), .A(n7325), .ZN(n7324) );
  INV_X1 U9383 ( .A(n9269), .ZN(n7328) );
  NAND2_X1 U9384 ( .A1(n7329), .A2(n7330), .ZN(n9217) );
  NAND3_X1 U9385 ( .A1(n9212), .A2(n6571), .A3(n9211), .ZN(n7329) );
  NAND3_X1 U9386 ( .A1(n7333), .A2(n8108), .A3(n8107), .ZN(n8503) );
  NAND2_X1 U9387 ( .A1(n8106), .A2(n8105), .ZN(n8108) );
  NAND2_X1 U9388 ( .A1(n8103), .A2(n10899), .ZN(n7333) );
  NAND2_X1 U9389 ( .A1(n8117), .A2(n8118), .ZN(n8522) );
  NAND3_X1 U9390 ( .A1(n9197), .A2(n9196), .A3(n7339), .ZN(n7337) );
  NAND2_X1 U9391 ( .A1(n7340), .A2(n7341), .ZN(n9284) );
  NAND3_X1 U9392 ( .A1(n9278), .A2(n9277), .A3(n6575), .ZN(n7340) );
  NAND2_X1 U9393 ( .A1(n9070), .A2(n7342), .ZN(n9068) );
  INV_X1 U9394 ( .A(n9068), .ZN(n9065) );
  NAND2_X1 U9395 ( .A1(n9068), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9063) );
  AOI21_X1 U9396 ( .B1(n7351), .B2(n10706), .A(n6559), .ZN(n7349) );
  INV_X1 U9397 ( .A(n10706), .ZN(n7350) );
  NAND2_X1 U9398 ( .A1(n10707), .A2(n10706), .ZN(n10705) );
  NAND2_X1 U9399 ( .A1(n6573), .A2(n7356), .ZN(n7355) );
  NAND2_X1 U9400 ( .A1(n13997), .A2(n7357), .ZN(n7356) );
  NAND2_X1 U9401 ( .A1(n12479), .A2(n12468), .ZN(n12474) );
  INV_X1 U9402 ( .A(n12856), .ZN(n13080) );
  INV_X1 U9403 ( .A(n8037), .ZN(P3_U3486) );
  NAND2_X1 U9404 ( .A1(n11142), .A2(n11141), .ZN(n11140) );
  NAND2_X1 U9405 ( .A1(n13886), .A2(n9176), .ZN(n9360) );
  XNOR2_X1 U9406 ( .A(n7498), .B(n7497), .ZN(n7955) );
  NAND2_X1 U9407 ( .A1(n12536), .A2(n15053), .ZN(n12537) );
  NOR2_X2 U9408 ( .A1(n13514), .A2(n13418), .ZN(n13409) );
  NAND2_X1 U9409 ( .A1(n12306), .A2(n12491), .ZN(n12333) );
  NAND2_X1 U9410 ( .A1(n13734), .A2(n13735), .ZN(n13733) );
  XNOR2_X1 U9411 ( .A(n10452), .B(n10453), .ZN(n10617) );
  XNOR2_X1 U9412 ( .A(n6480), .B(n11180), .ZN(n10452) );
  NAND2_X1 U9413 ( .A1(n13693), .A2(n13694), .ZN(n14393) );
  INV_X1 U9414 ( .A(n11114), .ZN(n11115) );
  INV_X1 U9415 ( .A(n12535), .ZN(n12538) );
  NAND2_X1 U9416 ( .A1(n13072), .A2(n15131), .ZN(n8000) );
  INV_X1 U9417 ( .A(n11070), .ZN(n10104) );
  NAND2_X1 U9418 ( .A1(n8681), .A2(n9475), .ZN(n14769) );
  NAND2_X1 U9419 ( .A1(n9449), .A2(n15131), .ZN(n9452) );
  INV_X1 U9420 ( .A(n11173), .ZN(n9643) );
  NAND2_X1 U9421 ( .A1(n8201), .A2(n9477), .ZN(n10970) );
  NAND2_X2 U9422 ( .A1(n13611), .A2(n12120), .ZN(n12262) );
  NAND2_X1 U9423 ( .A1(n9065), .A2(n9064), .ZN(n9151) );
  NAND2_X1 U9424 ( .A1(n12492), .A2(n12491), .ZN(n12499) );
  AOI21_X1 U9425 ( .B1(n12492), .B2(n12490), .A(n12529), .ZN(n12501) );
  NOR2_X1 U9426 ( .A1(n9129), .A2(n9128), .ZN(n9130) );
  INV_X1 U9427 ( .A(n9129), .ZN(n9124) );
  NAND2_X1 U9428 ( .A1(n7955), .A2(n10898), .ZN(n9958) );
  OR2_X1 U9429 ( .A1(n7542), .A2(n10329), .ZN(n7531) );
  NAND2_X1 U9430 ( .A1(n9371), .A2(n9076), .ZN(n9185) );
  AND2_X1 U9431 ( .A1(n10090), .A2(n10089), .ZN(n10091) );
  NAND2_X1 U9432 ( .A1(n13900), .A2(n9061), .ZN(n13922) );
  AOI21_X1 U9433 ( .B1(n8034), .B2(n15060), .A(n8033), .ZN(n12858) );
  NAND2_X1 U9434 ( .A1(n7070), .A2(n9097), .ZN(n9099) );
  NAND2_X1 U9435 ( .A1(n9403), .A2(n9404), .ZN(n9407) );
  NAND2_X1 U9436 ( .A1(n6475), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8051) );
  INV_X1 U9437 ( .A(n10341), .ZN(n7790) );
  NAND2_X1 U9438 ( .A1(n10341), .A2(n6706), .ZN(n7550) );
  NOR2_X1 U9439 ( .A1(n10719), .A2(n10718), .ZN(n10721) );
  INV_X1 U9440 ( .A(n13774), .ZN(n8741) );
  INV_X1 U9441 ( .A(n11674), .ZN(n14913) );
  OR2_X1 U9442 ( .A1(n12862), .A2(n13063), .ZN(n7362) );
  OR2_X1 U9443 ( .A1(n13075), .A2(n13063), .ZN(n7363) );
  INV_X2 U9444 ( .A(n15080), .ZN(n15082) );
  INV_X1 U9445 ( .A(n15131), .ZN(n9450) );
  AND2_X1 U9446 ( .A1(n9248), .A2(n9247), .ZN(n7364) );
  XNOR2_X1 U9447 ( .A(n12162), .B(n12163), .ZN(n13265) );
  OR2_X1 U9448 ( .A1(n9422), .A2(n9421), .ZN(n7365) );
  AND3_X1 U9449 ( .A1(n7510), .A2(n7509), .A3(n7508), .ZN(n14334) );
  OR2_X1 U9450 ( .A1(n12862), .A2(n13121), .ZN(n7366) );
  INV_X1 U9451 ( .A(SI_23_), .ZN(n11288) );
  AND2_X1 U9452 ( .A1(n6587), .A2(n9447), .ZN(n7367) );
  AND2_X1 U9453 ( .A1(n8683), .A2(n9665), .ZN(n7368) );
  AND2_X1 U9454 ( .A1(n13074), .A2(n13073), .ZN(n7369) );
  AND2_X1 U9455 ( .A1(n12178), .A2(n12177), .ZN(n7370) );
  AND2_X1 U9456 ( .A1(n13109), .A2(n12978), .ZN(n7371) );
  AND2_X1 U9457 ( .A1(n6586), .A2(n9451), .ZN(n7372) );
  AND2_X1 U9458 ( .A1(n12165), .A2(n12164), .ZN(n7373) );
  XOR2_X1 U9459 ( .A(n12335), .B(n12334), .Z(n7375) );
  AND2_X1 U9460 ( .A1(n8083), .A2(n8082), .ZN(n7376) );
  AND3_X1 U9461 ( .A1(n8715), .A2(n8714), .A3(n8713), .ZN(n7377) );
  OR2_X2 U9462 ( .A1(n8942), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n7378) );
  NAND2_X1 U9463 ( .A1(n11069), .A2(n11068), .ZN(n7379) );
  AND2_X1 U9464 ( .A1(n6476), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7381) );
  OR2_X1 U9465 ( .A1(n11504), .A2(n13297), .ZN(n7382) );
  BUF_X1 U9466 ( .A(n7495), .Z(n7715) );
  AND2_X1 U9467 ( .A1(n12526), .A2(n12467), .ZN(n7384) );
  NAND2_X1 U9468 ( .A1(n11074), .A2(n11075), .ZN(n7385) );
  INV_X1 U9469 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n7719) );
  INV_X1 U9470 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8386) );
  INV_X1 U9471 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n7684) );
  INV_X1 U9472 ( .A(n13890), .ZN(n9359) );
  INV_X1 U9473 ( .A(n14232), .ZN(n9158) );
  AND2_X1 U9474 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n7386) );
  OR2_X1 U9475 ( .A1(n9985), .A2(n9984), .ZN(n7387) );
  AND2_X1 U9476 ( .A1(n12185), .A2(n12184), .ZN(n7388) );
  INV_X1 U9477 ( .A(n14023), .ZN(n11860) );
  AND3_X1 U9478 ( .A1(n12502), .A2(n12487), .A3(n12328), .ZN(n7390) );
  INV_X1 U9479 ( .A(n12529), .ZN(n12331) );
  AND3_X1 U9480 ( .A1(n9658), .A2(n9626), .A3(n9625), .ZN(n7391) );
  AND4_X1 U9481 ( .A1(n9658), .A2(n9620), .A3(n9626), .A4(n9619), .ZN(n7392)
         );
  AND2_X1 U9482 ( .A1(n9407), .A2(n9406), .ZN(n7393) );
  INV_X1 U9483 ( .A(n9404), .ZN(n9364) );
  OR2_X1 U9484 ( .A1(n13557), .A2(n9648), .ZN(n7394) );
  INV_X1 U9485 ( .A(n9384), .ZN(n8899) );
  AND3_X1 U9486 ( .A1(n13948), .A2(n13960), .A3(n9392), .ZN(n7395) );
  AND2_X1 U9487 ( .A1(n11829), .A2(n15116), .ZN(n14354) );
  NAND2_X1 U9488 ( .A1(n7932), .A2(n12496), .ZN(n14339) );
  OR2_X1 U9489 ( .A1(n12844), .A2(n14354), .ZN(n7398) );
  NAND2_X1 U9490 ( .A1(n12898), .A2(n12897), .ZN(n12880) );
  AND2_X1 U9491 ( .A1(n10487), .A2(n10447), .ZN(n9476) );
  OAI211_X1 U9492 ( .C1(n9482), .C2(n9481), .A(n9480), .B(n9479), .ZN(n9485)
         );
  NAND2_X1 U9493 ( .A1(n9493), .A2(n9492), .ZN(n9494) );
  NAND2_X1 U9494 ( .A1(n9505), .A2(n9504), .ZN(n9506) );
  AOI21_X1 U9495 ( .B1(n9227), .B2(n9226), .A(n9225), .ZN(n9229) );
  INV_X1 U9496 ( .A(n9258), .ZN(n9259) );
  INV_X1 U9497 ( .A(n9285), .ZN(n9286) );
  MUX2_X1 U9498 ( .A(n13751), .B(n14212), .S(n9176), .Z(n9292) );
  INV_X1 U9499 ( .A(n9301), .ZN(n9302) );
  INV_X1 U9500 ( .A(n9307), .ZN(n6524) );
  OAI21_X1 U9501 ( .B1(n12471), .B2(n12470), .A(n12469), .ZN(n12472) );
  INV_X1 U9502 ( .A(n12472), .ZN(n12473) );
  NAND2_X1 U9503 ( .A1(n9393), .A2(n7395), .ZN(n9394) );
  NAND2_X1 U9504 ( .A1(n12474), .A2(n12473), .ZN(n12484) );
  NOR2_X1 U9505 ( .A1(n9394), .A2(n13932), .ZN(n9395) );
  AND2_X1 U9506 ( .A1(n13068), .A2(n12494), .ZN(n12495) );
  INV_X1 U9507 ( .A(n9621), .ZN(n9614) );
  NOR3_X1 U9508 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .A3(
        P2_IR_REG_20__SCAN_IN), .ZN(n8138) );
  OR2_X1 U9509 ( .A1(n13886), .A2(n9359), .ZN(n9361) );
  INV_X1 U9510 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7458) );
  INV_X1 U9511 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n7452) );
  INV_X1 U9512 ( .A(n13291), .ZN(n8486) );
  INV_X1 U9513 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n8128) );
  NAND2_X1 U9514 ( .A1(n9364), .A2(n9405), .ZN(n9406) );
  OR4_X1 U9515 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n9143) );
  INV_X1 U9516 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n9923) );
  AND2_X1 U9517 ( .A1(n7969), .A2(n7458), .ZN(n7459) );
  INV_X1 U9518 ( .A(n11106), .ZN(n11102) );
  AND2_X1 U9519 ( .A1(n8539), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n8545) );
  INV_X1 U9520 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8139) );
  AND2_X1 U9521 ( .A1(n8099), .A2(n8472), .ZN(n8100) );
  INV_X1 U9522 ( .A(n7835), .ZN(n7834) );
  INV_X1 U9523 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11610) );
  NAND2_X1 U9524 ( .A1(n7478), .A2(n9923), .ZN(n7820) );
  AND2_X1 U9525 ( .A1(n11908), .A2(n12692), .ZN(n7709) );
  INV_X1 U9526 ( .A(n13161), .ZN(n10467) );
  AND2_X1 U9527 ( .A1(n8545), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n8563) );
  NOR2_X1 U9528 ( .A1(n13543), .A2(n13292), .ZN(n8470) );
  AOI22_X1 U9529 ( .A1(n11076), .A2(n13774), .B1(n10085), .B2(n12282), .ZN(
        n10086) );
  INV_X1 U9530 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n8865) );
  INV_X1 U9531 ( .A(n12005), .ZN(n12006) );
  XNOR2_X1 U9532 ( .A(n9400), .B(n11860), .ZN(n9409) );
  AND2_X1 U9533 ( .A1(n8919), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8934) );
  AND2_X1 U9534 ( .A1(SI_20_), .A2(n8104), .ZN(n8105) );
  INV_X1 U9535 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n8929) );
  AND2_X1 U9536 ( .A1(n9678), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n9679) );
  NOR2_X1 U9537 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n9728), .ZN(n9688) );
  INV_X1 U9538 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n9795) );
  INV_X1 U9539 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n7750) );
  OR2_X1 U9540 ( .A1(n7820), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n7835) );
  NOR2_X1 U9541 ( .A1(n11674), .A2(n11610), .ZN(n11611) );
  INV_X1 U9542 ( .A(n11803), .ZN(n11811) );
  NAND2_X1 U9543 ( .A1(n8025), .A2(n12470), .ZN(n9444) );
  AOI21_X1 U9544 ( .B1(n12913), .B2(n7827), .A(n7826), .ZN(n12902) );
  INV_X1 U9545 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n11934) );
  INV_X1 U9546 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n7586) );
  INV_X1 U9547 ( .A(n12543), .ZN(n7960) );
  OR2_X1 U9548 ( .A1(n7954), .A2(n7953), .ZN(n10038) );
  AND2_X1 U9549 ( .A1(n8462), .A2(n8162), .ZN(n8491) );
  NOR2_X1 U9550 ( .A1(n8419), .A2(n13270), .ZN(n8418) );
  AND2_X1 U9551 ( .A1(n8565), .A2(n8548), .ZN(n13380) );
  INV_X1 U9552 ( .A(n9522), .ZN(n11332) );
  INV_X1 U9553 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8132) );
  AND2_X1 U9554 ( .A1(n13677), .A2(n12109), .ZN(n13613) );
  INV_X1 U9555 ( .A(n9010), .ZN(n9011) );
  OR2_X1 U9556 ( .A1(n8949), .A2(n8948), .ZN(n8962) );
  INV_X1 U9557 ( .A(n8992), .ZN(n8993) );
  INV_X1 U9558 ( .A(n10099), .ZN(n10233) );
  AND2_X1 U9559 ( .A1(n13921), .A2(n13928), .ZN(n9121) );
  INV_X1 U9560 ( .A(n11520), .ZN(n11743) );
  INV_X1 U9561 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n9687) );
  NAND2_X1 U9562 ( .A1(n7477), .A2(n9795), .ZN(n7807) );
  OR2_X1 U9563 ( .A1(n9969), .A2(n12700), .ZN(n9970) );
  INV_X1 U9564 ( .A(n12696), .ZN(n11388) );
  AND2_X1 U9565 ( .A1(n7720), .A2(n7719), .ZN(n7734) );
  INV_X1 U9566 ( .A(n9972), .ZN(n9973) );
  NAND2_X1 U9567 ( .A1(n10037), .A2(n15063), .ZN(n12665) );
  INV_X2 U9568 ( .A(n12496), .ZN(n12488) );
  INV_X1 U9569 ( .A(n14272), .ZN(n10347) );
  INV_X1 U9570 ( .A(n14930), .ZN(n11612) );
  INV_X1 U9571 ( .A(n14965), .ZN(n11615) );
  OR2_X1 U9572 ( .A1(n10353), .A2(n10352), .ZN(n10355) );
  OR2_X1 U9573 ( .A1(n14339), .A2(n9440), .ZN(n12833) );
  INV_X1 U9574 ( .A(n12964), .ZN(n12970) );
  AND2_X1 U9575 ( .A1(n7734), .A2(n11934), .ZN(n7751) );
  INV_X1 U9576 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n7655) );
  NAND2_X1 U9577 ( .A1(n12334), .A2(n10898), .ZN(n15073) );
  AND2_X1 U9578 ( .A1(n10043), .A2(n10660), .ZN(n10663) );
  OR2_X1 U9579 ( .A1(n15120), .A2(n9446), .ZN(n9447) );
  AND2_X1 U9580 ( .A1(n7434), .A2(n7433), .ZN(n7757) );
  AND2_X1 U9581 ( .A1(n7427), .A2(n7426), .ZN(n7701) );
  AND2_X1 U9582 ( .A1(n7419), .A2(n7418), .ZN(n7648) );
  NAND2_X1 U9583 ( .A1(n7408), .A2(n7407), .ZN(n7595) );
  NOR2_X1 U9584 ( .A1(n8527), .A2(n13155), .ZN(n8536) );
  INV_X1 U9585 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n13210) );
  INV_X1 U9586 ( .A(n13288), .ZN(n13180) );
  AND2_X1 U9587 ( .A1(n8574), .A2(n8573), .ZN(n13352) );
  AND2_X1 U9588 ( .A1(n8491), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n8514) );
  OR2_X1 U9589 ( .A1(n8450), .A2(n13210), .ZN(n8463) );
  INV_X1 U9590 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n11167) );
  OR2_X1 U9591 ( .A1(n10207), .A2(n10208), .ZN(n14595) );
  INV_X1 U9592 ( .A(n13287), .ZN(n13234) );
  INV_X1 U9593 ( .A(n13537), .ZN(n13464) );
  OR2_X1 U9594 ( .A1(n8324), .A2(n8161), .ZN(n8340) );
  NAND2_X1 U9595 ( .A1(n14733), .A2(n14719), .ZN(n13453) );
  INV_X1 U9596 ( .A(n10971), .ZN(n10968) );
  OR2_X1 U9597 ( .A1(n14769), .A2(n9666), .ZN(n10844) );
  NAND2_X1 U9598 ( .A1(n13339), .A2(n13338), .ZN(n13337) );
  INV_X1 U9599 ( .A(n9650), .ZN(n11713) );
  INV_X1 U9600 ( .A(n14725), .ZN(n13462) );
  INV_X1 U9601 ( .A(n13641), .ZN(n12017) );
  AND3_X1 U9602 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n8797) );
  NOR2_X1 U9603 ( .A1(n8970), .A2(n13688), .ZN(n8981) );
  INV_X1 U9604 ( .A(n13717), .ZN(n13633) );
  INV_X1 U9605 ( .A(n10107), .ZN(n10112) );
  NAND2_X1 U9606 ( .A1(n10181), .A2(n10108), .ZN(n10116) );
  INV_X1 U9607 ( .A(n10116), .ZN(n10651) );
  NAND2_X1 U9608 ( .A1(n8122), .A2(n8121), .ZN(n8560) );
  INV_X1 U9609 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9062) );
  NOR2_X1 U9610 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n9740), .ZN(n9692) );
  AOI21_X1 U9611 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n9714), .A(n9713), .ZN(
        n9718) );
  AND2_X1 U9612 ( .A1(n10037), .A2(n15062), .ZN(n12663) );
  AND2_X1 U9613 ( .A1(n10033), .A2(n12670), .ZN(n10034) );
  NAND2_X1 U9614 ( .A1(n10407), .A2(n12546), .ZN(n12678) );
  NAND2_X1 U9615 ( .A1(n13125), .A2(n10073), .ZN(n12541) );
  AND4_X1 U9616 ( .A1(n7911), .A2(n7910), .A3(n7909), .A4(n7908), .ZN(n12560)
         );
  XNOR2_X1 U9617 ( .A(n11613), .B(n11612), .ZN(n14924) );
  INV_X1 U9618 ( .A(n14985), .ZN(n14962) );
  INV_X1 U9619 ( .A(n14341), .ZN(n15062) );
  AND2_X1 U9620 ( .A1(n12408), .A2(n12407), .ZN(n12517) );
  INV_X1 U9621 ( .A(n12960), .ZN(n14346) );
  NOR2_X1 U9622 ( .A1(n10665), .A2(n15053), .ZN(n15036) );
  INV_X1 U9623 ( .A(n15009), .ZN(n15077) );
  AND3_X1 U9624 ( .A1(n8007), .A2(n7995), .A3(n8014), .ZN(n10662) );
  INV_X1 U9625 ( .A(n15116), .ZN(n15112) );
  INV_X1 U9626 ( .A(n14354), .ZN(n15100) );
  XNOR2_X1 U9627 ( .A(n7980), .B(n7979), .ZN(n10339) );
  INV_X1 U9628 ( .A(n13256), .ZN(n13172) );
  AND2_X1 U9629 ( .A1(n10479), .A2(n10478), .ZN(n13257) );
  AND4_X1 U9630 ( .A1(n8170), .A2(n8169), .A3(n8168), .A4(n8167), .ZN(n13146)
         );
  AND2_X1 U9631 ( .A1(n10209), .A2(n10208), .ZN(n14692) );
  OR2_X1 U9632 ( .A1(n10199), .A2(n10198), .ZN(n10202) );
  NAND2_X1 U9633 ( .A1(n8692), .A2(n8691), .ZN(n8693) );
  INV_X1 U9634 ( .A(n14724), .ZN(n14705) );
  AND2_X1 U9635 ( .A1(n14733), .A2(n14720), .ZN(n13473) );
  INV_X1 U9636 ( .A(n14715), .ZN(n13426) );
  AND2_X1 U9637 ( .A1(n14769), .A2(n10449), .ZN(n14817) );
  INV_X1 U9638 ( .A(n14817), .ZN(n14809) );
  AND2_X1 U9639 ( .A1(n10849), .A2(n14742), .ZN(n10857) );
  OR2_X1 U9640 ( .A1(n11942), .A2(n13594), .ZN(n8641) );
  INV_X1 U9641 ( .A(n9669), .ZN(n11533) );
  OR2_X1 U9642 ( .A1(n10117), .A2(n10116), .ZN(n13739) );
  INV_X1 U9643 ( .A(n14417), .ZN(n13742) );
  OR2_X1 U9644 ( .A1(n8768), .A2(n13924), .ZN(n9053) );
  AND4_X1 U9645 ( .A1(n8998), .A2(n8997), .A3(n8996), .A4(n8995), .ZN(n13634)
         );
  OR2_X1 U9646 ( .A1(n10377), .A2(n13888), .ZN(n13880) );
  INV_X1 U9647 ( .A(n13880), .ZN(n14462) );
  AND2_X1 U9648 ( .A1(n10391), .A2(n10390), .ZN(n13883) );
  INV_X1 U9649 ( .A(n9375), .ZN(n10758) );
  INV_X1 U9650 ( .A(n14491), .ZN(n14080) );
  INV_X1 U9651 ( .A(n11188), .ZN(n10730) );
  NAND2_X1 U9652 ( .A1(n9105), .A2(n9104), .ZN(n14526) );
  NAND2_X1 U9653 ( .A1(n9154), .A2(n9153), .ZN(n10232) );
  NOR2_X1 U9654 ( .A1(n8831), .A2(n8830), .ZN(n13834) );
  AND2_X1 U9655 ( .A1(n8790), .A2(n8803), .ZN(n10384) );
  AND2_X1 U9656 ( .A1(n10354), .A2(n10353), .ZN(n14969) );
  INV_X1 U9657 ( .A(n12670), .ZN(n12650) );
  INV_X1 U9658 ( .A(n14340), .ZN(n12692) );
  INV_X1 U9659 ( .A(n14969), .ZN(n15000) );
  INV_X1 U9660 ( .A(n14300), .ZN(n14991) );
  NAND2_X1 U9661 ( .A1(n10664), .A2(n15053), .ZN(n15009) );
  NAND2_X1 U9662 ( .A1(n15131), .A2(n15071), .ZN(n13063) );
  AND2_X2 U9663 ( .A1(n7996), .A2(n10662), .ZN(n15131) );
  INV_X1 U9664 ( .A(n7800), .ZN(n13105) );
  NAND2_X1 U9665 ( .A1(n15120), .A2(n15071), .ZN(n13121) );
  AND2_X2 U9666 ( .A1(n8017), .A2(n10029), .ZN(n15120) );
  NAND2_X1 U9667 ( .A1(n13125), .A2(n10168), .ZN(n10169) );
  OR2_X1 U9668 ( .A1(n10339), .A2(P3_U3151), .ZN(n12546) );
  INV_X1 U9669 ( .A(SI_18_), .ZN(n10546) );
  INV_X1 U9670 ( .A(SI_13_), .ZN(n10219) );
  INV_X1 U9671 ( .A(n11677), .ZN(n14947) );
  NAND2_X1 U9672 ( .A1(n10445), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13259) );
  INV_X1 U9673 ( .A(n13257), .ZN(n13272) );
  INV_X1 U9674 ( .A(n12171), .ZN(n13543) );
  INV_X1 U9675 ( .A(n12214), .ZN(n13281) );
  INV_X1 U9676 ( .A(n14685), .ZN(n14620) );
  INV_X1 U9677 ( .A(n14692), .ZN(n14652) );
  OR2_X1 U9678 ( .A1(n10202), .A2(P2_U3088), .ZN(n14647) );
  AND2_X1 U9679 ( .A1(n11315), .A2(n11314), .ZN(n14828) );
  NAND2_X1 U9680 ( .A1(n14733), .A2(n8686), .ZN(n14715) );
  INV_X1 U9681 ( .A(n14853), .ZN(n14850) );
  OR2_X1 U9682 ( .A1(n13545), .A2(n13544), .ZN(n13574) );
  AND2_X1 U9683 ( .A1(n14828), .A2(n14827), .ZN(n14852) );
  INV_X1 U9684 ( .A(n14831), .ZN(n14829) );
  AND2_X2 U9685 ( .A1(n10857), .A2(n14740), .ZN(n14831) );
  OR2_X1 U9686 ( .A1(n14743), .A2(n14737), .ZN(n14738) );
  INV_X1 U9687 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10402) );
  INV_X1 U9688 ( .A(n12069), .ZN(n14167) );
  NAND2_X1 U9689 ( .A1(n10110), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14417) );
  INV_X1 U9690 ( .A(n9170), .ZN(n13747) );
  INV_X1 U9691 ( .A(n12048), .ZN(n13759) );
  INV_X1 U9692 ( .A(n14465), .ZN(n13806) );
  INV_X1 U9693 ( .A(n13883), .ZN(n14468) );
  OR2_X1 U9694 ( .A1(n14491), .A2(n10713), .ZN(n14482) );
  AND2_X1 U9695 ( .A1(n14048), .A2(n14047), .ZN(n14160) );
  INV_X1 U9696 ( .A(n14080), .ZN(n14479) );
  OR2_X1 U9697 ( .A1(n14491), .A2(n10702), .ZN(n11414) );
  AND2_X2 U9698 ( .A1(n9162), .A2(n9161), .ZN(n14560) );
  INV_X1 U9699 ( .A(n14083), .ZN(n14228) );
  INV_X1 U9700 ( .A(n14549), .ZN(n14547) );
  AND2_X1 U9701 ( .A1(n10232), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10188) );
  INV_X1 U9702 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11149) );
  INV_X1 U9703 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10657) );
  XNOR2_X1 U9704 ( .A(n9954), .B(n9953), .ZN(n9955) );
  AND2_X2 U9705 ( .A1(n13125), .A2(n10074), .ZN(P3_U3897) );
  OR4_X1 U9706 ( .A1(n10072), .A2(n10071), .A3(n10070), .A4(n10069), .ZN(
        P3_U3174) );
  NAND2_X1 U9707 ( .A1(n9452), .A2(n7372), .ZN(P3_U3488) );
  NAND2_X1 U9708 ( .A1(n9448), .A2(n7367), .ZN(P3_U3456) );
  AND2_X1 U9709 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10199), .ZN(P2_U3947) );
  OAI21_X1 U9710 ( .B1(n13484), .B2(n14736), .A(n8695), .ZN(P2_U3236) );
  NOR2_X1 U9711 ( .A1(n10077), .A2(n10060), .ZN(P1_U4016) );
  XNOR2_X1 U9712 ( .A(n9956), .B(n9955), .ZN(SUB_1596_U4) );
  INV_X1 U9713 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10145) );
  NAND2_X1 U9714 ( .A1(n10145), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7399) );
  NAND2_X1 U9715 ( .A1(n7400), .A2(n7399), .ZN(n7549) );
  NAND2_X1 U9716 ( .A1(n10178), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7402) );
  INV_X1 U9717 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10131) );
  NAND2_X1 U9718 ( .A1(n10131), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7401) );
  AND2_X1 U9719 ( .A1(n7402), .A2(n7401), .ZN(n7548) );
  NAND2_X1 U9720 ( .A1(n7549), .A2(n7548), .ZN(n7547) );
  NAND2_X1 U9721 ( .A1(n10142), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7404) );
  INV_X1 U9722 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10129) );
  NAND2_X1 U9723 ( .A1(n10129), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7403) );
  NAND2_X1 U9724 ( .A1(n7564), .A2(n7563), .ZN(n7405) );
  NAND2_X1 U9725 ( .A1(n7405), .A2(n7404), .ZN(n7581) );
  NAND2_X1 U9726 ( .A1(n10139), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7407) );
  NAND2_X1 U9727 ( .A1(n10133), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n7406) );
  NAND2_X1 U9728 ( .A1(n7581), .A2(n7580), .ZN(n7408) );
  NAND2_X1 U9729 ( .A1(n10141), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n7410) );
  NAND2_X1 U9730 ( .A1(n10136), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n7409) );
  NAND2_X1 U9731 ( .A1(n7595), .A2(n7594), .ZN(n7411) );
  NAND2_X1 U9732 ( .A1(n7411), .A2(n7410), .ZN(n7615) );
  NAND2_X1 U9733 ( .A1(n10152), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7412) );
  NAND2_X1 U9734 ( .A1(n7615), .A2(n7412), .ZN(n7414) );
  NAND2_X1 U9735 ( .A1(n10180), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n7413) );
  NAND2_X1 U9736 ( .A1(n10165), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7417) );
  NAND2_X1 U9737 ( .A1(n10176), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n7415) );
  INV_X1 U9738 ( .A(n7627), .ZN(n7416) );
  NAND2_X1 U9739 ( .A1(n10171), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n7419) );
  NAND2_X1 U9740 ( .A1(n10174), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n7418) );
  NAND2_X1 U9741 ( .A1(n10192), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n7421) );
  NAND2_X1 U9742 ( .A1(n10191), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n7420) );
  NAND2_X1 U9743 ( .A1(n10221), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n7423) );
  NAND2_X1 U9744 ( .A1(n10223), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n7422) );
  NAND2_X1 U9745 ( .A1(n10237), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n7425) );
  NAND2_X1 U9746 ( .A1(n10236), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n7424) );
  NAND2_X1 U9747 ( .A1(n10323), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n7427) );
  NAND2_X1 U9748 ( .A1(n10322), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n7426) );
  NAND2_X1 U9749 ( .A1(n10597), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n7430) );
  NAND2_X1 U9750 ( .A1(n10599), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n7429) );
  NAND2_X1 U9751 ( .A1(n10657), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n7432) );
  NAND2_X1 U9752 ( .A1(n10656), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n7431) );
  NAND2_X1 U9753 ( .A1(n10571), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n7434) );
  NAND2_X1 U9754 ( .A1(n10570), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n7433) );
  NAND2_X1 U9755 ( .A1(n10673), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n7437) );
  NAND2_X1 U9756 ( .A1(n10672), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n7435) );
  NAND2_X1 U9757 ( .A1(n7437), .A2(n7435), .ZN(n7771) );
  INV_X1 U9758 ( .A(n7771), .ZN(n7436) );
  NAND2_X1 U9759 ( .A1(n10876), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n7439) );
  NAND2_X1 U9760 ( .A1(n10874), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n7438) );
  INV_X1 U9761 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10951) );
  NAND2_X1 U9762 ( .A1(n10951), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n7441) );
  INV_X1 U9763 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10950) );
  NAND2_X1 U9764 ( .A1(n10950), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n7440) );
  INV_X1 U9765 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11250) );
  NAND2_X1 U9766 ( .A1(n11250), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n7815) );
  INV_X1 U9767 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11268) );
  NAND2_X1 U9768 ( .A1(n11268), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n7443) );
  OR2_X1 U9769 ( .A1(n7445), .A2(n7444), .ZN(n7446) );
  NAND2_X1 U9770 ( .A1(n7816), .A2(n7446), .ZN(n10986) );
  NAND4_X1 U9771 ( .A1(n7450), .A2(n7449), .A3(n7448), .A4(n7629), .ZN(n7451)
         );
  NAND2_X1 U9772 ( .A1(n7462), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7464) );
  OR2_X1 U9773 ( .A1(n10986), .A2(n7804), .ZN(n7468) );
  INV_X1 U9774 ( .A(SI_21_), .ZN(n10985) );
  OR2_X1 U9775 ( .A1(n9431), .A2(n10985), .ZN(n7467) );
  NAND2_X1 U9776 ( .A1(n7471), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7472) );
  INV_X1 U9777 ( .A(n7473), .ZN(n13128) );
  NAND2_X1 U9778 ( .A1(n12315), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n7485) );
  AND2_X2 U9779 ( .A1(n7481), .A2(n7480), .ZN(n7529) );
  INV_X1 U9780 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n7476) );
  NOR2_X1 U9781 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7587) );
  NAND2_X1 U9782 ( .A1(n7587), .A2(n7586), .ZN(n7606) );
  NAND2_X1 U9783 ( .A1(n7476), .A2(n7779), .ZN(n7795) );
  INV_X1 U9784 ( .A(n7795), .ZN(n7477) );
  NAND2_X1 U9785 ( .A1(n7809), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n7479) );
  NAND2_X1 U9786 ( .A1(n7820), .A2(n7479), .ZN(n12929) );
  NAND2_X1 U9787 ( .A1(n7529), .A2(n12929), .ZN(n7484) );
  NAND2_X4 U9788 ( .A1(n7475), .A2(n13133), .ZN(n12314) );
  INV_X1 U9789 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13095) );
  OR2_X1 U9790 ( .A1(n12314), .A2(n13095), .ZN(n7483) );
  NAND2_X2 U9791 ( .A1(n7481), .A2(n13133), .ZN(n7542) );
  INV_X2 U9792 ( .A(n9435), .ZN(n12317) );
  INV_X1 U9793 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n12931) );
  OR2_X1 U9794 ( .A1(n12317), .A2(n12931), .ZN(n7482) );
  INV_X1 U9795 ( .A(n12940), .ZN(n12686) );
  NAND2_X1 U9796 ( .A1(n7795), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n7486) );
  NAND2_X1 U9797 ( .A1(n7807), .A2(n7486), .ZN(n12956) );
  NAND2_X1 U9798 ( .A1(n7529), .A2(n12956), .ZN(n7490) );
  NAND2_X1 U9799 ( .A1(n12315), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n7489) );
  INV_X1 U9800 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13103) );
  OR2_X1 U9801 ( .A1(n12314), .A2(n13103), .ZN(n7488) );
  INV_X1 U9802 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12812) );
  OR2_X1 U9803 ( .A1(n7542), .A2(n12812), .ZN(n7487) );
  OR2_X1 U9804 ( .A1(n7492), .A2(n7491), .ZN(n7493) );
  NAND2_X1 U9805 ( .A1(n7494), .A2(n7493), .ZN(n10688) );
  OR2_X1 U9806 ( .A1(n10688), .A2(n7804), .ZN(n7500) );
  NAND2_X1 U9807 ( .A1(n7761), .A2(n7496), .ZN(n7773) );
  OAI21_X2 U9808 ( .B1(n6510), .B2(P3_IR_REG_18__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7498) );
  AOI22_X1 U9809 ( .A1(n12312), .A2(SI_19_), .B1(n12334), .B2(n7790), .ZN(
        n7499) );
  NAND2_X1 U9810 ( .A1(n7500), .A2(n7499), .ZN(n7800) );
  OR2_X1 U9811 ( .A1(n7502), .A2(n7501), .ZN(n7503) );
  NAND2_X1 U9812 ( .A1(n7504), .A2(n7503), .ZN(n10162) );
  NAND2_X1 U9813 ( .A1(n12322), .A2(n10162), .ZN(n7510) );
  OR2_X1 U9814 ( .A1(n9431), .A2(SI_11_), .ZN(n7509) );
  NOR2_X1 U9815 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n7505) );
  NAND2_X1 U9816 ( .A1(n7630), .A2(n7505), .ZN(n7646) );
  OAI21_X1 U9817 ( .B1(n7685), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7507) );
  INV_X1 U9818 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n7506) );
  XNOR2_X1 U9819 ( .A(n7507), .B(n7506), .ZN(n11803) );
  OR2_X1 U9820 ( .A1(n10341), .A2(n11811), .ZN(n7508) );
  NAND2_X1 U9821 ( .A1(n9436), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n7516) );
  NAND2_X1 U9822 ( .A1(n12315), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n7515) );
  NAND2_X1 U9823 ( .A1(n7674), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7511) );
  NAND2_X1 U9824 ( .A1(n7693), .A2(n7511), .ZN(n14335) );
  NAND2_X1 U9825 ( .A1(n7926), .A2(n14335), .ZN(n7514) );
  INV_X1 U9826 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n7512) );
  OR2_X1 U9827 ( .A1(n12317), .A2(n7512), .ZN(n7513) );
  NAND2_X1 U9828 ( .A1(n7529), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n7520) );
  NAND2_X1 U9829 ( .A1(n7540), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7519) );
  NAND2_X1 U9830 ( .A1(n6471), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n7518) );
  INV_X1 U9831 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10326) );
  OR2_X1 U9832 ( .A1(n7542), .A2(n10326), .ZN(n7517) );
  NAND2_X1 U9833 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n7522) );
  INV_X1 U9834 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7521) );
  MUX2_X1 U9835 ( .A(n7522), .B(P3_IR_REG_31__SCAN_IN), .S(n7521), .Z(n7525)
         );
  INV_X1 U9836 ( .A(n10346), .ZN(n7524) );
  INV_X1 U9837 ( .A(SI_1_), .ZN(n10149) );
  OR2_X1 U9838 ( .A1(n7550), .A2(n10149), .ZN(n7528) );
  XNOR2_X1 U9839 ( .A(n7526), .B(n7537), .ZN(n10150) );
  INV_X1 U9840 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10329) );
  NAND2_X1 U9841 ( .A1(n7529), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n7530) );
  INV_X1 U9842 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n7532) );
  NAND2_X1 U9843 ( .A1(n7540), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n7533) );
  INV_X1 U9844 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8747) );
  NAND2_X1 U9845 ( .A1(n8747), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7536) );
  NAND2_X1 U9846 ( .A1(n7537), .A2(n7536), .ZN(n7538) );
  MUX2_X1 U9847 ( .A(n7538), .B(SI_0_), .S(n6706), .Z(n13143) );
  MUX2_X1 U9848 ( .A(n13142), .B(n13143), .S(n10341), .Z(n10668) );
  NAND2_X1 U9849 ( .A1(n15042), .A2(n7539), .ZN(n15043) );
  NAND2_X1 U9850 ( .A1(n15058), .A2(n15043), .ZN(n7556) );
  NAND2_X1 U9851 ( .A1(n7540), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7546) );
  NAND2_X1 U9852 ( .A1(n7529), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n7545) );
  INV_X1 U9853 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n7541) );
  OR2_X1 U9854 ( .A1(n12314), .A2(n7541), .ZN(n7544) );
  INV_X1 U9855 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10331) );
  OR2_X1 U9856 ( .A1(n7542), .A2(n10331), .ZN(n7543) );
  AND4_X2 U9857 ( .A1(n7546), .A2(n7545), .A3(n7544), .A4(n7543), .ZN(n10914)
         );
  OAI21_X1 U9858 ( .B1(n7549), .B2(n7548), .A(n7547), .ZN(n14269) );
  OR2_X1 U9859 ( .A1(n7804), .A2(n14269), .ZN(n7555) );
  OR2_X1 U9860 ( .A1(n7550), .A2(SI_2_), .ZN(n7554) );
  INV_X1 U9861 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7551) );
  OR2_X1 U9862 ( .A1(n10341), .A2(n10347), .ZN(n7553) );
  NAND2_X1 U9863 ( .A1(n10914), .A2(n10493), .ZN(n12346) );
  INV_X1 U9864 ( .A(n10493), .ZN(n15051) );
  NAND2_X1 U9865 ( .A1(n7556), .A2(n7935), .ZN(n15047) );
  NAND2_X1 U9866 ( .A1(n10914), .A2(n15051), .ZN(n7557) );
  NAND2_X1 U9867 ( .A1(n15047), .A2(n7557), .ZN(n10917) );
  INV_X1 U9868 ( .A(n10917), .ZN(n7571) );
  INV_X1 U9869 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n10920) );
  NAND2_X1 U9870 ( .A1(n7529), .A2(n10920), .ZN(n7562) );
  NAND2_X1 U9871 ( .A1(n12315), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n7561) );
  INV_X1 U9872 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n7558) );
  OR2_X1 U9873 ( .A1(n12314), .A2(n7558), .ZN(n7560) );
  INV_X1 U9874 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n11621) );
  OR2_X1 U9875 ( .A1(n12317), .A2(n11621), .ZN(n7559) );
  AND4_X2 U9876 ( .A1(n7562), .A2(n7561), .A3(n7560), .A4(n7559), .ZN(n15041)
         );
  OR2_X1 U9877 ( .A1(n9431), .A2(SI_3_), .ZN(n7569) );
  XNOR2_X1 U9878 ( .A(n7564), .B(n7563), .ZN(n10126) );
  OR2_X1 U9879 ( .A1(n7804), .A2(n10126), .ZN(n7568) );
  INV_X1 U9880 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n7566) );
  NAND2_X1 U9881 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n6525), .ZN(n7565) );
  XNOR2_X1 U9882 ( .A(n7566), .B(n7565), .ZN(n14861) );
  INV_X1 U9883 ( .A(n14861), .ZN(n11668) );
  OR2_X1 U9884 ( .A1(n10341), .A2(n11668), .ZN(n7567) );
  NAND2_X1 U9885 ( .A1(n15041), .A2(n10795), .ZN(n12352) );
  INV_X1 U9886 ( .A(n10795), .ZN(n12358) );
  NAND2_X1 U9887 ( .A1(n12701), .A2(n12358), .ZN(n12350) );
  NAND2_X1 U9888 ( .A1(n7571), .A2(n7570), .ZN(n10915) );
  NAND2_X1 U9889 ( .A1(n12701), .A2(n10795), .ZN(n7572) );
  NAND2_X1 U9890 ( .A1(n9436), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n7576) );
  OR2_X1 U9891 ( .A1(n7386), .A2(n7587), .ZN(n15035) );
  NAND2_X1 U9892 ( .A1(n7926), .A2(n15035), .ZN(n7575) );
  NAND2_X1 U9893 ( .A1(n12315), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7574) );
  INV_X1 U9894 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11627) );
  OR2_X1 U9895 ( .A1(n7542), .A2(n11627), .ZN(n7573) );
  NAND4_X1 U9896 ( .A1(n7576), .A2(n7575), .A3(n7574), .A4(n7573), .ZN(n12700)
         );
  NAND2_X1 U9897 ( .A1(n10346), .A2(n7577), .ZN(n7578) );
  NAND2_X1 U9898 ( .A1(n7578), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7579) );
  XNOR2_X1 U9899 ( .A(n7579), .B(n7447), .ZN(n14878) );
  INV_X1 U9900 ( .A(n14878), .ZN(n11670) );
  XNOR2_X1 U9901 ( .A(n7581), .B(n7580), .ZN(n10155) );
  OR2_X1 U9902 ( .A1(n7804), .A2(n10155), .ZN(n7583) );
  OR2_X1 U9903 ( .A1(n9431), .A2(SI_4_), .ZN(n7582) );
  OAI211_X1 U9904 ( .C1(n11670), .C2(n10341), .A(n7583), .B(n7582), .ZN(n15034) );
  XNOR2_X1 U9905 ( .A(n12700), .B(n15034), .ZN(n15027) );
  NAND2_X1 U9906 ( .A1(n15028), .A2(n15027), .ZN(n7585) );
  INV_X1 U9907 ( .A(n15034), .ZN(n10894) );
  NAND2_X1 U9908 ( .A1(n12700), .A2(n10894), .ZN(n7584) );
  OR2_X1 U9909 ( .A1(n7587), .A2(n7586), .ZN(n7588) );
  NAND2_X1 U9910 ( .A1(n7606), .A2(n7588), .ZN(n15021) );
  NAND2_X1 U9911 ( .A1(n7926), .A2(n15021), .ZN(n7593) );
  NAND2_X1 U9912 ( .A1(n12315), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7592) );
  INV_X1 U9913 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n11632) );
  OR2_X1 U9914 ( .A1(n12317), .A2(n11632), .ZN(n7591) );
  INV_X1 U9915 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n7589) );
  OR2_X1 U9916 ( .A1(n12314), .A2(n7589), .ZN(n7590) );
  OR2_X1 U9917 ( .A1(n9431), .A2(SI_5_), .ZN(n7602) );
  XNOR2_X1 U9918 ( .A(n7595), .B(n7594), .ZN(n10153) );
  OR2_X1 U9919 ( .A1(n7804), .A2(n10153), .ZN(n7601) );
  INV_X1 U9920 ( .A(n7630), .ZN(n7599) );
  NAND2_X1 U9921 ( .A1(n6645), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7597) );
  MUX2_X1 U9922 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7597), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n7598) );
  NAND2_X1 U9923 ( .A1(n7599), .A2(n7598), .ZN(n14895) );
  INV_X1 U9924 ( .A(n14895), .ZN(n11672) );
  OR2_X1 U9925 ( .A1(n10341), .A2(n11672), .ZN(n7600) );
  NAND2_X1 U9926 ( .A1(n15029), .A2(n15020), .ZN(n12369) );
  INV_X1 U9927 ( .A(n15029), .ZN(n12699) );
  INV_X1 U9928 ( .A(n15020), .ZN(n7604) );
  NAND2_X1 U9929 ( .A1(n12699), .A2(n7604), .ZN(n12364) );
  NAND2_X1 U9930 ( .A1(n15029), .A2(n7604), .ZN(n7605) );
  NAND2_X1 U9931 ( .A1(n7606), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7607) );
  NAND2_X1 U9932 ( .A1(n7620), .A2(n7607), .ZN(n11262) );
  NAND2_X1 U9933 ( .A1(n7926), .A2(n11262), .ZN(n7612) );
  NAND2_X1 U9934 ( .A1(n12315), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n7611) );
  INV_X1 U9935 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n7608) );
  OR2_X1 U9936 ( .A1(n12314), .A2(n7608), .ZN(n7610) );
  OR2_X1 U9937 ( .A1(n12317), .A2(n11610), .ZN(n7609) );
  OR2_X1 U9938 ( .A1(n7630), .A2(n7460), .ZN(n7613) );
  XNOR2_X1 U9939 ( .A(n7613), .B(P3_IR_REG_6__SCAN_IN), .ZN(n11674) );
  XNOR2_X1 U9940 ( .A(n10180), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n7614) );
  XNOR2_X1 U9941 ( .A(n7615), .B(n7614), .ZN(n10158) );
  OR2_X1 U9942 ( .A1(n7804), .A2(n10158), .ZN(n7617) );
  INV_X1 U9943 ( .A(SI_6_), .ZN(n10157) );
  OR2_X1 U9944 ( .A1(n9431), .A2(n10157), .ZN(n7616) );
  OAI211_X1 U9945 ( .C1(n10341), .C2(n14913), .A(n7617), .B(n7616), .ZN(n11261) );
  NAND2_X1 U9946 ( .A1(n15018), .A2(n11261), .ZN(n12371) );
  INV_X1 U9947 ( .A(n11261), .ZN(n7618) );
  NAND2_X1 U9948 ( .A1(n12698), .A2(n7618), .ZN(n12377) );
  NAND2_X1 U9949 ( .A1(n11255), .A2(n12507), .ZN(n11254) );
  NAND2_X1 U9950 ( .A1(n12698), .A2(n11261), .ZN(n7619) );
  NAND2_X1 U9951 ( .A1(n11254), .A2(n7619), .ZN(n11227) );
  AND2_X1 U9952 ( .A1(n7620), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7621) );
  OR2_X1 U9953 ( .A1(n7621), .A2(n7640), .ZN(n11234) );
  NAND2_X1 U9954 ( .A1(n7926), .A2(n11234), .ZN(n7626) );
  NAND2_X1 U9955 ( .A1(n12315), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n7625) );
  INV_X1 U9956 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n7622) );
  OR2_X1 U9957 ( .A1(n12314), .A2(n7622), .ZN(n7624) );
  INV_X1 U9958 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11642) );
  OR2_X1 U9959 ( .A1(n12317), .A2(n11642), .ZN(n7623) );
  XNOR2_X1 U9960 ( .A(n7628), .B(n7627), .ZN(n14266) );
  OR2_X1 U9961 ( .A1(n7804), .A2(n14266), .ZN(n7636) );
  OR2_X1 U9962 ( .A1(n9431), .A2(SI_7_), .ZN(n7635) );
  NAND2_X1 U9963 ( .A1(n7630), .A2(n7629), .ZN(n7631) );
  NAND2_X1 U9964 ( .A1(n7631), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7633) );
  INV_X1 U9965 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n7632) );
  XNOR2_X1 U9966 ( .A(n7633), .B(n7632), .ZN(n14930) );
  OR2_X1 U9967 ( .A1(n10341), .A2(n11612), .ZN(n7634) );
  NAND2_X1 U9968 ( .A1(n11354), .A2(n11233), .ZN(n12381) );
  INV_X1 U9969 ( .A(n11354), .ZN(n12697) );
  INV_X1 U9970 ( .A(n11233), .ZN(n12376) );
  NAND2_X1 U9971 ( .A1(n12697), .A2(n12376), .ZN(n7637) );
  NAND2_X1 U9972 ( .A1(n11227), .A2(n11226), .ZN(n7639) );
  NAND2_X1 U9973 ( .A1(n12697), .A2(n11233), .ZN(n7638) );
  NAND2_X1 U9974 ( .A1(n9436), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n7645) );
  NOR2_X1 U9975 ( .A1(n7640), .A2(n11273), .ZN(n7641) );
  OR2_X1 U9976 ( .A1(n7656), .A2(n7641), .ZN(n11269) );
  NAND2_X1 U9977 ( .A1(n7926), .A2(n11269), .ZN(n7644) );
  NAND2_X1 U9978 ( .A1(n12315), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7643) );
  INV_X1 U9979 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11648) );
  OR2_X1 U9980 ( .A1(n7542), .A2(n11648), .ZN(n7642) );
  NAND4_X1 U9981 ( .A1(n7645), .A2(n7644), .A3(n7643), .A4(n7642), .ZN(n12696)
         );
  NAND2_X1 U9982 ( .A1(n7646), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7647) );
  XNOR2_X1 U9983 ( .A(n7647), .B(P3_IR_REG_8__SCAN_IN), .ZN(n11677) );
  INV_X1 U9984 ( .A(SI_8_), .ZN(n10124) );
  OR2_X1 U9985 ( .A1(n9431), .A2(n10124), .ZN(n7653) );
  OR2_X1 U9986 ( .A1(n7649), .A2(n7648), .ZN(n7650) );
  NAND2_X1 U9987 ( .A1(n7651), .A2(n7650), .ZN(n10125) );
  OR2_X1 U9988 ( .A1(n7804), .A2(n10125), .ZN(n7652) );
  OAI211_X1 U9989 ( .C1(n10341), .C2(n14947), .A(n7653), .B(n7652), .ZN(n11360) );
  AND2_X1 U9990 ( .A1(n12696), .A2(n11360), .ZN(n7654) );
  NAND2_X1 U9991 ( .A1(n9436), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n7661) );
  NAND2_X1 U9992 ( .A1(n12315), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n7660) );
  OR2_X1 U9993 ( .A1(n7656), .A2(n7655), .ZN(n7657) );
  AND2_X1 U9994 ( .A1(n7672), .A2(n7657), .ZN(n15010) );
  INV_X1 U9995 ( .A(n15010), .ZN(n11390) );
  NAND2_X1 U9996 ( .A1(n7926), .A2(n11390), .ZN(n7659) );
  INV_X1 U9997 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11652) );
  OR2_X1 U9998 ( .A1(n12317), .A2(n11652), .ZN(n7658) );
  NAND4_X1 U9999 ( .A1(n7661), .A2(n7660), .A3(n7659), .A4(n7658), .ZN(n12695)
         );
  OR2_X1 U10000 ( .A1(n7663), .A2(n7662), .ZN(n7664) );
  AND2_X1 U10001 ( .A1(n7665), .A2(n7664), .ZN(n10159) );
  OR2_X1 U10002 ( .A1(n7804), .A2(n10159), .ZN(n7671) );
  OR2_X1 U10003 ( .A1(n9431), .A2(SI_9_), .ZN(n7670) );
  NAND2_X1 U10004 ( .A1(n7666), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7667) );
  MUX2_X1 U10005 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7667), .S(
        P3_IR_REG_9__SCAN_IN), .Z(n7668) );
  NAND2_X1 U10006 ( .A1(n7668), .A2(n7685), .ZN(n14965) );
  OR2_X1 U10007 ( .A1(n10341), .A2(n11615), .ZN(n7669) );
  XNOR2_X1 U10008 ( .A(n12695), .B(n15003), .ZN(n12511) );
  NAND2_X1 U10009 ( .A1(n7672), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7673) );
  NAND2_X1 U10010 ( .A1(n7674), .A2(n7673), .ZN(n11492) );
  NAND2_X1 U10011 ( .A1(n7926), .A2(n11492), .ZN(n7679) );
  NAND2_X1 U10012 ( .A1(n12315), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7678) );
  INV_X1 U10013 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11658) );
  OR2_X1 U10014 ( .A1(n7542), .A2(n11658), .ZN(n7677) );
  INV_X1 U10015 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n7675) );
  OR2_X1 U10016 ( .A1(n12314), .A2(n7675), .ZN(n7676) );
  OR2_X1 U10017 ( .A1(n7681), .A2(n7680), .ZN(n7682) );
  AND2_X1 U10018 ( .A1(n7683), .A2(n7682), .ZN(n10146) );
  OR2_X1 U10019 ( .A1(n7804), .A2(n10146), .ZN(n7689) );
  OR2_X1 U10020 ( .A1(n9431), .A2(SI_10_), .ZN(n7688) );
  NAND2_X1 U10021 ( .A1(n7685), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7686) );
  INV_X1 U10022 ( .A(n11665), .ZN(n14995) );
  OR2_X1 U10023 ( .A1(n10341), .A2(n14995), .ZN(n7687) );
  NAND2_X1 U10024 ( .A1(n14342), .A2(n11593), .ZN(n12395) );
  INV_X1 U10025 ( .A(n11593), .ZN(n15114) );
  NAND2_X1 U10026 ( .A1(n12694), .A2(n15114), .ZN(n7938) );
  NAND2_X1 U10027 ( .A1(n12395), .A2(n7938), .ZN(n12505) );
  NAND2_X1 U10028 ( .A1(n12694), .A2(n11593), .ZN(n7690) );
  OAI21_X1 U10029 ( .B1(n14334), .B2(n12693), .A(n14338), .ZN(n7692) );
  INV_X1 U10030 ( .A(n14334), .ZN(n9983) );
  NAND2_X1 U10031 ( .A1(n12693), .A2(n14334), .ZN(n7691) );
  AND2_X1 U10032 ( .A1(n7693), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7694) );
  OR2_X1 U10033 ( .A1(n7694), .A2(n7720), .ZN(n11898) );
  NAND2_X1 U10034 ( .A1(n7529), .A2(n11898), .ZN(n7700) );
  NAND2_X1 U10035 ( .A1(n12315), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n7699) );
  INV_X1 U10036 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n7695) );
  OR2_X1 U10037 ( .A1(n12314), .A2(n7695), .ZN(n7698) );
  INV_X1 U10038 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n7696) );
  OR2_X1 U10039 ( .A1(n7542), .A2(n7696), .ZN(n7697) );
  OR2_X1 U10040 ( .A1(n7702), .A2(n7701), .ZN(n7703) );
  NAND2_X1 U10041 ( .A1(n7704), .A2(n7703), .ZN(n10166) );
  OR2_X1 U10042 ( .A1(n10166), .A2(n7804), .ZN(n7708) );
  OR2_X1 U10043 ( .A1(n7705), .A2(n7460), .ZN(n7706) );
  XNOR2_X1 U10044 ( .A(n7706), .B(P3_IR_REG_12__SCAN_IN), .ZN(n12706) );
  AOI22_X1 U10045 ( .A1(n12312), .A2(SI_12_), .B1(n7790), .B2(n12706), .ZN(
        n7707) );
  NAND2_X1 U10046 ( .A1(n7708), .A2(n7707), .ZN(n11908) );
  NAND2_X1 U10047 ( .A1(n14340), .A2(n11908), .ZN(n12406) );
  INV_X1 U10048 ( .A(n11908), .ZN(n14359) );
  NAND2_X1 U10049 ( .A1(n12692), .A2(n14359), .ZN(n12404) );
  NAND2_X1 U10050 ( .A1(n12406), .A2(n12404), .ZN(n12514) );
  NAND2_X1 U10051 ( .A1(n7710), .A2(n10402), .ZN(n7711) );
  NAND2_X1 U10052 ( .A1(n7712), .A2(n7711), .ZN(n10218) );
  NAND2_X1 U10053 ( .A1(n10218), .A2(n12322), .ZN(n7718) );
  NAND2_X1 U10054 ( .A1(n7713), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7714) );
  MUX2_X1 U10055 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7714), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n7716) );
  NAND2_X1 U10056 ( .A1(n7716), .A2(n7715), .ZN(n12727) );
  AOI22_X1 U10057 ( .A1(n12312), .A2(n10219), .B1(n7790), .B2(n12727), .ZN(
        n7717) );
  NAND2_X1 U10058 ( .A1(n7718), .A2(n7717), .ZN(n14353) );
  NAND2_X1 U10059 ( .A1(n9436), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n7726) );
  NAND2_X1 U10060 ( .A1(n12315), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n7725) );
  NOR2_X1 U10061 ( .A1(n7720), .A2(n7719), .ZN(n7721) );
  OR2_X1 U10062 ( .A1(n7734), .A2(n7721), .ZN(n11913) );
  NAND2_X1 U10063 ( .A1(n7529), .A2(n11913), .ZN(n7724) );
  INV_X1 U10064 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n7722) );
  OR2_X1 U10065 ( .A1(n12317), .A2(n7722), .ZN(n7723) );
  NAND4_X1 U10066 ( .A1(n7726), .A2(n7725), .A3(n7724), .A4(n7723), .ZN(n12691) );
  OR2_X1 U10067 ( .A1(n14353), .A2(n12691), .ZN(n12408) );
  NAND2_X1 U10068 ( .A1(n14353), .A2(n12691), .ZN(n12407) );
  INV_X1 U10069 ( .A(n12691), .ZN(n14328) );
  OR2_X1 U10070 ( .A1(n7728), .A2(n7727), .ZN(n7729) );
  NAND2_X1 U10071 ( .A1(n7730), .A2(n7729), .ZN(n10278) );
  NAND2_X1 U10072 ( .A1(n10278), .A2(n12322), .ZN(n7733) );
  INV_X1 U10073 ( .A(SI_14_), .ZN(n10279) );
  NAND2_X1 U10074 ( .A1(n7715), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7731) );
  XNOR2_X1 U10075 ( .A(n7731), .B(n6634), .ZN(n12734) );
  AOI22_X1 U10076 ( .A1(n12312), .A2(n10279), .B1(n7790), .B2(n12734), .ZN(
        n7732) );
  NAND2_X1 U10077 ( .A1(n7733), .A2(n7732), .ZN(n14330) );
  NAND2_X1 U10078 ( .A1(n9436), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n7740) );
  NAND2_X1 U10079 ( .A1(n12315), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n7739) );
  NOR2_X1 U10080 ( .A1(n7734), .A2(n11934), .ZN(n7735) );
  OR2_X1 U10081 ( .A1(n7751), .A2(n7735), .ZN(n14331) );
  NAND2_X1 U10082 ( .A1(n7529), .A2(n14331), .ZN(n7738) );
  INV_X1 U10083 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n7736) );
  OR2_X1 U10084 ( .A1(n7542), .A2(n7736), .ZN(n7737) );
  NAND4_X1 U10085 ( .A1(n7740), .A2(n7739), .A3(n7738), .A4(n7737), .ZN(n12690) );
  OR2_X1 U10086 ( .A1(n14330), .A2(n12690), .ZN(n12412) );
  NAND2_X1 U10087 ( .A1(n14330), .A2(n12690), .ZN(n12413) );
  NAND2_X1 U10088 ( .A1(n12412), .A2(n12413), .ZN(n14325) );
  INV_X1 U10089 ( .A(n14330), .ZN(n9989) );
  OR2_X1 U10090 ( .A1(n7742), .A2(n7741), .ZN(n7743) );
  NAND2_X1 U10091 ( .A1(n7744), .A2(n7743), .ZN(n10319) );
  OR2_X1 U10092 ( .A1(n10319), .A2(n7804), .ZN(n7749) );
  NAND2_X1 U10093 ( .A1(n7745), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7747) );
  XNOR2_X1 U10094 ( .A(n7747), .B(n7746), .ZN(n12795) );
  INV_X1 U10095 ( .A(n12795), .ZN(n12774) );
  AOI22_X1 U10096 ( .A1(n12312), .A2(SI_15_), .B1(n7790), .B2(n12774), .ZN(
        n7748) );
  NAND2_X1 U10097 ( .A1(n7749), .A2(n7748), .ZN(n9993) );
  NAND2_X1 U10098 ( .A1(n12315), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n7756) );
  OR2_X1 U10099 ( .A1(n7751), .A2(n7750), .ZN(n7752) );
  NAND2_X1 U10100 ( .A1(n7765), .A2(n7752), .ZN(n13005) );
  NAND2_X1 U10101 ( .A1(n7529), .A2(n13005), .ZN(n7755) );
  INV_X1 U10102 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13119) );
  OR2_X1 U10103 ( .A1(n12314), .A2(n13119), .ZN(n7754) );
  INV_X1 U10104 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12754) );
  OR2_X1 U10105 ( .A1(n12317), .A2(n12754), .ZN(n7753) );
  OR2_X1 U10106 ( .A1(n9993), .A2(n14329), .ZN(n12417) );
  NAND2_X1 U10107 ( .A1(n9993), .A2(n14329), .ZN(n12422) );
  OR2_X1 U10108 ( .A1(n7758), .A2(n7757), .ZN(n7759) );
  NAND2_X1 U10109 ( .A1(n7760), .A2(n7759), .ZN(n10368) );
  OR2_X1 U10110 ( .A1(n10368), .A2(n7804), .ZN(n7764) );
  OR2_X1 U10111 ( .A1(n7761), .A2(n7460), .ZN(n7762) );
  XNOR2_X1 U10112 ( .A(n7762), .B(P3_IR_REG_16__SCAN_IN), .ZN(n14289) );
  AOI22_X1 U10113 ( .A1(n12312), .A2(SI_16_), .B1(n7790), .B2(n14289), .ZN(
        n7763) );
  NAND2_X1 U10114 ( .A1(n12315), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n7770) );
  NAND2_X1 U10115 ( .A1(n7765), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n7766) );
  NAND2_X1 U10116 ( .A1(n7778), .A2(n7766), .ZN(n12993) );
  NAND2_X1 U10117 ( .A1(n7529), .A2(n12993), .ZN(n7769) );
  INV_X1 U10118 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13115) );
  OR2_X1 U10119 ( .A1(n12314), .A2(n13115), .ZN(n7768) );
  INV_X1 U10120 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12784) );
  OR2_X1 U10121 ( .A1(n12317), .A2(n12784), .ZN(n7767) );
  OR2_X1 U10122 ( .A1(n12992), .A2(n13001), .ZN(n12424) );
  NAND2_X1 U10123 ( .A1(n12992), .A2(n13001), .ZN(n12423) );
  NAND2_X1 U10124 ( .A1(n12424), .A2(n12423), .ZN(n12986) );
  INV_X1 U10125 ( .A(n13001), .ZN(n12689) );
  XNOR2_X1 U10126 ( .A(n7772), .B(n7771), .ZN(n10438) );
  NAND2_X1 U10127 ( .A1(n10438), .A2(n12322), .ZN(n7777) );
  NAND2_X1 U10128 ( .A1(n7773), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7774) );
  MUX2_X1 U10129 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7774), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n7775) );
  NAND2_X1 U10130 ( .A1(n7775), .A2(n6510), .ZN(n12798) );
  INV_X1 U10131 ( .A(n12798), .ZN(n14312) );
  AOI22_X1 U10132 ( .A1(n12312), .A2(SI_17_), .B1(n7790), .B2(n14312), .ZN(
        n7776) );
  NAND2_X1 U10133 ( .A1(n7777), .A2(n7776), .ZN(n9998) );
  NAND2_X1 U10134 ( .A1(n7778), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n7780) );
  INV_X1 U10135 ( .A(n7779), .ZN(n7793) );
  NAND2_X1 U10136 ( .A1(n7780), .A2(n7793), .ZN(n12981) );
  NAND2_X1 U10137 ( .A1(n7529), .A2(n12981), .ZN(n7784) );
  NAND2_X1 U10138 ( .A1(n12315), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n7783) );
  INV_X1 U10139 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13111) );
  OR2_X1 U10140 ( .A1(n12314), .A2(n13111), .ZN(n7782) );
  INV_X1 U10141 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14309) );
  OR2_X1 U10142 ( .A1(n7542), .A2(n14309), .ZN(n7781) );
  OR2_X1 U10143 ( .A1(n9998), .A2(n12989), .ZN(n12430) );
  NAND2_X1 U10144 ( .A1(n9998), .A2(n12989), .ZN(n12427) );
  OR2_X1 U10145 ( .A1(n7786), .A2(n7785), .ZN(n7787) );
  NAND2_X1 U10146 ( .A1(n7788), .A2(n7787), .ZN(n10545) );
  OR2_X1 U10147 ( .A1(n10545), .A2(n7804), .ZN(n7792) );
  NAND2_X1 U10148 ( .A1(n6510), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7789) );
  XNOR2_X1 U10149 ( .A(n7789), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12824) );
  AOI22_X1 U10150 ( .A1(n12312), .A2(SI_18_), .B1(n7790), .B2(n12824), .ZN(
        n7791) );
  NAND2_X1 U10151 ( .A1(n7792), .A2(n7791), .ZN(n10005) );
  NAND2_X1 U10152 ( .A1(n12315), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n7799) );
  NAND2_X1 U10153 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(n7793), .ZN(n7794) );
  NAND2_X1 U10154 ( .A1(n7795), .A2(n7794), .ZN(n12971) );
  NAND2_X1 U10155 ( .A1(n7529), .A2(n12971), .ZN(n7798) );
  INV_X1 U10156 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13107) );
  OR2_X1 U10157 ( .A1(n12314), .A2(n13107), .ZN(n7797) );
  INV_X1 U10158 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12786) );
  OR2_X1 U10159 ( .A1(n12317), .A2(n12786), .ZN(n7796) );
  OR2_X1 U10160 ( .A1(n10005), .A2(n12978), .ZN(n12428) );
  NAND2_X1 U10161 ( .A1(n10005), .A2(n12978), .ZN(n12433) );
  OR2_X1 U10162 ( .A1(n7800), .A2(n12966), .ZN(n12438) );
  NAND2_X1 U10163 ( .A1(n7800), .A2(n12966), .ZN(n12439) );
  NAND2_X1 U10164 ( .A1(n12438), .A2(n12439), .ZN(n12951) );
  NAND2_X1 U10165 ( .A1(n7801), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7802) );
  NAND2_X1 U10166 ( .A1(n7803), .A2(n7802), .ZN(n10900) );
  OR2_X1 U10167 ( .A1(n10900), .A2(n7804), .ZN(n7806) );
  OR2_X1 U10168 ( .A1(n9431), .A2(n10899), .ZN(n7805) );
  NAND2_X1 U10169 ( .A1(n7807), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n7808) );
  NAND2_X1 U10170 ( .A1(n7809), .A2(n7808), .ZN(n12944) );
  NAND2_X1 U10171 ( .A1(n7529), .A2(n12944), .ZN(n7814) );
  NAND2_X1 U10172 ( .A1(n12315), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n7813) );
  INV_X1 U10173 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n7810) );
  OR2_X1 U10174 ( .A1(n7542), .A2(n7810), .ZN(n7812) );
  INV_X1 U10175 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13099) );
  OR2_X1 U10176 ( .A1(n12314), .A2(n13099), .ZN(n7811) );
  NAND2_X1 U10177 ( .A1(n12943), .A2(n12955), .ZN(n12443) );
  NAND2_X1 U10178 ( .A1(n12442), .A2(n12443), .ZN(n12937) );
  NAND2_X1 U10179 ( .A1(n13033), .A2(n12940), .ZN(n12447) );
  NAND2_X1 U10180 ( .A1(n12446), .A2(n12447), .ZN(n12933) );
  NAND2_X1 U10181 ( .A1(n12925), .A2(n12933), .ZN(n12924) );
  INV_X1 U10182 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7828) );
  XNOR2_X1 U10183 ( .A(n7828), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n7830) );
  XNOR2_X1 U10184 ( .A(n7831), .B(n7830), .ZN(n11063) );
  NAND2_X1 U10185 ( .A1(n11063), .A2(n12322), .ZN(n7819) );
  INV_X1 U10186 ( .A(SI_22_), .ZN(n7817) );
  OR2_X1 U10187 ( .A1(n9431), .A2(n7817), .ZN(n7818) );
  NAND2_X1 U10188 ( .A1(n9435), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n7825) );
  NAND2_X1 U10189 ( .A1(n7820), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n7821) );
  NAND2_X1 U10190 ( .A1(n7835), .A2(n7821), .ZN(n12919) );
  NAND2_X1 U10191 ( .A1(n7529), .A2(n12919), .ZN(n7824) );
  NAND2_X1 U10192 ( .A1(n12315), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n7823) );
  INV_X1 U10193 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13091) );
  OR2_X1 U10194 ( .A1(n12314), .A2(n13091), .ZN(n7822) );
  NAND4_X1 U10195 ( .A1(n7825), .A2(n7824), .A3(n7823), .A4(n7822), .ZN(n12927) );
  NAND2_X1 U10196 ( .A1(n12918), .A2(n12927), .ZN(n7827) );
  NOR2_X1 U10197 ( .A1(n12918), .A2(n12927), .ZN(n7826) );
  NAND2_X1 U10198 ( .A1(n7828), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n7829) );
  XNOR2_X1 U10199 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n7842) );
  XNOR2_X1 U10200 ( .A(n7843), .B(n7842), .ZN(n11286) );
  NAND2_X1 U10201 ( .A1(n11286), .A2(n12322), .ZN(n7833) );
  OR2_X1 U10202 ( .A1(n9431), .A2(n11288), .ZN(n7832) );
  NAND2_X1 U10203 ( .A1(n7835), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n7836) );
  NAND2_X1 U10204 ( .A1(n7849), .A2(n7836), .ZN(n12905) );
  NAND2_X1 U10205 ( .A1(n7529), .A2(n12905), .ZN(n7840) );
  NAND2_X1 U10206 ( .A1(n12315), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n7839) );
  INV_X1 U10207 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n12907) );
  OR2_X1 U10208 ( .A1(n7542), .A2(n12907), .ZN(n7838) );
  INV_X1 U10209 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13087) );
  OR2_X1 U10210 ( .A1(n12314), .A2(n13087), .ZN(n7837) );
  XNOR2_X1 U10211 ( .A(n13024), .B(n12915), .ZN(n12901) );
  NAND2_X1 U10212 ( .A1(n12902), .A2(n12901), .ZN(n12900) );
  NAND2_X1 U10213 ( .A1(n13024), .A2(n12685), .ZN(n7841) );
  INV_X1 U10214 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7844) );
  NAND2_X1 U10215 ( .A1(n7844), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7845) );
  INV_X1 U10216 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11943) );
  INV_X1 U10217 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11940) );
  XNOR2_X1 U10218 ( .A(n7858), .B(n11940), .ZN(n11466) );
  NAND2_X1 U10219 ( .A1(n11466), .A2(n12322), .ZN(n7848) );
  OR2_X1 U10220 ( .A1(n9431), .A2(n6810), .ZN(n7847) );
  NAND2_X2 U10221 ( .A1(n7848), .A2(n7847), .ZN(n13020) );
  NAND2_X1 U10222 ( .A1(n12315), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n7856) );
  NAND2_X1 U10223 ( .A1(n7849), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n7850) );
  NAND2_X1 U10224 ( .A1(n7864), .A2(n7850), .ZN(n12892) );
  NAND2_X1 U10225 ( .A1(n7926), .A2(n12892), .ZN(n7855) );
  INV_X1 U10226 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n7851) );
  OR2_X1 U10227 ( .A1(n12314), .A2(n7851), .ZN(n7854) );
  INV_X1 U10228 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n7852) );
  OR2_X1 U10229 ( .A1(n7542), .A2(n7852), .ZN(n7853) );
  NAND2_X1 U10230 ( .A1(n13020), .A2(n6647), .ZN(n7857) );
  INV_X1 U10231 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n11977) );
  XNOR2_X1 U10232 ( .A(n11977), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n7860) );
  XNOR2_X1 U10233 ( .A(n7872), .B(n7860), .ZN(n11690) );
  NAND2_X1 U10234 ( .A1(n11690), .A2(n12322), .ZN(n7862) );
  INV_X1 U10235 ( .A(SI_25_), .ZN(n11691) );
  NAND2_X1 U10236 ( .A1(n7864), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n7865) );
  NAND2_X1 U10237 ( .A1(n7891), .A2(n7865), .ZN(n12875) );
  NAND2_X1 U10238 ( .A1(n7926), .A2(n12875), .ZN(n7870) );
  NAND2_X1 U10239 ( .A1(n12315), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n7869) );
  INV_X1 U10240 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n7866) );
  OR2_X1 U10241 ( .A1(n7542), .A2(n7866), .ZN(n7868) );
  INV_X1 U10242 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13082) );
  OR2_X1 U10243 ( .A1(n12314), .A2(n13082), .ZN(n7867) );
  XNOR2_X1 U10244 ( .A(n12592), .B(n12885), .ZN(n12868) );
  INV_X1 U10245 ( .A(n12885), .ZN(n12684) );
  NAND2_X1 U10246 ( .A1(n12592), .A2(n12684), .ZN(n8002) );
  NAND2_X1 U10247 ( .A1(n11977), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n7871) );
  NAND2_X1 U10248 ( .A1(n7872), .A2(n7871), .ZN(n7874) );
  INV_X1 U10249 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n11978) );
  NAND2_X1 U10250 ( .A1(n11978), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n7873) );
  INV_X1 U10251 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7885) );
  XNOR2_X1 U10252 ( .A(n7885), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n7875) );
  XNOR2_X1 U10253 ( .A(n7884), .B(n7875), .ZN(n11768) );
  NAND2_X1 U10254 ( .A1(n11768), .A2(n12322), .ZN(n7877) );
  INV_X1 U10255 ( .A(SI_26_), .ZN(n11770) );
  OR2_X1 U10256 ( .A1(n9431), .A2(n11770), .ZN(n7876) );
  XNOR2_X1 U10257 ( .A(n7891), .B(P3_REG3_REG_26__SCAN_IN), .ZN(n12860) );
  NAND2_X1 U10258 ( .A1(n7926), .A2(n12860), .ZN(n7882) );
  NAND2_X1 U10259 ( .A1(n12315), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n7881) );
  INV_X1 U10260 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n8018) );
  OR2_X1 U10261 ( .A1(n12314), .A2(n8018), .ZN(n7880) );
  INV_X1 U10262 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n7878) );
  OR2_X1 U10263 ( .A1(n7542), .A2(n7878), .ZN(n7879) );
  NAND2_X1 U10264 ( .A1(n7949), .A2(n12870), .ZN(n7883) );
  AND2_X1 U10265 ( .A1(n8002), .A2(n7883), .ZN(n8026) );
  INV_X1 U10266 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14249) );
  NAND2_X1 U10267 ( .A1(n7885), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n7886) );
  XNOR2_X1 U10268 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n7887) );
  XNOR2_X1 U10269 ( .A(n7899), .B(n7887), .ZN(n11886) );
  NAND2_X1 U10270 ( .A1(n11886), .A2(n12322), .ZN(n7889) );
  INV_X1 U10271 ( .A(SI_27_), .ZN(n11887) );
  NAND2_X2 U10272 ( .A1(n7889), .A2(n7888), .ZN(n12856) );
  OAI21_X1 U10273 ( .B1(n7891), .B2(P3_REG3_REG_26__SCAN_IN), .A(
        P3_REG3_REG_27__SCAN_IN), .ZN(n7892) );
  INV_X1 U10274 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n9829) );
  INV_X1 U10275 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n9854) );
  NAND2_X1 U10276 ( .A1(n9829), .A2(n9854), .ZN(n7890) );
  NAND2_X1 U10277 ( .A1(n7892), .A2(n7905), .ZN(n12849) );
  NAND2_X1 U10278 ( .A1(n7926), .A2(n12849), .ZN(n7896) );
  NAND2_X1 U10279 ( .A1(n12315), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n7895) );
  INV_X1 U10280 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n13078) );
  OR2_X1 U10281 ( .A1(n12314), .A2(n13078), .ZN(n7894) );
  INV_X1 U10282 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n12851) );
  OR2_X1 U10283 ( .A1(n12317), .A2(n12851), .ZN(n7893) );
  OR2_X1 U10284 ( .A1(n12856), .A2(n12666), .ZN(n12477) );
  NAND2_X1 U10285 ( .A1(n12856), .A2(n12666), .ZN(n12470) );
  AND2_X2 U10286 ( .A1(n12477), .A2(n12470), .ZN(n12526) );
  INV_X1 U10287 ( .A(n12526), .ZN(n8030) );
  AND2_X1 U10288 ( .A1(n8026), .A2(n8030), .ZN(n7897) );
  NAND2_X1 U10289 ( .A1(n12862), .A2(n7948), .ZN(n8027) );
  NAND2_X1 U10290 ( .A1(n13080), .A2(n12666), .ZN(n7923) );
  NAND2_X1 U10291 ( .A1(n8029), .A2(n7923), .ZN(n7922) );
  INV_X1 U10292 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13590) );
  AND2_X1 U10293 ( .A1(n13590), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n7898) );
  INV_X1 U10294 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14246) );
  INV_X1 U10295 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9428) );
  XNOR2_X1 U10296 ( .A(n9428), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n7900) );
  XNOR2_X1 U10297 ( .A(n9427), .B(n7900), .ZN(n13136) );
  NAND2_X1 U10298 ( .A1(n13136), .A2(n12322), .ZN(n7902) );
  INV_X1 U10299 ( .A(SI_28_), .ZN(n13141) );
  OR2_X1 U10300 ( .A1(n9431), .A2(n13141), .ZN(n7901) );
  INV_X1 U10301 ( .A(n7905), .ZN(n7904) );
  INV_X1 U10302 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n7903) );
  NAND2_X1 U10303 ( .A1(n7904), .A2(n7903), .ZN(n12548) );
  NAND2_X1 U10304 ( .A1(n7905), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n7906) );
  NAND2_X1 U10305 ( .A1(n12548), .A2(n7906), .ZN(n12841) );
  NAND2_X1 U10306 ( .A1(n7926), .A2(n12841), .ZN(n7911) );
  NAND2_X1 U10307 ( .A1(n12315), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n7910) );
  INV_X1 U10308 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n12843) );
  OR2_X1 U10309 ( .A1(n7542), .A2(n12843), .ZN(n7909) );
  INV_X1 U10310 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n7907) );
  OR2_X1 U10311 ( .A1(n12314), .A2(n7907), .ZN(n7908) );
  NAND2_X1 U10312 ( .A1(n7997), .A2(n12560), .ZN(n12469) );
  NAND2_X1 U10313 ( .A1(n7978), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7914) );
  NAND2_X1 U10314 ( .A1(n12334), .A2(n12543), .ZN(n7921) );
  INV_X1 U10315 ( .A(n7915), .ZN(n7916) );
  NAND2_X1 U10316 ( .A1(n7916), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7917) );
  XNOR2_X2 U10317 ( .A(n7917), .B(P3_IR_REG_21__SCAN_IN), .ZN(n12337) );
  NAND2_X1 U10318 ( .A1(n7918), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7920) );
  INV_X1 U10319 ( .A(n10898), .ZN(n7959) );
  NAND2_X1 U10320 ( .A1(n12337), .A2(n7959), .ZN(n12336) );
  AOI21_X1 U10321 ( .B1(n7922), .B2(n12479), .A(n15045), .ZN(n7934) );
  INV_X1 U10322 ( .A(n12479), .ZN(n12527) );
  AND2_X1 U10323 ( .A1(n7923), .A2(n12527), .ZN(n7924) );
  NAND2_X1 U10324 ( .A1(n8029), .A2(n7924), .ZN(n9425) );
  INV_X1 U10325 ( .A(n12548), .ZN(n7925) );
  NAND2_X1 U10326 ( .A1(n7926), .A2(n7925), .ZN(n12321) );
  NAND2_X1 U10327 ( .A1(n9436), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n7929) );
  NAND2_X1 U10328 ( .A1(n12315), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n7928) );
  NAND2_X1 U10329 ( .A1(n9435), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n7927) );
  INV_X1 U10330 ( .A(n13139), .ZN(n10342) );
  NAND2_X1 U10331 ( .A1(n10342), .A2(n12820), .ZN(n10343) );
  NAND2_X1 U10332 ( .A1(n10341), .A2(n10343), .ZN(n7932) );
  AND2_X4 U10333 ( .A1(n12543), .A2(n12337), .ZN(n12496) );
  OAI22_X1 U10334 ( .A1(n11029), .A2(n14339), .B1(n12666), .B2(n14341), .ZN(
        n7933) );
  AOI21_X1 U10335 ( .B1(n7934), .B2(n9425), .A(n7933), .ZN(n12848) );
  INV_X1 U10336 ( .A(n10668), .ZN(n10600) );
  NOR2_X2 U10337 ( .A1(n10404), .A2(n10600), .ZN(n15067) );
  NAND2_X1 U10338 ( .A1(n10522), .A2(n12348), .ZN(n15040) );
  NAND2_X1 U10339 ( .A1(n15040), .A2(n15044), .ZN(n15039) );
  NAND2_X1 U10340 ( .A1(n10913), .A2(n12509), .ZN(n7936) );
  NAND2_X1 U10341 ( .A1(n7936), .A2(n12352), .ZN(n15026) );
  INV_X1 U10342 ( .A(n15027), .ZN(n15025) );
  NAND2_X1 U10343 ( .A1(n15026), .A2(n15025), .ZN(n15024) );
  NAND2_X1 U10344 ( .A1(n15017), .A2(n10894), .ZN(n12361) );
  NAND2_X1 U10345 ( .A1(n15011), .A2(n15015), .ZN(n7937) );
  INV_X1 U10346 ( .A(n12507), .ZN(n11252) );
  INV_X1 U10347 ( .A(n11226), .ZN(n12504) );
  NAND2_X1 U10348 ( .A1(n11228), .A2(n12381), .ZN(n11350) );
  NAND2_X1 U10349 ( .A1(n11388), .A2(n11360), .ZN(n12382) );
  INV_X1 U10350 ( .A(n11360), .ZN(n15108) );
  NAND2_X1 U10351 ( .A1(n12696), .A2(n15108), .ZN(n12383) );
  NAND2_X1 U10352 ( .A1(n11586), .A2(n7938), .ZN(n7939) );
  NAND2_X1 U10353 ( .A1(n11825), .A2(n14334), .ZN(n12397) );
  NAND2_X1 U10354 ( .A1(n12693), .A2(n9983), .ZN(n12402) );
  NAND2_X1 U10355 ( .A1(n14336), .A2(n14337), .ZN(n7940) );
  NAND2_X1 U10356 ( .A1(n7940), .A2(n12397), .ZN(n11828) );
  INV_X1 U10357 ( .A(n12514), .ZN(n11827) );
  INV_X1 U10358 ( .A(n12408), .ZN(n7941) );
  NAND2_X1 U10359 ( .A1(n13004), .A2(n13003), .ZN(n13002) );
  NAND2_X1 U10360 ( .A1(n13002), .A2(n12422), .ZN(n12991) );
  INV_X1 U10361 ( .A(n12986), .ZN(n12990) );
  NAND2_X1 U10362 ( .A1(n12991), .A2(n12990), .ZN(n7942) );
  NAND2_X1 U10363 ( .A1(n7942), .A2(n12423), .ZN(n12979) );
  NAND2_X1 U10364 ( .A1(n12979), .A2(n12980), .ZN(n7943) );
  NAND2_X1 U10365 ( .A1(n7944), .A2(n12438), .ZN(n7945) );
  NAND2_X1 U10366 ( .A1(n7945), .A2(n12439), .ZN(n12942) );
  INV_X1 U10367 ( .A(n12927), .ZN(n12588) );
  NAND2_X1 U10368 ( .A1(n12918), .A2(n12588), .ZN(n12452) );
  OR2_X1 U10369 ( .A1(n12918), .A2(n12588), .ZN(n12451) );
  NAND2_X1 U10370 ( .A1(n7946), .A2(n12451), .ZN(n12898) );
  INV_X1 U10371 ( .A(n12901), .ZN(n12897) );
  OR2_X1 U10372 ( .A1(n13024), .A2(n12915), .ZN(n12881) );
  NAND2_X1 U10373 ( .A1(n12880), .A2(n12463), .ZN(n12883) );
  NAND2_X1 U10374 ( .A1(n13020), .A2(n12601), .ZN(n12461) );
  NAND2_X1 U10375 ( .A1(n12883), .A2(n12461), .ZN(n12874) );
  NAND2_X1 U10376 ( .A1(n12874), .A2(n12873), .ZN(n7947) );
  NAND2_X1 U10377 ( .A1(n12592), .A2(n12885), .ZN(n12459) );
  NAND2_X1 U10378 ( .A1(n8001), .A2(n12467), .ZN(n7950) );
  NAND2_X1 U10379 ( .A1(n7949), .A2(n7948), .ZN(n12475) );
  NAND2_X1 U10380 ( .A1(n7950), .A2(n12475), .ZN(n8023) );
  NAND2_X1 U10381 ( .A1(n8023), .A2(n12526), .ZN(n8025) );
  XOR2_X1 U10382 ( .A(n12479), .B(n9444), .Z(n12844) );
  NAND2_X1 U10383 ( .A1(n12543), .A2(n10898), .ZN(n7951) );
  AOI21_X1 U10384 ( .B1(n12334), .B2(n7951), .A(n12337), .ZN(n7954) );
  NAND2_X1 U10385 ( .A1(n12342), .A2(n10898), .ZN(n7952) );
  AND2_X1 U10386 ( .A1(n7960), .A2(n7952), .ZN(n7953) );
  NAND2_X1 U10387 ( .A1(n10038), .A2(n15115), .ZN(n10513) );
  OR2_X1 U10388 ( .A1(n10513), .A2(n12542), .ZN(n7957) );
  AND2_X1 U10389 ( .A1(n12543), .A2(n7959), .ZN(n7956) );
  NAND2_X1 U10390 ( .A1(n12818), .A2(n7956), .ZN(n7958) );
  NAND2_X1 U10391 ( .A1(n12848), .A2(n7398), .ZN(n13072) );
  NAND2_X1 U10392 ( .A1(n12542), .A2(n12496), .ZN(n10043) );
  NAND2_X1 U10393 ( .A1(n7958), .A2(n12488), .ZN(n10660) );
  OAI22_X1 U10394 ( .A1(n12334), .A2(n7960), .B1(n7959), .B2(n15115), .ZN(
        n7961) );
  AOI21_X1 U10395 ( .B1(n7961), .B2(n12542), .A(n12496), .ZN(n7976) );
  NAND2_X1 U10396 ( .A1(n7963), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7962) );
  NAND2_X1 U10397 ( .A1(n7965), .A2(n7966), .ZN(n7977) );
  XNOR2_X1 U10398 ( .A(n7977), .B(P3_B_REG_SCAN_IN), .ZN(n7971) );
  MUX2_X1 U10399 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7967), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n7970) );
  NAND2_X1 U10400 ( .A1(n7968), .A2(n7969), .ZN(n7972) );
  NAND2_X1 U10401 ( .A1(n7971), .A2(n11693), .ZN(n7974) );
  NAND2_X1 U10402 ( .A1(n7972), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7973) );
  INV_X1 U10403 ( .A(n7983), .ZN(n11771) );
  NAND2_X1 U10404 ( .A1(n11771), .A2(n11693), .ZN(n7975) );
  MUX2_X1 U10405 ( .A(n10663), .B(n7976), .S(n10659), .Z(n7996) );
  INV_X1 U10406 ( .A(n7977), .ZN(n7982) );
  OAI22_X2 U10407 ( .A1(n10168), .A2(P3_D_REG_0__SCAN_IN), .B1(n7982), .B2(
        n7983), .ZN(n13124) );
  OR2_X1 U10408 ( .A1(n13124), .A2(n10659), .ZN(n8007) );
  INV_X1 U10409 ( .A(n11693), .ZN(n7981) );
  NAND3_X1 U10410 ( .A1(n7983), .A2(n7982), .A3(n7981), .ZN(n10073) );
  NOR2_X1 U10411 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .ZN(
        n7987) );
  NOR4_X1 U10412 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n7986) );
  NOR4_X1 U10413 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n7985) );
  NOR4_X1 U10414 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n7984) );
  NAND4_X1 U10415 ( .A1(n7987), .A2(n7986), .A3(n7985), .A4(n7984), .ZN(n7993)
         );
  NOR4_X1 U10416 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n7991) );
  NOR4_X1 U10417 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n7990) );
  NOR4_X1 U10418 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n7989) );
  NOR4_X1 U10419 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n7988) );
  NAND4_X1 U10420 ( .A1(n7991), .A2(n7990), .A3(n7989), .A4(n7988), .ZN(n7992)
         );
  NOR2_X1 U10421 ( .A1(n7993), .A2(n7992), .ZN(n7994) );
  NOR2_X1 U10422 ( .A1(n12541), .A2(n8013), .ZN(n7995) );
  NAND2_X1 U10423 ( .A1(n13124), .A2(n10659), .ZN(n8014) );
  INV_X1 U10424 ( .A(n7997), .ZN(n13075) );
  INV_X1 U10425 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n7998) );
  OR2_X1 U10426 ( .A1(n15131), .A2(n7998), .ZN(n7999) );
  XNOR2_X1 U10427 ( .A(n8001), .B(n12525), .ZN(n12864) );
  XOR2_X1 U10428 ( .A(n12525), .B(n8003), .Z(n8006) );
  OAI22_X1 U10429 ( .A1(n12885), .A2(n14341), .B1(n12666), .B2(n14339), .ZN(
        n8004) );
  AOI21_X1 U10430 ( .B1(n12864), .B2(n15070), .A(n8004), .ZN(n8005) );
  AOI21_X1 U10431 ( .B1(n15112), .B2(n12864), .A(n12859), .ZN(n8020) );
  INV_X1 U10432 ( .A(n8007), .ZN(n8009) );
  INV_X1 U10433 ( .A(n8013), .ZN(n8008) );
  NAND2_X1 U10434 ( .A1(n8009), .A2(n8008), .ZN(n10039) );
  INV_X1 U10435 ( .A(n12534), .ZN(n8010) );
  NAND2_X1 U10436 ( .A1(n8010), .A2(n12543), .ZN(n8011) );
  OR2_X1 U10437 ( .A1(n8011), .A2(n12818), .ZN(n10040) );
  OAI21_X1 U10438 ( .B1(n12542), .B2(n12488), .A(n10040), .ZN(n8012) );
  INV_X1 U10439 ( .A(n8012), .ZN(n8016) );
  OR2_X1 U10440 ( .A1(n8014), .A2(n8013), .ZN(n10046) );
  INV_X1 U10441 ( .A(n10038), .ZN(n8015) );
  OAI22_X1 U10442 ( .A1(n10039), .A2(n8016), .B1(n10046), .B2(n8015), .ZN(
        n8017) );
  INV_X1 U10443 ( .A(n12541), .ZN(n10029) );
  NAND2_X1 U10444 ( .A1(n8019), .A2(n7366), .ZN(P3_U3453) );
  INV_X1 U10445 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n8021) );
  NAND2_X1 U10446 ( .A1(n8022), .A2(n7362), .ZN(P3_U3485) );
  NAND2_X1 U10447 ( .A1(n12867), .A2(n8026), .ZN(n8028) );
  NAND2_X1 U10448 ( .A1(n8028), .A2(n8027), .ZN(n8031) );
  OAI21_X1 U10449 ( .B1(n8031), .B2(n8030), .A(n8029), .ZN(n8034) );
  INV_X1 U10450 ( .A(n12560), .ZN(n12682) );
  AOI22_X1 U10451 ( .A1(n15062), .A2(n12870), .B1(n12682), .B2(n15063), .ZN(
        n8032) );
  OAI21_X1 U10452 ( .B1(n12853), .B2(n15116), .A(n12858), .ZN(n13076) );
  INV_X1 U10453 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n8035) );
  AND2_X1 U10454 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n8038) );
  NAND2_X1 U10455 ( .A1(n8726), .A2(n8038), .ZN(n8750) );
  AND2_X1 U10456 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8039) );
  NAND2_X1 U10457 ( .A1(n8043), .A2(n8039), .ZN(n8188) );
  NAND2_X1 U10458 ( .A1(n8750), .A2(n8188), .ZN(n8198) );
  INV_X1 U10459 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10134) );
  NAND2_X1 U10460 ( .A1(n8043), .A2(n10145), .ZN(n8040) );
  NAND2_X1 U10461 ( .A1(n8198), .A2(n8199), .ZN(n8208) );
  INV_X1 U10462 ( .A(n8041), .ZN(n8042) );
  NAND2_X1 U10463 ( .A1(n8042), .A2(SI_1_), .ZN(n8207) );
  MUX2_X1 U10464 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n8043), .Z(n8209) );
  NAND2_X1 U10465 ( .A1(n8209), .A2(SI_2_), .ZN(n8044) );
  AND2_X1 U10466 ( .A1(n8207), .A2(n8044), .ZN(n8045) );
  NAND2_X1 U10467 ( .A1(n8208), .A2(n8045), .ZN(n8049) );
  INV_X1 U10468 ( .A(n8209), .ZN(n8047) );
  INV_X1 U10469 ( .A(SI_2_), .ZN(n8046) );
  NAND2_X1 U10470 ( .A1(n8047), .A2(n8046), .ZN(n8048) );
  NAND2_X1 U10471 ( .A1(n8049), .A2(n8048), .ZN(n8224) );
  INV_X1 U10472 ( .A(n8052), .ZN(n8053) );
  INV_X1 U10473 ( .A(SI_3_), .ZN(n10128) );
  MUX2_X1 U10474 ( .A(n10133), .B(n10139), .S(n6475), .Z(n8054) );
  XNOR2_X1 U10475 ( .A(n8054), .B(SI_4_), .ZN(n8243) );
  INV_X1 U10476 ( .A(n8054), .ZN(n8055) );
  NAND2_X1 U10477 ( .A1(n8055), .A2(SI_4_), .ZN(n8056) );
  MUX2_X1 U10478 ( .A(n10136), .B(n10141), .S(n6475), .Z(n8057) );
  XNOR2_X1 U10479 ( .A(n8057), .B(SI_5_), .ZN(n8258) );
  INV_X1 U10480 ( .A(n8057), .ZN(n8058) );
  NAND2_X1 U10481 ( .A1(n8058), .A2(SI_5_), .ZN(n8059) );
  MUX2_X1 U10482 ( .A(n10152), .B(n10180), .S(n6475), .Z(n8061) );
  XNOR2_X1 U10483 ( .A(n8061), .B(SI_6_), .ZN(n8270) );
  INV_X1 U10484 ( .A(n8061), .ZN(n8062) );
  NAND2_X1 U10485 ( .A1(n8062), .A2(SI_6_), .ZN(n8063) );
  MUX2_X1 U10486 ( .A(n10165), .B(n10176), .S(n6475), .Z(n8064) );
  XNOR2_X1 U10487 ( .A(n8064), .B(SI_7_), .ZN(n8287) );
  INV_X1 U10488 ( .A(n8064), .ZN(n8065) );
  MUX2_X1 U10489 ( .A(n10171), .B(n10174), .S(n6706), .Z(n8066) );
  XNOR2_X1 U10490 ( .A(n8066), .B(SI_8_), .ZN(n8305) );
  INV_X1 U10491 ( .A(n8066), .ZN(n8067) );
  MUX2_X1 U10492 ( .A(n10192), .B(n10191), .S(n6706), .Z(n8068) );
  INV_X1 U10493 ( .A(n8068), .ZN(n8069) );
  NAND2_X1 U10494 ( .A1(n8069), .A2(SI_9_), .ZN(n8070) );
  MUX2_X1 U10495 ( .A(n10221), .B(n10223), .S(n6706), .Z(n8073) );
  NAND2_X1 U10496 ( .A1(n8073), .A2(n10148), .ZN(n8072) );
  INV_X1 U10497 ( .A(n8073), .ZN(n8333) );
  NAND2_X1 U10498 ( .A1(n8333), .A2(SI_10_), .ZN(n8074) );
  MUX2_X1 U10499 ( .A(n10237), .B(n10236), .S(n6706), .Z(n8076) );
  NAND2_X1 U10500 ( .A1(n8076), .A2(n10163), .ZN(n8079) );
  INV_X1 U10501 ( .A(n8076), .ZN(n8077) );
  NAND2_X1 U10502 ( .A1(n8077), .A2(SI_11_), .ZN(n8078) );
  NAND2_X1 U10503 ( .A1(n8079), .A2(n8078), .ZN(n8346) );
  MUX2_X1 U10504 ( .A(n10323), .B(n10322), .S(n6706), .Z(n8080) );
  NAND2_X1 U10505 ( .A1(n8080), .A2(n10167), .ZN(n8083) );
  INV_X1 U10506 ( .A(n8080), .ZN(n8081) );
  NAND2_X1 U10507 ( .A1(n8081), .A2(SI_12_), .ZN(n8082) );
  MUX2_X1 U10508 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n6706), .Z(n8379) );
  INV_X1 U10509 ( .A(n8379), .ZN(n8084) );
  NAND2_X1 U10510 ( .A1(n8084), .A2(n10219), .ZN(n8085) );
  MUX2_X1 U10511 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n6706), .Z(n8394) );
  NAND2_X1 U10512 ( .A1(n8394), .A2(SI_14_), .ZN(n8087) );
  MUX2_X1 U10513 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n6706), .Z(n8411) );
  NAND2_X1 U10514 ( .A1(n8411), .A2(SI_15_), .ZN(n8090) );
  NOR2_X1 U10515 ( .A1(n8394), .A2(SI_14_), .ZN(n8091) );
  INV_X1 U10516 ( .A(n8411), .ZN(n8089) );
  AOI22_X1 U10517 ( .A1(n8091), .A2(n8090), .B1(n10320), .B2(n8089), .ZN(n8092) );
  MUX2_X1 U10518 ( .A(n10571), .B(n10570), .S(n6706), .Z(n8093) );
  XNOR2_X1 U10519 ( .A(n8093), .B(SI_16_), .ZN(n8428) );
  NAND2_X1 U10520 ( .A1(n8093), .A2(n10369), .ZN(n8094) );
  NAND2_X1 U10521 ( .A1(n8095), .A2(n8094), .ZN(n8444) );
  MUX2_X1 U10522 ( .A(n10673), .B(n10672), .S(n6706), .Z(n8096) );
  NAND2_X1 U10523 ( .A1(n8096), .A2(n10440), .ZN(n8097) );
  MUX2_X1 U10524 ( .A(n10876), .B(n10874), .S(n6706), .Z(n8457) );
  MUX2_X1 U10525 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n6706), .Z(n8101) );
  XNOR2_X1 U10526 ( .A(n8101), .B(SI_19_), .ZN(n8473) );
  INV_X1 U10527 ( .A(n8473), .ZN(n8099) );
  NAND2_X1 U10528 ( .A1(n8455), .A2(n8100), .ZN(n8106) );
  INV_X1 U10529 ( .A(n8101), .ZN(n8102) );
  NAND2_X1 U10530 ( .A1(n8102), .A2(n10689), .ZN(n8104) );
  NAND2_X1 U10531 ( .A1(n8106), .A2(n8104), .ZN(n8103) );
  MUX2_X1 U10532 ( .A(n11149), .B(n6950), .S(n6475), .Z(n8500) );
  NAND2_X1 U10533 ( .A1(n8503), .A2(n8108), .ZN(n8171) );
  MUX2_X1 U10534 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n6706), .Z(n8109) );
  OAI21_X1 U10535 ( .B1(SI_21_), .B2(n8109), .A(n8111), .ZN(n8172) );
  INV_X1 U10536 ( .A(n8172), .ZN(n8110) );
  NAND2_X1 U10537 ( .A1(n8171), .A2(n8110), .ZN(n8174) );
  NAND2_X1 U10538 ( .A1(n8174), .A2(n8111), .ZN(n8112) );
  MUX2_X1 U10539 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n6706), .Z(n8507) );
  MUX2_X1 U10540 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n6706), .Z(n8115) );
  INV_X1 U10541 ( .A(n8115), .ZN(n8114) );
  MUX2_X1 U10542 ( .A(n11940), .B(n11943), .S(n6706), .Z(n8533) );
  MUX2_X1 U10543 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n6475), .Z(n8119) );
  XNOR2_X1 U10544 ( .A(n8119), .B(SI_25_), .ZN(n8553) );
  INV_X1 U10545 ( .A(n8558), .ZN(n8122) );
  MUX2_X1 U10546 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n6706), .Z(n8120) );
  NAND2_X1 U10547 ( .A1(n8120), .A2(SI_26_), .ZN(n8123) );
  OAI21_X1 U10548 ( .B1(SI_26_), .B2(n8120), .A(n8123), .ZN(n8557) );
  INV_X1 U10549 ( .A(n8557), .ZN(n8121) );
  NAND2_X1 U10550 ( .A1(n8560), .A2(n8123), .ZN(n8581) );
  MUX2_X1 U10551 ( .A(n14246), .B(n13590), .S(n6706), .Z(n8125) );
  NAND2_X1 U10552 ( .A1(n8125), .A2(n11887), .ZN(n8124) );
  NAND2_X1 U10553 ( .A1(n8581), .A2(n8124), .ZN(n8127) );
  INV_X1 U10554 ( .A(n8125), .ZN(n8582) );
  NAND2_X1 U10555 ( .A1(n8582), .A2(SI_27_), .ZN(n8126) );
  MUX2_X1 U10556 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n6706), .Z(n8586) );
  XNOR2_X1 U10557 ( .A(n8586), .B(SI_28_), .ZN(n8587) );
  NOR2_X1 U10558 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n8131) );
  NAND4_X1 U10559 ( .A1(n8131), .A2(n8130), .A3(n8129), .A4(n8128), .ZN(n8363)
         );
  INV_X1 U10560 ( .A(n8363), .ZN(n8134) );
  NOR2_X1 U10561 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), 
        .ZN(n8137) );
  NOR2_X1 U10562 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), 
        .ZN(n8136) );
  NOR2_X1 U10563 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), 
        .ZN(n8135) );
  NOR2_X1 U10564 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), 
        .ZN(n8141) );
  NAND2_X1 U10565 ( .A1(n8150), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8142) );
  NAND2_X1 U10566 ( .A1(n12296), .A2(n9460), .ZN(n8148) );
  INV_X4 U10567 ( .A(n8225), .ZN(n9459) );
  NAND2_X1 U10568 ( .A1(n9459), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8147) );
  OR2_X1 U10569 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n8149) );
  INV_X1 U10570 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8151) );
  NAND2_X1 U10571 ( .A1(n8154), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n8157) );
  NAND2_X1 U10572 ( .A1(n9453), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8170) );
  NAND2_X2 U10573 ( .A1(n13579), .A2(n8160), .ZN(n9457) );
  NAND2_X1 U10574 ( .A1(n6482), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8169) );
  AND2_X1 U10575 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8236) );
  NAND2_X1 U10576 ( .A1(n8236), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8276) );
  INV_X1 U10577 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8275) );
  NOR2_X1 U10578 ( .A1(n8276), .A2(n8275), .ZN(n8274) );
  NAND2_X1 U10579 ( .A1(n8274), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8324) );
  NAND2_X1 U10580 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG3_REG_8__SCAN_IN), 
        .ZN(n8161) );
  NAND2_X1 U10581 ( .A1(n8352), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8387) );
  INV_X1 U10582 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n11039) );
  INV_X1 U10583 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n13270) );
  NAND2_X1 U10584 ( .A1(n8418), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8450) );
  INV_X1 U10585 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n13314) );
  AND2_X1 U10586 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(P2_REG3_REG_19__SCAN_IN), 
        .ZN(n8162) );
  INV_X1 U10587 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13155) );
  INV_X1 U10588 ( .A(n8688), .ZN(n8166) );
  INV_X1 U10589 ( .A(n8163), .ZN(n8574) );
  INV_X1 U10590 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8164) );
  NAND2_X1 U10591 ( .A1(n8574), .A2(n8164), .ZN(n8165) );
  NAND2_X1 U10592 ( .A1(n8575), .A2(n12212), .ZN(n8168) );
  NAND2_X1 U10593 ( .A1(n8576), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8167) );
  INV_X1 U10594 ( .A(n8171), .ZN(n8173) );
  NAND2_X1 U10595 ( .A1(n8173), .A2(n8172), .ZN(n8175) );
  NAND2_X1 U10596 ( .A1(n8175), .A2(n8174), .ZN(n11266) );
  OR2_X1 U10597 ( .A1(n11266), .A2(n8206), .ZN(n8177) );
  NAND2_X1 U10598 ( .A1(n9459), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8176) );
  INV_X1 U10599 ( .A(n13526), .ZN(n8687) );
  NOR2_X1 U10600 ( .A1(n8491), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n8178) );
  OR2_X1 U10601 ( .A1(n8514), .A2(n8178), .ZN(n13434) );
  INV_X2 U10602 ( .A(n8465), .ZN(n8591) );
  INV_X1 U10603 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8181) );
  NAND2_X1 U10604 ( .A1(n8576), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8180) );
  NAND2_X1 U10605 ( .A1(n9453), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8179) );
  OAI211_X1 U10606 ( .C1(n9457), .C2(n8181), .A(n8180), .B(n8179), .ZN(n8182)
         );
  INV_X1 U10607 ( .A(n8182), .ZN(n8183) );
  OAI21_X1 U10608 ( .B1(n13434), .B2(n8465), .A(n8183), .ZN(n13289) );
  INV_X1 U10609 ( .A(n13289), .ZN(n13235) );
  NAND2_X1 U10610 ( .A1(n8591), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8185) );
  NAND2_X1 U10611 ( .A1(n8278), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n8184) );
  INV_X1 U10612 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10226) );
  NAND2_X1 U10613 ( .A1(n6706), .A2(SI_0_), .ZN(n8187) );
  NAND2_X1 U10614 ( .A1(n8187), .A2(n8186), .ZN(n8189) );
  NAND2_X1 U10615 ( .A1(n8189), .A2(n8188), .ZN(n13597) );
  MUX2_X1 U10616 ( .A(n10226), .B(n13597), .S(n10196), .Z(n14721) );
  OR2_X1 U10617 ( .A1(n9457), .A2(n14834), .ZN(n8194) );
  NAND2_X1 U10618 ( .A1(n8575), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n8193) );
  NAND2_X1 U10619 ( .A1(n8278), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8192) );
  INV_X1 U10620 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n8190) );
  NAND2_X1 U10621 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8195) );
  MUX2_X1 U10622 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8195), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n8197) );
  INV_X1 U10623 ( .A(n8196), .ZN(n8212) );
  XNOR2_X1 U10624 ( .A(n8198), .B(n8199), .ZN(n10144) );
  XNOR2_X2 U10625 ( .A(n13308), .B(n11180), .ZN(n9474) );
  NAND2_X1 U10626 ( .A1(n11173), .A2(n9474), .ZN(n8201) );
  INV_X1 U10627 ( .A(n13308), .ZN(n8200) );
  NAND2_X1 U10628 ( .A1(n8200), .A2(n11180), .ZN(n9477) );
  NAND2_X1 U10629 ( .A1(n8278), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8205) );
  NAND2_X1 U10630 ( .A1(n6482), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8204) );
  NAND2_X1 U10631 ( .A1(n8576), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8203) );
  NAND2_X1 U10632 ( .A1(n8591), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n8202) );
  NAND2_X1 U10633 ( .A1(n8208), .A2(n8207), .ZN(n8211) );
  XNOR2_X1 U10634 ( .A(n8209), .B(SI_2_), .ZN(n8210) );
  XNOR2_X1 U10635 ( .A(n8211), .B(n8210), .ZN(n10130) );
  NAND2_X1 U10636 ( .A1(n9460), .A2(n10130), .ZN(n8218) );
  OR2_X1 U10637 ( .A1(n8225), .A2(n10178), .ZN(n8217) );
  NAND2_X1 U10638 ( .A1(n8212), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8213) );
  MUX2_X1 U10639 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8213), .S(
        P2_IR_REG_2__SCAN_IN), .Z(n8215) );
  INV_X1 U10640 ( .A(n8214), .ZN(n8227) );
  NAND2_X1 U10641 ( .A1(n8215), .A2(n8227), .ZN(n14562) );
  INV_X1 U10642 ( .A(n14562), .ZN(n10252) );
  NAND2_X1 U10643 ( .A1(n8477), .A2(n10252), .ZN(n8216) );
  NAND2_X1 U10644 ( .A1(n10863), .A2(n10864), .ZN(n8232) );
  NAND2_X1 U10645 ( .A1(n6482), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8222) );
  INV_X1 U10646 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8234) );
  NAND2_X1 U10647 ( .A1(n8575), .A2(n8234), .ZN(n8221) );
  NAND2_X1 U10648 ( .A1(n8278), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n8220) );
  NAND2_X1 U10649 ( .A1(n8576), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8219) );
  INV_X1 U10650 ( .A(n13307), .ZN(n8648) );
  XNOR2_X1 U10651 ( .A(n8224), .B(n8223), .ZN(n10143) );
  OR2_X1 U10652 ( .A1(n8225), .A2(n10142), .ZN(n8230) );
  NAND2_X1 U10653 ( .A1(n8227), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8226) );
  MUX2_X1 U10654 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8226), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n8228) );
  AND2_X1 U10655 ( .A1(n8228), .A2(n8260), .ZN(n10253) );
  NAND2_X1 U10656 ( .A1(n8477), .A2(n10253), .ZN(n8229) );
  OAI211_X2 U10657 ( .C1(n8206), .C2(n10143), .A(n8230), .B(n8229), .ZN(n14766) );
  NAND2_X1 U10658 ( .A1(n8648), .A2(n14766), .ZN(n10997) );
  NAND2_X1 U10659 ( .A1(n13307), .A2(n10869), .ZN(n8231) );
  INV_X1 U10660 ( .A(n8647), .ZN(n10861) );
  NAND2_X1 U10661 ( .A1(n10999), .A2(n10997), .ZN(n8249) );
  NAND2_X1 U10662 ( .A1(n6482), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8241) );
  INV_X1 U10663 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n8235) );
  NAND2_X1 U10664 ( .A1(n8235), .A2(n8234), .ZN(n8237) );
  INV_X1 U10665 ( .A(n8236), .ZN(n8251) );
  AND2_X1 U10666 ( .A1(n8237), .A2(n8251), .ZN(n10446) );
  NAND2_X1 U10667 ( .A1(n8591), .A2(n10446), .ZN(n8240) );
  NAND2_X1 U10668 ( .A1(n9453), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n8239) );
  NAND2_X1 U10669 ( .A1(n8576), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8238) );
  INV_X1 U10670 ( .A(n13306), .ZN(n10867) );
  XNOR2_X1 U10671 ( .A(n8242), .B(n7273), .ZN(n10132) );
  NAND2_X1 U10672 ( .A1(n10132), .A2(n9460), .ZN(n8246) );
  NAND2_X1 U10673 ( .A1(n8260), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8244) );
  XNOR2_X1 U10674 ( .A(n8244), .B(P2_IR_REG_4__SCAN_IN), .ZN(n14583) );
  AOI22_X1 U10675 ( .A1(n9459), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n8477), .B2(
        n14583), .ZN(n8245) );
  NAND2_X1 U10676 ( .A1(n8246), .A2(n8245), .ZN(n11008) );
  NAND2_X1 U10677 ( .A1(n10867), .A2(n11008), .ZN(n11131) );
  INV_X1 U10678 ( .A(n11008), .ZN(n14776) );
  NAND2_X1 U10679 ( .A1(n13306), .A2(n14776), .ZN(n8247) );
  NAND2_X1 U10680 ( .A1(n11131), .A2(n8247), .ZN(n10998) );
  INV_X1 U10681 ( .A(n10998), .ZN(n8248) );
  NAND2_X1 U10682 ( .A1(n8249), .A2(n8248), .ZN(n10996) );
  NAND2_X1 U10683 ( .A1(n10996), .A2(n11131), .ZN(n8269) );
  NAND2_X1 U10684 ( .A1(n6482), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8256) );
  INV_X1 U10685 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8250) );
  NAND2_X1 U10686 ( .A1(n8251), .A2(n8250), .ZN(n8252) );
  AND2_X1 U10687 ( .A1(n8276), .A2(n8252), .ZN(n11128) );
  NAND2_X1 U10688 ( .A1(n8575), .A2(n11128), .ZN(n8255) );
  NAND2_X1 U10689 ( .A1(n9453), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8254) );
  NAND2_X1 U10690 ( .A1(n8576), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8253) );
  NAND4_X1 U10691 ( .A1(n8256), .A2(n8255), .A3(n8254), .A4(n8253), .ZN(n13305) );
  INV_X1 U10692 ( .A(n13305), .ZN(n8266) );
  INV_X1 U10693 ( .A(n8258), .ZN(n8259) );
  XNOR2_X1 U10694 ( .A(n8257), .B(n8259), .ZN(n10135) );
  NAND2_X1 U10695 ( .A1(n10135), .A2(n9460), .ZN(n8265) );
  INV_X1 U10696 ( .A(n8260), .ZN(n8262) );
  INV_X1 U10697 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8261) );
  NAND2_X1 U10698 ( .A1(n8262), .A2(n8261), .ZN(n8364) );
  NAND2_X1 U10699 ( .A1(n8364), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8263) );
  XNOR2_X1 U10700 ( .A(n8263), .B(P2_IR_REG_5__SCAN_IN), .ZN(n14599) );
  AOI22_X1 U10701 ( .A1(n9459), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8477), .B2(
        n14599), .ZN(n8264) );
  NAND2_X1 U10702 ( .A1(n8265), .A2(n8264), .ZN(n11129) );
  NAND2_X1 U10703 ( .A1(n8266), .A2(n11129), .ZN(n10832) );
  INV_X1 U10704 ( .A(n11129), .ZN(n14783) );
  NAND2_X1 U10705 ( .A1(n14783), .A2(n13305), .ZN(n8267) );
  NAND2_X1 U10706 ( .A1(n10832), .A2(n8267), .ZN(n11132) );
  INV_X1 U10707 ( .A(n11132), .ZN(n8268) );
  NAND2_X1 U10708 ( .A1(n8269), .A2(n8268), .ZN(n10831) );
  NAND2_X1 U10709 ( .A1(n10831), .A2(n10832), .ZN(n8283) );
  XNOR2_X1 U10710 ( .A(n8271), .B(n7284), .ZN(n10151) );
  NAND2_X1 U10711 ( .A1(n10151), .A2(n9460), .ZN(n8273) );
  NAND2_X1 U10712 ( .A1(n8307), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8289) );
  XNOR2_X1 U10713 ( .A(n8289), .B(P2_IR_REG_6__SCAN_IN), .ZN(n10290) );
  AOI22_X1 U10714 ( .A1(n9459), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8477), .B2(
        n10290), .ZN(n8272) );
  NAND2_X1 U10715 ( .A1(n6482), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8282) );
  INV_X1 U10716 ( .A(n8274), .ZN(n8295) );
  NAND2_X1 U10717 ( .A1(n8276), .A2(n8275), .ZN(n8277) );
  AND2_X1 U10718 ( .A1(n8295), .A2(n8277), .ZN(n10839) );
  NAND2_X1 U10719 ( .A1(n8575), .A2(n10839), .ZN(n8281) );
  NAND2_X1 U10720 ( .A1(n9453), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n8280) );
  NAND2_X1 U10721 ( .A1(n8576), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8279) );
  NAND4_X1 U10722 ( .A1(n8282), .A2(n8281), .A3(n8280), .A4(n8279), .ZN(n13304) );
  XNOR2_X1 U10723 ( .A(n10911), .B(n13304), .ZN(n10826) );
  INV_X1 U10724 ( .A(n13304), .ZN(n8284) );
  NAND2_X1 U10725 ( .A1(n10911), .A2(n8284), .ZN(n8285) );
  XNOR2_X1 U10726 ( .A(n8286), .B(n7287), .ZN(n10164) );
  NAND2_X1 U10727 ( .A1(n10164), .A2(n9460), .ZN(n8293) );
  INV_X1 U10728 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8288) );
  NAND2_X1 U10729 ( .A1(n8289), .A2(n8288), .ZN(n8290) );
  NAND2_X1 U10730 ( .A1(n8290), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8291) );
  XNOR2_X1 U10731 ( .A(n8291), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10268) );
  AOI22_X1 U10732 ( .A1(n9459), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8477), .B2(
        n10268), .ZN(n8292) );
  NAND2_X1 U10733 ( .A1(n6482), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8300) );
  INV_X1 U10734 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8294) );
  NAND2_X1 U10735 ( .A1(n8295), .A2(n8294), .ZN(n8296) );
  AND2_X1 U10736 ( .A1(n8324), .A2(n8296), .ZN(n10782) );
  NAND2_X1 U10737 ( .A1(n8575), .A2(n10782), .ZN(n8299) );
  NAND2_X1 U10738 ( .A1(n9453), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8298) );
  NAND2_X1 U10739 ( .A1(n8576), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8297) );
  NAND4_X1 U10740 ( .A1(n8300), .A2(n8299), .A3(n8298), .A4(n8297), .ZN(n13303) );
  INV_X1 U10741 ( .A(n13303), .ZN(n8302) );
  OR2_X1 U10742 ( .A1(n14789), .A2(n8302), .ZN(n8301) );
  NAND2_X1 U10743 ( .A1(n14789), .A2(n8302), .ZN(n8303) );
  INV_X1 U10744 ( .A(n8305), .ZN(n8306) );
  XNOR2_X1 U10745 ( .A(n8304), .B(n8306), .ZN(n10170) );
  NAND2_X1 U10746 ( .A1(n10170), .A2(n9460), .ZN(n8312) );
  INV_X1 U10747 ( .A(n8307), .ZN(n8309) );
  NOR2_X1 U10748 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n8308) );
  NAND2_X1 U10749 ( .A1(n8309), .A2(n8308), .ZN(n8318) );
  NAND2_X1 U10750 ( .A1(n8318), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8310) );
  XNOR2_X1 U10751 ( .A(n8310), .B(P2_IR_REG_8__SCAN_IN), .ZN(n10585) );
  AOI22_X1 U10752 ( .A1(n9459), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8477), .B2(
        n10585), .ZN(n8311) );
  NAND2_X1 U10753 ( .A1(n6482), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8316) );
  XNOR2_X1 U10754 ( .A(n8324), .B(P2_REG3_REG_8__SCAN_IN), .ZN(n11153) );
  NAND2_X1 U10755 ( .A1(n8575), .A2(n11153), .ZN(n8315) );
  NAND2_X1 U10756 ( .A1(n9453), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8314) );
  NAND2_X1 U10757 ( .A1(n8576), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8313) );
  NAND4_X1 U10758 ( .A1(n8316), .A2(n8315), .A3(n8314), .A4(n8313), .ZN(n13302) );
  XNOR2_X1 U10759 ( .A(n11154), .B(n13302), .ZN(n11157) );
  NAND2_X1 U10760 ( .A1(n11156), .A2(n11157), .ZN(n14700) );
  XNOR2_X1 U10761 ( .A(n8317), .B(n6558), .ZN(n10190) );
  NAND2_X1 U10762 ( .A1(n10190), .A2(n9460), .ZN(n8321) );
  NAND2_X1 U10763 ( .A1(n8335), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8319) );
  XNOR2_X1 U10764 ( .A(n8319), .B(P2_IR_REG_9__SCAN_IN), .ZN(n14614) );
  AOI22_X1 U10765 ( .A1(n9459), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8477), .B2(
        n14614), .ZN(n8320) );
  NAND2_X1 U10766 ( .A1(n6482), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n8329) );
  INV_X1 U10767 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8323) );
  INV_X1 U10768 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8322) );
  OAI21_X1 U10769 ( .B1(n8324), .B2(n8323), .A(n8322), .ZN(n8325) );
  AND2_X1 U10770 ( .A1(n8325), .A2(n8340), .ZN(n14704) );
  NAND2_X1 U10771 ( .A1(n8591), .A2(n14704), .ZN(n8328) );
  NAND2_X1 U10772 ( .A1(n9453), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8327) );
  NAND2_X1 U10773 ( .A1(n8576), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8326) );
  NAND4_X1 U10774 ( .A1(n8329), .A2(n8328), .A3(n8327), .A4(n8326), .ZN(n13301) );
  INV_X1 U10775 ( .A(n13301), .ZN(n9523) );
  NAND2_X1 U10776 ( .A1(n14710), .A2(n9523), .ZN(n8330) );
  INV_X1 U10777 ( .A(n13302), .ZN(n11108) );
  NAND2_X1 U10778 ( .A1(n11154), .A2(n11108), .ZN(n14699) );
  AND2_X1 U10779 ( .A1(n8330), .A2(n14699), .ZN(n8331) );
  OR2_X1 U10780 ( .A1(n14710), .A2(n9523), .ZN(n8332) );
  XNOR2_X1 U10781 ( .A(n8333), .B(SI_10_), .ZN(n8334) );
  NAND2_X1 U10782 ( .A1(n10220), .A2(n9460), .ZN(n8338) );
  NAND2_X1 U10783 ( .A1(n8348), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8336) );
  XNOR2_X1 U10784 ( .A(n8336), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10588) );
  AOI22_X1 U10785 ( .A1(n9459), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n8477), 
        .B2(n10588), .ZN(n8337) );
  NAND2_X1 U10786 ( .A1(n6482), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8345) );
  INV_X1 U10787 ( .A(n8339), .ZN(n8354) );
  NAND2_X1 U10788 ( .A1(n8340), .A2(n11167), .ZN(n8341) );
  AND2_X1 U10789 ( .A1(n8354), .A2(n8341), .ZN(n11328) );
  NAND2_X1 U10790 ( .A1(n8591), .A2(n11328), .ZN(n8344) );
  NAND2_X1 U10791 ( .A1(n9453), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n8343) );
  NAND2_X1 U10792 ( .A1(n8576), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8342) );
  NAND4_X1 U10793 ( .A1(n8345), .A2(n8344), .A3(n8343), .A4(n8342), .ZN(n13300) );
  XNOR2_X1 U10794 ( .A(n14813), .B(n13300), .ZN(n9522) );
  INV_X1 U10795 ( .A(n13300), .ZN(n11107) );
  NAND2_X1 U10796 ( .A1(n14813), .A2(n11107), .ZN(n11307) );
  NAND2_X1 U10797 ( .A1(n11324), .A2(n11307), .ZN(n8360) );
  XNOR2_X1 U10798 ( .A(n8346), .B(n8347), .ZN(n10235) );
  NAND2_X1 U10799 ( .A1(n10235), .A2(n9460), .ZN(n8351) );
  OAI21_X1 U10800 ( .B1(n8348), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8349) );
  XNOR2_X1 U10801 ( .A(n8349), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11034) );
  AOI22_X1 U10802 ( .A1(n9459), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n11034), 
        .B2(n8477), .ZN(n8350) );
  INV_X1 U10803 ( .A(n8352), .ZN(n8369) );
  INV_X1 U10804 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8353) );
  NAND2_X1 U10805 ( .A1(n8354), .A2(n8353), .ZN(n8355) );
  AND2_X1 U10806 ( .A1(n8369), .A2(n8355), .ZN(n11376) );
  NAND2_X1 U10807 ( .A1(n8591), .A2(n11376), .ZN(n8359) );
  NAND2_X1 U10808 ( .A1(n6482), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8358) );
  NAND2_X1 U10809 ( .A1(n9453), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8357) );
  NAND2_X1 U10810 ( .A1(n8576), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n8356) );
  NAND4_X1 U10811 ( .A1(n8359), .A2(n8358), .A3(n8357), .A4(n8356), .ZN(n13299) );
  INV_X1 U10812 ( .A(n13299), .ZN(n11402) );
  XNOR2_X1 U10813 ( .A(n11382), .B(n11402), .ZN(n11308) );
  INV_X1 U10814 ( .A(n11308), .ZN(n11305) );
  NAND2_X1 U10815 ( .A1(n11382), .A2(n11402), .ZN(n8361) );
  NAND2_X1 U10816 ( .A1(n11310), .A2(n8361), .ZN(n11435) );
  XNOR2_X1 U10817 ( .A(n8362), .B(n7376), .ZN(n10321) );
  NAND2_X1 U10818 ( .A1(n10321), .A2(n9460), .ZN(n8367) );
  OAI21_X1 U10819 ( .B1(n8364), .B2(n8363), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8365) );
  XNOR2_X1 U10820 ( .A(n8365), .B(P2_IR_REG_12__SCAN_IN), .ZN(n14643) );
  AOI22_X1 U10821 ( .A1(n9459), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8477), 
        .B2(n14643), .ZN(n8366) );
  NAND2_X1 U10822 ( .A1(n6482), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8374) );
  INV_X1 U10823 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8368) );
  NAND2_X1 U10824 ( .A1(n8369), .A2(n8368), .ZN(n8370) );
  AND2_X1 U10825 ( .A1(n8387), .A2(n8370), .ZN(n11442) );
  NAND2_X1 U10826 ( .A1(n8591), .A2(n11442), .ZN(n8373) );
  NAND2_X1 U10827 ( .A1(n9453), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n8372) );
  NAND2_X1 U10828 ( .A1(n8576), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8371) );
  NAND4_X1 U10829 ( .A1(n8374), .A2(n8373), .A3(n8372), .A4(n8371), .ZN(n13298) );
  INV_X1 U10830 ( .A(n13298), .ZN(n8375) );
  NAND2_X1 U10831 ( .A1(n11435), .A2(n11443), .ZN(n8376) );
  XNOR2_X1 U10832 ( .A(n8379), .B(n10219), .ZN(n8380) );
  XNOR2_X1 U10833 ( .A(n8378), .B(n8380), .ZN(n10400) );
  NAND2_X1 U10834 ( .A1(n10400), .A2(n9460), .ZN(n8385) );
  NAND2_X1 U10835 ( .A1(n8381), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8382) );
  MUX2_X1 U10836 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8382), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n8383) );
  INV_X1 U10837 ( .A(n8601), .ZN(n8395) );
  AND2_X1 U10838 ( .A1(n8383), .A2(n8395), .ZN(n14657) );
  AOI22_X1 U10839 ( .A1(n9459), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8477), 
        .B2(n14657), .ZN(n8384) );
  NAND2_X1 U10840 ( .A1(n6482), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8392) );
  NAND2_X1 U10841 ( .A1(n8387), .A2(n8386), .ZN(n8388) );
  AND2_X1 U10842 ( .A1(n8399), .A2(n8388), .ZN(n11515) );
  NAND2_X1 U10843 ( .A1(n8575), .A2(n11515), .ZN(n8391) );
  NAND2_X1 U10844 ( .A1(n9453), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8390) );
  NAND2_X1 U10845 ( .A1(n8576), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n8389) );
  NAND4_X1 U10846 ( .A1(n8392), .A2(n8391), .A3(n8390), .A4(n8389), .ZN(n13297) );
  INV_X1 U10847 ( .A(n8394), .ZN(n8409) );
  XNOR2_X1 U10848 ( .A(n8410), .B(n8409), .ZN(n10596) );
  NAND2_X1 U10849 ( .A1(n10596), .A2(n9460), .ZN(n8398) );
  NAND2_X1 U10850 ( .A1(n8395), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8396) );
  XNOR2_X1 U10851 ( .A(n8396), .B(P2_IR_REG_14__SCAN_IN), .ZN(n12226) );
  AOI22_X1 U10852 ( .A1(n9459), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8477), 
        .B2(n12226), .ZN(n8397) );
  NAND2_X1 U10853 ( .A1(n6482), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8404) );
  NAND2_X1 U10854 ( .A1(n8399), .A2(n11039), .ZN(n8400) );
  AND2_X1 U10855 ( .A1(n8419), .A2(n8400), .ZN(n11761) );
  NAND2_X1 U10856 ( .A1(n8591), .A2(n11761), .ZN(n8403) );
  NAND2_X1 U10857 ( .A1(n9453), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8402) );
  NAND2_X1 U10858 ( .A1(n8576), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n8401) );
  NAND4_X1 U10859 ( .A1(n8404), .A2(n8403), .A3(n8402), .A4(n8401), .ZN(n13296) );
  INV_X1 U10860 ( .A(n13296), .ZN(n9648) );
  NAND2_X1 U10861 ( .A1(n8405), .A2(n7394), .ZN(n8407) );
  NAND2_X1 U10862 ( .A1(n13557), .A2(n9648), .ZN(n8406) );
  NAND2_X1 U10863 ( .A1(n8407), .A2(n8406), .ZN(n11711) );
  AND2_X1 U10864 ( .A1(n8393), .A2(n10279), .ZN(n8408) );
  AOI21_X1 U10865 ( .B1(n8410), .B2(n8409), .A(n8408), .ZN(n8413) );
  XNOR2_X1 U10866 ( .A(n8411), .B(SI_15_), .ZN(n8412) );
  XNOR2_X1 U10867 ( .A(n8413), .B(n8412), .ZN(n10655) );
  NAND2_X1 U10868 ( .A1(n10655), .A2(n9460), .ZN(n8417) );
  INV_X1 U10869 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n8414) );
  NAND2_X1 U10870 ( .A1(n8601), .A2(n8414), .ZN(n8429) );
  NAND2_X1 U10871 ( .A1(n8429), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8415) );
  XNOR2_X1 U10872 ( .A(n8415), .B(P2_IR_REG_15__SCAN_IN), .ZN(n14662) );
  AOI22_X1 U10873 ( .A1(n9459), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n8477), 
        .B2(n14662), .ZN(n8416) );
  NAND2_X1 U10874 ( .A1(n6482), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8424) );
  INV_X1 U10875 ( .A(n8418), .ZN(n8435) );
  NAND2_X1 U10876 ( .A1(n8419), .A2(n13270), .ZN(n8420) );
  AND2_X1 U10877 ( .A1(n8435), .A2(n8420), .ZN(n13275) );
  NAND2_X1 U10878 ( .A1(n8591), .A2(n13275), .ZN(n8423) );
  NAND2_X1 U10879 ( .A1(n9453), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8422) );
  NAND2_X1 U10880 ( .A1(n8576), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n8421) );
  NAND4_X1 U10881 ( .A1(n8424), .A2(n8423), .A3(n8422), .A4(n8421), .ZN(n13295) );
  INV_X1 U10882 ( .A(n13295), .ZN(n8425) );
  OR2_X1 U10883 ( .A1(n12161), .A2(n8425), .ZN(n8426) );
  XNOR2_X1 U10884 ( .A(n8427), .B(n8428), .ZN(n10569) );
  NAND2_X1 U10885 ( .A1(n10569), .A2(n9460), .ZN(n8434) );
  INV_X1 U10886 ( .A(n8429), .ZN(n8431) );
  INV_X1 U10887 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8430) );
  NAND2_X1 U10888 ( .A1(n8446), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8432) );
  XNOR2_X1 U10889 ( .A(n8432), .B(P2_IR_REG_16__SCAN_IN), .ZN(n12236) );
  AOI22_X1 U10890 ( .A1(n9459), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8477), 
        .B2(n12236), .ZN(n8433) );
  INV_X1 U10891 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n13197) );
  NAND2_X1 U10892 ( .A1(n8435), .A2(n13197), .ZN(n8436) );
  NAND2_X1 U10893 ( .A1(n8450), .A2(n8436), .ZN(n11889) );
  NAND2_X1 U10894 ( .A1(n6482), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8438) );
  NAND2_X1 U10895 ( .A1(n9453), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8437) );
  AND2_X1 U10896 ( .A1(n8438), .A2(n8437), .ZN(n8440) );
  NAND2_X1 U10897 ( .A1(n8576), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n8439) );
  OAI211_X1 U10898 ( .C1(n11889), .C2(n8465), .A(n8440), .B(n8439), .ZN(n13294) );
  INV_X1 U10899 ( .A(n13294), .ZN(n8441) );
  NAND2_X1 U10900 ( .A1(n13553), .A2(n8441), .ZN(n8442) );
  NAND2_X1 U10901 ( .A1(n8443), .A2(n8442), .ZN(n11959) );
  XNOR2_X1 U10902 ( .A(n8444), .B(n8445), .ZN(n10671) );
  NAND2_X1 U10903 ( .A1(n10671), .A2(n9460), .ZN(n8449) );
  NAND2_X1 U10904 ( .A1(n6591), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8447) );
  XNOR2_X1 U10905 ( .A(n8447), .B(P2_IR_REG_17__SCAN_IN), .ZN(n14686) );
  AOI22_X1 U10906 ( .A1(n9459), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8477), 
        .B2(n14686), .ZN(n8448) );
  NAND2_X1 U10907 ( .A1(n8450), .A2(n13210), .ZN(n8451) );
  NAND2_X1 U10908 ( .A1(n8463), .A2(n8451), .ZN(n11966) );
  AOI22_X1 U10909 ( .A1(n6482), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n9453), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n8453) );
  NAND2_X1 U10910 ( .A1(n8576), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8452) );
  OAI211_X1 U10911 ( .C1(n11966), .C2(n8465), .A(n8453), .B(n8452), .ZN(n13293) );
  INV_X1 U10912 ( .A(n13293), .ZN(n8454) );
  XNOR2_X1 U10913 ( .A(n13547), .B(n8454), .ZN(n11968) );
  NAND2_X1 U10914 ( .A1(n8456), .A2(n8457), .ZN(n8458) );
  NAND2_X1 U10915 ( .A1(n8455), .A2(n8458), .ZN(n10875) );
  OR2_X1 U10916 ( .A1(n10875), .A2(n8206), .ZN(n8461) );
  NAND2_X1 U10917 ( .A1(n8475), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8459) );
  XNOR2_X1 U10918 ( .A(n8459), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13318) );
  AOI22_X1 U10919 ( .A1(n13318), .A2(n8477), .B1(n9459), .B2(
        P1_DATAO_REG_18__SCAN_IN), .ZN(n8460) );
  INV_X1 U10920 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8468) );
  INV_X1 U10921 ( .A(n8462), .ZN(n8490) );
  NAND2_X1 U10922 ( .A1(n8463), .A2(n13314), .ZN(n8464) );
  NAND2_X1 U10923 ( .A1(n8490), .A2(n8464), .ZN(n11946) );
  OR2_X1 U10924 ( .A1(n11946), .A2(n8465), .ZN(n8467) );
  AOI22_X1 U10925 ( .A1(n6482), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n9453), .B2(
        P2_REG2_REG_18__SCAN_IN), .ZN(n8466) );
  OAI211_X1 U10926 ( .C1(n8469), .C2(n8468), .A(n8467), .B(n8466), .ZN(n13292)
         );
  NAND2_X1 U10927 ( .A1(n8455), .A2(n8472), .ZN(n8474) );
  XNOR2_X1 U10928 ( .A(n8474), .B(n8473), .ZN(n10949) );
  NAND2_X1 U10929 ( .A1(n10949), .A2(n9460), .ZN(n8479) );
  XNOR2_X1 U10930 ( .A(n8476), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8683) );
  AOI22_X1 U10931 ( .A1(n8683), .A2(n8477), .B1(n9459), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n8478) );
  XNOR2_X1 U10932 ( .A(n8490), .B(P2_REG3_REG_19__SCAN_IN), .ZN(n13468) );
  NAND2_X1 U10933 ( .A1(n13468), .A2(n8591), .ZN(n8485) );
  INV_X1 U10934 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8482) );
  NAND2_X1 U10935 ( .A1(n8576), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8481) );
  NAND2_X1 U10936 ( .A1(n9453), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8480) );
  OAI211_X1 U10937 ( .C1(n9457), .C2(n8482), .A(n8481), .B(n8480), .ZN(n8483)
         );
  INV_X1 U10938 ( .A(n8483), .ZN(n8484) );
  NAND2_X1 U10939 ( .A1(n8485), .A2(n8484), .ZN(n13291) );
  NAND2_X1 U10940 ( .A1(n13537), .A2(n8486), .ZN(n8487) );
  INV_X1 U10941 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8489) );
  INV_X1 U10942 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8488) );
  OAI21_X1 U10943 ( .B1(n8490), .B2(n8489), .A(n8488), .ZN(n8493) );
  INV_X1 U10944 ( .A(n8491), .ZN(n8492) );
  AND2_X1 U10945 ( .A1(n8493), .A2(n8492), .ZN(n13450) );
  NAND2_X1 U10946 ( .A1(n13450), .A2(n8591), .ZN(n8499) );
  INV_X1 U10947 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8496) );
  NAND2_X1 U10948 ( .A1(n9453), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8495) );
  NAND2_X1 U10949 ( .A1(n8576), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8494) );
  OAI211_X1 U10950 ( .C1(n8496), .C2(n9457), .A(n8495), .B(n8494), .ZN(n8497)
         );
  INV_X1 U10951 ( .A(n8497), .ZN(n8498) );
  NAND2_X1 U10952 ( .A1(n8499), .A2(n8498), .ZN(n13290) );
  NAND2_X1 U10953 ( .A1(n8501), .A2(n8500), .ZN(n8502) );
  NAND2_X1 U10954 ( .A1(n11148), .A2(n9460), .ZN(n8505) );
  NAND2_X1 U10955 ( .A1(n9459), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8504) );
  XOR2_X1 U10956 ( .A(n13290), .B(n13531), .Z(n13443) );
  INV_X1 U10957 ( .A(n13531), .ZN(n13454) );
  INV_X1 U10958 ( .A(n8506), .ZN(n8509) );
  INV_X1 U10959 ( .A(n8507), .ZN(n8508) );
  NAND2_X1 U10960 ( .A1(n8509), .A2(n8508), .ZN(n8510) );
  AND2_X1 U10961 ( .A1(n8511), .A2(n8510), .ZN(n11534) );
  NAND2_X1 U10962 ( .A1(n11534), .A2(n9460), .ZN(n8513) );
  NAND2_X1 U10963 ( .A1(n9459), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8512) );
  OR2_X1 U10964 ( .A1(n8514), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8515) );
  AND2_X1 U10965 ( .A1(n8515), .A2(n8527), .ZN(n13420) );
  NAND2_X1 U10966 ( .A1(n13420), .A2(n8591), .ZN(n8521) );
  INV_X1 U10967 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8518) );
  NAND2_X1 U10968 ( .A1(n8576), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8517) );
  NAND2_X1 U10969 ( .A1(n9453), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8516) );
  OAI211_X1 U10970 ( .C1(n9457), .C2(n8518), .A(n8517), .B(n8516), .ZN(n8519)
         );
  INV_X1 U10971 ( .A(n8519), .ZN(n8520) );
  NAND2_X1 U10972 ( .A1(n8521), .A2(n8520), .ZN(n13288) );
  XNOR2_X1 U10973 ( .A(n13518), .B(n13180), .ZN(n9653) );
  NAND2_X1 U10974 ( .A1(n8522), .A2(n11288), .ZN(n8523) );
  NAND2_X1 U10975 ( .A1(n11752), .A2(n9460), .ZN(n8526) );
  NAND2_X1 U10976 ( .A1(n9459), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8525) );
  NAND2_X1 U10977 ( .A1(n6482), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8531) );
  AOI21_X1 U10978 ( .B1(n13155), .B2(n8527), .A(n8536), .ZN(n13403) );
  NAND2_X1 U10979 ( .A1(n8591), .A2(n13403), .ZN(n8530) );
  NAND2_X1 U10980 ( .A1(n9453), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8529) );
  NAND2_X1 U10981 ( .A1(n8576), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8528) );
  NAND4_X1 U10982 ( .A1(n8531), .A2(n8530), .A3(n8529), .A4(n8528), .ZN(n13287) );
  NOR2_X1 U10983 ( .A1(n13514), .A2(n13234), .ZN(n8532) );
  INV_X1 U10984 ( .A(n13514), .ZN(n13411) );
  NAND2_X1 U10985 ( .A1(n9459), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8535) );
  NAND2_X1 U10986 ( .A1(n6482), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8544) );
  NAND2_X1 U10987 ( .A1(n9453), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8543) );
  INV_X1 U10988 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8538) );
  INV_X1 U10989 ( .A(n8536), .ZN(n8537) );
  NAND2_X1 U10990 ( .A1(n8538), .A2(n8537), .ZN(n8540) );
  INV_X1 U10991 ( .A(n8539), .ZN(n8547) );
  NAND2_X1 U10992 ( .A1(n8575), .A2(n13394), .ZN(n8542) );
  NAND2_X1 U10993 ( .A1(n8576), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8541) );
  INV_X1 U10994 ( .A(n13187), .ZN(n13286) );
  XNOR2_X1 U10995 ( .A(n13507), .B(n13286), .ZN(n13398) );
  NAND2_X1 U10996 ( .A1(n6482), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8552) );
  NAND2_X1 U10997 ( .A1(n9453), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8551) );
  INV_X1 U10998 ( .A(n8545), .ZN(n8565) );
  INV_X1 U10999 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8546) );
  NAND2_X1 U11000 ( .A1(n8547), .A2(n8546), .ZN(n8548) );
  NAND2_X1 U11001 ( .A1(n8591), .A2(n13380), .ZN(n8550) );
  NAND2_X1 U11002 ( .A1(n8576), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8549) );
  XNOR2_X1 U11003 ( .A(n8554), .B(n8553), .ZN(n11975) );
  NAND2_X1 U11004 ( .A1(n11975), .A2(n9460), .ZN(n8556) );
  NAND2_X1 U11005 ( .A1(n9459), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8555) );
  NAND2_X1 U11006 ( .A1(n8558), .A2(n8557), .ZN(n8559) );
  NAND2_X1 U11007 ( .A1(n13592), .A2(n9460), .ZN(n8562) );
  NAND2_X1 U11008 ( .A1(n9459), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8561) );
  NAND2_X1 U11009 ( .A1(n6482), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8570) );
  INV_X1 U11010 ( .A(n8563), .ZN(n8572) );
  INV_X1 U11011 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8564) );
  NAND2_X1 U11012 ( .A1(n8565), .A2(n8564), .ZN(n8566) );
  NAND2_X1 U11013 ( .A1(n8575), .A2(n13366), .ZN(n8569) );
  NAND2_X1 U11014 ( .A1(n9453), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8568) );
  NAND2_X1 U11015 ( .A1(n8576), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8567) );
  NAND4_X1 U11016 ( .A1(n8570), .A2(n8569), .A3(n8568), .A4(n8567), .ZN(n13284) );
  XNOR2_X1 U11017 ( .A(n13497), .B(n13284), .ZN(n13370) );
  INV_X1 U11018 ( .A(n13284), .ZN(n13188) );
  NAND2_X1 U11019 ( .A1(n6482), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8580) );
  INV_X1 U11020 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8571) );
  NAND2_X1 U11021 ( .A1(n8572), .A2(n8571), .ZN(n8573) );
  NAND2_X1 U11022 ( .A1(n8575), .A2(n13352), .ZN(n8579) );
  NAND2_X1 U11023 ( .A1(n9453), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8578) );
  NAND2_X1 U11024 ( .A1(n8576), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8577) );
  NAND4_X1 U11025 ( .A1(n8580), .A2(n8579), .A3(n8578), .A4(n8577), .ZN(n13283) );
  XNOR2_X1 U11026 ( .A(n8582), .B(SI_27_), .ZN(n8583) );
  NAND2_X1 U11027 ( .A1(n9459), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8584) );
  NAND2_X1 U11028 ( .A1(n13487), .A2(n13282), .ZN(n8678) );
  MUX2_X1 U11029 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n6475), .Z(n9324) );
  INV_X1 U11030 ( .A(SI_29_), .ZN(n13135) );
  XNOR2_X1 U11031 ( .A(n9324), .B(n13135), .ZN(n9322) );
  XNOR2_X1 U11032 ( .A(n9323), .B(n9322), .ZN(n13581) );
  NAND2_X1 U11033 ( .A1(n13581), .A2(n9460), .ZN(n8590) );
  NAND2_X1 U11034 ( .A1(n9459), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8589) );
  NAND2_X1 U11035 ( .A1(n9453), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8595) );
  NAND2_X1 U11036 ( .A1(n8576), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8594) );
  NAND2_X1 U11037 ( .A1(n8591), .A2(n8688), .ZN(n8593) );
  NAND2_X1 U11038 ( .A1(n6482), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8592) );
  AND4_X1 U11039 ( .A1(n8595), .A2(n8594), .A3(n8593), .A4(n8592), .ZN(n12214)
         );
  XNOR2_X1 U11040 ( .A(n13482), .B(n13281), .ZN(n9657) );
  NAND2_X1 U11041 ( .A1(n8597), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8598) );
  MUX2_X1 U11042 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8598), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n8599) );
  INV_X1 U11043 ( .A(n8623), .ZN(n8636) );
  NAND2_X1 U11044 ( .A1(n8683), .A2(n11533), .ZN(n8607) );
  NAND2_X1 U11045 ( .A1(n8601), .A2(n8600), .ZN(n8603) );
  XNOR2_X1 U11046 ( .A(n8602), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8682) );
  INV_X1 U11047 ( .A(n8681), .ZN(n9667) );
  NAND2_X1 U11048 ( .A1(n9666), .A2(n9667), .ZN(n8606) );
  INV_X1 U11049 ( .A(n8608), .ZN(n8609) );
  INV_X1 U11050 ( .A(n13588), .ZN(n10208) );
  NAND2_X1 U11051 ( .A1(n10473), .A2(n8608), .ZN(n13256) );
  AOI21_X1 U11052 ( .B1(n10208), .B2(P2_B_REG_SCAN_IN), .A(n13256), .ZN(n13324) );
  INV_X1 U11053 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8612) );
  NAND2_X1 U11054 ( .A1(n9453), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8611) );
  NAND2_X1 U11055 ( .A1(n8576), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8610) );
  OAI211_X1 U11056 ( .C1(n9457), .C2(n8612), .A(n8611), .B(n8610), .ZN(n13280)
         );
  AOI22_X1 U11057 ( .A1(n13282), .A2(n13171), .B1(n13324), .B2(n13280), .ZN(
        n8613) );
  NOR2_X1 U11058 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n8618) );
  NOR4_X1 U11059 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n8617) );
  NOR4_X1 U11060 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n8616) );
  NOR4_X1 U11061 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n8615) );
  NAND4_X1 U11062 ( .A1(n8618), .A2(n8617), .A3(n8616), .A4(n8615), .ZN(n8634)
         );
  NOR4_X1 U11063 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n8622) );
  NOR4_X1 U11064 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n8621) );
  NOR4_X1 U11065 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8620) );
  NOR4_X1 U11066 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n8619) );
  NAND4_X1 U11067 ( .A1(n8622), .A2(n8621), .A3(n8620), .A4(n8619), .ZN(n8633)
         );
  NAND2_X1 U11068 ( .A1(n8623), .A2(n8637), .ZN(n8625) );
  NAND2_X1 U11069 ( .A1(n8625), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8624) );
  MUX2_X1 U11070 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8624), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n8626) );
  INV_X1 U11071 ( .A(P2_B_REG_SCAN_IN), .ZN(n8627) );
  XNOR2_X1 U11072 ( .A(n11942), .B(n8627), .ZN(n8629) );
  NAND2_X1 U11073 ( .A1(n8630), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8628) );
  INV_X1 U11074 ( .A(n8639), .ZN(n11976) );
  NAND2_X1 U11075 ( .A1(n8629), .A2(n11976), .ZN(n8632) );
  AND2_X1 U11076 ( .A1(n8632), .A2(n13594), .ZN(n14737) );
  OAI21_X1 U11077 ( .B1(n8634), .B2(n8633), .A(n14737), .ZN(n10441) );
  INV_X1 U11078 ( .A(n10441), .ZN(n8635) );
  INV_X1 U11079 ( .A(n8683), .ZN(n14720) );
  NAND2_X1 U11080 ( .A1(n14720), .A2(n8681), .ZN(n10472) );
  AND2_X1 U11081 ( .A1(n10472), .A2(n10473), .ZN(n10443) );
  OR2_X1 U11082 ( .A1(n8635), .A2(n10443), .ZN(n10845) );
  INV_X1 U11083 ( .A(n10845), .ZN(n8643) );
  NAND3_X1 U11084 ( .A1(n13594), .A2(n11942), .A3(n8639), .ZN(n10059) );
  NAND2_X1 U11085 ( .A1(n8636), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8638) );
  XNOR2_X1 U11086 ( .A(n8638), .B(n8637), .ZN(n10195) );
  AND2_X1 U11087 ( .A1(n10059), .A2(n10195), .ZN(n10444) );
  INV_X1 U11088 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14744) );
  NOR2_X1 U11089 ( .A1(n13594), .A2(n8639), .ZN(n8640) );
  AOI21_X1 U11090 ( .B1(n14737), .B2(n14744), .A(n8640), .ZN(n10847) );
  INV_X1 U11091 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14739) );
  NAND2_X1 U11092 ( .A1(n14737), .A2(n14739), .ZN(n8642) );
  NAND2_X1 U11093 ( .A1(n8642), .A2(n8641), .ZN(n14740) );
  NAND4_X1 U11094 ( .A1(n8643), .A2(n14741), .A3(n10847), .A4(n14740), .ZN(
        n8644) );
  INV_X1 U11095 ( .A(n14741), .ZN(n14743) );
  INV_X1 U11096 ( .A(n13374), .ZN(n13385) );
  NAND2_X1 U11097 ( .A1(n10969), .A2(n10968), .ZN(n8646) );
  NAND2_X1 U11098 ( .A1(n10866), .A2(n14759), .ZN(n8645) );
  NAND2_X1 U11099 ( .A1(n8646), .A2(n8645), .ZN(n10862) );
  NAND2_X1 U11100 ( .A1(n10862), .A2(n8647), .ZN(n8650) );
  NAND2_X1 U11101 ( .A1(n8648), .A2(n10869), .ZN(n8649) );
  NAND2_X1 U11102 ( .A1(n8650), .A2(n8649), .ZN(n10995) );
  NAND2_X1 U11103 ( .A1(n10995), .A2(n10998), .ZN(n8652) );
  NAND2_X1 U11104 ( .A1(n10867), .A2(n14776), .ZN(n8651) );
  NOR2_X1 U11105 ( .A1(n11129), .A2(n13305), .ZN(n8653) );
  NAND2_X1 U11106 ( .A1(n11129), .A2(n13305), .ZN(n8654) );
  INV_X1 U11107 ( .A(n10826), .ZN(n10833) );
  NAND2_X1 U11108 ( .A1(n10911), .A2(n13304), .ZN(n8655) );
  OR2_X1 U11109 ( .A1(n14789), .A2(n13303), .ZN(n8657) );
  XNOR2_X1 U11110 ( .A(n14710), .B(n9523), .ZN(n14708) );
  NAND2_X1 U11111 ( .A1(n14710), .A2(n13301), .ZN(n8658) );
  NAND2_X1 U11112 ( .A1(n14813), .A2(n13300), .ZN(n8659) );
  OR2_X1 U11113 ( .A1(n11382), .A2(n13299), .ZN(n8660) );
  NAND2_X1 U11114 ( .A1(n11382), .A2(n13299), .ZN(n8661) );
  AND2_X1 U11115 ( .A1(n11443), .A2(n13298), .ZN(n8662) );
  NAND2_X1 U11116 ( .A1(n8663), .A2(n7382), .ZN(n8665) );
  NAND2_X1 U11117 ( .A1(n11504), .A2(n13297), .ZN(n8664) );
  AND2_X1 U11118 ( .A1(n13557), .A2(n13296), .ZN(n8667) );
  OR2_X1 U11119 ( .A1(n13557), .A2(n13296), .ZN(n8666) );
  XNOR2_X1 U11120 ( .A(n12161), .B(n13295), .ZN(n9650) );
  XNOR2_X1 U11121 ( .A(n13553), .B(n13294), .ZN(n11892) );
  NAND2_X1 U11122 ( .A1(n13553), .A2(n13294), .ZN(n8668) );
  NAND2_X1 U11123 ( .A1(n13547), .A2(n13293), .ZN(n8669) );
  XNOR2_X1 U11124 ( .A(n12171), .B(n13292), .ZN(n11951) );
  OR2_X1 U11125 ( .A1(n12171), .A2(n13292), .ZN(n8670) );
  NOR2_X1 U11126 ( .A1(n13537), .A2(n13291), .ZN(n8671) );
  AND2_X1 U11127 ( .A1(n13531), .A2(n13290), .ZN(n8673) );
  OR2_X1 U11128 ( .A1(n13531), .A2(n13290), .ZN(n8672) );
  XNOR2_X1 U11129 ( .A(n13526), .B(n13235), .ZN(n13436) );
  NAND2_X1 U11130 ( .A1(n8687), .A2(n13235), .ZN(n8674) );
  NAND2_X1 U11131 ( .A1(n13518), .A2(n13288), .ZN(n8675) );
  NAND2_X1 U11132 ( .A1(n13411), .A2(n13234), .ZN(n8677) );
  AND2_X1 U11133 ( .A1(n13514), .A2(n13287), .ZN(n8676) );
  INV_X1 U11134 ( .A(n13497), .ZN(n13368) );
  XNOR2_X1 U11135 ( .A(n8685), .B(n11533), .ZN(n8684) );
  OR2_X2 U11136 ( .A1(n8684), .A2(n8683), .ZN(n10449) );
  NAND2_X1 U11137 ( .A1(n8683), .A2(n10447), .ZN(n10828) );
  NAND2_X1 U11138 ( .A1(n10449), .A2(n10828), .ZN(n8686) );
  NOR2_X1 U11139 ( .A1(n13480), .A2(n14715), .ZN(n8694) );
  AND2_X1 U11140 ( .A1(n14755), .A2(n14721), .ZN(n11177) );
  NAND2_X1 U11141 ( .A1(n11177), .A2(n14759), .ZN(n10977) );
  NOR2_X1 U11142 ( .A1(n10977), .A2(n14766), .ZN(n11004) );
  NAND2_X1 U11143 ( .A1(n11004), .A2(n14776), .ZN(n11125) );
  OR2_X1 U11144 ( .A1(n11125), .A2(n11129), .ZN(n11126) );
  OR2_X1 U11145 ( .A1(n11126), .A2(n10911), .ZN(n10882) );
  INV_X1 U11146 ( .A(n11154), .ZN(n14797) );
  INV_X1 U11147 ( .A(n11382), .ZN(n14823) );
  INV_X1 U11148 ( .A(n11443), .ZN(n14385) );
  NAND2_X1 U11149 ( .A1(n11441), .A2(n14385), .ZN(n11456) );
  INV_X1 U11150 ( .A(n13547), .ZN(n13216) );
  AND2_X2 U11151 ( .A1(n11963), .A2(n13216), .ZN(n11964) );
  OR2_X2 U11152 ( .A1(n13518), .A2(n13431), .ZN(n13418) );
  AND2_X2 U11153 ( .A1(n13396), .A2(n13409), .ZN(n13392) );
  NOR2_X1 U11154 ( .A1(n13482), .A2(n13340), .ZN(n13329) );
  AOI211_X1 U11155 ( .C1(n13482), .C2(n13340), .A(n11505), .B(n13329), .ZN(
        n13481) );
  NAND2_X1 U11156 ( .A1(n14745), .A2(n9667), .ZN(n10475) );
  INV_X1 U11157 ( .A(n10475), .ZN(n14719) );
  AOI22_X1 U11158 ( .A1(n14736), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n8688), 
        .B2(n14705), .ZN(n8689) );
  OAI21_X1 U11159 ( .B1(n9458), .B2(n13453), .A(n8689), .ZN(n8690) );
  INV_X1 U11160 ( .A(n8690), .ZN(n8691) );
  INV_X2 U11161 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8728) );
  NOR2_X1 U11162 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n8699) );
  NOR2_X1 U11163 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), 
        .ZN(n8698) );
  NOR2_X1 U11164 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), 
        .ZN(n8697) );
  NOR2_X1 U11165 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .ZN(n8702) );
  NOR3_X1 U11166 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), 
        .A3(P1_IR_REG_26__SCAN_IN), .ZN(n8706) );
  NOR2_X1 U11167 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), 
        .ZN(n8705) );
  NOR2_X1 U11168 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n8704) );
  NAND2_X1 U11169 ( .A1(n8706), .A2(n9122), .ZN(n8721) );
  NOR2_X1 U11170 ( .A1(n8721), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n8707) );
  NAND2_X1 U11171 ( .A1(n8709), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8710) );
  AND2_X4 U11172 ( .A1(n6474), .A2(n8716), .ZN(n8766) );
  NAND2_X1 U11173 ( .A1(n8766), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n8715) );
  INV_X1 U11174 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n8711) );
  OR2_X1 U11175 ( .A1(n9109), .A2(n8711), .ZN(n8714) );
  NAND2_X1 U11176 ( .A1(n8767), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n8713) );
  INV_X1 U11177 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n13790) );
  OR2_X1 U11178 ( .A1(n8768), .A2(n13790), .ZN(n8718) );
  NAND2_X1 U11179 ( .A1(n8774), .A2(n10130), .ZN(n8732) );
  OR2_X1 U11180 ( .A1(n8759), .A2(n10131), .ZN(n8731) );
  OR2_X1 U11181 ( .A1(n8727), .A2(n14236), .ZN(n8729) );
  XNOR2_X1 U11182 ( .A(n8729), .B(n8728), .ZN(n13789) );
  OR2_X1 U11183 ( .A1(n8739), .A2(n13789), .ZN(n8730) );
  AND3_X4 U11184 ( .A1(n8732), .A2(n8731), .A3(n8730), .ZN(n14503) );
  NAND2_X1 U11185 ( .A1(n13773), .A2(n14503), .ZN(n8733) );
  INV_X1 U11186 ( .A(n10752), .ZN(n8752) );
  NAND2_X1 U11187 ( .A1(n8767), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n8737) );
  NAND2_X1 U11188 ( .A1(n8983), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n8736) );
  NAND4_X2 U11189 ( .A1(n8737), .A2(n8736), .A3(n8735), .A4(n8734), .ZN(n13774) );
  INV_X1 U11190 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n8738) );
  OR2_X1 U11191 ( .A1(n8739), .A2(n10379), .ZN(n8740) );
  NAND2_X1 U11192 ( .A1(n13774), .A2(n10087), .ZN(n9174) );
  NAND2_X1 U11193 ( .A1(n8983), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n8746) );
  NAND2_X1 U11194 ( .A1(n8766), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n8744) );
  NAND2_X1 U11195 ( .A1(n8767), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n8743) );
  INV_X1 U11196 ( .A(n14256), .ZN(n12152) );
  INV_X1 U11197 ( .A(SI_0_), .ZN(n8748) );
  OAI21_X1 U11198 ( .B1(n6706), .B2(n8748), .A(n8747), .ZN(n8749) );
  NAND2_X1 U11199 ( .A1(n8750), .A2(n8749), .ZN(n14255) );
  NAND2_X1 U11200 ( .A1(n8739), .A2(n14255), .ZN(n8751) );
  AND2_X1 U11201 ( .A1(n13776), .A2(n10730), .ZN(n10728) );
  NAND2_X1 U11202 ( .A1(n10693), .A2(n14503), .ZN(n8753) );
  NAND2_X1 U11203 ( .A1(n8754), .A2(n8753), .ZN(n10699) );
  NAND2_X1 U11204 ( .A1(n8767), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n8758) );
  NAND2_X1 U11205 ( .A1(n8742), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n8757) );
  NAND2_X1 U11206 ( .A1(n8766), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n8756) );
  OR2_X1 U11207 ( .A1(n8768), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n8755) );
  NAND2_X1 U11208 ( .A1(n8760), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8762) );
  INV_X1 U11209 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n8761) );
  XNOR2_X1 U11210 ( .A(n8762), .B(n8761), .ZN(n13812) );
  OR2_X1 U11211 ( .A1(n8739), .A2(n13812), .ZN(n8763) );
  NAND2_X1 U11212 ( .A1(n10699), .A2(n7350), .ZN(n8765) );
  INV_X1 U11213 ( .A(n13772), .ZN(n9193) );
  INV_X1 U11214 ( .A(n10714), .ZN(n14514) );
  NAND2_X1 U11215 ( .A1(n9193), .A2(n14514), .ZN(n8764) );
  NAND2_X1 U11216 ( .A1(n8766), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n8773) );
  INV_X1 U11217 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10381) );
  OR2_X1 U11218 ( .A1(n8991), .A2(n10381), .ZN(n8772) );
  XNOR2_X1 U11219 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n11123) );
  OR2_X1 U11220 ( .A1(n9107), .A2(n11123), .ZN(n8771) );
  INV_X1 U11221 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n8769) );
  OR2_X1 U11222 ( .A1(n9109), .A2(n8769), .ZN(n8770) );
  NAND2_X1 U11223 ( .A1(n10132), .A2(n8774), .ZN(n8777) );
  OR2_X1 U11224 ( .A1(n8760), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n8784) );
  NAND2_X1 U11225 ( .A1(n8784), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8775) );
  XNOR2_X1 U11226 ( .A(n8775), .B(P1_IR_REG_4__SCAN_IN), .ZN(n10382) );
  AOI22_X1 U11227 ( .A1(n8958), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n8957), .B2(
        n10382), .ZN(n8776) );
  AND2_X2 U11228 ( .A1(n8777), .A2(n8776), .ZN(n14520) );
  NAND2_X1 U11229 ( .A1(n11071), .A2(n14520), .ZN(n9373) );
  INV_X1 U11230 ( .A(n9373), .ZN(n8778) );
  INV_X1 U11231 ( .A(n11071), .ZN(n13771) );
  INV_X1 U11232 ( .A(n14520), .ZN(n11120) );
  NAND2_X1 U11233 ( .A1(n13771), .A2(n11120), .ZN(n9372) );
  NAND2_X1 U11234 ( .A1(n9334), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n8783) );
  NAND2_X1 U11235 ( .A1(n8742), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n8782) );
  AOI21_X1 U11236 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n8779) );
  NOR2_X1 U11237 ( .A1(n8779), .A2(n8797), .ZN(n11994) );
  NAND2_X1 U11238 ( .A1(n8983), .A2(n11994), .ZN(n8781) );
  NAND2_X1 U11239 ( .A1(n8766), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n8780) );
  NAND4_X1 U11240 ( .A1(n8783), .A2(n8782), .A3(n8781), .A4(n8780), .ZN(n13770) );
  NAND2_X1 U11241 ( .A1(n10135), .A2(n8774), .ZN(n8792) );
  INV_X1 U11242 ( .A(n8784), .ZN(n8785) );
  NAND2_X1 U11243 ( .A1(n8785), .A2(n6813), .ZN(n8787) );
  NAND2_X1 U11244 ( .A1(n8787), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8786) );
  MUX2_X1 U11245 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8786), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n8790) );
  INV_X1 U11246 ( .A(n8787), .ZN(n8789) );
  NAND2_X1 U11247 ( .A1(n8789), .A2(n8788), .ZN(n8803) );
  AOI22_X1 U11248 ( .A1(n8958), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n8957), .B2(
        n10384), .ZN(n8791) );
  XNOR2_X1 U11249 ( .A(n11078), .B(n11990), .ZN(n11981) );
  INV_X1 U11250 ( .A(n11981), .ZN(n11983) );
  OR2_X1 U11251 ( .A1(n13770), .A2(n11990), .ZN(n8793) );
  NAND2_X1 U11252 ( .A1(n11986), .A2(n8793), .ZN(n10759) );
  NAND2_X1 U11253 ( .A1(n10151), .A2(n8774), .ZN(n8796) );
  NAND2_X1 U11254 ( .A1(n8803), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8794) );
  XNOR2_X1 U11255 ( .A(n8794), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10385) );
  AOI22_X1 U11256 ( .A1(n8958), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n8957), .B2(
        n10385), .ZN(n8795) );
  NAND2_X1 U11257 ( .A1(n8796), .A2(n8795), .ZN(n14537) );
  NAND2_X1 U11258 ( .A1(n8766), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n8801) );
  NAND2_X1 U11259 ( .A1(n9334), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n8800) );
  NAND2_X1 U11260 ( .A1(n8742), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n8799) );
  NAND2_X1 U11261 ( .A1(n8797), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8820) );
  OAI21_X1 U11262 ( .B1(n8797), .B2(P1_REG3_REG_6__SCAN_IN), .A(n8820), .ZN(
        n11424) );
  OR2_X1 U11263 ( .A1(n9107), .A2(n11424), .ZN(n8798) );
  NAND4_X1 U11264 ( .A1(n8801), .A2(n8800), .A3(n8799), .A4(n8798), .ZN(n13769) );
  XNOR2_X1 U11265 ( .A(n14537), .B(n13769), .ZN(n9375) );
  NAND2_X1 U11266 ( .A1(n10759), .A2(n10758), .ZN(n10757) );
  OR2_X1 U11267 ( .A1(n14537), .A2(n13769), .ZN(n8802) );
  NAND2_X1 U11268 ( .A1(n10757), .A2(n8802), .ZN(n11195) );
  NAND2_X1 U11269 ( .A1(n10164), .A2(n8774), .ZN(n8806) );
  OAI21_X1 U11270 ( .B1(n8803), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8804) );
  XNOR2_X1 U11271 ( .A(n8804), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10429) );
  AOI22_X1 U11272 ( .A1(n8958), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n8957), .B2(
        n10429), .ZN(n8805) );
  NAND2_X1 U11273 ( .A1(n9334), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n8811) );
  NAND2_X1 U11274 ( .A1(n8742), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n8810) );
  INV_X1 U11275 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n8807) );
  XNOR2_X1 U11276 ( .A(n8820), .B(n8807), .ZN(n14476) );
  OR2_X1 U11277 ( .A1(n9107), .A2(n14476), .ZN(n8809) );
  NAND2_X1 U11278 ( .A1(n8766), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n8808) );
  NAND4_X1 U11279 ( .A1(n8811), .A2(n8810), .A3(n8809), .A4(n8808), .ZN(n13768) );
  XNOR2_X1 U11280 ( .A(n14475), .B(n13768), .ZN(n9376) );
  INV_X1 U11281 ( .A(n9376), .ZN(n11200) );
  NAND2_X1 U11282 ( .A1(n11195), .A2(n11200), .ZN(n11194) );
  OR2_X1 U11283 ( .A1(n14475), .A2(n13768), .ZN(n8812) );
  NAND2_X1 U11284 ( .A1(n10170), .A2(n8774), .ZN(n8817) );
  NAND2_X1 U11285 ( .A1(n8814), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8815) );
  XNOR2_X1 U11286 ( .A(n8815), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10549) );
  AOI22_X1 U11287 ( .A1(n8958), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n8957), .B2(
        n10549), .ZN(n8816) );
  NAND2_X1 U11288 ( .A1(n8817), .A2(n8816), .ZN(n11552) );
  NAND2_X1 U11289 ( .A1(n8766), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n8825) );
  NAND2_X1 U11290 ( .A1(n9334), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n8824) );
  NAND2_X1 U11291 ( .A1(n8742), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n8823) );
  INV_X1 U11292 ( .A(n8820), .ZN(n8818) );
  AOI21_X1 U11293 ( .B1(n8818), .B2(P1_REG3_REG_7__SCAN_IN), .A(
        P1_REG3_REG_8__SCAN_IN), .ZN(n8821) );
  NAND2_X1 U11294 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n8819) );
  NOR2_X1 U11295 ( .A1(n8820), .A2(n8819), .ZN(n8834) );
  OR2_X1 U11296 ( .A1(n8821), .A2(n8834), .ZN(n11559) );
  OR2_X1 U11297 ( .A1(n9107), .A2(n11559), .ZN(n8822) );
  NAND4_X1 U11298 ( .A1(n8825), .A2(n8824), .A3(n8823), .A4(n8822), .ZN(n13767) );
  XNOR2_X1 U11299 ( .A(n11552), .B(n13767), .ZN(n10953) );
  INV_X1 U11300 ( .A(n10953), .ZN(n10963) );
  OR2_X1 U11301 ( .A1(n11552), .A2(n13767), .ZN(n8826) );
  NAND2_X1 U11302 ( .A1(n10190), .A2(n8774), .ZN(n8833) );
  NOR2_X1 U11303 ( .A1(n8814), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n8829) );
  NOR2_X1 U11304 ( .A1(n8829), .A2(n14236), .ZN(n8827) );
  MUX2_X1 U11305 ( .A(n14236), .B(n8827), .S(P1_IR_REG_9__SCAN_IN), .Z(n8831)
         );
  INV_X1 U11306 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8828) );
  NAND2_X1 U11307 ( .A1(n8829), .A2(n8828), .ZN(n8848) );
  INV_X1 U11308 ( .A(n8848), .ZN(n8830) );
  AOI22_X1 U11309 ( .A1(n8958), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n8957), .B2(
        n13834), .ZN(n8832) );
  NAND2_X1 U11310 ( .A1(n8766), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n8839) );
  NAND2_X1 U11311 ( .A1(n9334), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n8838) );
  NAND2_X1 U11312 ( .A1(n8742), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n8837) );
  NAND2_X1 U11313 ( .A1(n8834), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n8854) );
  OR2_X1 U11314 ( .A1(n8834), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n8835) );
  NAND2_X1 U11315 ( .A1(n8854), .A2(n8835), .ZN(n11849) );
  OR2_X1 U11316 ( .A1(n9107), .A2(n11849), .ZN(n8836) );
  NAND4_X1 U11317 ( .A1(n8839), .A2(n8838), .A3(n8837), .A4(n8836), .ZN(n13766) );
  INV_X1 U11318 ( .A(n13766), .ZN(n10955) );
  XNOR2_X1 U11319 ( .A(n11851), .B(n10955), .ZN(n11059) );
  NAND2_X1 U11320 ( .A1(n10220), .A2(n8774), .ZN(n8842) );
  NAND2_X1 U11321 ( .A1(n8848), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8840) );
  XNOR2_X1 U11322 ( .A(n8840), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10677) );
  AOI22_X1 U11323 ( .A1(n8958), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n8957), 
        .B2(n10677), .ZN(n8841) );
  NAND2_X1 U11324 ( .A1(n8766), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8846) );
  NAND2_X1 U11325 ( .A1(n9334), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n8845) );
  NAND2_X1 U11326 ( .A1(n8742), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n8844) );
  XNOR2_X1 U11327 ( .A(n8854), .B(n8852), .ZN(n11881) );
  OR2_X1 U11328 ( .A1(n9107), .A2(n11881), .ZN(n8843) );
  NAND4_X1 U11329 ( .A1(n8846), .A2(n8845), .A3(n8844), .A4(n8843), .ZN(n13765) );
  XNOR2_X1 U11330 ( .A(n11883), .B(n13765), .ZN(n9379) );
  OR2_X1 U11331 ( .A1(n11883), .A2(n13765), .ZN(n8847) );
  NAND2_X1 U11332 ( .A1(n11245), .A2(n8847), .ZN(n11296) );
  NAND2_X1 U11333 ( .A1(n10235), .A2(n8774), .ZN(n8851) );
  NAND2_X1 U11334 ( .A1(n8861), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8849) );
  XNOR2_X1 U11335 ( .A(n8849), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10817) );
  AOI22_X1 U11336 ( .A1(n8958), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n8957), 
        .B2(n10817), .ZN(n8850) );
  NAND2_X1 U11337 ( .A1(n8742), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n8859) );
  INV_X1 U11338 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n8853) );
  OAI21_X1 U11339 ( .B1(n8854), .B2(n8852), .A(n8853), .ZN(n8855) );
  NAND2_X1 U11340 ( .A1(n8855), .A2(n8866), .ZN(n14416) );
  OR2_X1 U11341 ( .A1(n9107), .A2(n14416), .ZN(n8858) );
  INV_X1 U11342 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10678) );
  OR2_X1 U11343 ( .A1(n9338), .A2(n10678), .ZN(n8857) );
  INV_X1 U11344 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11299) );
  OR2_X1 U11345 ( .A1(n8991), .A2(n11299), .ZN(n8856) );
  XNOR2_X1 U11346 ( .A(n14413), .B(n13764), .ZN(n9380) );
  INV_X1 U11347 ( .A(n9380), .ZN(n11295) );
  NAND2_X1 U11348 ( .A1(n11296), .A2(n11295), .ZN(n11294) );
  NAND2_X1 U11349 ( .A1(n14426), .A2(n12007), .ZN(n8860) );
  NAND2_X1 U11350 ( .A1(n11294), .A2(n8860), .ZN(n11409) );
  NAND2_X1 U11351 ( .A1(n10321), .A2(n8774), .ZN(n8863) );
  OAI21_X1 U11352 ( .B1(n8861), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8875) );
  XNOR2_X1 U11353 ( .A(n8875), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11021) );
  AOI22_X1 U11354 ( .A1(n8958), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n8957), 
        .B2(n11021), .ZN(n8862) );
  INV_X1 U11355 ( .A(n13652), .ZN(n11418) );
  NAND2_X1 U11356 ( .A1(n8742), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n8872) );
  INV_X1 U11357 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n8864) );
  OR2_X1 U11358 ( .A1(n9338), .A2(n8864), .ZN(n8871) );
  INV_X1 U11359 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11416) );
  OR2_X1 U11360 ( .A1(n8991), .A2(n11416), .ZN(n8870) );
  INV_X1 U11361 ( .A(n8879), .ZN(n8868) );
  NAND2_X1 U11362 ( .A1(n8866), .A2(n8865), .ZN(n8867) );
  NAND2_X1 U11363 ( .A1(n8868), .A2(n8867), .ZN(n13645) );
  OR2_X1 U11364 ( .A1(n9107), .A2(n13645), .ZN(n8869) );
  XNOR2_X1 U11365 ( .A(n11418), .B(n13763), .ZN(n11411) );
  NAND2_X1 U11366 ( .A1(n11409), .A2(n7347), .ZN(n11408) );
  NAND2_X1 U11367 ( .A1(n13652), .A2(n12016), .ZN(n8873) );
  NAND2_X1 U11368 ( .A1(n11408), .A2(n8873), .ZN(n11469) );
  NAND2_X1 U11369 ( .A1(n10400), .A2(n8774), .ZN(n8878) );
  INV_X1 U11370 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n8874) );
  NAND2_X1 U11371 ( .A1(n8875), .A2(n8874), .ZN(n8876) );
  NAND2_X1 U11372 ( .A1(n8876), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8887) );
  XNOR2_X1 U11373 ( .A(n8887), .B(P1_IR_REG_13__SCAN_IN), .ZN(n11212) );
  AOI22_X1 U11374 ( .A1(n8958), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n11212), 
        .B2(n8957), .ZN(n8877) );
  NAND2_X1 U11375 ( .A1(n9334), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n8884) );
  NAND2_X1 U11376 ( .A1(n8742), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n8883) );
  NAND2_X1 U11377 ( .A1(n8766), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n8882) );
  NAND2_X1 U11378 ( .A1(n8879), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8893) );
  OR2_X1 U11379 ( .A1(n8879), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8880) );
  NAND2_X1 U11380 ( .A1(n8893), .A2(n8880), .ZN(n13695) );
  OR2_X1 U11381 ( .A1(n9107), .A2(n13695), .ZN(n8881) );
  NAND4_X1 U11382 ( .A1(n8884), .A2(n8883), .A3(n8882), .A4(n8881), .ZN(n13762) );
  INV_X1 U11383 ( .A(n13762), .ZN(n12022) );
  XNOR2_X1 U11384 ( .A(n12024), .B(n12022), .ZN(n11474) );
  NAND2_X1 U11385 ( .A1(n11469), .A2(n11474), .ZN(n11468) );
  OR2_X1 U11386 ( .A1(n12024), .A2(n13762), .ZN(n8885) );
  NAND2_X1 U11387 ( .A1(n10596), .A2(n8774), .ZN(n8891) );
  INV_X1 U11388 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8886) );
  NAND2_X1 U11389 ( .A1(n8887), .A2(n8886), .ZN(n8888) );
  NAND2_X1 U11390 ( .A1(n8888), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8889) );
  XNOR2_X1 U11391 ( .A(n8889), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11695) );
  AOI22_X1 U11392 ( .A1(n11695), .A2(n8957), .B1(n8958), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n8890) );
  NAND2_X1 U11393 ( .A1(n8742), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n8898) );
  INV_X1 U11394 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8892) );
  NAND2_X1 U11395 ( .A1(n8893), .A2(n8892), .ZN(n8894) );
  NAND2_X1 U11396 ( .A1(n8906), .A2(n8894), .ZN(n14402) );
  OR2_X1 U11397 ( .A1(n8768), .A2(n14402), .ZN(n8897) );
  INV_X1 U11398 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11216) );
  OR2_X1 U11399 ( .A1(n8991), .A2(n11216), .ZN(n8896) );
  INV_X1 U11400 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11210) );
  OR2_X1 U11401 ( .A1(n9338), .A2(n11210), .ZN(n8895) );
  NAND2_X1 U11402 ( .A1(n14419), .A2(n12029), .ZN(n9241) );
  INV_X1 U11403 ( .A(n12029), .ZN(n13761) );
  NAND2_X1 U11404 ( .A1(n14419), .A2(n13761), .ZN(n8900) );
  NAND2_X1 U11405 ( .A1(n10655), .A2(n8774), .ZN(n8904) );
  OR2_X1 U11406 ( .A1(n8901), .A2(n14236), .ZN(n8902) );
  XNOR2_X1 U11407 ( .A(n8902), .B(P1_IR_REG_15__SCAN_IN), .ZN(n14464) );
  AOI22_X1 U11408 ( .A1(n8958), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n8957), 
        .B2(n14464), .ZN(n8903) );
  NAND2_X1 U11409 ( .A1(n8742), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n8911) );
  INV_X1 U11410 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n11742) );
  OR2_X1 U11411 ( .A1(n8991), .A2(n11742), .ZN(n8910) );
  INV_X1 U11412 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14460) );
  OR2_X1 U11413 ( .A1(n9338), .A2(n14460), .ZN(n8909) );
  INV_X1 U11414 ( .A(n8919), .ZN(n8921) );
  NAND2_X1 U11415 ( .A1(n8906), .A2(n8905), .ZN(n8907) );
  NAND2_X1 U11416 ( .A1(n8921), .A2(n8907), .ZN(n11739) );
  OR2_X1 U11417 ( .A1(n9107), .A2(n11739), .ZN(n8908) );
  NAND2_X1 U11418 ( .A1(n12041), .A2(n11523), .ZN(n9252) );
  NAND2_X1 U11419 ( .A1(n9251), .A2(n9252), .ZN(n9386) );
  INV_X1 U11420 ( .A(n9386), .ZN(n8912) );
  INV_X1 U11421 ( .A(n11523), .ZN(n13760) );
  OR2_X1 U11422 ( .A1(n12041), .A2(n13760), .ZN(n8913) );
  NAND2_X1 U11423 ( .A1(n8914), .A2(n8913), .ZN(n11863) );
  NAND2_X1 U11424 ( .A1(n10569), .A2(n8774), .ZN(n8918) );
  AND2_X1 U11425 ( .A1(n8901), .A2(n8915), .ZN(n8930) );
  OR2_X1 U11426 ( .A1(n8930), .A2(n14236), .ZN(n8916) );
  XNOR2_X1 U11427 ( .A(n8916), .B(P1_IR_REG_16__SCAN_IN), .ZN(n13847) );
  AOI22_X1 U11428 ( .A1(n8958), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n8957), 
        .B2(n13847), .ZN(n8917) );
  NAND2_X1 U11429 ( .A1(n8742), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n8927) );
  INV_X1 U11430 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11864) );
  OR2_X1 U11431 ( .A1(n8991), .A2(n11864), .ZN(n8926) );
  INV_X1 U11432 ( .A(n8934), .ZN(n8936) );
  INV_X1 U11433 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8920) );
  NAND2_X1 U11434 ( .A1(n8921), .A2(n8920), .ZN(n8922) );
  NAND2_X1 U11435 ( .A1(n8936), .A2(n8922), .ZN(n13655) );
  OR2_X1 U11436 ( .A1(n8768), .A2(n13655), .ZN(n8925) );
  INV_X1 U11437 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n8923) );
  OR2_X1 U11438 ( .A1(n9338), .A2(n8923), .ZN(n8924) );
  XNOR2_X1 U11439 ( .A(n14189), .B(n13759), .ZN(n11856) );
  INV_X1 U11440 ( .A(n11856), .ZN(n11862) );
  NAND2_X1 U11441 ( .A1(n12049), .A2(n12048), .ZN(n8928) );
  NAND2_X1 U11442 ( .A1(n10671), .A2(n8774), .ZN(n8933) );
  NAND2_X1 U11443 ( .A1(n8930), .A2(n8929), .ZN(n8942) );
  NAND2_X1 U11444 ( .A1(n8942), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8931) );
  XNOR2_X1 U11445 ( .A(n8931), .B(P1_IR_REG_17__SCAN_IN), .ZN(n13855) );
  AOI22_X1 U11446 ( .A1(n8958), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n8957), 
        .B2(n13855), .ZN(n8932) );
  NAND2_X1 U11447 ( .A1(n8766), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n8941) );
  INV_X1 U11448 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8935) );
  NAND2_X1 U11449 ( .A1(n8936), .A2(n8935), .ZN(n8937) );
  NAND2_X1 U11450 ( .A1(n8949), .A2(n8937), .ZN(n13668) );
  OR2_X1 U11451 ( .A1(n8768), .A2(n13668), .ZN(n8940) );
  NAND2_X1 U11452 ( .A1(n9334), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8939) );
  NAND2_X1 U11453 ( .A1(n8742), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n8938) );
  NAND4_X1 U11454 ( .A1(n8941), .A2(n8940), .A3(n8939), .A4(n8938), .ZN(n13758) );
  OR2_X1 U11455 ( .A1(n13670), .A2(n13758), .ZN(n9369) );
  OR2_X1 U11456 ( .A1(n10875), .A2(n8978), .ZN(n8945) );
  NAND2_X1 U11457 ( .A1(n7378), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8943) );
  XNOR2_X1 U11458 ( .A(n8943), .B(P1_IR_REG_18__SCAN_IN), .ZN(n13875) );
  AOI22_X1 U11459 ( .A1(n8958), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n8957), 
        .B2(n13875), .ZN(n8944) );
  NAND2_X1 U11460 ( .A1(n9334), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8947) );
  INV_X1 U11461 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n14177) );
  OR2_X1 U11462 ( .A1(n9338), .A2(n14177), .ZN(n8946) );
  AND2_X1 U11463 ( .A1(n8947), .A2(n8946), .ZN(n8953) );
  INV_X1 U11464 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8948) );
  NAND2_X1 U11465 ( .A1(n8949), .A2(n8948), .ZN(n8950) );
  NAND2_X1 U11466 ( .A1(n8962), .A2(n8950), .ZN(n14078) );
  OR2_X1 U11467 ( .A1(n14078), .A2(n9107), .ZN(n8952) );
  NAND2_X1 U11468 ( .A1(n8742), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n8951) );
  INV_X1 U11469 ( .A(n13625), .ZN(n13757) );
  NAND2_X1 U11470 ( .A1(n14083), .A2(n13757), .ZN(n8954) );
  NAND2_X1 U11471 ( .A1(n10949), .A2(n8774), .ZN(n8960) );
  OAI21_X2 U11472 ( .B1(n7378), .B2(P1_IR_REG_18__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8956) );
  AOI22_X1 U11473 ( .A1(n8958), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14023), 
        .B2(n8957), .ZN(n8959) );
  INV_X1 U11474 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8961) );
  NAND2_X1 U11475 ( .A1(n8962), .A2(n8961), .ZN(n8963) );
  NAND2_X1 U11476 ( .A1(n8970), .A2(n8963), .ZN(n14066) );
  AOI22_X1 U11477 ( .A1(n8766), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n9334), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n8965) );
  NAND2_X1 U11478 ( .A1(n8742), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8964) );
  OAI211_X1 U11479 ( .C1(n14066), .C2(n9107), .A(n8965), .B(n8964), .ZN(n13756) );
  INV_X1 U11480 ( .A(n13756), .ZN(n8966) );
  OR2_X1 U11481 ( .A1(n12069), .A2(n8966), .ZN(n9265) );
  NAND2_X1 U11482 ( .A1(n12069), .A2(n8966), .ZN(n9266) );
  OR2_X1 U11483 ( .A1(n12069), .A2(n13756), .ZN(n8967) );
  NAND2_X1 U11484 ( .A1(n11148), .A2(n8774), .ZN(n8969) );
  OR2_X1 U11485 ( .A1(n8759), .A2(n11149), .ZN(n8968) );
  INV_X1 U11486 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13688) );
  AND2_X1 U11487 ( .A1(n8970), .A2(n13688), .ZN(n8971) );
  OR2_X1 U11488 ( .A1(n8971), .A2(n8981), .ZN(n14055) );
  INV_X1 U11489 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n8974) );
  NAND2_X1 U11490 ( .A1(n9334), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8973) );
  NAND2_X1 U11491 ( .A1(n8742), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n8972) );
  OAI211_X1 U11492 ( .C1(n8974), .C2(n9338), .A(n8973), .B(n8972), .ZN(n8975)
         );
  INV_X1 U11493 ( .A(n8975), .ZN(n8976) );
  OAI21_X1 U11494 ( .B1(n14055), .B2(n9107), .A(n8976), .ZN(n13755) );
  INV_X1 U11495 ( .A(n13755), .ZN(n9093) );
  XNOR2_X1 U11496 ( .A(n14222), .B(n9093), .ZN(n14043) );
  INV_X1 U11497 ( .A(n14043), .ZN(n14049) );
  NAND2_X1 U11498 ( .A1(n14222), .A2(n13755), .ZN(n8977) );
  OR2_X1 U11499 ( .A1(n11266), .A2(n8978), .ZN(n8980) );
  OR2_X1 U11500 ( .A1(n8759), .A2(n11250), .ZN(n8979) );
  OR2_X1 U11501 ( .A1(n8981), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8982) );
  NAND2_X1 U11502 ( .A1(n8981), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8992) );
  AND2_X1 U11503 ( .A1(n8982), .A2(n8992), .ZN(n14035) );
  NAND2_X1 U11504 ( .A1(n14035), .A2(n8983), .ZN(n8989) );
  INV_X1 U11505 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n8986) );
  NAND2_X1 U11506 ( .A1(n8742), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8985) );
  NAND2_X1 U11507 ( .A1(n9334), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8984) );
  OAI211_X1 U11508 ( .C1(n9338), .C2(n8986), .A(n8985), .B(n8984), .ZN(n8987)
         );
  INV_X1 U11509 ( .A(n8987), .ZN(n8988) );
  NAND2_X1 U11510 ( .A1(n8989), .A2(n8988), .ZN(n13754) );
  XNOR2_X1 U11511 ( .A(n14155), .B(n13754), .ZN(n14030) );
  NAND2_X1 U11512 ( .A1(n8506), .A2(n8726), .ZN(n8990) );
  XNOR2_X1 U11513 ( .A(n8990), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14254) );
  NAND2_X1 U11514 ( .A1(n8766), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n8998) );
  INV_X1 U11515 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n14012) );
  OR2_X1 U11516 ( .A1(n8991), .A2(n14012), .ZN(n8997) );
  NAND2_X1 U11517 ( .A1(n8993), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9001) );
  OAI21_X1 U11518 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n8993), .A(n9001), .ZN(
        n14011) );
  OR2_X1 U11519 ( .A1(n8768), .A2(n14011), .ZN(n8996) );
  INV_X1 U11520 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n8994) );
  OR2_X1 U11521 ( .A1(n9109), .A2(n8994), .ZN(n8995) );
  XNOR2_X1 U11522 ( .A(n14218), .B(n13634), .ZN(n9390) );
  NAND2_X1 U11523 ( .A1(n11752), .A2(n8774), .ZN(n9000) );
  INV_X1 U11524 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11755) );
  OR2_X1 U11525 ( .A1(n8759), .A2(n11755), .ZN(n8999) );
  NAND2_X2 U11526 ( .A1(n9000), .A2(n8999), .ZN(n14142) );
  NAND2_X1 U11527 ( .A1(n8766), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n9006) );
  NAND2_X1 U11528 ( .A1(n9334), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n9005) );
  NAND2_X1 U11529 ( .A1(n8742), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n9004) );
  NAND2_X1 U11530 ( .A1(n9002), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n9010) );
  OAI21_X1 U11531 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n9002), .A(n9010), .ZN(
        n14000) );
  OR2_X1 U11532 ( .A1(n8768), .A2(n14000), .ZN(n9003) );
  NAND4_X1 U11533 ( .A1(n9006), .A2(n9005), .A3(n9004), .A4(n9003), .ZN(n13752) );
  XNOR2_X1 U11534 ( .A(n14142), .B(n13752), .ZN(n13997) );
  NAND2_X1 U11535 ( .A1(n14142), .A2(n13752), .ZN(n9007) );
  OR2_X1 U11536 ( .A1(n8759), .A2(n11940), .ZN(n9008) );
  NAND2_X1 U11537 ( .A1(n9334), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n9015) );
  NAND2_X1 U11538 ( .A1(n8742), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n9014) );
  NAND2_X1 U11539 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(n9011), .ZN(n9021) );
  OAI21_X1 U11540 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n9011), .A(n9021), .ZN(
        n13987) );
  OR2_X1 U11541 ( .A1(n8768), .A2(n13987), .ZN(n9013) );
  NAND2_X1 U11542 ( .A1(n8766), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n9012) );
  NAND4_X1 U11543 ( .A1(n9015), .A2(n9014), .A3(n9013), .A4(n9012), .ZN(n13751) );
  INV_X1 U11544 ( .A(n13751), .ZN(n12113) );
  XNOR2_X1 U11545 ( .A(n14212), .B(n12113), .ZN(n13979) );
  OR2_X1 U11546 ( .A1(n14212), .A2(n13751), .ZN(n9016) );
  NAND2_X1 U11547 ( .A1(n11975), .A2(n8774), .ZN(n9018) );
  OR2_X1 U11548 ( .A1(n8759), .A2(n11978), .ZN(n9017) );
  NAND2_X1 U11549 ( .A1(n8766), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n9026) );
  NAND2_X1 U11550 ( .A1(n9334), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n9025) );
  NAND2_X1 U11551 ( .A1(n8742), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n9024) );
  INV_X1 U11552 ( .A(n9021), .ZN(n9019) );
  NAND2_X1 U11553 ( .A1(n9019), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n9031) );
  INV_X1 U11554 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9020) );
  NAND2_X1 U11555 ( .A1(n9021), .A2(n9020), .ZN(n9022) );
  NAND2_X1 U11556 ( .A1(n9031), .A2(n9022), .ZN(n13969) );
  OR2_X1 U11557 ( .A1(n8768), .A2(n13969), .ZN(n9023) );
  NAND4_X1 U11558 ( .A1(n9026), .A2(n9025), .A3(n9024), .A4(n9023), .ZN(n13750) );
  XNOR2_X1 U11559 ( .A(n14208), .B(n13750), .ZN(n13960) );
  INV_X1 U11560 ( .A(n13960), .ZN(n13963) );
  NAND2_X1 U11561 ( .A1(n13592), .A2(n8774), .ZN(n9028) );
  OR2_X1 U11562 ( .A1(n8759), .A2(n14249), .ZN(n9027) );
  NAND2_X1 U11563 ( .A1(n8766), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n9036) );
  NAND2_X1 U11564 ( .A1(n8767), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n9035) );
  NAND2_X1 U11565 ( .A1(n8742), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n9034) );
  INV_X1 U11566 ( .A(n9031), .ZN(n9029) );
  NAND2_X1 U11567 ( .A1(n9029), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n9042) );
  INV_X1 U11568 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9030) );
  NAND2_X1 U11569 ( .A1(n9031), .A2(n9030), .ZN(n9032) );
  NAND2_X1 U11570 ( .A1(n9042), .A2(n9032), .ZN(n13950) );
  OR2_X1 U11571 ( .A1(n8768), .A2(n13950), .ZN(n9033) );
  NAND4_X1 U11572 ( .A1(n9036), .A2(n9035), .A3(n9034), .A4(n9033), .ZN(n13749) );
  XNOR2_X1 U11573 ( .A(n14117), .B(n13749), .ZN(n13948) );
  INV_X1 U11574 ( .A(n13948), .ZN(n13945) );
  NAND2_X1 U11575 ( .A1(n14117), .A2(n13749), .ZN(n9037) );
  NAND2_X1 U11576 ( .A1(n13587), .A2(n8774), .ZN(n9039) );
  OR2_X1 U11577 ( .A1(n8759), .A2(n14246), .ZN(n9038) );
  NAND2_X1 U11578 ( .A1(n9334), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n9047) );
  NAND2_X1 U11579 ( .A1(n8742), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n9046) );
  NAND2_X1 U11580 ( .A1(n8766), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n9045) );
  INV_X1 U11581 ( .A(n9042), .ZN(n9040) );
  NAND2_X1 U11582 ( .A1(n9040), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n9051) );
  INV_X1 U11583 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9041) );
  NAND2_X1 U11584 ( .A1(n9042), .A2(n9041), .ZN(n9043) );
  NAND2_X1 U11585 ( .A1(n9051), .A2(n9043), .ZN(n13939) );
  OR2_X1 U11586 ( .A1(n8768), .A2(n13939), .ZN(n9044) );
  NAND4_X1 U11587 ( .A1(n9047), .A2(n9046), .A3(n9045), .A4(n9044), .ZN(n13748) );
  INV_X1 U11588 ( .A(n13748), .ZN(n9102) );
  XNOR2_X1 U11589 ( .A(n14203), .B(n9102), .ZN(n13932) );
  INV_X1 U11590 ( .A(n13932), .ZN(n13936) );
  INV_X1 U11591 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12297) );
  OR2_X1 U11592 ( .A1(n8759), .A2(n12297), .ZN(n9048) );
  NAND2_X1 U11593 ( .A1(n8766), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n9056) );
  NAND2_X1 U11594 ( .A1(n9334), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n9055) );
  NAND2_X1 U11595 ( .A1(n8742), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n9054) );
  INV_X1 U11596 ( .A(n9051), .ZN(n9050) );
  NAND2_X1 U11597 ( .A1(n9050), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n13911) );
  INV_X1 U11598 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n12290) );
  NAND2_X1 U11599 ( .A1(n9051), .A2(n12290), .ZN(n9052) );
  NAND2_X1 U11600 ( .A1(n13911), .A2(n9052), .ZN(n13924) );
  NAND4_X1 U11601 ( .A1(n9056), .A2(n9055), .A3(n9054), .A4(n9053), .ZN(n13914) );
  OR2_X1 U11602 ( .A1(n13926), .A2(n13914), .ZN(n9057) );
  NAND2_X1 U11603 ( .A1(n13926), .A2(n13914), .ZN(n13899) );
  INV_X1 U11604 ( .A(n9393), .ZN(n9058) );
  NAND2_X1 U11605 ( .A1(n9059), .A2(n9058), .ZN(n13900) );
  INV_X1 U11606 ( .A(n9059), .ZN(n9060) );
  NAND2_X1 U11607 ( .A1(n9060), .A2(n9393), .ZN(n9061) );
  MUX2_X1 U11608 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9067), .S(
        P1_IR_REG_21__SCAN_IN), .Z(n9069) );
  NAND2_X1 U11609 ( .A1(n9071), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9072) );
  MUX2_X1 U11610 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9072), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n9073) );
  INV_X1 U11611 ( .A(n10075), .ZN(n10076) );
  AOI21_X1 U11612 ( .B1(n14253), .B2(n10075), .A(n14023), .ZN(n9074) );
  NAND2_X1 U11613 ( .A1(n12066), .A2(n9074), .ZN(n10726) );
  NAND2_X1 U11614 ( .A1(n9167), .A2(n11150), .ZN(n9365) );
  INV_X1 U11615 ( .A(n9365), .ZN(n9075) );
  NAND2_X1 U11616 ( .A1(n9075), .A2(n14023), .ZN(n14541) );
  NAND2_X1 U11617 ( .A1(n11071), .A2(n11120), .ZN(n9077) );
  NAND2_X1 U11618 ( .A1(n11078), .A2(n11990), .ZN(n9078) );
  NAND2_X1 U11619 ( .A1(n9079), .A2(n9078), .ZN(n10756) );
  NAND2_X1 U11620 ( .A1(n10756), .A2(n9375), .ZN(n9082) );
  INV_X1 U11621 ( .A(n13769), .ZN(n9080) );
  NAND2_X1 U11622 ( .A1(n14537), .A2(n9080), .ZN(n9081) );
  INV_X1 U11623 ( .A(n13768), .ZN(n11542) );
  AND2_X1 U11624 ( .A1(n14475), .A2(n11542), .ZN(n9083) );
  OR2_X1 U11625 ( .A1(n14475), .A2(n11542), .ZN(n9084) );
  INV_X1 U11626 ( .A(n13767), .ZN(n11050) );
  INV_X1 U11627 ( .A(n11059), .ZN(n11047) );
  INV_X1 U11628 ( .A(n13765), .ZN(n11049) );
  NAND2_X1 U11629 ( .A1(n14426), .A2(n13764), .ZN(n9085) );
  NAND2_X1 U11630 ( .A1(n13652), .A2(n13763), .ZN(n9087) );
  INV_X1 U11631 ( .A(n11474), .ZN(n9088) );
  NAND2_X1 U11632 ( .A1(n11530), .A2(n9384), .ZN(n9089) );
  INV_X1 U11633 ( .A(n13758), .ZN(n9091) );
  OR2_X1 U11634 ( .A1(n13670), .A2(n9091), .ZN(n9090) );
  NAND2_X1 U11635 ( .A1(n13670), .A2(n9091), .ZN(n9092) );
  OR2_X1 U11636 ( .A1(n14083), .A2(n13625), .ZN(n9260) );
  NAND2_X1 U11637 ( .A1(n14083), .A2(n13625), .ZN(n9261) );
  INV_X1 U11638 ( .A(n14088), .ZN(n9387) );
  OR2_X1 U11639 ( .A1(n14222), .A2(n9093), .ZN(n9094) );
  INV_X1 U11640 ( .A(n14155), .ZN(n14038) );
  NAND2_X1 U11641 ( .A1(n14038), .A2(n13754), .ZN(n9095) );
  INV_X1 U11642 ( .A(n13634), .ZN(n13753) );
  OR2_X1 U11643 ( .A1(n14218), .A2(n13753), .ZN(n9096) );
  INV_X1 U11644 ( .A(n13752), .ZN(n12103) );
  INV_X1 U11645 ( .A(n13978), .ZN(n9097) );
  NAND2_X1 U11646 ( .A1(n14212), .A2(n12113), .ZN(n9098) );
  NAND2_X1 U11647 ( .A1(n9099), .A2(n9098), .ZN(n13959) );
  INV_X1 U11648 ( .A(n13750), .ZN(n12126) );
  NAND2_X1 U11649 ( .A1(n14208), .A2(n12126), .ZN(n9100) );
  INV_X1 U11650 ( .A(n13749), .ZN(n9101) );
  NAND2_X1 U11651 ( .A1(n14203), .A2(n9102), .ZN(n9103) );
  XNOR2_X1 U11652 ( .A(n13904), .B(n9393), .ZN(n9117) );
  NAND2_X1 U11653 ( .A1(n14253), .A2(n14023), .ZN(n9105) );
  NAND2_X1 U11654 ( .A1(n9343), .A2(n10111), .ZN(n9104) );
  NAND2_X1 U11655 ( .A1(n8767), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9113) );
  INV_X1 U11656 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n9106) );
  OR2_X1 U11657 ( .A1(n9338), .A2(n9106), .ZN(n9112) );
  OR2_X1 U11658 ( .A1(n9107), .A2(n13911), .ZN(n9111) );
  INV_X1 U11659 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n9108) );
  OR2_X1 U11660 ( .A1(n9109), .A2(n9108), .ZN(n9110) );
  AND4_X1 U11661 ( .A1(n9113), .A2(n9112), .A3(n9111), .A4(n9110), .ZN(n9170)
         );
  NAND2_X1 U11662 ( .A1(n14253), .A2(n9343), .ZN(n10099) );
  INV_X1 U11663 ( .A(n6483), .ZN(n9115) );
  NOR2_X2 U11664 ( .A1(n10099), .A2(n9115), .ZN(n13717) );
  NAND2_X1 U11665 ( .A1(n10233), .A2(n9115), .ZN(n13624) );
  AOI22_X1 U11666 ( .A1(n13747), .A2(n13717), .B1(n13913), .B2(n13748), .ZN(
        n12291) );
  INV_X1 U11667 ( .A(n12291), .ZN(n9116) );
  INV_X1 U11668 ( .A(n14117), .ZN(n13952) );
  AND2_X1 U11669 ( .A1(n10087), .A2(n11188), .ZN(n10748) );
  NAND2_X1 U11670 ( .A1(n10748), .A2(n14503), .ZN(n10747) );
  NOR2_X2 U11671 ( .A1(n11197), .A2(n14475), .ZN(n11196) );
  INV_X1 U11672 ( .A(n11552), .ZN(n11565) );
  NAND2_X1 U11673 ( .A1(n11196), .A2(n11565), .ZN(n11052) );
  NOR2_X2 U11674 ( .A1(n11241), .A2(n11883), .ZN(n11298) );
  NAND2_X1 U11675 ( .A1(n11415), .A2(n13652), .ZN(n11472) );
  OR2_X2 U11676 ( .A1(n11472), .A2(n12024), .ZN(n11519) );
  NOR2_X2 U11677 ( .A1(n11519), .A2(n14419), .ZN(n11520) );
  NAND2_X1 U11678 ( .A1(n14218), .A2(n14032), .ZN(n14015) );
  OR2_X2 U11679 ( .A1(n14203), .A2(n13949), .ZN(n13938) );
  NAND2_X1 U11680 ( .A1(n13926), .A2(n13938), .ZN(n9119) );
  NAND2_X2 U11681 ( .A1(n9118), .A2(n11150), .ZN(n14119) );
  NAND2_X1 U11682 ( .A1(n9119), .A2(n14493), .ZN(n9120) );
  OR2_X1 U11683 ( .A1(n9120), .A2(n13908), .ZN(n13928) );
  OAI21_X1 U11684 ( .B1(n13922), .B2(n14521), .A(n9121), .ZN(n9163) );
  INV_X1 U11685 ( .A(n9122), .ZN(n9123) );
  NAND2_X1 U11686 ( .A1(n9124), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9125) );
  MUX2_X1 U11687 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9125), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n9126) );
  NAND2_X1 U11688 ( .A1(n9126), .A2(n9133), .ZN(n11980) );
  NAND2_X1 U11689 ( .A1(n11980), .A2(P1_B_REG_SCAN_IN), .ZN(n9132) );
  MUX2_X1 U11690 ( .A(P1_B_REG_SCAN_IN), .B(n9132), .S(n11941), .Z(n9137) );
  INV_X1 U11691 ( .A(n14252), .ZN(n9136) );
  NAND2_X1 U11692 ( .A1(n9137), .A2(n9136), .ZN(n10182) );
  NOR4_X1 U11693 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n9146) );
  NOR4_X1 U11694 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n9145) );
  NOR4_X1 U11695 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n9141) );
  NOR4_X1 U11696 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n9140) );
  NOR4_X1 U11697 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9139) );
  NOR4_X1 U11698 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n9138) );
  NAND4_X1 U11699 ( .A1(n9141), .A2(n9140), .A3(n9139), .A4(n9138), .ZN(n9142)
         );
  NOR4_X1 U11700 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n9143), .A4(n9142), .ZN(n9144) );
  AND3_X1 U11701 ( .A1(n9146), .A2(n9145), .A3(n9144), .ZN(n9147) );
  NOR2_X1 U11702 ( .A1(n10182), .A2(n9147), .ZN(n10095) );
  NAND2_X1 U11703 ( .A1(n14493), .A2(n14023), .ZN(n10107) );
  NOR2_X1 U11704 ( .A1(n10095), .A2(n10112), .ZN(n9148) );
  NAND2_X1 U11705 ( .A1(n14252), .A2(n11980), .ZN(n10183) );
  OAI21_X1 U11706 ( .B1(n10182), .B2(P1_D_REG_1__SCAN_IN), .A(n10183), .ZN(
        n10096) );
  AND2_X1 U11707 ( .A1(n9148), .A2(n10096), .ZN(n9162) );
  NAND2_X1 U11708 ( .A1(n11941), .A2(n14252), .ZN(n10186) );
  NOR2_X1 U11709 ( .A1(n14252), .A2(n11980), .ZN(n9150) );
  INV_X1 U11710 ( .A(n11941), .ZN(n9149) );
  NAND2_X1 U11711 ( .A1(n9150), .A2(n9149), .ZN(n10077) );
  NAND2_X1 U11712 ( .A1(n9151), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9152) );
  MUX2_X1 U11713 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9152), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n9154) );
  NAND2_X1 U11714 ( .A1(n11860), .A2(n11150), .ZN(n9157) );
  NAND2_X1 U11715 ( .A1(n10233), .A2(n9157), .ZN(n10108) );
  AND2_X1 U11716 ( .A1(n10097), .A2(n10651), .ZN(n10700) );
  INV_X1 U11717 ( .A(n9155), .ZN(n9160) );
  INV_X1 U11718 ( .A(n13926), .ZN(n9156) );
  INV_X1 U11719 ( .A(n14528), .ZN(n14538) );
  NAND2_X1 U11720 ( .A1(n14549), .A2(n14538), .ZN(n14232) );
  NAND2_X1 U11721 ( .A1(n13926), .A2(n9158), .ZN(n9159) );
  NAND2_X1 U11722 ( .A1(n9160), .A2(n9159), .ZN(P1_U3524) );
  NOR2_X1 U11723 ( .A1(n10097), .A2(n10116), .ZN(n9161) );
  NAND2_X1 U11724 ( .A1(n14560), .A2(n14538), .ZN(n14186) );
  OAI21_X1 U11725 ( .B1(n14186), .B2(n9156), .A(n9164), .ZN(P1_U3556) );
  NAND2_X1 U11726 ( .A1(n13581), .A2(n8774), .ZN(n9166) );
  INV_X1 U11727 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14242) );
  OR2_X1 U11728 ( .A1(n8759), .A2(n14242), .ZN(n9165) );
  MUX2_X1 U11729 ( .A(n11150), .B(n9343), .S(n9341), .Z(n9169) );
  INV_X2 U11730 ( .A(n9176), .ZN(n9345) );
  MUX2_X1 U11731 ( .A(n9170), .B(n14106), .S(n9345), .Z(n9320) );
  INV_X1 U11732 ( .A(n9320), .ZN(n9321) );
  NOR2_X1 U11733 ( .A1(n13762), .A2(n9176), .ZN(n9172) );
  NOR2_X1 U11734 ( .A1(n12024), .A2(n9345), .ZN(n9171) );
  MUX2_X1 U11735 ( .A(n13762), .B(n12024), .S(n9345), .Z(n9233) );
  NAND2_X1 U11736 ( .A1(n13776), .A2(n11188), .ZN(n9370) );
  NAND2_X1 U11737 ( .A1(n9370), .A2(n10075), .ZN(n9173) );
  NAND2_X1 U11738 ( .A1(n9173), .A2(n9371), .ZN(n9175) );
  NAND2_X1 U11739 ( .A1(n9175), .A2(n9174), .ZN(n9184) );
  MUX2_X1 U11740 ( .A(n13774), .B(n10085), .S(n9169), .Z(n9178) );
  NAND2_X1 U11741 ( .A1(n13774), .A2(n10085), .ZN(n9177) );
  NAND2_X1 U11742 ( .A1(n9178), .A2(n9177), .ZN(n9188) );
  INV_X1 U11743 ( .A(n9185), .ZN(n9180) );
  NAND2_X1 U11744 ( .A1(n13773), .A2(n7066), .ZN(n9179) );
  AOI21_X1 U11745 ( .B1(n9180), .B2(n9176), .A(n9179), .ZN(n9181) );
  OAI211_X1 U11746 ( .C1(n9184), .C2(n9176), .A(n9188), .B(n9181), .ZN(n9192)
         );
  NAND3_X1 U11747 ( .A1(n9169), .A2(n14503), .A3(n13773), .ZN(n9182) );
  INV_X1 U11748 ( .A(n9183), .ZN(n9191) );
  NAND3_X1 U11749 ( .A1(n9184), .A2(n14503), .A3(n9169), .ZN(n9187) );
  NAND3_X1 U11750 ( .A1(n9185), .A2(n9176), .A3(n10693), .ZN(n9186) );
  NAND2_X1 U11751 ( .A1(n9187), .A2(n9186), .ZN(n9189) );
  NAND2_X1 U11752 ( .A1(n9189), .A2(n9188), .ZN(n9190) );
  NAND4_X1 U11753 ( .A1(n9192), .A2(n9191), .A3(n10706), .A4(n9190), .ZN(n9197) );
  NAND2_X1 U11754 ( .A1(n9176), .A2(n13772), .ZN(n9195) );
  NAND2_X1 U11755 ( .A1(n9193), .A2(n9169), .ZN(n9194) );
  MUX2_X1 U11756 ( .A(n9195), .B(n9194), .S(n10714), .Z(n9196) );
  MUX2_X1 U11757 ( .A(n14520), .B(n11071), .S(n9169), .Z(n9199) );
  MUX2_X1 U11758 ( .A(n11120), .B(n13771), .S(n9176), .Z(n9198) );
  MUX2_X1 U11759 ( .A(n11990), .B(n13770), .S(n9176), .Z(n9202) );
  MUX2_X1 U11760 ( .A(n13770), .B(n11990), .S(n9176), .Z(n9200) );
  NAND2_X1 U11761 ( .A1(n9201), .A2(n9200), .ZN(n9204) );
  NAND2_X1 U11762 ( .A1(n6549), .A2(n7336), .ZN(n9203) );
  NAND2_X1 U11763 ( .A1(n9204), .A2(n9203), .ZN(n9207) );
  MUX2_X1 U11764 ( .A(n13769), .B(n14537), .S(n9176), .Z(n9208) );
  NAND2_X1 U11765 ( .A1(n9207), .A2(n9208), .ZN(n9206) );
  MUX2_X1 U11766 ( .A(n13769), .B(n14537), .S(n9345), .Z(n9205) );
  NAND2_X1 U11767 ( .A1(n9206), .A2(n9205), .ZN(n9212) );
  INV_X1 U11768 ( .A(n9207), .ZN(n9210) );
  INV_X1 U11769 ( .A(n9208), .ZN(n9209) );
  NAND2_X1 U11770 ( .A1(n9210), .A2(n9209), .ZN(n9211) );
  MUX2_X1 U11771 ( .A(n13768), .B(n14475), .S(n9345), .Z(n9214) );
  MUX2_X1 U11772 ( .A(n13768), .B(n14475), .S(n9176), .Z(n9213) );
  MUX2_X1 U11773 ( .A(n13767), .B(n11552), .S(n9176), .Z(n9218) );
  NAND2_X1 U11774 ( .A1(n9217), .A2(n9218), .ZN(n9216) );
  MUX2_X1 U11775 ( .A(n13767), .B(n11552), .S(n9345), .Z(n9215) );
  NAND2_X1 U11776 ( .A1(n9216), .A2(n9215), .ZN(n9222) );
  INV_X1 U11777 ( .A(n9217), .ZN(n9220) );
  INV_X1 U11778 ( .A(n9218), .ZN(n9219) );
  NAND2_X1 U11779 ( .A1(n9220), .A2(n9219), .ZN(n9221) );
  MUX2_X1 U11780 ( .A(n13766), .B(n11851), .S(n9345), .Z(n9224) );
  MUX2_X1 U11781 ( .A(n13766), .B(n11851), .S(n9176), .Z(n9223) );
  MUX2_X1 U11782 ( .A(n13765), .B(n11883), .S(n9176), .Z(n9226) );
  INV_X1 U11783 ( .A(n11883), .ZN(n11346) );
  MUX2_X1 U11784 ( .A(n11049), .B(n11346), .S(n9345), .Z(n9225) );
  NOR2_X1 U11785 ( .A1(n9227), .A2(n9226), .ZN(n9228) );
  MUX2_X1 U11786 ( .A(n12007), .B(n14426), .S(n9176), .Z(n9231) );
  MUX2_X1 U11787 ( .A(n13764), .B(n14413), .S(n9345), .Z(n9230) );
  OAI22_X1 U11788 ( .A1(n9229), .A2(n9228), .B1(n9231), .B2(n9230), .ZN(n9236)
         );
  MUX2_X1 U11789 ( .A(n12016), .B(n13652), .S(n9176), .Z(n9238) );
  MUX2_X1 U11790 ( .A(n13763), .B(n11418), .S(n9345), .Z(n9237) );
  AOI22_X1 U11791 ( .A1(n9238), .A2(n9237), .B1(n9231), .B2(n9230), .ZN(n9235)
         );
  INV_X1 U11792 ( .A(n12024), .ZN(n13702) );
  NAND2_X1 U11793 ( .A1(n9345), .A2(n13762), .ZN(n9232) );
  OAI211_X1 U11794 ( .C1(n13702), .C2(n9345), .A(n9233), .B(n9232), .ZN(n9234)
         );
  AND2_X1 U11795 ( .A1(n9384), .A2(n9234), .ZN(n9244) );
  NAND3_X1 U11796 ( .A1(n9236), .A2(n9235), .A3(n9244), .ZN(n9249) );
  INV_X1 U11797 ( .A(n9237), .ZN(n9240) );
  INV_X1 U11798 ( .A(n9238), .ZN(n9239) );
  AND2_X1 U11799 ( .A1(n9240), .A2(n9239), .ZN(n9243) );
  NAND2_X1 U11800 ( .A1(n9252), .A2(n9241), .ZN(n9242) );
  AOI22_X1 U11801 ( .A1(n9244), .A2(n9243), .B1(n9176), .B2(n9242), .ZN(n9248)
         );
  NAND2_X1 U11802 ( .A1(n9251), .A2(n9245), .ZN(n9246) );
  NAND2_X1 U11803 ( .A1(n9246), .A2(n9345), .ZN(n9247) );
  NAND3_X1 U11804 ( .A1(n9250), .A2(n9249), .A3(n7364), .ZN(n9254) );
  MUX2_X1 U11805 ( .A(n9252), .B(n9251), .S(n9176), .Z(n9253) );
  NAND2_X1 U11806 ( .A1(n9254), .A2(n9253), .ZN(n9257) );
  MUX2_X1 U11807 ( .A(n12048), .B(n12049), .S(n9176), .Z(n9256) );
  MUX2_X1 U11808 ( .A(n13759), .B(n14189), .S(n9345), .Z(n9255) );
  MUX2_X1 U11809 ( .A(n13758), .B(n13670), .S(n9176), .Z(n9258) );
  MUX2_X1 U11810 ( .A(n9261), .B(n9260), .S(n9345), .Z(n9262) );
  NAND2_X1 U11811 ( .A1(n9263), .A2(n9262), .ZN(n9264) );
  NAND2_X1 U11812 ( .A1(n9264), .A2(n14064), .ZN(n9268) );
  MUX2_X1 U11813 ( .A(n9266), .B(n9265), .S(n9345), .Z(n9267) );
  MUX2_X1 U11814 ( .A(n14222), .B(n13755), .S(n9345), .Z(n9270) );
  MUX2_X1 U11815 ( .A(n13755), .B(n14222), .S(n9345), .Z(n9269) );
  MUX2_X1 U11816 ( .A(n13754), .B(n14155), .S(n9345), .Z(n9274) );
  NAND2_X1 U11817 ( .A1(n9273), .A2(n9274), .ZN(n9272) );
  MUX2_X1 U11818 ( .A(n14155), .B(n13754), .S(n9345), .Z(n9271) );
  NAND2_X1 U11819 ( .A1(n9272), .A2(n9271), .ZN(n9278) );
  INV_X1 U11820 ( .A(n9273), .ZN(n9276) );
  INV_X1 U11821 ( .A(n9274), .ZN(n9275) );
  NAND2_X1 U11822 ( .A1(n9276), .A2(n9275), .ZN(n9277) );
  MUX2_X1 U11823 ( .A(n14218), .B(n13634), .S(n9345), .Z(n9279) );
  INV_X1 U11824 ( .A(n9279), .ZN(n9281) );
  MUX2_X1 U11825 ( .A(n13634), .B(n14218), .S(n9345), .Z(n9280) );
  MUX2_X1 U11826 ( .A(n13752), .B(n14142), .S(n9345), .Z(n9285) );
  NAND2_X1 U11827 ( .A1(n9284), .A2(n9285), .ZN(n9283) );
  MUX2_X1 U11828 ( .A(n14142), .B(n13752), .S(n9345), .Z(n9282) );
  NAND2_X1 U11829 ( .A1(n9283), .A2(n9282), .ZN(n9289) );
  INV_X1 U11830 ( .A(n9284), .ZN(n9287) );
  NAND2_X1 U11831 ( .A1(n9287), .A2(n9286), .ZN(n9288) );
  MUX2_X1 U11832 ( .A(n13751), .B(n14212), .S(n9345), .Z(n9290) );
  NAND2_X1 U11833 ( .A1(n9291), .A2(n9290), .ZN(n9297) );
  INV_X1 U11834 ( .A(n9292), .ZN(n9295) );
  INV_X1 U11835 ( .A(n9293), .ZN(n9294) );
  NAND2_X1 U11836 ( .A1(n9295), .A2(n9294), .ZN(n9296) );
  NAND2_X1 U11837 ( .A1(n9297), .A2(n9296), .ZN(n9300) );
  MUX2_X1 U11838 ( .A(n14208), .B(n13750), .S(n9176), .Z(n9301) );
  NAND2_X1 U11839 ( .A1(n9300), .A2(n9301), .ZN(n9299) );
  MUX2_X1 U11840 ( .A(n14208), .B(n13750), .S(n9345), .Z(n9298) );
  NAND2_X1 U11841 ( .A1(n9299), .A2(n9298), .ZN(n9305) );
  INV_X1 U11842 ( .A(n9300), .ZN(n9303) );
  NAND2_X1 U11843 ( .A1(n9303), .A2(n9302), .ZN(n9304) );
  MUX2_X1 U11844 ( .A(n14117), .B(n13749), .S(n9345), .Z(n9307) );
  MUX2_X1 U11845 ( .A(n13749), .B(n14117), .S(n9345), .Z(n9306) );
  MUX2_X1 U11846 ( .A(n14203), .B(n13748), .S(n9345), .Z(n9308) );
  NAND2_X1 U11847 ( .A1(n9309), .A2(n9308), .ZN(n9315) );
  INV_X1 U11848 ( .A(n9310), .ZN(n9313) );
  INV_X1 U11849 ( .A(n9311), .ZN(n9312) );
  NAND2_X1 U11850 ( .A1(n9313), .A2(n9312), .ZN(n9314) );
  NAND2_X1 U11851 ( .A1(n9315), .A2(n9314), .ZN(n9317) );
  MUX2_X1 U11852 ( .A(n13914), .B(n13926), .S(n9176), .Z(n9318) );
  MUX2_X1 U11853 ( .A(n13914), .B(n13926), .S(n9345), .Z(n9316) );
  MUX2_X1 U11854 ( .A(n9368), .B(n13747), .S(n9345), .Z(n9319) );
  INV_X1 U11855 ( .A(n9348), .ZN(n9351) );
  INV_X1 U11856 ( .A(n9324), .ZN(n9325) );
  MUX2_X1 U11857 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n6706), .Z(n9326) );
  NAND2_X1 U11858 ( .A1(n9326), .A2(SI_30_), .ZN(n9352) );
  OAI21_X1 U11859 ( .B1(SI_30_), .B2(n9326), .A(n9352), .ZN(n9327) );
  NAND2_X1 U11860 ( .A1(n9328), .A2(n9327), .ZN(n9329) );
  NAND2_X1 U11861 ( .A1(n12257), .A2(n8774), .ZN(n9331) );
  INV_X1 U11862 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12301) );
  OR2_X1 U11863 ( .A1(n8759), .A2(n12301), .ZN(n9330) );
  INV_X1 U11864 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n14096) );
  NAND2_X1 U11865 ( .A1(n8767), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n9333) );
  NAND2_X1 U11866 ( .A1(n8742), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n9332) );
  OAI211_X1 U11867 ( .C1(n9338), .C2(n14096), .A(n9333), .B(n9332), .ZN(n13890) );
  INV_X1 U11868 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9337) );
  NAND2_X1 U11869 ( .A1(n9334), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9336) );
  NAND2_X1 U11870 ( .A1(n8742), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n9335) );
  OAI211_X1 U11871 ( .C1(n9338), .C2(n9337), .A(n9336), .B(n9335), .ZN(n13910)
         );
  OAI21_X1 U11872 ( .B1(n13890), .B2(n11150), .A(n13910), .ZN(n9339) );
  INV_X1 U11873 ( .A(n9339), .ZN(n9340) );
  MUX2_X1 U11874 ( .A(n14198), .B(n9340), .S(n9345), .Z(n9347) );
  INV_X1 U11875 ( .A(n9347), .ZN(n9350) );
  INV_X1 U11876 ( .A(n9341), .ZN(n9342) );
  NAND2_X1 U11877 ( .A1(n9176), .A2(n13890), .ZN(n9362) );
  OAI21_X1 U11878 ( .B1(n9343), .B2(n9342), .A(n9362), .ZN(n9344) );
  AOI22_X1 U11879 ( .A1(n14198), .A2(n9345), .B1(n13910), .B2(n9344), .ZN(
        n9346) );
  AOI21_X1 U11880 ( .B1(n9348), .B2(n9347), .A(n9346), .ZN(n9349) );
  AOI21_X2 U11881 ( .B1(n9351), .B2(n9350), .A(n9349), .ZN(n9416) );
  INV_X1 U11882 ( .A(n9416), .ZN(n9413) );
  MUX2_X1 U11883 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n6706), .Z(n9354) );
  XNOR2_X1 U11884 ( .A(n9354), .B(SI_31_), .ZN(n9355) );
  NAND2_X1 U11885 ( .A1(n12219), .A2(n8774), .ZN(n9358) );
  INV_X1 U11886 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9356) );
  OR2_X1 U11887 ( .A1(n8759), .A2(n9356), .ZN(n9357) );
  NAND2_X1 U11888 ( .A1(n9361), .A2(n9360), .ZN(n9363) );
  NAND2_X1 U11889 ( .A1(n10099), .A2(n9365), .ZN(n9366) );
  NAND2_X1 U11890 ( .A1(n10075), .A2(n14023), .ZN(n10702) );
  NAND2_X1 U11891 ( .A1(n9366), .A2(n10702), .ZN(n9414) );
  NAND2_X1 U11892 ( .A1(n11251), .A2(n10111), .ZN(n9408) );
  NAND2_X1 U11893 ( .A1(n9414), .A2(n9408), .ZN(n9401) );
  INV_X1 U11894 ( .A(n9401), .ZN(n9367) );
  XNOR2_X1 U11895 ( .A(n13886), .B(n9359), .ZN(n9415) );
  INV_X1 U11896 ( .A(n9415), .ZN(n9402) );
  XOR2_X1 U11897 ( .A(n13910), .B(n14198), .Z(n9398) );
  NAND2_X1 U11898 ( .A1(n9369), .A2(n6547), .ZN(n11922) );
  AND2_X1 U11899 ( .A1(n9371), .A2(n9370), .ZN(n11193) );
  NAND2_X1 U11900 ( .A1(n9373), .A2(n9372), .ZN(n10806) );
  NAND4_X1 U11901 ( .A1(n10752), .A2(n11193), .A3(n10734), .A4(n10806), .ZN(
        n9374) );
  NOR3_X1 U11902 ( .A1(n9374), .A2(n11981), .A3(n7350), .ZN(n9377) );
  NAND4_X1 U11903 ( .A1(n10953), .A2(n9377), .A3(n9376), .A4(n9375), .ZN(n9378) );
  NOR2_X1 U11904 ( .A1(n11059), .A2(n9378), .ZN(n9381) );
  NAND4_X1 U11905 ( .A1(n11411), .A2(n9381), .A3(n9380), .A4(n9379), .ZN(n9382) );
  NOR2_X1 U11906 ( .A1(n11474), .A2(n9382), .ZN(n9383) );
  NAND4_X1 U11907 ( .A1(n9384), .A2(n11922), .A3(n9383), .A4(n11856), .ZN(
        n9385) );
  OR4_X1 U11908 ( .A1(n9387), .A2(n14061), .A3(n9386), .A4(n9385), .ZN(n9388)
         );
  NOR2_X1 U11909 ( .A1(n14043), .A2(n9388), .ZN(n9389) );
  NAND4_X1 U11910 ( .A1(n13997), .A2(n9390), .A3(n9389), .A4(n14030), .ZN(
        n9391) );
  NOR2_X1 U11911 ( .A1(n13979), .A2(n9391), .ZN(n9392) );
  NAND2_X1 U11912 ( .A1(n9396), .A2(n9395), .ZN(n9397) );
  NOR2_X1 U11913 ( .A1(n9402), .A2(n9401), .ZN(n9403) );
  INV_X1 U11914 ( .A(n9414), .ZN(n9405) );
  OAI21_X1 U11915 ( .B1(n9409), .B2(n9408), .A(n7393), .ZN(n9410) );
  INV_X1 U11916 ( .A(n9410), .ZN(n9411) );
  OAI21_X2 U11917 ( .B1(n9413), .B2(n9412), .A(n9411), .ZN(n9420) );
  NOR3_X1 U11918 ( .A1(n9416), .A2(n9415), .A3(n9414), .ZN(n9419) );
  INV_X1 U11919 ( .A(n10232), .ZN(n9417) );
  NAND2_X1 U11920 ( .A1(n9417), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11753) );
  INV_X1 U11921 ( .A(n11753), .ZN(n9418) );
  OAI21_X1 U11922 ( .B1(n9420), .B2(n9419), .A(n9418), .ZN(n9423) );
  NOR3_X1 U11923 ( .A1(n10116), .A2(n14248), .A3(n13624), .ZN(n9422) );
  OAI21_X1 U11924 ( .B1(n11753), .B2(n14253), .A(P1_B_REG_SCAN_IN), .ZN(n9421)
         );
  NAND2_X1 U11925 ( .A1(n9423), .A2(n7365), .ZN(P1_U3242) );
  NAND2_X1 U11926 ( .A1(n7997), .A2(n12682), .ZN(n9424) );
  NAND2_X1 U11927 ( .A1(n9425), .A2(n9424), .ZN(n9434) );
  AND2_X1 U11928 ( .A1(n12297), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9426) );
  NAND2_X1 U11929 ( .A1(n9428), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9429) );
  XNOR2_X1 U11930 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n12298) );
  NAND2_X1 U11931 ( .A1(n13132), .A2(n12322), .ZN(n9433) );
  OR2_X1 U11932 ( .A1(n9431), .A2(n13135), .ZN(n9432) );
  NAND2_X1 U11933 ( .A1(n9445), .A2(n11029), .ZN(n12487) );
  XNOR2_X1 U11934 ( .A(n9434), .B(n12485), .ZN(n9442) );
  NAND2_X1 U11935 ( .A1(n9435), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n9439) );
  NAND2_X1 U11936 ( .A1(n9436), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9438) );
  NAND2_X1 U11937 ( .A1(n12315), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n9437) );
  AND2_X1 U11938 ( .A1(n10342), .A2(P3_B_REG_SCAN_IN), .ZN(n9440) );
  OAI22_X1 U11939 ( .A1(n12494), .A2(n12833), .B1(n12560), .B2(n14341), .ZN(
        n9441) );
  INV_X1 U11940 ( .A(n12469), .ZN(n9443) );
  NAND2_X1 U11941 ( .A1(n9449), .A2(n15120), .ZN(n9448) );
  INV_X1 U11942 ( .A(n9445), .ZN(n12549) );
  INV_X1 U11943 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n9446) );
  NAND2_X1 U11944 ( .A1(n9450), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n9451) );
  INV_X1 U11945 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9456) );
  NAND2_X1 U11946 ( .A1(n9453), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9455) );
  NAND2_X1 U11947 ( .A1(n8576), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9454) );
  OAI211_X1 U11948 ( .C1(n9457), .C2(n9456), .A(n9455), .B(n9454), .ZN(n13325)
         );
  NAND2_X1 U11949 ( .A1(n9475), .A2(n10447), .ZN(n9496) );
  MUX2_X1 U11950 ( .A(n13341), .B(n13146), .S(n9567), .Z(n9620) );
  MUX2_X1 U11951 ( .A(n12214), .B(n9458), .S(n9472), .Z(n9466) );
  MUX2_X1 U11952 ( .A(n13281), .B(n13482), .S(n9496), .Z(n9465) );
  NAND2_X1 U11953 ( .A1(n9466), .A2(n9465), .ZN(n9626) );
  MUX2_X1 U11954 ( .A(n13282), .B(n13487), .S(n9567), .Z(n9619) );
  INV_X1 U11955 ( .A(n13325), .ZN(n9636) );
  NOR2_X1 U11956 ( .A1(n9636), .A2(n9567), .ZN(n9462) );
  MUX2_X1 U11957 ( .A(n9636), .B(n9462), .S(n9634), .Z(n9470) );
  OAI211_X1 U11958 ( .C1(n9667), .C2(n9669), .A(n10472), .B(n9666), .ZN(n9461)
         );
  OAI21_X1 U11959 ( .B1(n9462), .B2(n9461), .A(n13280), .ZN(n9463) );
  OAI21_X1 U11960 ( .B1(n13479), .B2(n9496), .A(n9463), .ZN(n9630) );
  INV_X1 U11961 ( .A(n13280), .ZN(n9464) );
  MUX2_X1 U11962 ( .A(n9464), .B(n13479), .S(n9635), .Z(n9631) );
  INV_X1 U11963 ( .A(n9465), .ZN(n9468) );
  INV_X1 U11964 ( .A(n9466), .ZN(n9467) );
  AOI22_X1 U11965 ( .A1(n9630), .A2(n9631), .B1(n9468), .B2(n9467), .ZN(n9469)
         );
  NOR2_X1 U11966 ( .A1(n9470), .A2(n9469), .ZN(n9471) );
  NOR2_X1 U11967 ( .A1(n7392), .A2(n9471), .ZN(n9629) );
  MUX2_X1 U11968 ( .A(n13287), .B(n13514), .S(n9635), .Z(n9597) );
  MUX2_X1 U11969 ( .A(n13526), .B(n13289), .S(n9635), .Z(n9586) );
  OAI21_X1 U11970 ( .B1(n13308), .B2(n9635), .A(n11180), .ZN(n9473) );
  INV_X1 U11971 ( .A(n9473), .ZN(n9482) );
  AOI21_X1 U11972 ( .B1(n13308), .B2(n9635), .A(n11180), .ZN(n9481) );
  NAND2_X1 U11973 ( .A1(n13310), .A2(n14721), .ZN(n10487) );
  NAND3_X1 U11974 ( .A1(n9476), .A2(n9474), .A3(n9475), .ZN(n9480) );
  INV_X1 U11975 ( .A(n9476), .ZN(n9478) );
  NAND4_X1 U11976 ( .A1(n9478), .A2(n9643), .A3(n9477), .A4(n9635), .ZN(n9479)
         );
  MUX2_X1 U11977 ( .A(n10866), .B(n14759), .S(n9635), .Z(n9484) );
  MUX2_X1 U11978 ( .A(n10981), .B(n6995), .S(n9635), .Z(n9483) );
  OAI21_X1 U11979 ( .B1(n9485), .B2(n9484), .A(n9483), .ZN(n9487) );
  NAND2_X1 U11980 ( .A1(n9485), .A2(n9484), .ZN(n9486) );
  NAND2_X1 U11981 ( .A1(n9487), .A2(n9486), .ZN(n9490) );
  MUX2_X1 U11982 ( .A(n13307), .B(n14766), .S(n9472), .Z(n9491) );
  NAND2_X1 U11983 ( .A1(n9490), .A2(n9491), .ZN(n9489) );
  MUX2_X1 U11984 ( .A(n13307), .B(n14766), .S(n9635), .Z(n9488) );
  NAND2_X1 U11985 ( .A1(n9489), .A2(n9488), .ZN(n9495) );
  INV_X1 U11986 ( .A(n9490), .ZN(n9493) );
  INV_X1 U11987 ( .A(n9491), .ZN(n9492) );
  MUX2_X1 U11988 ( .A(n13306), .B(n11008), .S(n9635), .Z(n9498) );
  MUX2_X1 U11989 ( .A(n13306), .B(n11008), .S(n9567), .Z(n9497) );
  INV_X1 U11990 ( .A(n9498), .ZN(n9499) );
  MUX2_X1 U11991 ( .A(n11129), .B(n13305), .S(n9635), .Z(n9503) );
  NAND2_X1 U11992 ( .A1(n9502), .A2(n9503), .ZN(n9501) );
  MUX2_X1 U11993 ( .A(n13305), .B(n11129), .S(n9635), .Z(n9500) );
  NAND2_X1 U11994 ( .A1(n9501), .A2(n9500), .ZN(n9507) );
  INV_X1 U11995 ( .A(n9502), .ZN(n9505) );
  INV_X1 U11996 ( .A(n9503), .ZN(n9504) );
  MUX2_X1 U11997 ( .A(n13304), .B(n10911), .S(n9635), .Z(n9509) );
  MUX2_X1 U11998 ( .A(n13304), .B(n10911), .S(n9567), .Z(n9508) );
  INV_X1 U11999 ( .A(n9509), .ZN(n9510) );
  MUX2_X1 U12000 ( .A(n13303), .B(n14789), .S(n9567), .Z(n9514) );
  NAND2_X1 U12001 ( .A1(n9513), .A2(n9514), .ZN(n9512) );
  MUX2_X1 U12002 ( .A(n13303), .B(n14789), .S(n9496), .Z(n9511) );
  NAND2_X1 U12003 ( .A1(n9512), .A2(n9511), .ZN(n9518) );
  INV_X1 U12004 ( .A(n9513), .ZN(n9516) );
  INV_X1 U12005 ( .A(n9514), .ZN(n9515) );
  NAND2_X1 U12006 ( .A1(n9516), .A2(n9515), .ZN(n9517) );
  MUX2_X1 U12007 ( .A(n13302), .B(n11154), .S(n9635), .Z(n9520) );
  MUX2_X1 U12008 ( .A(n13302), .B(n11154), .S(n9567), .Z(n9519) );
  INV_X1 U12009 ( .A(n9520), .ZN(n9521) );
  MUX2_X1 U12010 ( .A(n13301), .B(n14710), .S(n9567), .Z(n9525) );
  OAI21_X1 U12011 ( .B1(n9526), .B2(n9525), .A(n9522), .ZN(n9528) );
  INV_X1 U12012 ( .A(n14710), .ZN(n14805) );
  MUX2_X1 U12013 ( .A(n9523), .B(n14805), .S(n9635), .Z(n9524) );
  AOI21_X1 U12014 ( .B1(n9526), .B2(n9525), .A(n9524), .ZN(n9527) );
  OR2_X1 U12015 ( .A1(n9528), .A2(n9527), .ZN(n9532) );
  AND2_X1 U12016 ( .A1(n13300), .A2(n9635), .ZN(n9530) );
  OAI21_X1 U12017 ( .B1(n13300), .B2(n9635), .A(n14813), .ZN(n9529) );
  OAI21_X1 U12018 ( .B1(n9530), .B2(n14813), .A(n9529), .ZN(n9531) );
  NAND2_X1 U12019 ( .A1(n9532), .A2(n9531), .ZN(n9534) );
  MUX2_X1 U12020 ( .A(n13299), .B(n11382), .S(n9472), .Z(n9535) );
  MUX2_X1 U12021 ( .A(n13299), .B(n11382), .S(n9635), .Z(n9533) );
  MUX2_X1 U12022 ( .A(n13298), .B(n11443), .S(n9635), .Z(n9538) );
  MUX2_X1 U12023 ( .A(n13298), .B(n11443), .S(n9567), .Z(n9536) );
  NAND2_X1 U12024 ( .A1(n9537), .A2(n9536), .ZN(n9541) );
  MUX2_X1 U12025 ( .A(n13297), .B(n11504), .S(n9567), .Z(n9543) );
  MUX2_X1 U12026 ( .A(n13297), .B(n11504), .S(n9635), .Z(n9542) );
  INV_X1 U12027 ( .A(n9543), .ZN(n9544) );
  MUX2_X1 U12028 ( .A(n13296), .B(n13557), .S(n9635), .Z(n9548) );
  NAND2_X1 U12029 ( .A1(n9547), .A2(n9548), .ZN(n9546) );
  MUX2_X1 U12030 ( .A(n13296), .B(n13557), .S(n9567), .Z(n9545) );
  NAND2_X1 U12031 ( .A1(n9546), .A2(n9545), .ZN(n9552) );
  INV_X1 U12032 ( .A(n9547), .ZN(n9550) );
  INV_X1 U12033 ( .A(n9548), .ZN(n9549) );
  NAND2_X1 U12034 ( .A1(n9550), .A2(n9549), .ZN(n9551) );
  MUX2_X1 U12035 ( .A(n13295), .B(n12161), .S(n9567), .Z(n9554) );
  MUX2_X1 U12036 ( .A(n13295), .B(n12161), .S(n9635), .Z(n9553) );
  INV_X1 U12037 ( .A(n9554), .ZN(n9555) );
  MUX2_X1 U12038 ( .A(n13294), .B(n13553), .S(n9635), .Z(n9559) );
  NAND2_X1 U12039 ( .A1(n9558), .A2(n9559), .ZN(n9557) );
  MUX2_X1 U12040 ( .A(n13294), .B(n13553), .S(n9567), .Z(n9556) );
  NAND2_X1 U12041 ( .A1(n9557), .A2(n9556), .ZN(n9563) );
  INV_X1 U12042 ( .A(n9558), .ZN(n9561) );
  INV_X1 U12043 ( .A(n9559), .ZN(n9560) );
  NAND2_X1 U12044 ( .A1(n9561), .A2(n9560), .ZN(n9562) );
  MUX2_X1 U12045 ( .A(n13293), .B(n13547), .S(n9472), .Z(n9565) );
  MUX2_X1 U12046 ( .A(n13293), .B(n13547), .S(n9635), .Z(n9564) );
  INV_X1 U12047 ( .A(n9565), .ZN(n9566) );
  MUX2_X1 U12048 ( .A(n13292), .B(n12171), .S(n9496), .Z(n9571) );
  NAND2_X1 U12049 ( .A1(n9570), .A2(n9571), .ZN(n9569) );
  MUX2_X1 U12050 ( .A(n13292), .B(n12171), .S(n9567), .Z(n9568) );
  NAND2_X1 U12051 ( .A1(n9569), .A2(n9568), .ZN(n9575) );
  INV_X1 U12052 ( .A(n9570), .ZN(n9573) );
  INV_X1 U12053 ( .A(n9571), .ZN(n9572) );
  NAND2_X1 U12054 ( .A1(n9573), .A2(n9572), .ZN(n9574) );
  MUX2_X1 U12055 ( .A(n13291), .B(n13537), .S(n9567), .Z(n9577) );
  MUX2_X1 U12056 ( .A(n13291), .B(n13537), .S(n9635), .Z(n9576) );
  INV_X1 U12057 ( .A(n9577), .ZN(n9578) );
  MUX2_X1 U12058 ( .A(n13531), .B(n13290), .S(n9472), .Z(n9582) );
  NAND2_X1 U12059 ( .A1(n9581), .A2(n9582), .ZN(n9580) );
  MUX2_X1 U12060 ( .A(n13531), .B(n13290), .S(n9496), .Z(n9579) );
  INV_X1 U12061 ( .A(n9581), .ZN(n9584) );
  INV_X1 U12062 ( .A(n9582), .ZN(n9583) );
  MUX2_X1 U12063 ( .A(n13289), .B(n13526), .S(n9635), .Z(n9585) );
  MUX2_X1 U12064 ( .A(n13288), .B(n13518), .S(n9635), .Z(n9590) );
  NAND2_X1 U12065 ( .A1(n9589), .A2(n9590), .ZN(n9588) );
  MUX2_X1 U12066 ( .A(n13518), .B(n13288), .S(n9635), .Z(n9587) );
  NAND2_X1 U12067 ( .A1(n9588), .A2(n9587), .ZN(n9594) );
  INV_X1 U12068 ( .A(n9590), .ZN(n9591) );
  NAND2_X1 U12069 ( .A1(n9594), .A2(n9593), .ZN(n9595) );
  MUX2_X1 U12070 ( .A(n13514), .B(n13287), .S(n9635), .Z(n9596) );
  MUX2_X1 U12071 ( .A(n13187), .B(n13396), .S(n9635), .Z(n9599) );
  MUX2_X1 U12072 ( .A(n13507), .B(n13286), .S(n9496), .Z(n9598) );
  MUX2_X1 U12073 ( .A(n13497), .B(n13284), .S(n9635), .Z(n9611) );
  INV_X1 U12074 ( .A(n9611), .ZN(n9600) );
  MUX2_X1 U12075 ( .A(n13284), .B(n13497), .S(n9635), .Z(n9605) );
  NAND2_X1 U12076 ( .A1(n9600), .A2(n9605), .ZN(n9606) );
  MUX2_X1 U12077 ( .A(n13502), .B(n13285), .S(n9496), .Z(n9607) );
  INV_X1 U12078 ( .A(n9607), .ZN(n9602) );
  MUX2_X1 U12079 ( .A(n13255), .B(n13382), .S(n9635), .Z(n9608) );
  INV_X1 U12080 ( .A(n9608), .ZN(n9601) );
  NAND2_X1 U12081 ( .A1(n9602), .A2(n9601), .ZN(n9603) );
  NAND3_X1 U12082 ( .A1(n9604), .A2(n9606), .A3(n9603), .ZN(n9618) );
  INV_X1 U12083 ( .A(n9605), .ZN(n9612) );
  INV_X1 U12084 ( .A(n9606), .ZN(n9609) );
  NOR3_X1 U12085 ( .A1(n9609), .A2(n9602), .A3(n9601), .ZN(n9610) );
  AOI21_X1 U12086 ( .B1(n9612), .B2(n9611), .A(n9610), .ZN(n9616) );
  MUX2_X1 U12087 ( .A(n13492), .B(n13283), .S(n9635), .Z(n9613) );
  INV_X1 U12088 ( .A(n9613), .ZN(n9622) );
  MUX2_X1 U12089 ( .A(n13492), .B(n13283), .S(n9567), .Z(n9621) );
  NAND2_X1 U12090 ( .A1(n9613), .A2(n9614), .ZN(n9615) );
  INV_X1 U12091 ( .A(n9619), .ZN(n9624) );
  INV_X1 U12092 ( .A(n9620), .ZN(n9623) );
  AOI22_X1 U12093 ( .A1(n9624), .A2(n9623), .B1(n9622), .B2(n9621), .ZN(n9625)
         );
  NAND2_X1 U12094 ( .A1(n9627), .A2(n7391), .ZN(n9628) );
  NAND2_X1 U12095 ( .A1(n9629), .A2(n9628), .ZN(n9642) );
  INV_X1 U12096 ( .A(n9630), .ZN(n9633) );
  INV_X1 U12097 ( .A(n9631), .ZN(n9632) );
  NAND2_X1 U12098 ( .A1(n9633), .A2(n9632), .ZN(n9641) );
  INV_X1 U12099 ( .A(n9634), .ZN(n9637) );
  NOR3_X1 U12100 ( .A1(n9637), .A2(n9636), .A3(n9635), .ZN(n9639) );
  NOR3_X1 U12101 ( .A1(n9634), .A2(n9472), .A3(n13325), .ZN(n9638) );
  INV_X1 U12102 ( .A(n9673), .ZN(n9663) );
  XOR2_X1 U12103 ( .A(n8486), .B(n13537), .Z(n13459) );
  AND2_X1 U12104 ( .A1(n9643), .A2(n10487), .ZN(n14749) );
  NAND4_X1 U12105 ( .A1(n10971), .A2(n9474), .A3(n14749), .A4(n9667), .ZN(
        n9644) );
  NOR4_X1 U12106 ( .A1(n11132), .A2(n9644), .A3(n10998), .A4(n8647), .ZN(n9645) );
  XNOR2_X1 U12107 ( .A(n14789), .B(n13303), .ZN(n10878) );
  NAND4_X1 U12108 ( .A1(n9645), .A2(n11157), .A3(n10878), .A4(n10826), .ZN(
        n9646) );
  NOR4_X1 U12109 ( .A1(n11308), .A2(n11332), .A3(n14708), .A4(n9646), .ZN(
        n9647) );
  XNOR2_X1 U12110 ( .A(n11504), .B(n13297), .ZN(n11454) );
  XNOR2_X1 U12111 ( .A(n11443), .B(n13298), .ZN(n11438) );
  NAND4_X1 U12112 ( .A1(n11892), .A2(n9647), .A3(n11454), .A4(n11438), .ZN(
        n9649) );
  XNOR2_X1 U12113 ( .A(n13557), .B(n9648), .ZN(n11763) );
  NOR3_X1 U12114 ( .A1(n11968), .A2(n9649), .A3(n11763), .ZN(n9651) );
  NAND4_X1 U12115 ( .A1(n13459), .A2(n9651), .A3(n9650), .A4(n11951), .ZN(
        n9652) );
  NOR4_X1 U12116 ( .A1(n9653), .A2(n13436), .A3(n13443), .A4(n9652), .ZN(n9654) );
  XNOR2_X1 U12117 ( .A(n13514), .B(n13287), .ZN(n13405) );
  NAND4_X1 U12118 ( .A1(n13370), .A2(n9654), .A3(n13398), .A4(n13405), .ZN(
        n9655) );
  XOR2_X1 U12119 ( .A(n13280), .B(n13479), .Z(n9656) );
  NAND4_X1 U12120 ( .A1(n9659), .A2(n9658), .A3(n9657), .A4(n9656), .ZN(n9660)
         );
  INV_X1 U12121 ( .A(n10195), .ZN(n10058) );
  NAND2_X1 U12122 ( .A1(n10058), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11749) );
  OR2_X1 U12123 ( .A1(n11749), .A2(n9666), .ZN(n9661) );
  OAI21_X1 U12124 ( .B1(n9663), .B2(n9667), .A(n9662), .ZN(n9676) );
  INV_X1 U12125 ( .A(n10472), .ZN(n10478) );
  NAND4_X1 U12126 ( .A1(n14741), .A2(n10208), .A3(n10478), .A4(n13171), .ZN(
        n9664) );
  OAI211_X1 U12127 ( .C1(n11533), .C2(n11749), .A(n9664), .B(P2_B_REG_SCAN_IN), 
        .ZN(n9675) );
  MUX2_X1 U12128 ( .A(n11533), .B(n9666), .S(n9667), .Z(n9665) );
  INV_X1 U12129 ( .A(n9666), .ZN(n11267) );
  AOI21_X1 U12130 ( .B1(n9667), .B2(n11267), .A(n8683), .ZN(n9668) );
  AOI21_X1 U12131 ( .B1(n10447), .B2(n9669), .A(n9668), .ZN(n9670) );
  NAND2_X1 U12132 ( .A1(n9673), .A2(n9670), .ZN(n9672) );
  INV_X1 U12133 ( .A(n11749), .ZN(n9671) );
  OAI211_X1 U12134 ( .C1(n9673), .C2(n7368), .A(n9672), .B(n9671), .ZN(n9674)
         );
  NAND3_X1 U12135 ( .A1(n9676), .A2(n9675), .A3(n9674), .ZN(P2_U3328) );
  INV_X1 U12136 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14315) );
  INV_X1 U12137 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9717) );
  XOR2_X1 U12138 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n9717), .Z(n9770) );
  INV_X1 U12139 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n9714) );
  XOR2_X1 U12140 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .Z(n9721) );
  INV_X1 U12141 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9711) );
  INV_X1 U12142 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9708) );
  INV_X1 U12143 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9703) );
  INV_X1 U12144 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9701) );
  INV_X1 U12145 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9695) );
  NAND2_X1 U12146 ( .A1(P3_ADDR_REG_0__SCAN_IN), .A2(n9734), .ZN(n9733) );
  AOI21_X2 U12147 ( .B1(n9681), .B2(n9680), .A(n9679), .ZN(n9682) );
  NOR2_X1 U12148 ( .A1(n9682), .A2(n9683), .ZN(n9685) );
  XNOR2_X1 U12149 ( .A(n9683), .B(n9682), .ZN(n9729) );
  NOR2_X1 U12150 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(n9729), .ZN(n9684) );
  NOR2_X1 U12151 ( .A1(n9686), .A2(n9687), .ZN(n9689) );
  NOR2_X1 U12152 ( .A1(n9690), .A2(n9691), .ZN(n9693) );
  XOR2_X1 U12153 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), .Z(
        n9744) );
  NOR2_X1 U12154 ( .A1(n9696), .A2(n9697), .ZN(n9699) );
  XNOR2_X1 U12155 ( .A(n9697), .B(n9696), .ZN(n9750) );
  XOR2_X1 U12156 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(P3_ADDR_REG_8__SCAN_IN), .Z(
        n9752) );
  XOR2_X1 U12157 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(P3_ADDR_REG_9__SCAN_IN), .Z(
        n9726) );
  NOR2_X1 U12158 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n9704), .ZN(n9706) );
  XNOR2_X1 U12159 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(n9704), .ZN(n9725) );
  INV_X1 U12160 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n14999) );
  INV_X1 U12161 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n9707) );
  XNOR2_X1 U12162 ( .A(P1_ADDR_REG_11__SCAN_IN), .B(n9707), .ZN(n9761) );
  INV_X1 U12163 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n9709) );
  XNOR2_X1 U12164 ( .A(P1_ADDR_REG_12__SCAN_IN), .B(n9709), .ZN(n9763) );
  INV_X1 U12165 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n9722) );
  AND2_X1 U12166 ( .A1(n9722), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n9712) );
  INV_X1 U12167 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n12763) );
  NAND2_X1 U12168 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n12763), .ZN(n9715) );
  INV_X1 U12169 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14474) );
  NAND2_X1 U12170 ( .A1(n9770), .A2(n9769), .ZN(n9716) );
  XNOR2_X1 U12171 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n9772), .ZN(n9773) );
  XOR2_X1 U12172 ( .A(n14315), .B(n9773), .Z(n14286) );
  XOR2_X1 U12173 ( .A(n14474), .B(P3_ADDR_REG_15__SCAN_IN), .Z(n9719) );
  XOR2_X1 U12174 ( .A(n9719), .B(n9718), .Z(n14451) );
  XNOR2_X1 U12175 ( .A(n9721), .B(n9720), .ZN(n14447) );
  XOR2_X1 U12176 ( .A(P1_ADDR_REG_13__SCAN_IN), .B(n9722), .Z(n9724) );
  XNOR2_X1 U12177 ( .A(n9724), .B(n9723), .ZN(n14443) );
  XOR2_X1 U12178 ( .A(n14999), .B(n9725), .Z(n14283) );
  XOR2_X1 U12179 ( .A(n9727), .B(n9726), .Z(n9757) );
  INV_X1 U12180 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n14589) );
  NOR2_X1 U12181 ( .A1(n9738), .A2(n14589), .ZN(n9739) );
  XOR2_X1 U12182 ( .A(n9729), .B(P1_ADDR_REG_3__SCAN_IN), .Z(n15144) );
  XOR2_X1 U12183 ( .A(n9731), .B(n9730), .Z(n14264) );
  INV_X1 U12184 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10200) );
  NOR2_X1 U12185 ( .A1(n9735), .A2(n10200), .ZN(n9736) );
  OAI21_X1 U12186 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n9734), .A(n9733), .ZN(
        n15138) );
  NAND2_X1 U12187 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15138), .ZN(n15148) );
  NOR2_X1 U12188 ( .A1(n15148), .A2(n15147), .ZN(n15146) );
  NAND2_X1 U12189 ( .A1(n14264), .A2(n14263), .ZN(n14262) );
  NAND2_X1 U12190 ( .A1(n15144), .A2(n15143), .ZN(n9737) );
  AOI21_X1 U12191 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n9737), .A(n15142), .ZN(
        n15134) );
  NOR2_X1 U12192 ( .A1(n15134), .A2(n15133), .ZN(n15132) );
  NAND2_X1 U12193 ( .A1(n9741), .A2(n9742), .ZN(n9743) );
  INV_X1 U12194 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15136) );
  NOR2_X1 U12195 ( .A1(n9746), .A2(n6876), .ZN(n9747) );
  XOR2_X1 U12196 ( .A(n9745), .B(n9744), .Z(n14275) );
  INV_X1 U12197 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n9748) );
  NAND2_X1 U12198 ( .A1(n9749), .A2(n9748), .ZN(n9751) );
  XOR2_X1 U12199 ( .A(n9750), .B(P1_ADDR_REG_7__SCAN_IN), .Z(n15140) );
  NAND2_X1 U12200 ( .A1(n15141), .A2(n15140), .ZN(n15139) );
  XOR2_X1 U12201 ( .A(n9753), .B(n9752), .Z(n9755) );
  INV_X1 U12202 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14277) );
  NAND2_X1 U12203 ( .A1(n9755), .A2(n9754), .ZN(n9756) );
  NOR2_X1 U12204 ( .A1(n9757), .A2(n9758), .ZN(n9759) );
  INV_X1 U12205 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14618) );
  NAND2_X1 U12206 ( .A1(n14283), .A2(n14282), .ZN(n9760) );
  XOR2_X1 U12207 ( .A(n9762), .B(n9761), .Z(n14436) );
  XOR2_X1 U12208 ( .A(n9764), .B(n9763), .Z(n9766) );
  INV_X1 U12209 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n14648) );
  NAND2_X1 U12210 ( .A1(n9766), .A2(n9765), .ZN(n9767) );
  NAND2_X1 U12211 ( .A1(n14443), .A2(n14442), .ZN(n14441) );
  NAND2_X1 U12212 ( .A1(n14447), .A2(n14446), .ZN(n14445) );
  NAND2_X1 U12213 ( .A1(n14451), .A2(n14450), .ZN(n9768) );
  XNOR2_X1 U12214 ( .A(n9770), .B(n9769), .ZN(n14454) );
  NAND2_X1 U12215 ( .A1(n14455), .A2(n14454), .ZN(n9771) );
  NAND2_X1 U12216 ( .A1(n14286), .A2(n14287), .ZN(n14285) );
  INV_X1 U12217 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n9779) );
  XOR2_X1 U12218 ( .A(n9779), .B(P1_ADDR_REG_18__SCAN_IN), .Z(n9776) );
  NOR2_X1 U12219 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n9772), .ZN(n9775) );
  NOR2_X1 U12220 ( .A1(n14315), .A2(n9773), .ZN(n9774) );
  NOR2_X1 U12221 ( .A1(n9775), .A2(n9774), .ZN(n9778) );
  XNOR2_X1 U12222 ( .A(n9776), .B(n9778), .ZN(n14259) );
  AND2_X1 U12223 ( .A1(n9779), .A2(P1_ADDR_REG_18__SCAN_IN), .ZN(n9777) );
  OAI22_X1 U12224 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n9779), .B1(n9778), .B2(
        n9777), .ZN(n9780) );
  INV_X1 U12225 ( .A(n9780), .ZN(n9954) );
  OAI22_X1 U12226 ( .A1(P3_REG3_REG_2__SCAN_IN), .A2(keyinput_f59), .B1(SI_14_), .B2(keyinput_f18), .ZN(n9781) );
  AOI221_X1 U12227 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(keyinput_f59), .C1(
        keyinput_f18), .C2(SI_14_), .A(n9781), .ZN(n9798) );
  OAI22_X1 U12228 ( .A1(P3_REG3_REG_28__SCAN_IN), .A2(keyinput_f42), .B1(
        keyinput_f52), .B2(P3_REG3_REG_4__SCAN_IN), .ZN(n9782) );
  AOI221_X1 U12229 ( .B1(P3_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .C1(
        P3_REG3_REG_4__SCAN_IN), .C2(keyinput_f52), .A(n9782), .ZN(n9797) );
  AOI22_X1 U12230 ( .A1(SI_7_), .A2(keyinput_f25), .B1(P3_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .ZN(n9783) );
  OAI221_X1 U12231 ( .B1(SI_7_), .B2(keyinput_f25), .C1(
        P3_REG3_REG_18__SCAN_IN), .C2(keyinput_f60), .A(n9783), .ZN(n9790) );
  AOI22_X1 U12232 ( .A1(SI_21_), .A2(keyinput_f11), .B1(
        P3_REG3_REG_21__SCAN_IN), .B2(keyinput_f45), .ZN(n9784) );
  OAI221_X1 U12233 ( .B1(SI_21_), .B2(keyinput_f11), .C1(
        P3_REG3_REG_21__SCAN_IN), .C2(keyinput_f45), .A(n9784), .ZN(n9789) );
  AOI22_X1 U12234 ( .A1(SI_30_), .A2(keyinput_f2), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(keyinput_f40), .ZN(n9785) );
  OAI221_X1 U12235 ( .B1(SI_30_), .B2(keyinput_f2), .C1(P3_REG3_REG_3__SCAN_IN), .C2(keyinput_f40), .A(n9785), .ZN(n9788) );
  AOI22_X1 U12236 ( .A1(SI_2_), .A2(keyinput_f30), .B1(P3_REG3_REG_14__SCAN_IN), .B2(keyinput_f37), .ZN(n9786) );
  OAI221_X1 U12237 ( .B1(SI_2_), .B2(keyinput_f30), .C1(
        P3_REG3_REG_14__SCAN_IN), .C2(keyinput_f37), .A(n9786), .ZN(n9787) );
  NOR4_X1 U12238 ( .A1(n9790), .A2(n9789), .A3(n9788), .A4(n9787), .ZN(n9793)
         );
  OAI22_X1 U12239 ( .A1(SI_11_), .A2(keyinput_f21), .B1(SI_31_), .B2(
        keyinput_f1), .ZN(n9791) );
  AOI221_X1 U12240 ( .B1(SI_11_), .B2(keyinput_f21), .C1(keyinput_f1), .C2(
        SI_31_), .A(n9791), .ZN(n9792) );
  OAI211_X1 U12241 ( .C1(n9795), .C2(keyinput_f41), .A(n9793), .B(n9792), .ZN(
        n9794) );
  AOI21_X1 U12242 ( .B1(n9795), .B2(keyinput_f41), .A(n9794), .ZN(n9796) );
  NAND3_X1 U12243 ( .A1(n9798), .A2(n9797), .A3(n9796), .ZN(n9862) );
  INV_X1 U12244 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n10990) );
  INV_X1 U12245 ( .A(P3_WR_REG_SCAN_IN), .ZN(n9800) );
  AOI22_X1 U12246 ( .A1(n10990), .A2(keyinput_f61), .B1(keyinput_f0), .B2(
        n9800), .ZN(n9799) );
  OAI221_X1 U12247 ( .B1(n10990), .B2(keyinput_f61), .C1(n9800), .C2(
        keyinput_f0), .A(n9799), .ZN(n9808) );
  INV_X1 U12248 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n9922) );
  AOI22_X1 U12249 ( .A1(n9922), .A2(keyinput_f55), .B1(keyinput_f3), .B2(
        n13135), .ZN(n9801) );
  OAI221_X1 U12250 ( .B1(n9922), .B2(keyinput_f55), .C1(n13135), .C2(
        keyinput_f3), .A(n9801), .ZN(n9807) );
  XNOR2_X1 U12251 ( .A(SI_22_), .B(keyinput_f10), .ZN(n9805) );
  XNOR2_X1 U12252 ( .A(SI_5_), .B(keyinput_f27), .ZN(n9804) );
  XNOR2_X1 U12253 ( .A(SI_3_), .B(keyinput_f29), .ZN(n9803) );
  XNOR2_X1 U12254 ( .A(SI_4_), .B(keyinput_f28), .ZN(n9802) );
  NAND4_X1 U12255 ( .A1(n9805), .A2(n9804), .A3(n9803), .A4(n9802), .ZN(n9806)
         );
  NOR3_X1 U12256 ( .A1(n9808), .A2(n9807), .A3(n9806), .ZN(n9839) );
  INV_X1 U12257 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n9810) );
  AOI22_X1 U12258 ( .A1(n9810), .A2(keyinput_f48), .B1(keyinput_f6), .B2(
        n11770), .ZN(n9809) );
  OAI221_X1 U12259 ( .B1(n9810), .B2(keyinput_f48), .C1(n11770), .C2(
        keyinput_f6), .A(n9809), .ZN(n9817) );
  INV_X1 U12260 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n11496) );
  INV_X1 U12261 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n11143) );
  AOI22_X1 U12262 ( .A1(n11496), .A2(keyinput_f39), .B1(keyinput_f35), .B2(
        n11143), .ZN(n9811) );
  OAI221_X1 U12263 ( .B1(n11496), .B2(keyinput_f39), .C1(n11143), .C2(
        keyinput_f35), .A(n9811), .ZN(n9816) );
  INV_X1 U12264 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10666) );
  INV_X1 U12265 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n9925) );
  AOI22_X1 U12266 ( .A1(n10666), .A2(keyinput_f54), .B1(n9925), .B2(
        keyinput_f47), .ZN(n9812) );
  OAI221_X1 U12267 ( .B1(n10666), .B2(keyinput_f54), .C1(n9925), .C2(
        keyinput_f47), .A(n9812), .ZN(n9815) );
  AOI22_X1 U12268 ( .A1(n13141), .A2(keyinput_f4), .B1(keyinput_f17), .B2(
        n10320), .ZN(n9813) );
  OAI221_X1 U12269 ( .B1(n13141), .B2(keyinput_f4), .C1(n10320), .C2(
        keyinput_f17), .A(n9813), .ZN(n9814) );
  NOR4_X1 U12270 ( .A1(n9817), .A2(n9816), .A3(n9815), .A4(n9814), .ZN(n9838)
         );
  INV_X1 U12271 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11683) );
  AOI22_X1 U12272 ( .A1(n7750), .A2(keyinput_f63), .B1(keyinput_f58), .B2(
        n11683), .ZN(n9818) );
  OAI221_X1 U12273 ( .B1(n7750), .B2(keyinput_f63), .C1(n11683), .C2(
        keyinput_f58), .A(n9818), .ZN(n9826) );
  INV_X1 U12274 ( .A(P3_RD_REG_SCAN_IN), .ZN(n10122) );
  AOI22_X1 U12275 ( .A1(n10440), .A2(keyinput_f15), .B1(keyinput_f33), .B2(
        n10122), .ZN(n9819) );
  OAI221_X1 U12276 ( .B1(n10440), .B2(keyinput_f15), .C1(n10122), .C2(
        keyinput_f33), .A(n9819), .ZN(n9825) );
  INV_X1 U12277 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n9895) );
  AOI22_X1 U12278 ( .A1(n7719), .A2(keyinput_f56), .B1(n9895), .B2(
        keyinput_f57), .ZN(n9820) );
  OAI221_X1 U12279 ( .B1(n7719), .B2(keyinput_f56), .C1(n9895), .C2(
        keyinput_f57), .A(n9820), .ZN(n9824) );
  INV_X1 U12280 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10502) );
  INV_X1 U12281 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n9822) );
  AOI22_X1 U12282 ( .A1(n10502), .A2(keyinput_f44), .B1(n9822), .B2(
        keyinput_f50), .ZN(n9821) );
  OAI221_X1 U12283 ( .B1(n10502), .B2(keyinput_f44), .C1(n9822), .C2(
        keyinput_f50), .A(n9821), .ZN(n9823) );
  NOR4_X1 U12284 ( .A1(n9826), .A2(n9825), .A3(n9824), .A4(n9823), .ZN(n9837)
         );
  AOI22_X1 U12285 ( .A1(n11288), .A2(keyinput_f9), .B1(n7586), .B2(
        keyinput_f49), .ZN(n9827) );
  OAI221_X1 U12286 ( .B1(n11288), .B2(keyinput_f9), .C1(n7586), .C2(
        keyinput_f49), .A(n9827), .ZN(n9835) );
  AOI22_X1 U12287 ( .A1(n10219), .A2(keyinput_f19), .B1(n9829), .B2(
        keyinput_f36), .ZN(n9828) );
  OAI221_X1 U12288 ( .B1(n10219), .B2(keyinput_f19), .C1(n9829), .C2(
        keyinput_f36), .A(n9828), .ZN(n9834) );
  INV_X1 U12289 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n12630) );
  AOI22_X1 U12290 ( .A1(n10689), .A2(keyinput_f13), .B1(n12630), .B2(
        keyinput_f51), .ZN(n9830) );
  OAI221_X1 U12291 ( .B1(n10689), .B2(keyinput_f13), .C1(n12630), .C2(
        keyinput_f51), .A(n9830), .ZN(n9833) );
  AOI22_X1 U12292 ( .A1(n11273), .A2(keyinput_f43), .B1(keyinput_f14), .B2(
        n10546), .ZN(n9831) );
  OAI221_X1 U12293 ( .B1(n11273), .B2(keyinput_f43), .C1(n10546), .C2(
        keyinput_f14), .A(n9831), .ZN(n9832) );
  NOR4_X1 U12294 ( .A1(n9835), .A2(n9834), .A3(n9833), .A4(n9832), .ZN(n9836)
         );
  NAND4_X1 U12295 ( .A1(n9839), .A2(n9838), .A3(n9837), .A4(n9836), .ZN(n9861)
         );
  OAI22_X1 U12296 ( .A1(P3_REG3_REG_9__SCAN_IN), .A2(keyinput_f53), .B1(
        keyinput_f12), .B2(SI_20_), .ZN(n9840) );
  AOI221_X1 U12297 ( .B1(P3_REG3_REG_9__SCAN_IN), .B2(keyinput_f53), .C1(
        SI_20_), .C2(keyinput_f12), .A(n9840), .ZN(n9847) );
  OAI22_X1 U12298 ( .A1(P3_STATE_REG_SCAN_IN), .A2(keyinput_f34), .B1(SI_9_), 
        .B2(keyinput_f23), .ZN(n9841) );
  AOI221_X1 U12299 ( .B1(P3_STATE_REG_SCAN_IN), .B2(keyinput_f34), .C1(
        keyinput_f23), .C2(SI_9_), .A(n9841), .ZN(n9846) );
  OAI22_X1 U12300 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(keyinput_f46), .B1(
        keyinput_f5), .B2(SI_27_), .ZN(n9842) );
  AOI221_X1 U12301 ( .B1(P3_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .C1(
        SI_27_), .C2(keyinput_f5), .A(n9842), .ZN(n9845) );
  OAI22_X1 U12302 ( .A1(SI_6_), .A2(keyinput_f26), .B1(SI_0_), .B2(
        keyinput_f32), .ZN(n9843) );
  AOI221_X1 U12303 ( .B1(SI_6_), .B2(keyinput_f26), .C1(keyinput_f32), .C2(
        SI_0_), .A(n9843), .ZN(n9844) );
  NAND4_X1 U12304 ( .A1(n9847), .A2(n9846), .A3(n9845), .A4(n9844), .ZN(n9851)
         );
  XNOR2_X1 U12305 ( .A(SI_10_), .B(keyinput_f22), .ZN(n9849) );
  XNOR2_X1 U12306 ( .A(SI_1_), .B(keyinput_f31), .ZN(n9848) );
  NAND2_X1 U12307 ( .A1(n9849), .A2(n9848), .ZN(n9850) );
  NOR2_X1 U12308 ( .A1(n9851), .A2(n9850), .ZN(n9859) );
  OAI22_X1 U12309 ( .A1(P3_REG3_REG_23__SCAN_IN), .A2(keyinput_f38), .B1(
        keyinput_f20), .B2(SI_12_), .ZN(n9852) );
  AOI221_X1 U12310 ( .B1(P3_REG3_REG_23__SCAN_IN), .B2(keyinput_f38), .C1(
        SI_12_), .C2(keyinput_f20), .A(n9852), .ZN(n9858) );
  OAI22_X1 U12311 ( .A1(n9854), .A2(keyinput_f62), .B1(keyinput_f8), .B2(
        SI_24_), .ZN(n9853) );
  AOI221_X1 U12312 ( .B1(n9854), .B2(keyinput_f62), .C1(SI_24_), .C2(
        keyinput_f8), .A(n9853), .ZN(n9857) );
  OAI22_X1 U12313 ( .A1(SI_16_), .A2(keyinput_f16), .B1(keyinput_f7), .B2(
        SI_25_), .ZN(n9855) );
  AOI221_X1 U12314 ( .B1(SI_16_), .B2(keyinput_f16), .C1(SI_25_), .C2(
        keyinput_f7), .A(n9855), .ZN(n9856) );
  NAND4_X1 U12315 ( .A1(n9859), .A2(n9858), .A3(n9857), .A4(n9856), .ZN(n9860)
         );
  NOR3_X1 U12316 ( .A1(n9862), .A2(n9861), .A3(n9860), .ZN(n9864) );
  INV_X1 U12317 ( .A(keyinput_g24), .ZN(n9863) );
  OAI211_X1 U12318 ( .C1(n9864), .C2(keyinput_f24), .A(n9863), .B(n10124), 
        .ZN(n9949) );
  INV_X1 U12319 ( .A(keyinput_f24), .ZN(n9865) );
  OAI211_X1 U12320 ( .C1(n9865), .C2(n9864), .A(SI_8_), .B(keyinput_g24), .ZN(
        n9948) );
  AOI22_X1 U12321 ( .A1(P3_WR_REG_SCAN_IN), .A2(keyinput_g0), .B1(SI_23_), 
        .B2(keyinput_g9), .ZN(n9866) );
  OAI221_X1 U12322 ( .B1(P3_WR_REG_SCAN_IN), .B2(keyinput_g0), .C1(SI_23_), 
        .C2(keyinput_g9), .A(n9866), .ZN(n9873) );
  AOI22_X1 U12323 ( .A1(SI_19_), .A2(keyinput_g13), .B1(
        P3_REG3_REG_28__SCAN_IN), .B2(keyinput_g42), .ZN(n9867) );
  OAI221_X1 U12324 ( .B1(SI_19_), .B2(keyinput_g13), .C1(
        P3_REG3_REG_28__SCAN_IN), .C2(keyinput_g42), .A(n9867), .ZN(n9872) );
  AOI22_X1 U12325 ( .A1(SI_24_), .A2(keyinput_g8), .B1(n10985), .B2(
        keyinput_g11), .ZN(n9868) );
  OAI221_X1 U12326 ( .B1(SI_24_), .B2(keyinput_g8), .C1(n10985), .C2(
        keyinput_g11), .A(n9868), .ZN(n9871) );
  AOI22_X1 U12327 ( .A1(SI_29_), .A2(keyinput_g3), .B1(P3_REG3_REG_14__SCAN_IN), .B2(keyinput_g37), .ZN(n9869) );
  OAI221_X1 U12328 ( .B1(SI_29_), .B2(keyinput_g3), .C1(
        P3_REG3_REG_14__SCAN_IN), .C2(keyinput_g37), .A(n9869), .ZN(n9870) );
  NOR4_X1 U12329 ( .A1(n9873), .A2(n9872), .A3(n9871), .A4(n9870), .ZN(n9905)
         );
  AOI22_X1 U12330 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(keyinput_g48), .B1(
        P3_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .ZN(n9874) );
  OAI221_X1 U12331 ( .B1(P3_REG3_REG_16__SCAN_IN), .B2(keyinput_g48), .C1(
        P3_REG3_REG_18__SCAN_IN), .C2(keyinput_g60), .A(n9874), .ZN(n9881) );
  AOI22_X1 U12332 ( .A1(SI_30_), .A2(keyinput_g2), .B1(SI_2_), .B2(
        keyinput_g30), .ZN(n9875) );
  OAI221_X1 U12333 ( .B1(SI_30_), .B2(keyinput_g2), .C1(SI_2_), .C2(
        keyinput_g30), .A(n9875), .ZN(n9880) );
  AOI22_X1 U12334 ( .A1(SI_6_), .A2(keyinput_g26), .B1(SI_22_), .B2(
        keyinput_g10), .ZN(n9876) );
  OAI221_X1 U12335 ( .B1(SI_6_), .B2(keyinput_g26), .C1(SI_22_), .C2(
        keyinput_g10), .A(n9876), .ZN(n9879) );
  AOI22_X1 U12336 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(keyinput_g39), .B1(
        P3_REG3_REG_27__SCAN_IN), .B2(keyinput_g36), .ZN(n9877) );
  OAI221_X1 U12337 ( .B1(P3_REG3_REG_10__SCAN_IN), .B2(keyinput_g39), .C1(
        P3_REG3_REG_27__SCAN_IN), .C2(keyinput_g36), .A(n9877), .ZN(n9878) );
  NOR4_X1 U12338 ( .A1(n9881), .A2(n9880), .A3(n9879), .A4(n9878), .ZN(n9904)
         );
  INV_X1 U12339 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n10892) );
  AOI22_X1 U12340 ( .A1(n11683), .A2(keyinput_g58), .B1(keyinput_g52), .B2(
        n10892), .ZN(n9882) );
  OAI221_X1 U12341 ( .B1(n11683), .B2(keyinput_g58), .C1(n10892), .C2(
        keyinput_g52), .A(n9882), .ZN(n9891) );
  AOI22_X1 U12342 ( .A1(n7586), .A2(keyinput_g49), .B1(n10990), .B2(
        keyinput_g61), .ZN(n9883) );
  OAI221_X1 U12343 ( .B1(n7586), .B2(keyinput_g49), .C1(n10990), .C2(
        keyinput_g61), .A(n9883), .ZN(n9890) );
  INV_X1 U12344 ( .A(SI_9_), .ZN(n10161) );
  AOI22_X1 U12345 ( .A1(n10122), .A2(keyinput_g33), .B1(n10161), .B2(
        keyinput_g23), .ZN(n9884) );
  OAI221_X1 U12346 ( .B1(n10122), .B2(keyinput_g33), .C1(n10161), .C2(
        keyinput_g23), .A(n9884), .ZN(n9889) );
  INV_X1 U12347 ( .A(SI_31_), .ZN(n9885) );
  XOR2_X1 U12348 ( .A(n9885), .B(keyinput_g1), .Z(n9887) );
  XNOR2_X1 U12349 ( .A(SI_1_), .B(keyinput_g31), .ZN(n9886) );
  NAND2_X1 U12350 ( .A1(n9887), .A2(n9886), .ZN(n9888) );
  NOR4_X1 U12351 ( .A1(n9891), .A2(n9890), .A3(n9889), .A4(n9888), .ZN(n9903)
         );
  INV_X1 U12352 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n9893) );
  AOI22_X1 U12353 ( .A1(n9893), .A2(keyinput_g38), .B1(keyinput_g44), .B2(
        n10502), .ZN(n9892) );
  OAI221_X1 U12354 ( .B1(n9893), .B2(keyinput_g38), .C1(n10502), .C2(
        keyinput_g44), .A(n9892), .ZN(n9901) );
  AOI22_X1 U12355 ( .A1(n9895), .A2(keyinput_g57), .B1(keyinput_g35), .B2(
        n11143), .ZN(n9894) );
  OAI221_X1 U12356 ( .B1(n9895), .B2(keyinput_g57), .C1(n11143), .C2(
        keyinput_g35), .A(n9894), .ZN(n9900) );
  AOI22_X1 U12357 ( .A1(n7719), .A2(keyinput_g56), .B1(keyinput_g20), .B2(
        n10167), .ZN(n9896) );
  OAI221_X1 U12358 ( .B1(n7719), .B2(keyinput_g56), .C1(n10167), .C2(
        keyinput_g20), .A(n9896), .ZN(n9899) );
  AOI22_X1 U12359 ( .A1(n11691), .A2(keyinput_g7), .B1(n10666), .B2(
        keyinput_g54), .ZN(n9897) );
  OAI221_X1 U12360 ( .B1(n11691), .B2(keyinput_g7), .C1(n10666), .C2(
        keyinput_g54), .A(n9897), .ZN(n9898) );
  NOR4_X1 U12361 ( .A1(n9901), .A2(n9900), .A3(n9899), .A4(n9898), .ZN(n9902)
         );
  NAND4_X1 U12362 ( .A1(n9905), .A2(n9904), .A3(n9903), .A4(n9902), .ZN(n9946)
         );
  AOI22_X1 U12363 ( .A1(SI_26_), .A2(keyinput_g6), .B1(P3_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .ZN(n9906) );
  OAI221_X1 U12364 ( .B1(SI_26_), .B2(keyinput_g6), .C1(
        P3_REG3_REG_19__SCAN_IN), .C2(keyinput_g41), .A(n9906), .ZN(n9913) );
  AOI22_X1 U12365 ( .A1(SI_16_), .A2(keyinput_g16), .B1(P3_REG3_REG_9__SCAN_IN), .B2(keyinput_g53), .ZN(n9907) );
  OAI221_X1 U12366 ( .B1(SI_16_), .B2(keyinput_g16), .C1(
        P3_REG3_REG_9__SCAN_IN), .C2(keyinput_g53), .A(n9907), .ZN(n9912) );
  AOI22_X1 U12367 ( .A1(SI_17_), .A2(keyinput_g15), .B1(
        P3_REG3_REG_26__SCAN_IN), .B2(keyinput_g62), .ZN(n9908) );
  OAI221_X1 U12368 ( .B1(SI_17_), .B2(keyinput_g15), .C1(
        P3_REG3_REG_26__SCAN_IN), .C2(keyinput_g62), .A(n9908), .ZN(n9911) );
  AOI22_X1 U12369 ( .A1(SI_3_), .A2(keyinput_g29), .B1(P3_REG3_REG_12__SCAN_IN), .B2(keyinput_g46), .ZN(n9909) );
  OAI221_X1 U12370 ( .B1(SI_3_), .B2(keyinput_g29), .C1(
        P3_REG3_REG_12__SCAN_IN), .C2(keyinput_g46), .A(n9909), .ZN(n9910) );
  NOR4_X1 U12371 ( .A1(n9913), .A2(n9912), .A3(n9911), .A4(n9910), .ZN(n9944)
         );
  XNOR2_X1 U12372 ( .A(n11273), .B(keyinput_g43), .ZN(n9920) );
  AOI22_X1 U12373 ( .A1(P3_REG3_REG_2__SCAN_IN), .A2(keyinput_g59), .B1(
        P3_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .ZN(n9914) );
  OAI221_X1 U12374 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .C1(
        P3_REG3_REG_15__SCAN_IN), .C2(keyinput_g63), .A(n9914), .ZN(n9919) );
  AOI22_X1 U12375 ( .A1(SI_15_), .A2(keyinput_g17), .B1(SI_0_), .B2(
        keyinput_g32), .ZN(n9915) );
  OAI221_X1 U12376 ( .B1(SI_15_), .B2(keyinput_g17), .C1(SI_0_), .C2(
        keyinput_g32), .A(n9915), .ZN(n9918) );
  AOI22_X1 U12377 ( .A1(SI_14_), .A2(keyinput_g18), .B1(SI_7_), .B2(
        keyinput_g25), .ZN(n9916) );
  OAI221_X1 U12378 ( .B1(SI_14_), .B2(keyinput_g18), .C1(SI_7_), .C2(
        keyinput_g25), .A(n9916), .ZN(n9917) );
  NOR4_X1 U12379 ( .A1(n9920), .A2(n9919), .A3(n9918), .A4(n9917), .ZN(n9943)
         );
  AOI22_X1 U12380 ( .A1(n9923), .A2(keyinput_g45), .B1(keyinput_g55), .B2(
        n9922), .ZN(n9921) );
  OAI221_X1 U12381 ( .B1(n9923), .B2(keyinput_g45), .C1(n9922), .C2(
        keyinput_g55), .A(n9921), .ZN(n9931) );
  AOI22_X1 U12382 ( .A1(n10546), .A2(keyinput_g14), .B1(n9925), .B2(
        keyinput_g47), .ZN(n9924) );
  OAI221_X1 U12383 ( .B1(n10546), .B2(keyinput_g14), .C1(n9925), .C2(
        keyinput_g47), .A(n9924), .ZN(n9930) );
  AOI22_X1 U12384 ( .A1(n10920), .A2(keyinput_g40), .B1(keyinput_g19), .B2(
        n10219), .ZN(n9926) );
  OAI221_X1 U12385 ( .B1(n10920), .B2(keyinput_g40), .C1(n10219), .C2(
        keyinput_g19), .A(n9926), .ZN(n9929) );
  AOI22_X1 U12386 ( .A1(n10899), .A2(keyinput_g12), .B1(n13141), .B2(
        keyinput_g4), .ZN(n9927) );
  OAI221_X1 U12387 ( .B1(n10899), .B2(keyinput_g12), .C1(n13141), .C2(
        keyinput_g4), .A(n9927), .ZN(n9928) );
  NOR4_X1 U12388 ( .A1(n9931), .A2(n9930), .A3(n9929), .A4(n9928), .ZN(n9942)
         );
  AOI22_X1 U12389 ( .A1(P3_U3151), .A2(keyinput_g34), .B1(keyinput_g5), .B2(
        n11887), .ZN(n9932) );
  OAI221_X1 U12390 ( .B1(P3_U3151), .B2(keyinput_g34), .C1(n11887), .C2(
        keyinput_g5), .A(n9932), .ZN(n9940) );
  AOI22_X1 U12391 ( .A1(n10148), .A2(keyinput_g22), .B1(n10163), .B2(
        keyinput_g21), .ZN(n9933) );
  OAI221_X1 U12392 ( .B1(n10148), .B2(keyinput_g22), .C1(n10163), .C2(
        keyinput_g21), .A(n9933), .ZN(n9939) );
  XNOR2_X1 U12393 ( .A(SI_4_), .B(keyinput_g28), .ZN(n9937) );
  XNOR2_X1 U12394 ( .A(P3_REG3_REG_24__SCAN_IN), .B(keyinput_g51), .ZN(n9936)
         );
  XNOR2_X1 U12395 ( .A(P3_REG3_REG_17__SCAN_IN), .B(keyinput_g50), .ZN(n9935)
         );
  XNOR2_X1 U12396 ( .A(SI_5_), .B(keyinput_g27), .ZN(n9934) );
  NAND4_X1 U12397 ( .A1(n9937), .A2(n9936), .A3(n9935), .A4(n9934), .ZN(n9938)
         );
  NOR3_X1 U12398 ( .A1(n9940), .A2(n9939), .A3(n9938), .ZN(n9941) );
  NAND4_X1 U12399 ( .A1(n9944), .A2(n9943), .A3(n9942), .A4(n9941), .ZN(n9945)
         );
  NOR2_X1 U12400 ( .A1(n9946), .A2(n9945), .ZN(n9947) );
  AOI21_X1 U12401 ( .B1(n9949), .B2(n9948), .A(n9947), .ZN(n9952) );
  XNOR2_X1 U12402 ( .A(P3_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n9950) );
  XNOR2_X1 U12403 ( .A(n7466), .B(n9950), .ZN(n9951) );
  XNOR2_X1 U12404 ( .A(n9952), .B(n9951), .ZN(n9953) );
  NAND2_X1 U12405 ( .A1(n12337), .A2(n10898), .ZN(n9957) );
  XNOR2_X1 U12406 ( .A(n15003), .B(n10521), .ZN(n9979) );
  XNOR2_X1 U12407 ( .A(n11360), .B(n10521), .ZN(n9978) );
  XNOR2_X1 U12408 ( .A(n10795), .B(n10521), .ZN(n9967) );
  INV_X1 U12409 ( .A(n9967), .ZN(n9968) );
  INV_X1 U12410 ( .A(n10522), .ZN(n9964) );
  OAI21_X1 U12411 ( .B1(n15059), .B2(n10521), .A(n15042), .ZN(n9962) );
  OAI22_X1 U12412 ( .A1(n15059), .A2(n15042), .B1(n10519), .B2(n15072), .ZN(
        n9961) );
  AOI21_X1 U12413 ( .B1(n15072), .B2(n9962), .A(n9961), .ZN(n9963) );
  XNOR2_X1 U12414 ( .A(n10493), .B(n10521), .ZN(n9965) );
  XNOR2_X1 U12415 ( .A(n9965), .B(n10914), .ZN(n10492) );
  INV_X1 U12416 ( .A(n9965), .ZN(n9966) );
  OAI22_X1 U12417 ( .A1(n10491), .A2(n10492), .B1(n15064), .B2(n9966), .ZN(
        n10791) );
  XNOR2_X1 U12418 ( .A(n9967), .B(n15041), .ZN(n10792) );
  AOI21_X1 U12419 ( .B1(n12701), .B2(n9968), .A(n10790), .ZN(n10889) );
  INV_X2 U12420 ( .A(n10519), .ZN(n10028) );
  XNOR2_X1 U12421 ( .A(n15034), .B(n10028), .ZN(n9969) );
  XNOR2_X1 U12422 ( .A(n15017), .B(n9969), .ZN(n10890) );
  NAND2_X1 U12423 ( .A1(n10889), .A2(n10890), .ZN(n10888) );
  XNOR2_X1 U12424 ( .A(n15020), .B(n10521), .ZN(n9971) );
  XNOR2_X1 U12425 ( .A(n12699), .B(n9971), .ZN(n10944) );
  NAND2_X1 U12426 ( .A1(n15029), .A2(n9971), .ZN(n9972) );
  XNOR2_X1 U12427 ( .A(n11261), .B(n10521), .ZN(n9974) );
  XNOR2_X1 U12428 ( .A(n12698), .B(n9974), .ZN(n10988) );
  INV_X1 U12429 ( .A(n9974), .ZN(n9975) );
  NAND2_X1 U12430 ( .A1(n9975), .A2(n12698), .ZN(n9976) );
  XNOR2_X1 U12431 ( .A(n11226), .B(n10519), .ZN(n11141) );
  NAND2_X1 U12432 ( .A1(n11140), .A2(n9977), .ZN(n11272) );
  XNOR2_X1 U12433 ( .A(n12696), .B(n9978), .ZN(n11271) );
  XNOR2_X1 U12434 ( .A(n12387), .B(n9979), .ZN(n11387) );
  XNOR2_X1 U12435 ( .A(n11593), .B(n10521), .ZN(n9980) );
  XNOR2_X1 U12436 ( .A(n12694), .B(n9980), .ZN(n11494) );
  INV_X1 U12437 ( .A(n9980), .ZN(n9981) );
  NAND2_X1 U12438 ( .A1(n9981), .A2(n12694), .ZN(n9982) );
  NAND2_X1 U12439 ( .A1(n11493), .A2(n9982), .ZN(n9985) );
  XNOR2_X1 U12440 ( .A(n9983), .B(n10521), .ZN(n9984) );
  NAND2_X1 U12441 ( .A1(n9985), .A2(n9984), .ZN(n11779) );
  NAND2_X1 U12442 ( .A1(n11779), .A2(n11825), .ZN(n9986) );
  XNOR2_X1 U12443 ( .A(n14359), .B(n10521), .ZN(n11902) );
  NOR2_X1 U12444 ( .A1(n11902), .A2(n12692), .ZN(n9987) );
  XNOR2_X1 U12445 ( .A(n14353), .B(n10028), .ZN(n9988) );
  NOR2_X1 U12446 ( .A1(n9988), .A2(n12691), .ZN(n10061) );
  NAND2_X1 U12447 ( .A1(n9988), .A2(n12691), .ZN(n10062) );
  XNOR2_X1 U12448 ( .A(n9989), .B(n10521), .ZN(n9990) );
  XNOR2_X1 U12449 ( .A(n9990), .B(n12690), .ZN(n11932) );
  INV_X1 U12450 ( .A(n9990), .ZN(n9991) );
  NAND2_X1 U12451 ( .A1(n9991), .A2(n12690), .ZN(n9992) );
  NAND2_X1 U12452 ( .A1(n11931), .A2(n9992), .ZN(n12673) );
  XNOR2_X1 U12453 ( .A(n9993), .B(n10028), .ZN(n9994) );
  XOR2_X1 U12454 ( .A(n14329), .B(n9994), .Z(n12672) );
  INV_X1 U12455 ( .A(n9994), .ZN(n9995) );
  NAND2_X1 U12456 ( .A1(n9995), .A2(n7255), .ZN(n9996) );
  XNOR2_X1 U12457 ( .A(n12992), .B(n10521), .ZN(n9999) );
  XNOR2_X1 U12458 ( .A(n9999), .B(n13001), .ZN(n12607) );
  XNOR2_X1 U12459 ( .A(n9998), .B(n10028), .ZN(n10002) );
  XNOR2_X1 U12460 ( .A(n10002), .B(n12989), .ZN(n12615) );
  INV_X1 U12461 ( .A(n12615), .ZN(n10000) );
  NAND2_X1 U12462 ( .A1(n9999), .A2(n13001), .ZN(n12613) );
  AND2_X1 U12463 ( .A1(n10000), .A2(n12613), .ZN(n10001) );
  INV_X1 U12464 ( .A(n10002), .ZN(n10003) );
  INV_X1 U12465 ( .A(n12989), .ZN(n12688) );
  NAND2_X1 U12466 ( .A1(n10003), .A2(n12688), .ZN(n10004) );
  NAND2_X1 U12467 ( .A1(n12617), .A2(n10004), .ZN(n12654) );
  XNOR2_X1 U12468 ( .A(n10005), .B(n10521), .ZN(n10006) );
  XOR2_X1 U12469 ( .A(n12978), .B(n10006), .Z(n12653) );
  NAND2_X1 U12470 ( .A1(n12654), .A2(n12653), .ZN(n12652) );
  INV_X1 U12471 ( .A(n10006), .ZN(n10007) );
  INV_X1 U12472 ( .A(n12978), .ZN(n12952) );
  NAND2_X1 U12473 ( .A1(n10007), .A2(n12952), .ZN(n10008) );
  NAND2_X1 U12474 ( .A1(n12652), .A2(n10008), .ZN(n12576) );
  XNOR2_X1 U12475 ( .A(n13105), .B(n10028), .ZN(n12574) );
  INV_X1 U12476 ( .A(n12966), .ZN(n12687) );
  XNOR2_X1 U12477 ( .A(n12943), .B(n10028), .ZN(n10009) );
  XNOR2_X1 U12478 ( .A(n10009), .B(n12926), .ZN(n12635) );
  INV_X1 U12479 ( .A(n10009), .ZN(n10010) );
  NAND2_X1 U12480 ( .A1(n10010), .A2(n12926), .ZN(n10011) );
  XNOR2_X1 U12481 ( .A(n13033), .B(n10521), .ZN(n10012) );
  NAND2_X1 U12482 ( .A1(n10012), .A2(n12940), .ZN(n10014) );
  OAI21_X1 U12483 ( .B1(n10012), .B2(n12940), .A(n10014), .ZN(n12585) );
  INV_X1 U12484 ( .A(n12585), .ZN(n10013) );
  NAND2_X1 U12485 ( .A1(n7013), .A2(n10013), .ZN(n12582) );
  NAND2_X1 U12486 ( .A1(n12582), .A2(n10014), .ZN(n10016) );
  XNOR2_X1 U12487 ( .A(n12918), .B(n10028), .ZN(n10015) );
  NAND2_X1 U12488 ( .A1(n12642), .A2(n10017), .ZN(n12565) );
  XNOR2_X1 U12489 ( .A(n10519), .B(n13024), .ZN(n12566) );
  NOR2_X1 U12490 ( .A1(n12566), .A2(n12685), .ZN(n10020) );
  XNOR2_X1 U12491 ( .A(n13020), .B(n10028), .ZN(n10018) );
  NAND2_X1 U12492 ( .A1(n10018), .A2(n12601), .ZN(n12594) );
  OAI21_X1 U12493 ( .B1(n10018), .B2(n12601), .A(n12594), .ZN(n12623) );
  AOI21_X1 U12494 ( .B1(n12566), .B2(n12685), .A(n12623), .ZN(n10019) );
  NAND2_X1 U12495 ( .A1(n12593), .A2(n12594), .ZN(n10024) );
  XNOR2_X1 U12496 ( .A(n12592), .B(n10521), .ZN(n10021) );
  NAND2_X1 U12497 ( .A1(n10021), .A2(n12885), .ZN(n10025) );
  INV_X1 U12498 ( .A(n10021), .ZN(n10022) );
  NAND2_X1 U12499 ( .A1(n10022), .A2(n12684), .ZN(n10023) );
  NAND2_X1 U12500 ( .A1(n10024), .A2(n12595), .ZN(n12597) );
  XNOR2_X1 U12501 ( .A(n12862), .B(n10028), .ZN(n10026) );
  NOR2_X1 U12502 ( .A1(n10026), .A2(n12870), .ZN(n10027) );
  AOI21_X1 U12503 ( .B1(n10026), .B2(n12870), .A(n10027), .ZN(n12661) );
  XNOR2_X1 U12504 ( .A(n12856), .B(n10519), .ZN(n10051) );
  NOR2_X1 U12505 ( .A1(n10051), .A2(n12683), .ZN(n10031) );
  AOI21_X1 U12506 ( .B1(n10051), .B2(n12683), .A(n10031), .ZN(n12555) );
  XNOR2_X1 U12507 ( .A(n12479), .B(n10028), .ZN(n10033) );
  INV_X1 U12508 ( .A(n10033), .ZN(n10052) );
  OAI22_X1 U12509 ( .A1(n10039), .A2(n10513), .B1(n10046), .B2(n10040), .ZN(
        n10030) );
  INV_X1 U12510 ( .A(n10031), .ZN(n10032) );
  NAND3_X1 U12511 ( .A1(n10052), .A2(n12670), .A3(n10032), .ZN(n10057) );
  NAND2_X1 U12512 ( .A1(n12558), .A2(n10034), .ZN(n10056) );
  NAND2_X1 U12513 ( .A1(n10039), .A2(n15073), .ZN(n10035) );
  NAND2_X1 U12514 ( .A1(n10035), .A2(n10664), .ZN(n12681) );
  OR2_X1 U12515 ( .A1(n12541), .A2(n12542), .ZN(n10036) );
  NOR2_X1 U12516 ( .A1(n10046), .A2(n10036), .ZN(n10037) );
  AOI22_X1 U12517 ( .A1(n12683), .A2(n12663), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n10050) );
  NAND2_X1 U12518 ( .A1(n10039), .A2(n10038), .ZN(n10044) );
  INV_X1 U12519 ( .A(n10040), .ZN(n10041) );
  NAND2_X1 U12520 ( .A1(n10046), .A2(n10041), .ZN(n10042) );
  NAND4_X1 U12521 ( .A1(n10044), .A2(n10073), .A3(n10043), .A4(n10042), .ZN(
        n10048) );
  NOR2_X1 U12522 ( .A1(n12541), .A2(n12488), .ZN(n10045) );
  AND2_X1 U12523 ( .A1(n10046), .A2(n10045), .ZN(n10047) );
  AOI21_X1 U12524 ( .B1(n10048), .B2(P3_STATE_REG_SCAN_IN), .A(n10047), .ZN(
        n10407) );
  NAND2_X1 U12525 ( .A1(n12678), .A2(n12841), .ZN(n10049) );
  OAI211_X1 U12526 ( .C1(n11029), .C2(n12665), .A(n10050), .B(n10049), .ZN(
        n10054) );
  NOR4_X1 U12527 ( .A1(n10052), .A2(n10051), .A3(n12683), .A4(n12650), .ZN(
        n10053) );
  AOI211_X1 U12528 ( .C1(n12648), .C2(n7997), .A(n10054), .B(n10053), .ZN(
        n10055) );
  OAI211_X1 U12529 ( .C1(n12558), .C2(n10057), .A(n10056), .B(n10055), .ZN(
        P3_U3160) );
  NOR2_X1 U12530 ( .A1(n10059), .A2(n10058), .ZN(n10199) );
  INV_X1 U12531 ( .A(n10188), .ZN(n10060) );
  INV_X1 U12532 ( .A(n10061), .ZN(n10063) );
  NAND2_X1 U12533 ( .A1(n10063), .A2(n10062), .ZN(n10064) );
  XNOR2_X1 U12534 ( .A(n10065), .B(n10064), .ZN(n10066) );
  NOR2_X1 U12535 ( .A1(n10066), .A2(n12650), .ZN(n10072) );
  NOR2_X1 U12536 ( .A1(n14353), .A2(n12681), .ZN(n10071) );
  AND2_X1 U12537 ( .A1(n12678), .A2(n11913), .ZN(n10070) );
  INV_X1 U12538 ( .A(n12663), .ZN(n12676) );
  INV_X1 U12539 ( .A(n12665), .ZN(n12674) );
  NAND2_X1 U12540 ( .A1(n12674), .A2(n12690), .ZN(n10068) );
  NOR2_X1 U12541 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n7719), .ZN(n12715) );
  INV_X1 U12542 ( .A(n12715), .ZN(n10067) );
  OAI211_X1 U12543 ( .C1(n12676), .C2(n14340), .A(n10068), .B(n10067), .ZN(
        n10069) );
  INV_X1 U12544 ( .A(n10073), .ZN(n10074) );
  AND2_X4 U12545 ( .A1(n10077), .A2(n10076), .ZN(n12282) );
  AOI22_X1 U12546 ( .A1(n12275), .A2(n13772), .B1(n12282), .B2(n10714), .ZN(
        n10078) );
  XNOR2_X1 U12547 ( .A(n10078), .B(n12066), .ZN(n11066) );
  AND2_X4 U12548 ( .A1(n12282), .A2(n14119), .ZN(n12284) );
  AOI22_X1 U12549 ( .A1(n12284), .A2(n13772), .B1(n12285), .B2(n10714), .ZN(
        n11067) );
  XNOR2_X1 U12550 ( .A(n11066), .B(n11067), .ZN(n10106) );
  NAND2_X1 U12551 ( .A1(n12284), .A2(n13776), .ZN(n10080) );
  INV_X1 U12552 ( .A(n10077), .ZN(n10081) );
  AOI22_X1 U12553 ( .A1(n11076), .A2(n10730), .B1(n10081), .B2(n14256), .ZN(
        n10079) );
  NAND2_X1 U12554 ( .A1(n10080), .A2(n10079), .ZN(n10719) );
  NAND2_X1 U12555 ( .A1(n13776), .A2(n11076), .ZN(n10084) );
  NAND2_X1 U12556 ( .A1(n10081), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10083) );
  NAND2_X1 U12557 ( .A1(n12282), .A2(n10730), .ZN(n10082) );
  AND3_X1 U12558 ( .A1(n10084), .A2(n10083), .A3(n10082), .ZN(n10718) );
  XNOR2_X1 U12559 ( .A(n12066), .B(n10086), .ZN(n10090) );
  NOR2_X1 U12560 ( .A1(n12092), .A2(n10087), .ZN(n10088) );
  AOI21_X1 U12561 ( .B1(n12284), .B2(n13774), .A(n10088), .ZN(n10089) );
  XNOR2_X1 U12562 ( .A(n10090), .B(n10089), .ZN(n10690) );
  NOR2_X1 U12563 ( .A1(n10692), .A2(n10690), .ZN(n10691) );
  NOR2_X1 U12564 ( .A1(n10691), .A2(n10091), .ZN(n10646) );
  OAI22_X1 U12565 ( .A1(n10693), .A2(n12092), .B1(n14503), .B2(n12090), .ZN(
        n10092) );
  XNOR2_X1 U12566 ( .A(n10092), .B(n12066), .ZN(n10094) );
  OAI22_X1 U12567 ( .A1(n12125), .A2(n10693), .B1(n14503), .B2(n12092), .ZN(
        n10093) );
  XNOR2_X1 U12568 ( .A(n10094), .B(n10093), .ZN(n10647) );
  OAI22_X1 U12569 ( .A1(n10646), .A2(n10647), .B1(n10094), .B2(n10093), .ZN(
        n10105) );
  NOR2_X1 U12570 ( .A1(n10096), .A2(n10095), .ZN(n10701) );
  INV_X1 U12571 ( .A(n10097), .ZN(n10098) );
  NAND2_X1 U12572 ( .A1(n10701), .A2(n10098), .ZN(n10117) );
  INV_X1 U12573 ( .A(n10181), .ZN(n10231) );
  OR2_X1 U12574 ( .A1(n10117), .A2(n10231), .ZN(n10113) );
  INV_X1 U12575 ( .A(n10113), .ZN(n10101) );
  AND2_X1 U12576 ( .A1(n14528), .A2(n10099), .ZN(n10100) );
  INV_X1 U12577 ( .A(n10105), .ZN(n10103) );
  NAND2_X1 U12578 ( .A1(n10103), .A2(n10102), .ZN(n11070) );
  AOI211_X1 U12579 ( .C1(n10106), .C2(n10105), .A(n13731), .B(n10104), .ZN(
        n10121) );
  NAND2_X1 U12580 ( .A1(n10117), .A2(n10107), .ZN(n10652) );
  AND3_X1 U12581 ( .A1(n10077), .A2(n10108), .A3(n10232), .ZN(n10109) );
  NAND2_X1 U12582 ( .A1(n10652), .A2(n10109), .ZN(n10110) );
  MUX2_X1 U12583 ( .A(n13742), .B(P1_U3086), .S(P1_REG3_REG_3__SCAN_IN), .Z(
        n10120) );
  NAND2_X1 U12584 ( .A1(n9118), .A2(n10111), .ZN(n10713) );
  INV_X1 U12585 ( .A(n6468), .ZN(n13745) );
  NOR2_X1 U12586 ( .A1(n11071), .A2(n13633), .ZN(n10115) );
  NOR2_X1 U12587 ( .A1(n10693), .A2(n13624), .ZN(n10114) );
  OR2_X1 U12588 ( .A1(n10115), .A2(n10114), .ZN(n10708) );
  INV_X1 U12589 ( .A(n10708), .ZN(n10118) );
  OAI22_X1 U12590 ( .A1(n13745), .A2(n14514), .B1(n10118), .B2(n13739), .ZN(
        n10119) );
  OR3_X1 U12591 ( .A1(n10121), .A2(n10120), .A3(n10119), .ZN(P1_U3218) );
  MUX2_X1 U12592 ( .A(P2_RD_REG_SCAN_IN), .B(n7465), .S(P1_RD_REG_SCAN_IN), 
        .Z(n10123) );
  NAND2_X1 U12593 ( .A1(n10123), .A2(n10122), .ZN(U29) );
  OAI222_X1 U12594 ( .A1(n13138), .A2(n10125), .B1(n12303), .B2(n10124), .C1(
        P3_U3151), .C2(n14947), .ZN(P3_U3287) );
  INV_X1 U12595 ( .A(n10126), .ZN(n10127) );
  OAI222_X1 U12596 ( .A1(P3_U3151), .A2(n14861), .B1(n12303), .B2(n10128), 
        .C1(n13138), .C2(n10127), .ZN(P3_U3292) );
  AND2_X1 U12597 ( .A1(n6706), .A2(P1_U3086), .ZN(n14239) );
  INV_X2 U12598 ( .A(n14239), .ZN(n14245) );
  AND2_X1 U12599 ( .A1(n8726), .A2(P1_U3086), .ZN(n11751) );
  INV_X2 U12600 ( .A(n11751), .ZN(n14251) );
  OAI222_X1 U12601 ( .A1(n14245), .A2(n10129), .B1(n14251), .B2(n10143), .C1(
        P1_U3086), .C2(n13812), .ZN(P1_U3352) );
  INV_X1 U12602 ( .A(n10130), .ZN(n10177) );
  OAI222_X1 U12603 ( .A1(n14245), .A2(n10131), .B1(n14251), .B2(n10177), .C1(
        n13789), .C2(P1_U3086), .ZN(P1_U3353) );
  INV_X1 U12604 ( .A(n10132), .ZN(n10138) );
  INV_X1 U12605 ( .A(n10382), .ZN(n12143) );
  OAI222_X1 U12606 ( .A1(n14245), .A2(n10133), .B1(n14251), .B2(n10138), .C1(
        n12143), .C2(P1_U3086), .ZN(P1_U3351) );
  OAI222_X1 U12607 ( .A1(n10379), .A2(P1_U3086), .B1(n14251), .B2(n10144), 
        .C1(n10134), .C2(n14245), .ZN(P1_U3354) );
  INV_X1 U12608 ( .A(n10384), .ZN(n10544) );
  INV_X1 U12609 ( .A(n10135), .ZN(n10140) );
  OAI222_X1 U12610 ( .A1(n10544), .A2(P1_U3086), .B1(n14251), .B2(n10140), 
        .C1(n10136), .C2(n14245), .ZN(P1_U3350) );
  NOR2_X1 U12611 ( .A1(n6475), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13593) );
  INV_X1 U12612 ( .A(n13593), .ZN(n13591) );
  NAND2_X1 U12613 ( .A1(n6706), .A2(P2_U3088), .ZN(n13596) );
  INV_X1 U12614 ( .A(n14583), .ZN(n10137) );
  OAI222_X1 U12615 ( .A1(n13591), .A2(n10139), .B1(n13596), .B2(n10138), .C1(
        P2_U3088), .C2(n10137), .ZN(P2_U3323) );
  INV_X1 U12616 ( .A(n14599), .ZN(n10254) );
  OAI222_X1 U12617 ( .A1(n13591), .A2(n10141), .B1(n13596), .B2(n10140), .C1(
        P2_U3088), .C2(n10254), .ZN(P2_U3322) );
  INV_X1 U12618 ( .A(n10253), .ZN(n10318) );
  OAI222_X1 U12619 ( .A1(P2_U3088), .A2(n10318), .B1(n13596), .B2(n10143), 
        .C1(n10142), .C2(n13591), .ZN(P2_U3324) );
  OAI222_X1 U12620 ( .A1(n13591), .A2(n10145), .B1(n13596), .B2(n10144), .C1(
        P2_U3088), .C2(n10217), .ZN(P2_U3326) );
  INV_X1 U12621 ( .A(n10146), .ZN(n10147) );
  OAI222_X1 U12622 ( .A1(P3_U3151), .A2(n11665), .B1(n12303), .B2(n10148), 
        .C1(n13138), .C2(n10147), .ZN(P3_U3285) );
  OAI222_X1 U12623 ( .A1(n13138), .A2(n10150), .B1(n12303), .B2(n10149), .C1(
        P3_U3151), .C2(n10345), .ZN(P3_U3294) );
  INV_X1 U12624 ( .A(n10385), .ZN(n10420) );
  INV_X1 U12625 ( .A(n10151), .ZN(n10179) );
  OAI222_X1 U12626 ( .A1(n10420), .A2(P1_U3086), .B1(n14251), .B2(n10179), 
        .C1(n10152), .C2(n14245), .ZN(P1_U3349) );
  INV_X1 U12627 ( .A(n13138), .ZN(n14270) );
  INV_X1 U12628 ( .A(n12303), .ZN(n14268) );
  AOI222_X1 U12629 ( .A1(n10153), .A2(n14270), .B1(n11672), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_5_), .C2(n14268), .ZN(n10154) );
  INV_X1 U12630 ( .A(n10154), .ZN(P3_U3290) );
  AOI222_X1 U12631 ( .A1(n10155), .A2(n14270), .B1(SI_4_), .B2(n14268), .C1(
        n11670), .C2(P3_STATE_REG_SCAN_IN), .ZN(n10156) );
  INV_X1 U12632 ( .A(n10156), .ZN(P3_U3291) );
  OAI222_X1 U12633 ( .A1(n14913), .A2(P3_U3151), .B1(n13138), .B2(n10158), 
        .C1(n10157), .C2(n12303), .ZN(P3_U3289) );
  INV_X1 U12634 ( .A(n10159), .ZN(n10160) );
  OAI222_X1 U12635 ( .A1(P3_U3151), .A2(n14965), .B1(n12303), .B2(n10161), 
        .C1(n13138), .C2(n10160), .ZN(P3_U3286) );
  OAI222_X1 U12636 ( .A1(P3_U3151), .A2(n11803), .B1(n12303), .B2(n10163), 
        .C1(n13138), .C2(n10162), .ZN(P3_U3284) );
  INV_X1 U12637 ( .A(n10429), .ZN(n10397) );
  INV_X1 U12638 ( .A(n10164), .ZN(n10175) );
  OAI222_X1 U12639 ( .A1(n10397), .A2(P1_U3086), .B1(n14251), .B2(n10175), 
        .C1(n10165), .C2(n14245), .ZN(P1_U3348) );
  OAI222_X1 U12640 ( .A1(P3_U3151), .A2(n12708), .B1(n12303), .B2(n10167), 
        .C1(n13138), .C2(n10166), .ZN(P3_U3283) );
  AND2_X1 U12641 ( .A1(n10169), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U12642 ( .A1(n10169), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U12643 ( .A1(n10169), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U12644 ( .A1(n10169), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U12645 ( .A1(n10169), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U12646 ( .A1(n10169), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U12647 ( .A1(n10169), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U12648 ( .A1(n10169), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U12649 ( .A1(n10169), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U12650 ( .A1(n10169), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U12651 ( .A1(n10169), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U12652 ( .A1(n10169), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U12653 ( .A1(n10169), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U12654 ( .A1(n10169), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U12655 ( .A1(n10169), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U12656 ( .A1(n10169), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U12657 ( .A1(n10169), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U12658 ( .A1(n10169), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U12659 ( .A1(n10169), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U12660 ( .A1(n10169), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U12661 ( .A1(n10169), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U12662 ( .A1(n10169), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U12663 ( .A1(n10169), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U12664 ( .A1(n10169), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U12665 ( .A1(n10169), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U12666 ( .A1(n10169), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U12667 ( .A1(n10169), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U12668 ( .A1(n10169), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U12669 ( .A1(n10169), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U12670 ( .A1(n10169), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  INV_X1 U12671 ( .A(n10549), .ZN(n10554) );
  INV_X1 U12672 ( .A(n10170), .ZN(n10173) );
  OAI222_X1 U12673 ( .A1(n10554), .A2(P1_U3086), .B1(n14251), .B2(n10173), 
        .C1(n10171), .C2(n14245), .ZN(P1_U3347) );
  INV_X1 U12674 ( .A(n13596), .ZN(n12220) );
  INV_X1 U12675 ( .A(n12220), .ZN(n13589) );
  INV_X1 U12676 ( .A(n10585), .ZN(n10172) );
  OAI222_X1 U12677 ( .A1(n13591), .A2(n10174), .B1(n13589), .B2(n10173), .C1(
        P2_U3088), .C2(n10172), .ZN(P2_U3319) );
  INV_X1 U12678 ( .A(n10268), .ZN(n10263) );
  OAI222_X1 U12679 ( .A1(n13591), .A2(n10176), .B1(n13589), .B2(n10175), .C1(
        P2_U3088), .C2(n10263), .ZN(P2_U3320) );
  OAI222_X1 U12680 ( .A1(n13591), .A2(n10178), .B1(n13589), .B2(n10177), .C1(
        P2_U3088), .C2(n14562), .ZN(P2_U3325) );
  INV_X1 U12681 ( .A(n10290), .ZN(n10304) );
  OAI222_X1 U12682 ( .A1(n13591), .A2(n10180), .B1(n13589), .B2(n10179), .C1(
        P2_U3088), .C2(n10304), .ZN(P2_U3321) );
  NAND2_X1 U12683 ( .A1(n10182), .A2(n10181), .ZN(n14492) );
  INV_X1 U12684 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10185) );
  INV_X1 U12685 ( .A(n10183), .ZN(n10184) );
  AOI22_X1 U12686 ( .A1(n14492), .A2(n10185), .B1(n10188), .B2(n10184), .ZN(
        P1_U3446) );
  INV_X1 U12687 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10189) );
  INV_X1 U12688 ( .A(n10186), .ZN(n10187) );
  AOI22_X1 U12689 ( .A1(n14492), .A2(n10189), .B1(n10188), .B2(n10187), .ZN(
        P1_U3445) );
  INV_X1 U12690 ( .A(n10190), .ZN(n10193) );
  INV_X1 U12691 ( .A(n14614), .ZN(n10586) );
  OAI222_X1 U12692 ( .A1(n13591), .A2(n10191), .B1(n13589), .B2(n10193), .C1(
        P2_U3088), .C2(n10586), .ZN(P2_U3318) );
  INV_X1 U12693 ( .A(n13834), .ZN(n10194) );
  OAI222_X1 U12694 ( .A1(n10194), .A2(P1_U3086), .B1(n14251), .B2(n10193), 
        .C1(n10192), .C2(n14245), .ZN(P1_U3346) );
  NAND2_X1 U12695 ( .A1(n10473), .A2(n10195), .ZN(n10197) );
  AND2_X1 U12696 ( .A1(n10197), .A2(n10196), .ZN(n10198) );
  AND2_X1 U12697 ( .A1(n10202), .A2(n8608), .ZN(n14561) );
  AND2_X1 U12698 ( .A1(n14561), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14685) );
  NOR2_X1 U12699 ( .A1(n14647), .A2(n10200), .ZN(n10206) );
  NAND2_X1 U12700 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n10204) );
  INV_X1 U12701 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n14834) );
  MUX2_X1 U12702 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n14834), .S(n10217), .Z(
        n10203) );
  INV_X1 U12703 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10201) );
  NOR3_X1 U12704 ( .A1(n10203), .A2(n10226), .A3(n10201), .ZN(n10250) );
  NOR2_X1 U12705 ( .A1(n8608), .A2(P2_U3088), .ZN(n13584) );
  NAND2_X1 U12706 ( .A1(n10202), .A2(n13584), .ZN(n10207) );
  AOI211_X1 U12707 ( .C1(n10204), .C2(n10203), .A(n10250), .B(n14595), .ZN(
        n10205) );
  AOI211_X1 U12708 ( .C1(P2_REG3_REG_1__SCAN_IN), .C2(P2_U3088), .A(n10206), 
        .B(n10205), .ZN(n10216) );
  INV_X1 U12709 ( .A(n10207), .ZN(n10209) );
  INV_X1 U12710 ( .A(n10217), .ZN(n10251) );
  NAND2_X1 U12711 ( .A1(n10251), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10240) );
  INV_X1 U12712 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10212) );
  NAND2_X1 U12713 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n10210) );
  AOI21_X1 U12714 ( .B1(n10217), .B2(n10212), .A(n10210), .ZN(n10211) );
  NAND2_X1 U12715 ( .A1(n10240), .A2(n10211), .ZN(n10241) );
  INV_X1 U12716 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n14735) );
  MUX2_X1 U12717 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n10212), .S(n10217), .Z(
        n10213) );
  OAI21_X1 U12718 ( .B1(n14735), .B2(n10226), .A(n10213), .ZN(n10214) );
  NAND3_X1 U12719 ( .A1(n14692), .A2(n10241), .A3(n10214), .ZN(n10215) );
  OAI211_X1 U12720 ( .C1(n14620), .C2(n10217), .A(n10216), .B(n10215), .ZN(
        P2_U3215) );
  OAI222_X1 U12721 ( .A1(P3_U3151), .A2(n12727), .B1(n12303), .B2(n10219), 
        .C1(n13138), .C2(n10218), .ZN(P3_U3282) );
  INV_X1 U12722 ( .A(n10677), .ZN(n10562) );
  INV_X1 U12723 ( .A(n10220), .ZN(n10222) );
  OAI222_X1 U12724 ( .A1(n10562), .A2(P1_U3086), .B1(n14251), .B2(n10222), 
        .C1(n10221), .C2(n14245), .ZN(P1_U3345) );
  INV_X1 U12725 ( .A(n10588), .ZN(n14619) );
  OAI222_X1 U12726 ( .A1(n13591), .A2(n10223), .B1(n13596), .B2(n10222), .C1(
        P2_U3088), .C2(n14619), .ZN(P2_U3317) );
  NAND2_X1 U12727 ( .A1(n14692), .A2(n14735), .ZN(n10224) );
  OAI211_X1 U12728 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n14595), .A(n14620), .B(
        n10224), .ZN(n10225) );
  INV_X1 U12729 ( .A(n10225), .ZN(n10228) );
  INV_X1 U12730 ( .A(n14595), .ZN(n14688) );
  AOI22_X1 U12731 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(n14688), .B1(n14692), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n10227) );
  MUX2_X1 U12732 ( .A(n10228), .B(n10227), .S(n10226), .Z(n10230) );
  INV_X1 U12733 ( .A(n14647), .ZN(n14684) );
  AOI22_X1 U12734 ( .A1(n14684), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n10229) );
  NAND2_X1 U12735 ( .A1(n10230), .A2(n10229), .ZN(P2_U3214) );
  NAND2_X1 U12736 ( .A1(n10231), .A2(n11753), .ZN(n10282) );
  NAND2_X1 U12737 ( .A1(n10233), .A2(n10232), .ZN(n10234) );
  NAND2_X1 U12738 ( .A1(n10234), .A2(n8739), .ZN(n10280) );
  NAND2_X1 U12739 ( .A1(n10282), .A2(n10280), .ZN(n14473) );
  INV_X1 U12740 ( .A(n14473), .ZN(n13827) );
  CLKBUF_X2 U12741 ( .A(P1_U4016), .Z(n13775) );
  NOR2_X1 U12742 ( .A1(n13827), .A2(n13775), .ZN(P1_U3085) );
  INV_X1 U12743 ( .A(n10235), .ZN(n10238) );
  INV_X1 U12744 ( .A(n11034), .ZN(n10582) );
  OAI222_X1 U12745 ( .A1(n13591), .A2(n10236), .B1(n13596), .B2(n10238), .C1(
        P2_U3088), .C2(n10582), .ZN(P2_U3316) );
  INV_X1 U12746 ( .A(n10817), .ZN(n10682) );
  OAI222_X1 U12747 ( .A1(n10682), .A2(P1_U3086), .B1(n14251), .B2(n10238), 
        .C1(n10237), .C2(n14245), .ZN(P1_U3344) );
  INV_X1 U12748 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10239) );
  MUX2_X1 U12749 ( .A(n10239), .B(P2_REG2_REG_3__SCAN_IN), .S(n10253), .Z(
        n10307) );
  XNOR2_X1 U12750 ( .A(n14562), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n14564) );
  NAND2_X1 U12751 ( .A1(n10241), .A2(n10240), .ZN(n14565) );
  AOI22_X1 U12752 ( .A1(n14564), .A2(n14565), .B1(n10252), .B2(
        P2_REG2_REG_2__SCAN_IN), .ZN(n10308) );
  OR2_X1 U12753 ( .A1(n10307), .A2(n10308), .ZN(n14578) );
  NAND2_X1 U12754 ( .A1(n10253), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n14577) );
  INV_X1 U12755 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11006) );
  MUX2_X1 U12756 ( .A(n11006), .B(P2_REG2_REG_4__SCAN_IN), .S(n14583), .Z(
        n14576) );
  AOI21_X1 U12757 ( .B1(n14578), .B2(n14577), .A(n14576), .ZN(n14580) );
  AOI21_X1 U12758 ( .B1(n14583), .B2(P2_REG2_REG_4__SCAN_IN), .A(n14580), .ZN(
        n14602) );
  INV_X1 U12759 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10242) );
  MUX2_X1 U12760 ( .A(n10242), .B(P2_REG2_REG_5__SCAN_IN), .S(n14599), .Z(
        n14601) );
  AOI21_X1 U12761 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n14599), .A(n14600), .ZN(
        n10298) );
  INV_X1 U12762 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10244) );
  MUX2_X1 U12763 ( .A(n10244), .B(P2_REG2_REG_6__SCAN_IN), .S(n10290), .Z(
        n10297) );
  INV_X1 U12764 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10243) );
  MUX2_X1 U12765 ( .A(n10243), .B(P2_REG2_REG_7__SCAN_IN), .S(n10268), .Z(
        n10246) );
  NOR2_X1 U12766 ( .A1(n10304), .A2(n10244), .ZN(n10248) );
  INV_X1 U12767 ( .A(n10248), .ZN(n10245) );
  NAND2_X1 U12768 ( .A1(n10246), .A2(n10245), .ZN(n10249) );
  MUX2_X1 U12769 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10243), .S(n10268), .Z(
        n10247) );
  OAI21_X1 U12770 ( .B1(n10296), .B2(n10248), .A(n10247), .ZN(n10272) );
  OAI211_X1 U12771 ( .C1(n10296), .C2(n10249), .A(n10272), .B(n14692), .ZN(
        n10262) );
  NAND2_X1 U12772 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n10786) );
  INV_X1 U12773 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10860) );
  AOI21_X1 U12774 ( .B1(n10251), .B2(P2_REG1_REG_1__SCAN_IN), .A(n10250), .ZN(
        n14568) );
  INV_X1 U12775 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n14836) );
  MUX2_X1 U12776 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n14836), .S(n14562), .Z(
        n14567) );
  OR2_X1 U12777 ( .A1(n14568), .A2(n14567), .ZN(n14570) );
  NAND2_X1 U12778 ( .A1(n10252), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10313) );
  INV_X1 U12779 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n14838) );
  MUX2_X1 U12780 ( .A(n14838), .B(P2_REG1_REG_3__SCAN_IN), .S(n10253), .Z(
        n10312) );
  AOI21_X1 U12781 ( .B1(P2_REG1_REG_3__SCAN_IN), .B2(n10253), .A(n10311), .ZN(
        n14585) );
  INV_X1 U12782 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n14840) );
  MUX2_X1 U12783 ( .A(n14840), .B(P2_REG1_REG_4__SCAN_IN), .S(n14583), .Z(
        n14584) );
  OR2_X1 U12784 ( .A1(n14585), .A2(n14584), .ZN(n14593) );
  NAND2_X1 U12785 ( .A1(n14583), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n14592) );
  INV_X1 U12786 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n14842) );
  MUX2_X1 U12787 ( .A(n14842), .B(P2_REG1_REG_5__SCAN_IN), .S(n14599), .Z(
        n14591) );
  NOR2_X1 U12788 ( .A1(n10254), .A2(n14842), .ZN(n10291) );
  MUX2_X1 U12789 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10860), .S(n10290), .Z(
        n10255) );
  OAI21_X1 U12790 ( .B1(n14596), .B2(n10291), .A(n10255), .ZN(n10294) );
  OAI21_X1 U12791 ( .B1(n10860), .B2(n10304), .A(n10294), .ZN(n10258) );
  INV_X1 U12792 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10256) );
  MUX2_X1 U12793 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10256), .S(n10268), .Z(
        n10257) );
  NAND2_X1 U12794 ( .A1(n10258), .A2(n10257), .ZN(n10266) );
  OAI211_X1 U12795 ( .C1(n10258), .C2(n10257), .A(n14688), .B(n10266), .ZN(
        n10259) );
  NAND2_X1 U12796 ( .A1(n10786), .A2(n10259), .ZN(n10260) );
  AOI21_X1 U12797 ( .B1(n14684), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n10260), .ZN(
        n10261) );
  OAI211_X1 U12798 ( .C1(n14620), .C2(n10263), .A(n10262), .B(n10261), .ZN(
        P2_U3221) );
  NAND2_X1 U12799 ( .A1(n10268), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10265) );
  INV_X1 U12800 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n14845) );
  MUX2_X1 U12801 ( .A(n14845), .B(P2_REG1_REG_8__SCAN_IN), .S(n10585), .Z(
        n10264) );
  NAND3_X1 U12802 ( .A1(n10266), .A2(n10265), .A3(n10264), .ZN(n10267) );
  NAND2_X1 U12803 ( .A1(n10267), .A2(n14688), .ZN(n10277) );
  NAND2_X1 U12804 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n10938) );
  OAI21_X1 U12805 ( .B1(n14647), .B2(n14277), .A(n10938), .ZN(n10275) );
  NAND2_X1 U12806 ( .A1(n10268), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10271) );
  INV_X1 U12807 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10269) );
  MUX2_X1 U12808 ( .A(n10269), .B(P2_REG2_REG_8__SCAN_IN), .S(n10585), .Z(
        n10270) );
  AOI21_X1 U12809 ( .B1(n10272), .B2(n10271), .A(n10270), .ZN(n10574) );
  AND3_X1 U12810 ( .A1(n10272), .A2(n10271), .A3(n10270), .ZN(n10273) );
  NOR3_X1 U12811 ( .A1(n10574), .A2(n10273), .A3(n14652), .ZN(n10274) );
  AOI211_X1 U12812 ( .C1(n14685), .C2(n10585), .A(n10275), .B(n10274), .ZN(
        n10276) );
  OAI21_X1 U12813 ( .B1(n10584), .B2(n10277), .A(n10276), .ZN(P2_U3222) );
  OAI222_X1 U12814 ( .A1(P3_U3151), .A2(n12734), .B1(n12303), .B2(n10279), 
        .C1(n13138), .C2(n10278), .ZN(P3_U3281) );
  INV_X1 U12815 ( .A(n10280), .ZN(n10281) );
  NAND2_X1 U12816 ( .A1(n10282), .A2(n10281), .ZN(n10377) );
  INV_X1 U12817 ( .A(n14248), .ZN(n13888) );
  NOR2_X1 U12818 ( .A1(n14248), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n10283) );
  OR2_X1 U12819 ( .A1(n6483), .A2(n10283), .ZN(n12153) );
  INV_X1 U12820 ( .A(n12153), .ZN(n10284) );
  OAI21_X1 U12821 ( .B1(n13888), .B2(P1_REG1_REG_0__SCAN_IN), .A(n10284), .ZN(
        n10285) );
  MUX2_X1 U12822 ( .A(n10285), .B(n10284), .S(n14256), .Z(n10286) );
  INV_X1 U12823 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n11186) );
  OAI22_X1 U12824 ( .A1(n10377), .A2(n10286), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11186), .ZN(n10288) );
  NOR3_X1 U12825 ( .A1(n13880), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n12152), .ZN(
        n10287) );
  AOI211_X1 U12826 ( .C1(n13827), .C2(P1_ADDR_REG_0__SCAN_IN), .A(n10288), .B(
        n10287), .ZN(n10289) );
  INV_X1 U12827 ( .A(n10289), .ZN(P1_U3243) );
  MUX2_X1 U12828 ( .A(n10860), .B(P2_REG1_REG_6__SCAN_IN), .S(n10290), .Z(
        n10293) );
  INV_X1 U12829 ( .A(n10291), .ZN(n10292) );
  NAND2_X1 U12830 ( .A1(n10293), .A2(n10292), .ZN(n10295) );
  OAI211_X1 U12831 ( .C1(n14596), .C2(n10295), .A(n10294), .B(n14688), .ZN(
        n10303) );
  NAND2_X1 U12832 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n10903) );
  AOI211_X1 U12833 ( .C1(n10298), .C2(n10297), .A(n10296), .B(n14652), .ZN(
        n10299) );
  INV_X1 U12834 ( .A(n10299), .ZN(n10300) );
  NAND2_X1 U12835 ( .A1(n10903), .A2(n10300), .ZN(n10301) );
  AOI21_X1 U12836 ( .B1(n14684), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n10301), .ZN(
        n10302) );
  OAI211_X1 U12837 ( .C1(n14620), .C2(n10304), .A(n10303), .B(n10302), .ZN(
        P2_U3220) );
  INV_X1 U12838 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10305) );
  NOR2_X1 U12839 ( .A1(n14647), .A2(n10305), .ZN(n10310) );
  INV_X1 U12840 ( .A(n14578), .ZN(n10306) );
  AOI211_X1 U12841 ( .C1(n10308), .C2(n10307), .A(n10306), .B(n14652), .ZN(
        n10309) );
  AOI211_X1 U12842 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(P2_U3088), .A(n10310), 
        .B(n10309), .ZN(n10317) );
  INV_X1 U12843 ( .A(n10311), .ZN(n10315) );
  NAND3_X1 U12844 ( .A1(n14570), .A2(n10313), .A3(n10312), .ZN(n10314) );
  NAND3_X1 U12845 ( .A1(n14688), .A2(n10315), .A3(n10314), .ZN(n10316) );
  OAI211_X1 U12846 ( .C1(n14620), .C2(n10318), .A(n10317), .B(n10316), .ZN(
        P2_U3217) );
  OAI222_X1 U12847 ( .A1(P3_U3151), .A2(n12795), .B1(n12303), .B2(n10320), 
        .C1(n13138), .C2(n10319), .ZN(P3_U3280) );
  INV_X1 U12848 ( .A(n14643), .ZN(n11035) );
  INV_X1 U12849 ( .A(n10321), .ZN(n10324) );
  OAI222_X1 U12850 ( .A1(P2_U3088), .A2(n11035), .B1(n13596), .B2(n10324), 
        .C1(n10322), .C2(n13591), .ZN(P2_U3315) );
  INV_X1 U12851 ( .A(n11021), .ZN(n10821) );
  OAI222_X1 U12852 ( .A1(P1_U3086), .A2(n10821), .B1(n14251), .B2(n10324), 
        .C1(n10323), .C2(n14245), .ZN(P1_U3343) );
  INV_X1 U12853 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10325) );
  MUX2_X1 U12854 ( .A(n10326), .B(n10325), .S(n7931), .Z(n10327) );
  INV_X1 U12855 ( .A(n10345), .ZN(n10509) );
  NAND2_X1 U12856 ( .A1(n10327), .A2(n10509), .ZN(n10330) );
  OAI21_X1 U12857 ( .B1(n10327), .B2(n10509), .A(n10330), .ZN(n10499) );
  INV_X1 U12858 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10328) );
  MUX2_X1 U12859 ( .A(n10329), .B(n10328), .S(n6473), .Z(n10603) );
  NAND2_X1 U12860 ( .A1(n10603), .A2(n13142), .ZN(n10614) );
  INV_X1 U12861 ( .A(n10330), .ZN(n10336) );
  INV_X1 U12862 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10356) );
  MUX2_X1 U12863 ( .A(n10331), .B(n10356), .S(n12776), .Z(n10332) );
  NAND2_X1 U12864 ( .A1(n10332), .A2(n10347), .ZN(n14857) );
  INV_X1 U12865 ( .A(n10332), .ZN(n10333) );
  NAND2_X1 U12866 ( .A1(n10333), .A2(n6476), .ZN(n10334) );
  AND2_X1 U12867 ( .A1(n14857), .A2(n10334), .ZN(n10335) );
  OAI21_X1 U12868 ( .B1(n10498), .B2(n10336), .A(n10335), .ZN(n14858) );
  INV_X1 U12869 ( .A(n14858), .ZN(n10338) );
  NOR3_X1 U12870 ( .A1(n10498), .A2(n10336), .A3(n10335), .ZN(n10337) );
  NAND2_X1 U12871 ( .A1(P3_U3897), .A2(n13139), .ZN(n14985) );
  OAI21_X1 U12872 ( .B1(n10338), .B2(n10337), .A(n14962), .ZN(n10367) );
  NAND2_X1 U12873 ( .A1(n12496), .A2(n10339), .ZN(n10340) );
  NAND2_X1 U12874 ( .A1(n10341), .A2(n10340), .ZN(n10353) );
  AND2_X1 U12875 ( .A1(n12541), .A2(n12546), .ZN(n10352) );
  INV_X1 U12876 ( .A(P3_U3897), .ZN(n12702) );
  MUX2_X1 U12877 ( .A(n10355), .B(n12702), .S(n10342), .Z(n14966) );
  INV_X1 U12878 ( .A(n14966), .ZN(n14996) );
  NOR2_X1 U12879 ( .A1(n13142), .A2(n10329), .ZN(n10608) );
  NAND2_X1 U12880 ( .A1(n10346), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10344) );
  OAI21_X1 U12881 ( .B1(n10345), .B2(n10608), .A(n10344), .ZN(n10504) );
  NOR2_X1 U12882 ( .A1(n10326), .A2(n10504), .ZN(n10503) );
  AOI21_X1 U12883 ( .B1(P3_REG2_REG_0__SCAN_IN), .B2(n10346), .A(n10503), .ZN(
        n10349) );
  AOI22_X1 U12884 ( .A1(n10347), .A2(P3_REG2_REG_2__SCAN_IN), .B1(n10331), 
        .B2(n6476), .ZN(n10348) );
  NOR2_X1 U12885 ( .A1(n10349), .A2(n10348), .ZN(n11605) );
  AOI21_X1 U12886 ( .B1(n10349), .B2(n10348), .A(n11605), .ZN(n10350) );
  INV_X1 U12887 ( .A(n10350), .ZN(n10351) );
  NAND2_X1 U12888 ( .A1(n14300), .A2(n10351), .ZN(n10364) );
  INV_X1 U12889 ( .A(n10352), .ZN(n10354) );
  AOI22_X1 U12890 ( .A1(n14969), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10363) );
  NOR2_X1 U12891 ( .A1(n10328), .A2(n13142), .ZN(n10607) );
  INV_X1 U12892 ( .A(n10607), .ZN(n10358) );
  NOR2_X1 U12893 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n10358), .ZN(n10357) );
  NAND2_X1 U12894 ( .A1(P3_REG1_REG_1__SCAN_IN), .A2(n10501), .ZN(n10500) );
  OAI21_X1 U12895 ( .B1(P3_IR_REG_1__SCAN_IN), .B2(n10358), .A(n10500), .ZN(
        n10359) );
  NAND2_X1 U12896 ( .A1(n10360), .A2(n10359), .ZN(n11666) );
  OAI21_X1 U12897 ( .B1(n10360), .B2(n10359), .A(n11666), .ZN(n10361) );
  NAND2_X1 U12898 ( .A1(n6467), .A2(n10361), .ZN(n10362) );
  NAND3_X1 U12899 ( .A1(n10364), .A2(n10363), .A3(n10362), .ZN(n10365) );
  AOI21_X1 U12900 ( .B1(n10347), .B2(n14996), .A(n10365), .ZN(n10366) );
  NAND2_X1 U12901 ( .A1(n10367), .A2(n10366), .ZN(P3_U3184) );
  INV_X1 U12902 ( .A(n14289), .ZN(n12793) );
  OAI222_X1 U12903 ( .A1(n12303), .A2(n10369), .B1(n13138), .B2(n10368), .C1(
        n12793), .C2(P3_U3151), .ZN(P3_U3279) );
  INV_X1 U12904 ( .A(n13812), .ZN(n10371) );
  INV_X1 U12905 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10370) );
  OAI21_X1 U12906 ( .B1(n10370), .B2(n10379), .A(n13780), .ZN(n13799) );
  INV_X1 U12907 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n14551) );
  MUX2_X1 U12908 ( .A(n14551), .B(P1_REG1_REG_2__SCAN_IN), .S(n13789), .Z(
        n13800) );
  NAND2_X1 U12909 ( .A1(n13799), .A2(n13800), .ZN(n13798) );
  OAI21_X1 U12910 ( .B1(n13789), .B2(n14551), .A(n13798), .ZN(n13809) );
  INV_X1 U12911 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n14553) );
  MUX2_X1 U12912 ( .A(n14553), .B(P1_REG1_REG_3__SCAN_IN), .S(n13812), .Z(
        n13810) );
  INV_X1 U12913 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10372) );
  MUX2_X1 U12914 ( .A(n10372), .B(P1_REG1_REG_4__SCAN_IN), .S(n10382), .Z(
        n12145) );
  XOR2_X1 U12915 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10384), .Z(n10534) );
  NAND2_X1 U12916 ( .A1(n10533), .A2(n10534), .ZN(n10532) );
  OAI21_X1 U12917 ( .B1(n10384), .B2(P1_REG1_REG_5__SCAN_IN), .A(n10532), .ZN(
        n10413) );
  INV_X1 U12918 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10373) );
  MUX2_X1 U12919 ( .A(n10373), .B(P1_REG1_REG_6__SCAN_IN), .S(n10385), .Z(
        n10414) );
  NOR2_X1 U12920 ( .A1(n10413), .A2(n10414), .ZN(n10412) );
  INV_X1 U12921 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10374) );
  MUX2_X1 U12922 ( .A(n10374), .B(P1_REG1_REG_7__SCAN_IN), .S(n10429), .Z(
        n10375) );
  AOI211_X1 U12923 ( .C1(n10376), .C2(n10375), .A(n13880), .B(n10428), .ZN(
        n10399) );
  INV_X1 U12924 ( .A(n10377), .ZN(n10391) );
  NAND2_X1 U12925 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n11598) );
  INV_X1 U12926 ( .A(n11598), .ZN(n10378) );
  AOI21_X1 U12927 ( .B1(n13827), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n10378), .ZN(
        n10396) );
  INV_X1 U12928 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n13813) );
  INV_X1 U12929 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10742) );
  MUX2_X1 U12930 ( .A(n10742), .B(P1_REG2_REG_1__SCAN_IN), .S(n10379), .Z(
        n13784) );
  NAND3_X1 U12931 ( .A1(n13784), .A2(P1_REG2_REG_0__SCAN_IN), .A3(n14256), 
        .ZN(n13795) );
  INV_X1 U12932 ( .A(n10379), .ZN(n13779) );
  NAND2_X1 U12933 ( .A1(n13779), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n13794) );
  INV_X1 U12934 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10746) );
  MUX2_X1 U12935 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n10746), .S(n13789), .Z(
        n13796) );
  AOI21_X1 U12936 ( .B1(n13795), .B2(n13794), .A(n13796), .ZN(n13793) );
  NOR2_X1 U12937 ( .A1(n13789), .A2(n10746), .ZN(n13811) );
  MUX2_X1 U12938 ( .A(n13813), .B(P1_REG2_REG_3__SCAN_IN), .S(n13812), .Z(
        n10380) );
  OAI21_X1 U12939 ( .B1(n13793), .B2(n13811), .A(n10380), .ZN(n13818) );
  OAI21_X1 U12940 ( .B1(n13813), .B2(n13812), .A(n13818), .ZN(n12139) );
  MUX2_X1 U12941 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10381), .S(n10382), .Z(
        n12140) );
  AOI22_X1 U12942 ( .A1(n12139), .A2(n12140), .B1(n10382), .B2(
        P1_REG2_REG_4__SCAN_IN), .ZN(n10538) );
  INV_X1 U12943 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10383) );
  MUX2_X1 U12944 ( .A(n10383), .B(P1_REG2_REG_5__SCAN_IN), .S(n10384), .Z(
        n10537) );
  OR2_X1 U12945 ( .A1(n10538), .A2(n10537), .ZN(n10535) );
  NAND2_X1 U12946 ( .A1(n10384), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10416) );
  INV_X1 U12947 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10386) );
  MUX2_X1 U12948 ( .A(n10386), .B(P1_REG2_REG_6__SCAN_IN), .S(n10385), .Z(
        n10415) );
  AOI21_X1 U12949 ( .B1(n10535), .B2(n10416), .A(n10415), .ZN(n10418) );
  NOR2_X1 U12950 ( .A1(n10420), .A2(n10386), .ZN(n10393) );
  INV_X1 U12951 ( .A(n10393), .ZN(n10389) );
  INV_X1 U12952 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10387) );
  MUX2_X1 U12953 ( .A(n10387), .B(P1_REG2_REG_7__SCAN_IN), .S(n10429), .Z(
        n10388) );
  NAND2_X1 U12954 ( .A1(n10389), .A2(n10388), .ZN(n10394) );
  NOR2_X1 U12955 ( .A1(n6483), .A2(n14248), .ZN(n10390) );
  MUX2_X1 U12956 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10387), .S(n10429), .Z(
        n10392) );
  OAI21_X1 U12957 ( .B1(n10418), .B2(n10393), .A(n10392), .ZN(n10426) );
  OAI211_X1 U12958 ( .C1(n10418), .C2(n10394), .A(n13883), .B(n10426), .ZN(
        n10395) );
  OAI211_X1 U12959 ( .C1(n13806), .C2(n10397), .A(n10396), .B(n10395), .ZN(
        n10398) );
  OR2_X1 U12960 ( .A1(n10399), .A2(n10398), .ZN(P1_U3250) );
  INV_X1 U12961 ( .A(n10400), .ZN(n10403) );
  INV_X1 U12962 ( .A(n11212), .ZN(n11218) );
  OAI222_X1 U12963 ( .A1(n14245), .A2(n10401), .B1(n14251), .B2(n10403), .C1(
        P1_U3086), .C2(n11218), .ZN(P1_U3342) );
  INV_X1 U12964 ( .A(n14657), .ZN(n11036) );
  OAI222_X1 U12965 ( .A1(P2_U3088), .A2(n11036), .B1(n13596), .B2(n10403), 
        .C1(n10402), .C2(n13591), .ZN(P2_U3314) );
  NAND2_X1 U12966 ( .A1(n10404), .A2(n10600), .ZN(n12339) );
  INV_X1 U12967 ( .A(n12339), .ZN(n10405) );
  NOR2_X1 U12968 ( .A1(n15067), .A2(n10405), .ZN(n12508) );
  AOI22_X1 U12969 ( .A1(n10406), .A2(n12674), .B1(n12648), .B2(n10668), .ZN(
        n10409) );
  NAND2_X1 U12970 ( .A1(n10407), .A2(n13125), .ZN(n10529) );
  NAND2_X1 U12971 ( .A1(n10529), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10408) );
  OAI211_X1 U12972 ( .C1(n12508), .C2(n12650), .A(n10409), .B(n10408), .ZN(
        P3_U3172) );
  NAND2_X1 U12973 ( .A1(n13774), .A2(n13717), .ZN(n11187) );
  INV_X1 U12974 ( .A(n11187), .ZN(n10723) );
  AOI21_X1 U12975 ( .B1(n14521), .B2(n14534), .A(n11193), .ZN(n10410) );
  AOI211_X1 U12976 ( .C1(n9118), .C2(n10730), .A(n10723), .B(n10410), .ZN(
        n10566) );
  NAND2_X1 U12977 ( .A1(n14558), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10411) );
  OAI21_X1 U12978 ( .B1(n10566), .B2(n14558), .A(n10411), .ZN(P1_U3528) );
  AOI211_X1 U12979 ( .C1(n10414), .C2(n10413), .A(n13880), .B(n10412), .ZN(
        n10423) );
  AND3_X1 U12980 ( .A1(n10535), .A2(n10416), .A3(n10415), .ZN(n10417) );
  NOR3_X1 U12981 ( .A1(n14468), .A2(n10418), .A3(n10417), .ZN(n10422) );
  NAND2_X1 U12982 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n11423) );
  NAND2_X1 U12983 ( .A1(n13827), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n10419) );
  OAI211_X1 U12984 ( .C1(n13806), .C2(n10420), .A(n11423), .B(n10419), .ZN(
        n10421) );
  OR3_X1 U12985 ( .A1(n10423), .A2(n10422), .A3(n10421), .ZN(P1_U3249) );
  NAND2_X1 U12986 ( .A1(n10429), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10425) );
  INV_X1 U12987 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10553) );
  MUX2_X1 U12988 ( .A(n10553), .B(P1_REG2_REG_8__SCAN_IN), .S(n10549), .Z(
        n10424) );
  AOI21_X1 U12989 ( .B1(n10426), .B2(n10425), .A(n10424), .ZN(n13833) );
  NAND3_X1 U12990 ( .A1(n10426), .A2(n10425), .A3(n10424), .ZN(n10427) );
  NAND2_X1 U12991 ( .A1(n13883), .A2(n10427), .ZN(n10437) );
  INV_X1 U12992 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10430) );
  MUX2_X1 U12993 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10430), .S(n10549), .Z(
        n10431) );
  OAI21_X1 U12994 ( .B1(n10432), .B2(n10431), .A(n10548), .ZN(n10433) );
  NAND2_X1 U12995 ( .A1(n10433), .A2(n14462), .ZN(n10436) );
  AND2_X1 U12996 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n11561) );
  NOR2_X1 U12997 ( .A1(n13806), .A2(n10554), .ZN(n10434) );
  AOI211_X1 U12998 ( .C1(n13827), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n11561), .B(
        n10434), .ZN(n10435) );
  OAI211_X1 U12999 ( .C1(n13833), .C2(n10437), .A(n10436), .B(n10435), .ZN(
        P1_U3251) );
  INV_X1 U13000 ( .A(n10438), .ZN(n10439) );
  OAI222_X1 U13001 ( .A1(n12303), .A2(n10440), .B1(n13138), .B2(n10439), .C1(
        P3_U3151), .C2(n12798), .ZN(P3_U3278) );
  NAND2_X1 U13002 ( .A1(n10847), .A2(n10441), .ZN(n10442) );
  OR2_X1 U13003 ( .A1(n10442), .A2(n14740), .ZN(n10471) );
  AOI21_X1 U13004 ( .B1(n10471), .B2(n10844), .A(n10443), .ZN(n10485) );
  NAND2_X1 U13005 ( .A1(n10485), .A2(n10444), .ZN(n10445) );
  INV_X1 U13006 ( .A(n10446), .ZN(n11005) );
  INV_X1 U13007 ( .A(n10447), .ZN(n10448) );
  NAND2_X4 U13008 ( .A1(n10449), .A2(n10448), .ZN(n12209) );
  NAND2_X1 U13009 ( .A1(n13308), .A2(n6477), .ZN(n10453) );
  NAND2_X1 U13010 ( .A1(n13310), .A2(n12193), .ZN(n10450) );
  NAND2_X1 U13011 ( .A1(n10450), .A2(n14746), .ZN(n10486) );
  NAND2_X1 U13012 ( .A1(n12209), .A2(n14721), .ZN(n10451) );
  NAND2_X1 U13013 ( .A1(n10486), .A2(n10451), .ZN(n10618) );
  NAND2_X1 U13014 ( .A1(n10617), .A2(n10618), .ZN(n10456) );
  INV_X1 U13015 ( .A(n10452), .ZN(n10454) );
  NAND2_X1 U13016 ( .A1(n10454), .A2(n10453), .ZN(n10455) );
  NAND2_X1 U13017 ( .A1(n10456), .A2(n10455), .ZN(n10622) );
  XNOR2_X1 U13018 ( .A(n10981), .B(n12209), .ZN(n10457) );
  XNOR2_X1 U13019 ( .A(n10457), .B(n10459), .ZN(n10623) );
  NAND2_X1 U13020 ( .A1(n10622), .A2(n10623), .ZN(n10461) );
  INV_X1 U13021 ( .A(n10457), .ZN(n10458) );
  NAND2_X1 U13022 ( .A1(n10459), .A2(n10458), .ZN(n10460) );
  NAND2_X1 U13023 ( .A1(n10461), .A2(n10460), .ZN(n13160) );
  INV_X1 U13024 ( .A(n13160), .ZN(n10468) );
  XNOR2_X1 U13025 ( .A(n12209), .B(n14766), .ZN(n10464) );
  INV_X1 U13026 ( .A(n10464), .ZN(n10463) );
  AND2_X1 U13027 ( .A1(n13307), .A2(n12193), .ZN(n10465) );
  INV_X1 U13028 ( .A(n10465), .ZN(n10462) );
  NAND2_X1 U13029 ( .A1(n10463), .A2(n10462), .ZN(n10466) );
  NAND2_X1 U13030 ( .A1(n10465), .A2(n10464), .ZN(n10469) );
  NAND2_X1 U13031 ( .A1(n10466), .A2(n10469), .ZN(n13161) );
  XNOR2_X1 U13032 ( .A(n12209), .B(n11008), .ZN(n10630) );
  NAND2_X1 U13033 ( .A1(n13306), .A2(n12193), .ZN(n10631) );
  XNOR2_X1 U13034 ( .A(n10630), .B(n10631), .ZN(n10470) );
  OAI21_X1 U13035 ( .B1(n6610), .B2(n10470), .A(n10636), .ZN(n10474) );
  NOR2_X1 U13036 ( .A1(n10471), .A2(n14743), .ZN(n10479) );
  INV_X1 U13037 ( .A(n10479), .ZN(n10476) );
  INV_X1 U13038 ( .A(n13267), .ZN(n13241) );
  NAND2_X1 U13039 ( .A1(n10474), .A2(n13241), .ZN(n10484) );
  OR2_X1 U13040 ( .A1(n10476), .A2(n10475), .ZN(n10477) );
  NAND2_X1 U13041 ( .A1(n13305), .A2(n13172), .ZN(n10481) );
  NAND2_X1 U13042 ( .A1(n13307), .A2(n13171), .ZN(n10480) );
  AND2_X1 U13043 ( .A1(n10481), .A2(n10480), .ZN(n11002) );
  NAND2_X1 U13044 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n14575) );
  OAI21_X1 U13045 ( .B1(n13272), .B2(n11002), .A(n14575), .ZN(n10482) );
  AOI21_X1 U13046 ( .B1(n11008), .B2(n13262), .A(n10482), .ZN(n10483) );
  OAI211_X1 U13047 ( .C1(n13259), .C2(n11005), .A(n10484), .B(n10483), .ZN(
        P2_U3202) );
  NAND2_X1 U13048 ( .A1(n13308), .A2(n13172), .ZN(n14727) );
  NAND2_X1 U13049 ( .A1(n10485), .A2(n14741), .ZN(n10627) );
  AOI22_X1 U13050 ( .A1(n13262), .A2(n14746), .B1(n10627), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n10490) );
  OAI21_X1 U13051 ( .B1(n10487), .B2(n11440), .A(n10486), .ZN(n10488) );
  NAND2_X1 U13052 ( .A1(n13241), .A2(n10488), .ZN(n10489) );
  OAI211_X1 U13053 ( .C1(n14727), .C2(n13272), .A(n10490), .B(n10489), .ZN(
        P2_U3204) );
  XOR2_X1 U13054 ( .A(n10491), .B(n10492), .Z(n10497) );
  AOI22_X1 U13055 ( .A1(n10406), .A2(n12663), .B1(n10493), .B2(n12648), .ZN(
        n10494) );
  OAI21_X1 U13056 ( .B1(n15041), .B2(n12665), .A(n10494), .ZN(n10495) );
  AOI21_X1 U13057 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n10529), .A(n10495), .ZN(
        n10496) );
  OAI21_X1 U13058 ( .B1(n10497), .B2(n12650), .A(n10496), .ZN(P3_U3177) );
  AOI21_X1 U13059 ( .B1(n10614), .B2(n10499), .A(n10498), .ZN(n10512) );
  OAI21_X1 U13060 ( .B1(n10501), .B2(P3_REG1_REG_1__SCAN_IN), .A(n10500), .ZN(
        n10508) );
  OAI22_X1 U13061 ( .A1(n15000), .A2(n6753), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10502), .ZN(n10507) );
  AOI21_X1 U13062 ( .B1(n10504), .B2(n10326), .A(n10503), .ZN(n10505) );
  NOR2_X1 U13063 ( .A1(n14991), .A2(n10505), .ZN(n10506) );
  AOI211_X1 U13064 ( .C1(n6467), .C2(n10508), .A(n10507), .B(n10506), .ZN(
        n10511) );
  NAND2_X1 U13065 ( .A1(n14996), .A2(n10509), .ZN(n10510) );
  OAI211_X1 U13066 ( .C1(n10512), .C2(n14985), .A(n10511), .B(n10510), .ZN(
        P3_U3183) );
  AOI21_X1 U13067 ( .B1(n15045), .B2(n10513), .A(n12508), .ZN(n10514) );
  AOI21_X1 U13068 ( .B1(n15063), .B2(n10406), .A(n10514), .ZN(n10670) );
  OAI22_X1 U13069 ( .A1(n13063), .A2(n10600), .B1(n15131), .B2(n10328), .ZN(
        n10515) );
  INV_X1 U13070 ( .A(n10515), .ZN(n10516) );
  OAI21_X1 U13071 ( .B1(n10670), .B2(n9450), .A(n10516), .ZN(P3_U3459) );
  INV_X1 U13072 ( .A(n15059), .ZN(n10526) );
  MUX2_X1 U13073 ( .A(n12348), .B(n15043), .S(n10519), .Z(n10518) );
  NAND3_X1 U13074 ( .A1(n10406), .A2(n10519), .A3(n15072), .ZN(n10517) );
  NAND2_X1 U13075 ( .A1(n10518), .A2(n10517), .ZN(n10525) );
  INV_X1 U13076 ( .A(n15068), .ZN(n10520) );
  NOR3_X1 U13077 ( .A1(n10520), .A2(n15067), .A3(n10519), .ZN(n10524) );
  AOI211_X1 U13078 ( .C1(n10522), .C2(n10521), .A(n10526), .B(n10525), .ZN(
        n10523) );
  AOI211_X1 U13079 ( .C1(n10526), .C2(n10525), .A(n10524), .B(n10523), .ZN(
        n10531) );
  AOI22_X1 U13080 ( .A1(n12663), .A2(n10404), .B1(n12648), .B2(n15072), .ZN(
        n10527) );
  OAI21_X1 U13081 ( .B1(n10914), .B2(n12665), .A(n10527), .ZN(n10528) );
  AOI21_X1 U13082 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(n10529), .A(n10528), .ZN(
        n10530) );
  OAI21_X1 U13083 ( .B1(n10531), .B2(n12650), .A(n10530), .ZN(P3_U3162) );
  OAI21_X1 U13084 ( .B1(n10534), .B2(n10533), .A(n10532), .ZN(n10540) );
  INV_X1 U13085 ( .A(n10535), .ZN(n10536) );
  AOI211_X1 U13086 ( .C1(n10538), .C2(n10537), .A(n10536), .B(n14468), .ZN(
        n10539) );
  AOI21_X1 U13087 ( .B1(n14462), .B2(n10540), .A(n10539), .ZN(n10543) );
  NAND2_X1 U13088 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n11080) );
  INV_X1 U13089 ( .A(n11080), .ZN(n10541) );
  AOI21_X1 U13090 ( .B1(n13827), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n10541), .ZN(
        n10542) );
  OAI211_X1 U13091 ( .C1(n10544), .C2(n13806), .A(n10543), .B(n10542), .ZN(
        P1_U3248) );
  INV_X1 U13092 ( .A(n12824), .ZN(n12814) );
  OAI222_X1 U13093 ( .A1(P3_U3151), .A2(n12814), .B1(n12303), .B2(n10546), 
        .C1(n13138), .C2(n10545), .ZN(P3_U3277) );
  INV_X1 U13094 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10547) );
  MUX2_X1 U13095 ( .A(n10547), .B(P1_REG1_REG_10__SCAN_IN), .S(n10677), .Z(
        n10552) );
  OAI21_X1 U13096 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n10549), .A(n10548), .ZN(
        n13823) );
  INV_X1 U13097 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10550) );
  MUX2_X1 U13098 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10550), .S(n13834), .Z(
        n13824) );
  NAND2_X1 U13099 ( .A1(n13823), .A2(n13824), .ZN(n13822) );
  OAI21_X1 U13100 ( .B1(n13834), .B2(P1_REG1_REG_9__SCAN_IN), .A(n13822), .ZN(
        n10551) );
  NOR2_X1 U13101 ( .A1(n10551), .A2(n10552), .ZN(n10676) );
  AOI211_X1 U13102 ( .C1(n10552), .C2(n10551), .A(n13880), .B(n10676), .ZN(
        n10565) );
  NOR2_X1 U13103 ( .A1(n10554), .A2(n10553), .ZN(n13828) );
  INV_X1 U13104 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n11055) );
  MUX2_X1 U13105 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n11055), .S(n13834), .Z(
        n10555) );
  OAI21_X1 U13106 ( .B1(n13833), .B2(n13828), .A(n10555), .ZN(n13831) );
  NAND2_X1 U13107 ( .A1(n13834), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10558) );
  INV_X1 U13108 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10556) );
  MUX2_X1 U13109 ( .A(n10556), .B(P1_REG2_REG_10__SCAN_IN), .S(n10677), .Z(
        n10557) );
  AOI21_X1 U13110 ( .B1(n13831), .B2(n10558), .A(n10557), .ZN(n10675) );
  AND3_X1 U13111 ( .A1(n13831), .A2(n10558), .A3(n10557), .ZN(n10559) );
  NOR3_X1 U13112 ( .A1(n10675), .A2(n10559), .A3(n14468), .ZN(n10564) );
  AND2_X1 U13113 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10560) );
  AOI21_X1 U13114 ( .B1(n13827), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n10560), 
        .ZN(n10561) );
  OAI21_X1 U13115 ( .B1(n13806), .B2(n10562), .A(n10561), .ZN(n10563) );
  OR3_X1 U13116 ( .A1(n10565), .A2(n10564), .A3(n10563), .ZN(P1_U3253) );
  INV_X1 U13117 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10568) );
  OR2_X1 U13118 ( .A1(n10566), .A2(n14547), .ZN(n10567) );
  OAI21_X1 U13119 ( .B1(n14549), .B2(n10568), .A(n10567), .ZN(P1_U3459) );
  INV_X1 U13120 ( .A(n12236), .ZN(n14671) );
  INV_X1 U13121 ( .A(n10569), .ZN(n10572) );
  OAI222_X1 U13122 ( .A1(P2_U3088), .A2(n14671), .B1(n13596), .B2(n10572), 
        .C1(n10570), .C2(n13591), .ZN(P2_U3311) );
  INV_X1 U13123 ( .A(n13847), .ZN(n10573) );
  OAI222_X1 U13124 ( .A1(P1_U3086), .A2(n10573), .B1(n14251), .B2(n10572), 
        .C1(n10571), .C2(n14245), .ZN(P1_U3339) );
  AOI21_X1 U13125 ( .B1(n10585), .B2(P2_REG2_REG_8__SCAN_IN), .A(n10574), .ZN(
        n14612) );
  INV_X1 U13126 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10575) );
  MUX2_X1 U13127 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n10575), .S(n14614), .Z(
        n14611) );
  NAND2_X1 U13128 ( .A1(n14612), .A2(n14611), .ZN(n14610) );
  OAI21_X1 U13129 ( .B1(n14614), .B2(P2_REG2_REG_9__SCAN_IN), .A(n14610), .ZN(
        n14627) );
  INV_X1 U13130 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10576) );
  MUX2_X1 U13131 ( .A(n10576), .B(P2_REG2_REG_10__SCAN_IN), .S(n10588), .Z(
        n14628) );
  NOR2_X1 U13132 ( .A1(n14627), .A2(n14628), .ZN(n14626) );
  AOI21_X1 U13133 ( .B1(n10588), .B2(P2_REG2_REG_10__SCAN_IN), .A(n14626), 
        .ZN(n10579) );
  INV_X1 U13134 ( .A(n10579), .ZN(n10581) );
  INV_X1 U13135 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10577) );
  MUX2_X1 U13136 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n10577), .S(n11034), .Z(
        n10578) );
  INV_X1 U13137 ( .A(n10578), .ZN(n10580) );
  AOI21_X1 U13138 ( .B1(n10581), .B2(n10580), .A(n14639), .ZN(n10595) );
  AND2_X1 U13139 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n11377) );
  NOR2_X1 U13140 ( .A1(n14620), .A2(n10582), .ZN(n10583) );
  AOI211_X1 U13141 ( .C1(n14684), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n11377), 
        .B(n10583), .ZN(n10594) );
  INV_X1 U13142 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n14847) );
  AOI21_X1 U13143 ( .B1(n10585), .B2(P2_REG1_REG_8__SCAN_IN), .A(n10584), .ZN(
        n14609) );
  MUX2_X1 U13144 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n14847), .S(n14614), .Z(
        n14608) );
  AND2_X1 U13145 ( .A1(n14609), .A2(n14608), .ZN(n14606) );
  INV_X1 U13146 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10587) );
  MUX2_X1 U13147 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n10587), .S(n10588), .Z(
        n14624) );
  NAND2_X1 U13148 ( .A1(n14625), .A2(n14624), .ZN(n14623) );
  NAND2_X1 U13149 ( .A1(n10588), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10590) );
  INV_X1 U13150 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n14851) );
  MUX2_X1 U13151 ( .A(n14851), .B(P2_REG1_REG_11__SCAN_IN), .S(n11034), .Z(
        n10589) );
  AOI21_X1 U13152 ( .B1(n14623), .B2(n10590), .A(n10589), .ZN(n11033) );
  INV_X1 U13153 ( .A(n11033), .ZN(n10592) );
  NAND3_X1 U13154 ( .A1(n14623), .A2(n10590), .A3(n10589), .ZN(n10591) );
  NAND3_X1 U13155 ( .A1(n10592), .A2(n14688), .A3(n10591), .ZN(n10593) );
  OAI211_X1 U13156 ( .C1(n10595), .C2(n14652), .A(n10594), .B(n10593), .ZN(
        P2_U3225) );
  INV_X1 U13157 ( .A(n11695), .ZN(n11704) );
  INV_X1 U13158 ( .A(n10596), .ZN(n10598) );
  OAI222_X1 U13159 ( .A1(P1_U3086), .A2(n11704), .B1(n14251), .B2(n10598), 
        .C1(n10597), .C2(n14245), .ZN(P1_U3341) );
  INV_X1 U13160 ( .A(n12226), .ZN(n12239) );
  OAI222_X1 U13161 ( .A1(n13591), .A2(n10599), .B1(n13596), .B2(n10598), .C1(
        n12239), .C2(P2_U3088), .ZN(P2_U3313) );
  INV_X1 U13162 ( .A(n15120), .ZN(n15121) );
  OAI22_X1 U13163 ( .A1(n13121), .A2(n10600), .B1(n15120), .B2(n7532), .ZN(
        n10601) );
  INV_X1 U13164 ( .A(n10601), .ZN(n10602) );
  OAI21_X1 U13165 ( .B1(n10670), .B2(n15121), .A(n10602), .ZN(P3_U3390) );
  NOR3_X1 U13166 ( .A1(n14300), .A2(n6467), .A3(n14962), .ZN(n10615) );
  INV_X1 U13167 ( .A(n10603), .ZN(n10605) );
  INV_X1 U13168 ( .A(n13142), .ZN(n10604) );
  NAND3_X1 U13169 ( .A1(n14962), .A2(n10605), .A3(n10604), .ZN(n10606) );
  OAI21_X1 U13170 ( .B1(P3_STATE_REG_SCAN_IN), .B2(n10666), .A(n10606), .ZN(
        n10611) );
  AOI22_X1 U13171 ( .A1(n14300), .A2(n10608), .B1(n6467), .B2(n10607), .ZN(
        n10609) );
  INV_X1 U13172 ( .A(n10609), .ZN(n10610) );
  AOI211_X1 U13173 ( .C1(n14969), .C2(P3_ADDR_REG_0__SCAN_IN), .A(n10611), .B(
        n10610), .ZN(n10613) );
  NAND2_X1 U13174 ( .A1(n14996), .A2(n13142), .ZN(n10612) );
  OAI211_X1 U13175 ( .C1(n10615), .C2(n10614), .A(n10613), .B(n10612), .ZN(
        P3_U3182) );
  INV_X1 U13176 ( .A(n13262), .ZN(n13278) );
  OAI22_X1 U13177 ( .A1(n10616), .A2(n13254), .B1(n10866), .B2(n13256), .ZN(
        n11174) );
  AOI22_X1 U13178 ( .A1(n13257), .A2(n11174), .B1(n10627), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n10621) );
  XNOR2_X1 U13179 ( .A(n10617), .B(n10618), .ZN(n10619) );
  NAND2_X1 U13180 ( .A1(n10619), .A2(n13241), .ZN(n10620) );
  OAI211_X1 U13181 ( .C1(n14755), .C2(n13278), .A(n10621), .B(n10620), .ZN(
        P2_U3194) );
  XNOR2_X1 U13182 ( .A(n10623), .B(n10622), .ZN(n10624) );
  NAND2_X1 U13183 ( .A1(n10624), .A2(n13241), .ZN(n10629) );
  NAND2_X1 U13184 ( .A1(n13307), .A2(n13172), .ZN(n10626) );
  NAND2_X1 U13185 ( .A1(n13308), .A2(n13171), .ZN(n10625) );
  NAND2_X1 U13186 ( .A1(n10626), .A2(n10625), .ZN(n10972) );
  AOI22_X1 U13187 ( .A1(n13257), .A2(n10972), .B1(n10627), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n10628) );
  OAI211_X1 U13188 ( .C1(n14759), .C2(n13278), .A(n10629), .B(n10628), .ZN(
        P2_U3209) );
  INV_X1 U13189 ( .A(n10636), .ZN(n10634) );
  INV_X1 U13190 ( .A(n10630), .ZN(n10632) );
  NAND2_X1 U13191 ( .A1(n10632), .A2(n10631), .ZN(n10635) );
  INV_X1 U13192 ( .A(n10635), .ZN(n10633) );
  XNOR2_X1 U13193 ( .A(n11129), .B(n12209), .ZN(n10769) );
  NAND2_X1 U13194 ( .A1(n13305), .A2(n12193), .ZN(n10770) );
  XNOR2_X1 U13195 ( .A(n10769), .B(n10770), .ZN(n10637) );
  NOR3_X1 U13196 ( .A1(n10634), .A2(n10633), .A3(n10637), .ZN(n10640) );
  NAND2_X1 U13197 ( .A1(n10638), .A2(n10637), .ZN(n10773) );
  INV_X1 U13198 ( .A(n10773), .ZN(n10639) );
  OAI21_X1 U13199 ( .B1(n10640), .B2(n10639), .A(n13241), .ZN(n10645) );
  INV_X1 U13200 ( .A(n13259), .ZN(n13274) );
  NAND2_X1 U13201 ( .A1(n13304), .A2(n13172), .ZN(n10642) );
  NAND2_X1 U13202 ( .A1(n13306), .A2(n13171), .ZN(n10641) );
  AND2_X1 U13203 ( .A1(n10642), .A2(n10641), .ZN(n11135) );
  NAND2_X1 U13204 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n14590) );
  OAI21_X1 U13205 ( .B1(n13272), .B2(n11135), .A(n14590), .ZN(n10643) );
  AOI21_X1 U13206 ( .B1(n11128), .B2(n13274), .A(n10643), .ZN(n10644) );
  OAI211_X1 U13207 ( .C1(n14783), .C2(n13278), .A(n10645), .B(n10644), .ZN(
        P2_U3199) );
  XNOR2_X1 U13208 ( .A(n10646), .B(n10647), .ZN(n10648) );
  NAND2_X1 U13209 ( .A1(n10648), .A2(n14409), .ZN(n10654) );
  NAND2_X1 U13210 ( .A1(n13774), .A2(n13913), .ZN(n10650) );
  NAND2_X1 U13211 ( .A1(n13772), .A2(n13717), .ZN(n10649) );
  NAND2_X1 U13212 ( .A1(n10650), .A2(n10649), .ZN(n14500) );
  NAND2_X1 U13213 ( .A1(n10652), .A2(n10651), .ZN(n10722) );
  AOI22_X1 U13214 ( .A1(n14411), .A2(n14500), .B1(n10722), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n10653) );
  OAI211_X1 U13215 ( .C1(n14503), .C2(n13745), .A(n10654), .B(n10653), .ZN(
        P1_U3237) );
  INV_X1 U13216 ( .A(n14662), .ZN(n12241) );
  INV_X1 U13217 ( .A(n10655), .ZN(n10658) );
  OAI222_X1 U13218 ( .A1(P2_U3088), .A2(n12241), .B1(n13596), .B2(n10658), 
        .C1(n10656), .C2(n13591), .ZN(P2_U3312) );
  INV_X1 U13219 ( .A(n14464), .ZN(n11697) );
  OAI222_X1 U13220 ( .A1(P1_U3086), .A2(n11697), .B1(n14251), .B2(n10658), 
        .C1(n10657), .C2(n14245), .ZN(P1_U3340) );
  INV_X1 U13221 ( .A(n10659), .ZN(n13123) );
  NAND2_X1 U13222 ( .A1(n13123), .A2(n10660), .ZN(n10661) );
  OAI22_X1 U13223 ( .A1(n15080), .A2(n10329), .B1(n10666), .B2(n15009), .ZN(
        n10667) );
  AOI21_X1 U13224 ( .B1(n15004), .B2(n10668), .A(n10667), .ZN(n10669) );
  OAI21_X1 U13225 ( .B1(n10670), .B2(n15082), .A(n10669), .ZN(P3_U3233) );
  INV_X1 U13226 ( .A(n10671), .ZN(n10674) );
  INV_X1 U13227 ( .A(n14686), .ZN(n12245) );
  OAI222_X1 U13228 ( .A1(n13591), .A2(n10672), .B1(n13589), .B2(n10674), .C1(
        n12245), .C2(P2_U3088), .ZN(P2_U3310) );
  INV_X1 U13229 ( .A(n13855), .ZN(n13862) );
  OAI222_X1 U13230 ( .A1(P1_U3086), .A2(n13862), .B1(n14251), .B2(n10674), 
        .C1(n10673), .C2(n14245), .ZN(P1_U3338) );
  AOI21_X1 U13231 ( .B1(n10677), .B2(P1_REG2_REG_10__SCAN_IN), .A(n10675), 
        .ZN(n10811) );
  MUX2_X1 U13232 ( .A(n11299), .B(P1_REG2_REG_11__SCAN_IN), .S(n10817), .Z(
        n10810) );
  XNOR2_X1 U13233 ( .A(n10811), .B(n10810), .ZN(n10687) );
  MUX2_X1 U13234 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10678), .S(n10817), .Z(
        n10679) );
  OAI21_X1 U13235 ( .B1(n10680), .B2(n10679), .A(n10816), .ZN(n10681) );
  NAND2_X1 U13236 ( .A1(n10681), .A2(n14462), .ZN(n10686) );
  NAND2_X1 U13237 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14414)
         );
  INV_X1 U13238 ( .A(n14414), .ZN(n10684) );
  NOR2_X1 U13239 ( .A1(n13806), .A2(n10682), .ZN(n10683) );
  AOI211_X1 U13240 ( .C1(n13827), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n10684), 
        .B(n10683), .ZN(n10685) );
  OAI211_X1 U13241 ( .C1(n14468), .C2(n10687), .A(n10686), .B(n10685), .ZN(
        P1_U3254) );
  OAI222_X1 U13242 ( .A1(n12303), .A2(n10689), .B1(P3_U3151), .B2(n12818), 
        .C1(n13138), .C2(n10688), .ZN(P3_U3276) );
  AOI21_X1 U13243 ( .B1(n10692), .B2(n10690), .A(n10691), .ZN(n10698) );
  INV_X1 U13244 ( .A(n10722), .ZN(n10695) );
  INV_X1 U13245 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n13777) );
  NOR2_X1 U13246 ( .A1(n10693), .A2(n13633), .ZN(n10740) );
  AOI21_X1 U13247 ( .B1(n13913), .B2(n13776), .A(n10740), .ZN(n10694) );
  OAI22_X1 U13248 ( .A1(n10695), .A2(n13777), .B1(n10694), .B2(n13739), .ZN(
        n10696) );
  AOI21_X1 U13249 ( .B1(n10085), .B2(n6468), .A(n10696), .ZN(n10697) );
  OAI21_X1 U13250 ( .B1(n10698), .B2(n13731), .A(n10697), .ZN(P1_U3222) );
  XNOR2_X1 U13251 ( .A(n7350), .B(n10699), .ZN(n14510) );
  INV_X1 U13252 ( .A(n14510), .ZN(n10717) );
  NAND2_X1 U13253 ( .A1(n10701), .A2(n10700), .ZN(n13912) );
  NAND2_X1 U13254 ( .A1(n10747), .A2(n10714), .ZN(n10703) );
  NAND2_X1 U13255 ( .A1(n10703), .A2(n14493), .ZN(n10704) );
  NOR2_X1 U13256 ( .A1(n10799), .A2(n10704), .ZN(n14511) );
  INV_X1 U13257 ( .A(n10726), .ZN(n14546) );
  NAND2_X1 U13258 ( .A1(n14510), .A2(n14546), .ZN(n10711) );
  OAI21_X1 U13259 ( .B1(n10707), .B2(n10706), .A(n10705), .ZN(n10709) );
  AOI21_X1 U13260 ( .B1(n10709), .B2(n14526), .A(n10708), .ZN(n10710) );
  NAND2_X1 U13261 ( .A1(n10711), .A2(n10710), .ZN(n14516) );
  AOI21_X1 U13262 ( .B1(n14511), .B2(n11860), .A(n14516), .ZN(n10712) );
  MUX2_X1 U13263 ( .A(n13813), .B(n10712), .S(n14080), .Z(n10716) );
  INV_X1 U13264 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n13805) );
  INV_X1 U13265 ( .A(n14477), .ZN(n14034) );
  AOI22_X1 U13266 ( .A1(n14082), .A2(n10714), .B1(n13805), .B2(n14034), .ZN(
        n10715) );
  OAI211_X1 U13267 ( .C1(n10717), .C2(n11414), .A(n10716), .B(n10715), .ZN(
        P1_U3290) );
  AND2_X1 U13268 ( .A1(n10719), .A2(n10718), .ZN(n10720) );
  NOR2_X1 U13269 ( .A1(n10721), .A2(n10720), .ZN(n12150) );
  AOI22_X1 U13270 ( .A1(n14411), .A2(n10723), .B1(n10722), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n10725) );
  NAND2_X1 U13271 ( .A1(n6468), .A2(n10730), .ZN(n10724) );
  OAI211_X1 U13272 ( .C1(n12150), .C2(n13731), .A(n10725), .B(n10724), .ZN(
        P1_U3232) );
  OR2_X1 U13273 ( .A1(n14491), .A2(n10726), .ZN(n10727) );
  XOR2_X1 U13274 ( .A(n10728), .B(n10734), .Z(n14497) );
  INV_X1 U13275 ( .A(n13912), .ZN(n10729) );
  NAND2_X1 U13276 ( .A1(n14485), .A2(n14493), .ZN(n13956) );
  INV_X1 U13277 ( .A(n10748), .ZN(n10732) );
  NAND2_X1 U13278 ( .A1(n10085), .A2(n10730), .ZN(n10731) );
  NAND2_X1 U13279 ( .A1(n10732), .A2(n10731), .ZN(n10736) );
  OAI22_X1 U13280 ( .A1(n13956), .A2(n10736), .B1(n13777), .B2(n14477), .ZN(
        n10733) );
  AOI21_X1 U13281 ( .B1(n14082), .B2(n10085), .A(n10733), .ZN(n10744) );
  INV_X1 U13282 ( .A(n13776), .ZN(n10735) );
  OAI21_X1 U13283 ( .B1(n6685), .B2(n10735), .A(n14526), .ZN(n10739) );
  INV_X1 U13284 ( .A(n10736), .ZN(n14494) );
  XOR2_X1 U13285 ( .A(n13774), .B(n14494), .Z(n10737) );
  AOI21_X1 U13286 ( .B1(n10737), .B2(n14526), .A(n13776), .ZN(n10738) );
  AOI21_X1 U13287 ( .B1(n13624), .B2(n10739), .A(n10738), .ZN(n10741) );
  NOR2_X1 U13288 ( .A1(n10741), .A2(n10740), .ZN(n14496) );
  MUX2_X1 U13289 ( .A(n10742), .B(n14496), .S(n14080), .Z(n10743) );
  OAI211_X1 U13290 ( .C1(n14073), .C2(n14497), .A(n10744), .B(n10743), .ZN(
        P1_U3292) );
  XNOR2_X1 U13291 ( .A(n10752), .B(n10745), .ZN(n14507) );
  NOR2_X1 U13292 ( .A1(n14080), .A2(n10746), .ZN(n10750) );
  OAI211_X1 U13293 ( .C1(n10748), .C2(n14503), .A(n14493), .B(n10747), .ZN(
        n14501) );
  OAI22_X1 U13294 ( .A1(n14085), .A2(n14501), .B1(n13790), .B2(n14477), .ZN(
        n10749) );
  AOI211_X1 U13295 ( .C1(n14080), .C2(n14500), .A(n10750), .B(n10749), .ZN(
        n10755) );
  OR2_X1 U13296 ( .A1(n14491), .A2(n14534), .ZN(n14042) );
  INV_X1 U13297 ( .A(n14042), .ZN(n14071) );
  OAI21_X1 U13298 ( .B1(n10753), .B2(n10752), .A(n10751), .ZN(n14505) );
  AOI22_X1 U13299 ( .A1(n14071), .A2(n14505), .B1(n14082), .B2(n7066), .ZN(
        n10754) );
  OAI211_X1 U13300 ( .C1(n14073), .C2(n14507), .A(n10755), .B(n10754), .ZN(
        P1_U3291) );
  XNOR2_X1 U13301 ( .A(n10756), .B(n10758), .ZN(n14535) );
  OAI21_X1 U13302 ( .B1(n10759), .B2(n10758), .A(n10757), .ZN(n14545) );
  NAND2_X1 U13303 ( .A1(n14545), .A2(n14092), .ZN(n10768) );
  AOI21_X1 U13304 ( .B1(n11992), .B2(n14537), .A(n14119), .ZN(n10760) );
  NAND2_X1 U13305 ( .A1(n10760), .A2(n11197), .ZN(n14539) );
  NOR2_X1 U13306 ( .A1(n14085), .A2(n14539), .ZN(n10766) );
  NAND2_X1 U13307 ( .A1(n13768), .A2(n13717), .ZN(n10762) );
  NAND2_X1 U13308 ( .A1(n13770), .A2(n13913), .ZN(n10761) );
  NAND2_X1 U13309 ( .A1(n10762), .A2(n10761), .ZN(n14536) );
  INV_X1 U13310 ( .A(n14536), .ZN(n10763) );
  MUX2_X1 U13311 ( .A(n10763), .B(n10386), .S(n14491), .Z(n10764) );
  OAI21_X1 U13312 ( .B1(n14477), .B2(n11424), .A(n10764), .ZN(n10765) );
  AOI211_X1 U13313 ( .C1(n14082), .C2(n14537), .A(n10766), .B(n10765), .ZN(
        n10767) );
  OAI211_X1 U13314 ( .C1(n14535), .C2(n14042), .A(n10768), .B(n10767), .ZN(
        P1_U3287) );
  INV_X1 U13315 ( .A(n10769), .ZN(n10771) );
  NAND2_X1 U13316 ( .A1(n10771), .A2(n10770), .ZN(n10772) );
  NAND2_X1 U13317 ( .A1(n10773), .A2(n10772), .ZN(n10907) );
  XNOR2_X1 U13318 ( .A(n10911), .B(n12209), .ZN(n10774) );
  AND2_X1 U13319 ( .A1(n13304), .A2(n12193), .ZN(n10775) );
  NAND2_X1 U13320 ( .A1(n10774), .A2(n10775), .ZN(n10779) );
  INV_X1 U13321 ( .A(n10774), .ZN(n10777) );
  INV_X1 U13322 ( .A(n10775), .ZN(n10776) );
  NAND2_X1 U13323 ( .A1(n10777), .A2(n10776), .ZN(n10778) );
  NAND2_X1 U13324 ( .A1(n10779), .A2(n10778), .ZN(n10908) );
  XNOR2_X1 U13325 ( .A(n14789), .B(n12209), .ZN(n10930) );
  INV_X1 U13326 ( .A(n12193), .ZN(n11457) );
  NAND2_X1 U13327 ( .A1(n13303), .A2(n12193), .ZN(n10928) );
  XNOR2_X1 U13328 ( .A(n10930), .B(n10928), .ZN(n10780) );
  OAI211_X1 U13329 ( .C1(n10781), .C2(n10780), .A(n10932), .B(n13241), .ZN(
        n10789) );
  INV_X1 U13330 ( .A(n10782), .ZN(n10883) );
  NAND2_X1 U13331 ( .A1(n13302), .A2(n13172), .ZN(n10784) );
  NAND2_X1 U13332 ( .A1(n13304), .A2(n13171), .ZN(n10783) );
  NAND2_X1 U13333 ( .A1(n10784), .A2(n10783), .ZN(n10880) );
  NAND2_X1 U13334 ( .A1(n13257), .A2(n10880), .ZN(n10785) );
  OAI211_X1 U13335 ( .C1(n13259), .C2(n10883), .A(n10786), .B(n10785), .ZN(
        n10787) );
  AOI21_X1 U13336 ( .B1(n14789), .B2(n13262), .A(n10787), .ZN(n10788) );
  NAND2_X1 U13337 ( .A1(n10789), .A2(n10788), .ZN(P2_U3185) );
  INV_X1 U13338 ( .A(n12678), .ZN(n11500) );
  AOI211_X1 U13339 ( .C1(n10792), .C2(n10791), .A(n12650), .B(n10790), .ZN(
        n10793) );
  INV_X1 U13340 ( .A(n10793), .ZN(n10797) );
  NOR2_X1 U13341 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10920), .ZN(n14863) );
  OAI22_X1 U13342 ( .A1(n10914), .A2(n12676), .B1(n15017), .B2(n12665), .ZN(
        n10794) );
  AOI211_X1 U13343 ( .C1(n12648), .C2(n10795), .A(n14863), .B(n10794), .ZN(
        n10796) );
  OAI211_X1 U13344 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n11500), .A(n10797), .B(
        n10796), .ZN(P3_U3158) );
  XNOR2_X1 U13345 ( .A(n10798), .B(n10806), .ZN(n14522) );
  OAI211_X1 U13346 ( .C1(n10799), .C2(n14520), .A(n14493), .B(n11991), .ZN(
        n14519) );
  INV_X1 U13347 ( .A(n14519), .ZN(n10805) );
  NAND2_X1 U13348 ( .A1(n13770), .A2(n13717), .ZN(n10801) );
  NAND2_X1 U13349 ( .A1(n13772), .A2(n13913), .ZN(n10800) );
  AND2_X1 U13350 ( .A1(n10801), .A2(n10800), .ZN(n14518) );
  INV_X1 U13351 ( .A(n14518), .ZN(n10802) );
  MUX2_X1 U13352 ( .A(n10802), .B(P1_REG2_REG_4__SCAN_IN), .S(n14491), .Z(
        n10804) );
  OAI22_X1 U13353 ( .A1(n14482), .A2(n14520), .B1(n11123), .B2(n14477), .ZN(
        n10803) );
  AOI211_X1 U13354 ( .C1(n10805), .C2(n14485), .A(n10804), .B(n10803), .ZN(
        n10809) );
  XNOR2_X1 U13355 ( .A(n10807), .B(n10806), .ZN(n14525) );
  NAND2_X1 U13356 ( .A1(n14525), .A2(n14071), .ZN(n10808) );
  OAI211_X1 U13357 ( .C1(n14073), .C2(n14522), .A(n10809), .B(n10808), .ZN(
        P1_U3289) );
  AOI22_X1 U13358 ( .A1(n11021), .A2(n11416), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n10821), .ZN(n10815) );
  NAND2_X1 U13359 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n10817), .ZN(n10813) );
  OR2_X1 U13360 ( .A1(n10811), .A2(n10810), .ZN(n10812) );
  NAND2_X1 U13361 ( .A1(n10813), .A2(n10812), .ZN(n10814) );
  NOR2_X1 U13362 ( .A1(n10815), .A2(n10814), .ZN(n11023) );
  AOI21_X1 U13363 ( .B1(n10815), .B2(n10814), .A(n11023), .ZN(n10825) );
  AOI22_X1 U13364 ( .A1(n11021), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n8864), 
        .B2(n10821), .ZN(n10819) );
  OAI21_X1 U13365 ( .B1(n10819), .B2(n10818), .A(n11015), .ZN(n10823) );
  NAND2_X1 U13366 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n13646)
         );
  NAND2_X1 U13367 ( .A1(n13827), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n10820) );
  OAI211_X1 U13368 ( .C1(n13806), .C2(n10821), .A(n13646), .B(n10820), .ZN(
        n10822) );
  AOI21_X1 U13369 ( .B1(n10823), .B2(n14462), .A(n10822), .ZN(n10824) );
  OAI21_X1 U13370 ( .B1(n10825), .B2(n14468), .A(n10824), .ZN(P1_U3255) );
  XNOR2_X1 U13371 ( .A(n10827), .B(n10826), .ZN(n10837) );
  INV_X1 U13372 ( .A(n10837), .ZN(n10853) );
  INV_X1 U13373 ( .A(n10828), .ZN(n14732) );
  NAND2_X1 U13374 ( .A1(n14733), .A2(n14732), .ZN(n10976) );
  INV_X1 U13375 ( .A(n10449), .ZN(n14801) );
  NAND2_X1 U13376 ( .A1(n13303), .A2(n13172), .ZN(n10830) );
  NAND2_X1 U13377 ( .A1(n13305), .A2(n13171), .ZN(n10829) );
  NAND2_X1 U13378 ( .A1(n10830), .A2(n10829), .ZN(n10901) );
  NAND3_X1 U13379 ( .A1(n10831), .A2(n10833), .A3(n10832), .ZN(n10834) );
  AOI21_X1 U13380 ( .B1(n10835), .B2(n10834), .A(n13462), .ZN(n10836) );
  AOI211_X1 U13381 ( .C1(n14801), .C2(n10837), .A(n10901), .B(n10836), .ZN(
        n10852) );
  MUX2_X1 U13382 ( .A(n10244), .B(n10852), .S(n14733), .Z(n10843) );
  INV_X1 U13383 ( .A(n10882), .ZN(n10838) );
  AOI211_X1 U13384 ( .C1(n10911), .C2(n11126), .A(n11505), .B(n10838), .ZN(
        n10850) );
  INV_X1 U13385 ( .A(n10911), .ZN(n10840) );
  INV_X1 U13386 ( .A(n10839), .ZN(n10904) );
  OAI22_X1 U13387 ( .A1(n13453), .A2(n10840), .B1(n14724), .B2(n10904), .ZN(
        n10841) );
  AOI21_X1 U13388 ( .B1(n10850), .B2(n13473), .A(n10841), .ZN(n10842) );
  OAI211_X1 U13389 ( .C1(n10853), .C2(n10976), .A(n10843), .B(n10842), .ZN(
        P2_U3259) );
  INV_X1 U13390 ( .A(n10844), .ZN(n10846) );
  NOR2_X1 U13391 ( .A1(n10846), .A2(n10845), .ZN(n10849) );
  INV_X1 U13392 ( .A(n10847), .ZN(n10848) );
  AND2_X1 U13393 ( .A1(n10848), .A2(n14741), .ZN(n14742) );
  INV_X1 U13394 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10855) );
  AOI21_X1 U13395 ( .B1(n14814), .B2(n10911), .A(n10850), .ZN(n10851) );
  OAI211_X1 U13396 ( .C1(n10853), .C2(n14769), .A(n10852), .B(n10851), .ZN(
        n10858) );
  NAND2_X1 U13397 ( .A1(n10858), .A2(n14831), .ZN(n10854) );
  OAI21_X1 U13398 ( .B1(n14831), .B2(n10855), .A(n10854), .ZN(P2_U3448) );
  INV_X1 U13399 ( .A(n14740), .ZN(n10856) );
  NAND2_X1 U13400 ( .A1(n10858), .A2(n14853), .ZN(n10859) );
  OAI21_X1 U13401 ( .B1(n14853), .B2(n10860), .A(n10859), .ZN(P2_U3505) );
  XNOR2_X1 U13402 ( .A(n10862), .B(n10861), .ZN(n14770) );
  NAND3_X1 U13403 ( .A1(n10863), .A2(n8647), .A3(n10864), .ZN(n10865) );
  AOI21_X1 U13404 ( .B1(n10999), .B2(n10865), .A(n13462), .ZN(n10868) );
  OAI22_X1 U13405 ( .A1(n10867), .A2(n13256), .B1(n10866), .B2(n13254), .ZN(
        n13164) );
  NOR2_X1 U13406 ( .A1(n10868), .A2(n13164), .ZN(n14768) );
  MUX2_X1 U13407 ( .A(n10239), .B(n14768), .S(n14733), .Z(n10872) );
  AOI211_X1 U13408 ( .C1(n14766), .C2(n10977), .A(n11505), .B(n11004), .ZN(
        n14765) );
  OAI22_X1 U13409 ( .A1(n13453), .A2(n10869), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n14724), .ZN(n10870) );
  AOI21_X1 U13410 ( .B1(n14765), .B2(n13473), .A(n10870), .ZN(n10871) );
  OAI211_X1 U13411 ( .C1(n14715), .C2(n14770), .A(n10872), .B(n10871), .ZN(
        P2_U3262) );
  INV_X1 U13412 ( .A(n13318), .ZN(n10873) );
  OAI222_X1 U13413 ( .A1(n13591), .A2(n10874), .B1(n13589), .B2(n10875), .C1(
        n10873), .C2(P2_U3088), .ZN(P2_U3309) );
  INV_X1 U13414 ( .A(n13875), .ZN(n13868) );
  OAI222_X1 U13415 ( .A1(n14245), .A2(n10876), .B1(n14251), .B2(n10875), .C1(
        P1_U3086), .C2(n13868), .ZN(P1_U3337) );
  XOR2_X1 U13416 ( .A(n10878), .B(n10877), .Z(n14792) );
  XNOR2_X1 U13417 ( .A(n10879), .B(n10878), .ZN(n10881) );
  AOI21_X1 U13418 ( .B1(n10881), .B2(n14725), .A(n10880), .ZN(n14791) );
  MUX2_X1 U13419 ( .A(n10243), .B(n14791), .S(n14733), .Z(n10887) );
  AOI211_X1 U13420 ( .C1(n14789), .C2(n10882), .A(n11505), .B(n11152), .ZN(
        n14788) );
  INV_X1 U13421 ( .A(n14789), .ZN(n10884) );
  OAI22_X1 U13422 ( .A1(n13453), .A2(n10884), .B1(n10883), .B2(n14724), .ZN(
        n10885) );
  AOI21_X1 U13423 ( .B1(n14788), .B2(n13473), .A(n10885), .ZN(n10886) );
  OAI211_X1 U13424 ( .C1(n14792), .C2(n14715), .A(n10887), .B(n10886), .ZN(
        P2_U3258) );
  INV_X1 U13425 ( .A(n15035), .ZN(n10897) );
  OAI21_X1 U13426 ( .B1(n10890), .B2(n10889), .A(n10888), .ZN(n10891) );
  NAND2_X1 U13427 ( .A1(n10891), .A2(n12670), .ZN(n10896) );
  NOR2_X1 U13428 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10892), .ZN(n14880) );
  OAI22_X1 U13429 ( .A1(n15041), .A2(n12676), .B1(n15029), .B2(n12665), .ZN(
        n10893) );
  AOI211_X1 U13430 ( .C1(n12648), .C2(n10894), .A(n14880), .B(n10893), .ZN(
        n10895) );
  OAI211_X1 U13431 ( .C1(n10897), .C2(n11500), .A(n10896), .B(n10895), .ZN(
        P3_U3170) );
  OAI222_X1 U13432 ( .A1(n13138), .A2(n10900), .B1(n12303), .B2(n10899), .C1(
        P3_U3151), .C2(n10898), .ZN(P3_U3275) );
  NAND2_X1 U13433 ( .A1(n13257), .A2(n10901), .ZN(n10902) );
  OAI211_X1 U13434 ( .C1(n13259), .C2(n10904), .A(n10903), .B(n10902), .ZN(
        n10910) );
  INV_X1 U13435 ( .A(n10905), .ZN(n10906) );
  AOI211_X1 U13436 ( .C1(n10908), .C2(n10907), .A(n13267), .B(n10906), .ZN(
        n10909) );
  AOI211_X1 U13437 ( .C1(n10911), .C2(n13262), .A(n10910), .B(n10909), .ZN(
        n10912) );
  INV_X1 U13438 ( .A(n10912), .ZN(P2_U3211) );
  XNOR2_X1 U13439 ( .A(n10913), .B(n12509), .ZN(n15093) );
  INV_X1 U13440 ( .A(n15093), .ZN(n10923) );
  OR2_X1 U13441 ( .A1(n15073), .A2(n12342), .ZN(n15054) );
  INV_X1 U13442 ( .A(n15054), .ZN(n15033) );
  NAND2_X1 U13443 ( .A1(n15080), .A2(n15033), .ZN(n12852) );
  OAI22_X1 U13444 ( .A1(n15017), .A2(n14339), .B1(n10914), .B2(n14341), .ZN(
        n10919) );
  INV_X1 U13445 ( .A(n10915), .ZN(n10916) );
  AOI211_X1 U13446 ( .C1(n12509), .C2(n10917), .A(n15045), .B(n10916), .ZN(
        n10918) );
  AOI211_X1 U13447 ( .C1(n15093), .C2(n15070), .A(n10919), .B(n10918), .ZN(
        n15090) );
  MUX2_X1 U13448 ( .A(n11621), .B(n15090), .S(n15080), .Z(n10922) );
  NOR2_X1 U13449 ( .A1(n12358), .A2(n15115), .ZN(n15092) );
  AOI22_X1 U13450 ( .A1(n15092), .A2(n15036), .B1(n15077), .B2(n10920), .ZN(
        n10921) );
  OAI211_X1 U13451 ( .C1(n10923), .C2(n12852), .A(n10922), .B(n10921), .ZN(
        P3_U3230) );
  XNOR2_X1 U13452 ( .A(n11154), .B(n12199), .ZN(n10924) );
  NAND2_X1 U13453 ( .A1(n13302), .A2(n12193), .ZN(n10925) );
  NAND2_X1 U13454 ( .A1(n10924), .A2(n10925), .ZN(n11098) );
  INV_X1 U13455 ( .A(n10924), .ZN(n10927) );
  INV_X1 U13456 ( .A(n10925), .ZN(n10926) );
  NAND2_X1 U13457 ( .A1(n10927), .A2(n10926), .ZN(n11100) );
  NAND2_X1 U13458 ( .A1(n11098), .A2(n11100), .ZN(n10933) );
  INV_X1 U13459 ( .A(n10928), .ZN(n10929) );
  NAND2_X1 U13460 ( .A1(n10930), .A2(n10929), .ZN(n10931) );
  NAND2_X1 U13461 ( .A1(n10932), .A2(n10931), .ZN(n11099) );
  XOR2_X1 U13462 ( .A(n10933), .B(n11099), .Z(n10942) );
  INV_X1 U13463 ( .A(n11153), .ZN(n10939) );
  NAND2_X1 U13464 ( .A1(n13301), .A2(n13172), .ZN(n10935) );
  NAND2_X1 U13465 ( .A1(n13303), .A2(n13171), .ZN(n10934) );
  AND2_X1 U13466 ( .A1(n10935), .A2(n10934), .ZN(n11158) );
  INV_X1 U13467 ( .A(n11158), .ZN(n10936) );
  NAND2_X1 U13468 ( .A1(n13257), .A2(n10936), .ZN(n10937) );
  OAI211_X1 U13469 ( .C1(n13259), .C2(n10939), .A(n10938), .B(n10937), .ZN(
        n10940) );
  AOI21_X1 U13470 ( .B1(n11154), .B2(n13262), .A(n10940), .ZN(n10941) );
  OAI21_X1 U13471 ( .B1(n10942), .B2(n13267), .A(n10941), .ZN(P2_U3193) );
  XOR2_X1 U13472 ( .A(n10944), .B(n10943), .Z(n10948) );
  NOR2_X1 U13473 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n7586), .ZN(n14897) );
  OAI22_X1 U13474 ( .A1(n15017), .A2(n12676), .B1(n15018), .B2(n12665), .ZN(
        n10945) );
  AOI211_X1 U13475 ( .C1(n12648), .C2(n15020), .A(n14897), .B(n10945), .ZN(
        n10947) );
  NAND2_X1 U13476 ( .A1(n12678), .A2(n15021), .ZN(n10946) );
  OAI211_X1 U13477 ( .C1(n10948), .C2(n12650), .A(n10947), .B(n10946), .ZN(
        P3_U3167) );
  INV_X1 U13478 ( .A(n10949), .ZN(n10952) );
  OAI222_X1 U13479 ( .A1(n13591), .A2(n10950), .B1(n13589), .B2(n10952), .C1(
        n14720), .C2(P2_U3088), .ZN(P2_U3308) );
  OAI222_X1 U13480 ( .A1(P1_U3086), .A2(n11860), .B1(n14251), .B2(n10952), 
        .C1(n10951), .C2(n14245), .ZN(P1_U3336) );
  INV_X1 U13481 ( .A(n11559), .ZN(n10958) );
  XNOR2_X1 U13482 ( .A(n10954), .B(n10953), .ZN(n10957) );
  OAI22_X1 U13483 ( .A1(n11542), .A2(n13624), .B1(n10955), .B2(n13633), .ZN(
        n11562) );
  INV_X1 U13484 ( .A(n11562), .ZN(n10956) );
  OAI21_X1 U13485 ( .B1(n10957), .B2(n14534), .A(n10956), .ZN(n11085) );
  AOI21_X1 U13486 ( .B1(n10958), .B2(n14034), .A(n11085), .ZN(n10967) );
  INV_X1 U13487 ( .A(n11196), .ZN(n10960) );
  INV_X1 U13488 ( .A(n11052), .ZN(n10959) );
  AOI211_X1 U13489 ( .C1(n11552), .C2(n10960), .A(n14119), .B(n10959), .ZN(
        n11086) );
  OAI22_X1 U13490 ( .A1(n11565), .A2(n14482), .B1(n14080), .B2(n10553), .ZN(
        n10961) );
  AOI21_X1 U13491 ( .B1(n11086), .B2(n14485), .A(n10961), .ZN(n10966) );
  OAI21_X1 U13492 ( .B1(n10964), .B2(n10963), .A(n10962), .ZN(n11087) );
  NAND2_X1 U13493 ( .A1(n11087), .A2(n14092), .ZN(n10965) );
  OAI211_X1 U13494 ( .C1(n10967), .C2(n14479), .A(n10966), .B(n10965), .ZN(
        P1_U3285) );
  XNOR2_X1 U13495 ( .A(n10969), .B(n10968), .ZN(n14761) );
  NAND2_X1 U13496 ( .A1(n14761), .A2(n14801), .ZN(n10975) );
  OAI21_X1 U13497 ( .B1(n10971), .B2(n10970), .A(n10863), .ZN(n10973) );
  AOI21_X1 U13498 ( .B1(n10973), .B2(n14725), .A(n10972), .ZN(n10974) );
  AND2_X1 U13499 ( .A1(n10975), .A2(n10974), .ZN(n14763) );
  INV_X1 U13500 ( .A(n10976), .ZN(n11320) );
  OAI211_X1 U13501 ( .C1(n11177), .C2(n14759), .A(n11440), .B(n10977), .ZN(
        n14758) );
  INV_X1 U13502 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10979) );
  INV_X1 U13503 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10978) );
  OAI22_X1 U13504 ( .A1(n14733), .A2(n10979), .B1(n10978), .B2(n14724), .ZN(
        n10980) );
  AOI21_X1 U13505 ( .B1(n14706), .B2(n10981), .A(n10980), .ZN(n10982) );
  OAI21_X1 U13506 ( .B1(n14714), .B2(n14758), .A(n10982), .ZN(n10983) );
  AOI21_X1 U13507 ( .B1(n11320), .B2(n14761), .A(n10983), .ZN(n10984) );
  OAI21_X1 U13508 ( .B1(n14736), .B2(n14763), .A(n10984), .ZN(P2_U3263) );
  OAI222_X1 U13509 ( .A1(n13138), .A2(n10986), .B1(n12303), .B2(n10985), .C1(
        P3_U3151), .C2(n12342), .ZN(P3_U3274) );
  INV_X1 U13510 ( .A(n11262), .ZN(n10994) );
  OAI211_X1 U13511 ( .C1(n10989), .C2(n10988), .A(n10987), .B(n12670), .ZN(
        n10993) );
  NOR2_X1 U13512 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10990), .ZN(n14915) );
  OAI22_X1 U13513 ( .A1(n15029), .A2(n12676), .B1(n11354), .B2(n12665), .ZN(
        n10991) );
  AOI211_X1 U13514 ( .C1(n12648), .C2(n11261), .A(n14915), .B(n10991), .ZN(
        n10992) );
  OAI211_X1 U13515 ( .C1(n10994), .C2(n11500), .A(n10993), .B(n10992), .ZN(
        P3_U3179) );
  XNOR2_X1 U13516 ( .A(n10995), .B(n10998), .ZN(n14774) );
  INV_X1 U13517 ( .A(n14774), .ZN(n11012) );
  NAND3_X1 U13518 ( .A1(n10999), .A2(n10998), .A3(n10997), .ZN(n11000) );
  NAND2_X1 U13519 ( .A1(n10996), .A2(n11000), .ZN(n11001) );
  NAND2_X1 U13520 ( .A1(n11001), .A2(n14725), .ZN(n11003) );
  NAND2_X1 U13521 ( .A1(n11003), .A2(n11002), .ZN(n14778) );
  OAI211_X1 U13522 ( .C1(n11004), .C2(n14776), .A(n11440), .B(n11125), .ZN(
        n14775) );
  OAI22_X1 U13523 ( .A1(n14733), .A2(n11006), .B1(n11005), .B2(n14724), .ZN(
        n11007) );
  AOI21_X1 U13524 ( .B1(n14706), .B2(n11008), .A(n11007), .ZN(n11009) );
  OAI21_X1 U13525 ( .B1(n14714), .B2(n14775), .A(n11009), .ZN(n11010) );
  AOI21_X1 U13526 ( .B1(n14778), .B2(n14733), .A(n11010), .ZN(n11011) );
  OAI21_X1 U13527 ( .B1(n11012), .B2(n14715), .A(n11011), .ZN(P2_U3261) );
  NAND2_X1 U13528 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n13696)
         );
  INV_X1 U13529 ( .A(n13696), .ZN(n11013) );
  AOI21_X1 U13530 ( .B1(n13827), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n11013), 
        .ZN(n11014) );
  INV_X1 U13531 ( .A(n11014), .ZN(n11020) );
  OAI21_X1 U13532 ( .B1(n11021), .B2(P1_REG1_REG_12__SCAN_IN), .A(n11015), 
        .ZN(n11018) );
  INV_X1 U13533 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n11016) );
  MUX2_X1 U13534 ( .A(n11016), .B(P1_REG1_REG_13__SCAN_IN), .S(n11212), .Z(
        n11017) );
  NOR2_X1 U13535 ( .A1(n11018), .A2(n11017), .ZN(n11211) );
  AOI211_X1 U13536 ( .C1(n11018), .C2(n11017), .A(n11211), .B(n13880), .ZN(
        n11019) );
  AOI211_X1 U13537 ( .C1(n14465), .C2(n11212), .A(n11020), .B(n11019), .ZN(
        n11027) );
  NOR2_X1 U13538 ( .A1(n11021), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n11022) );
  NOR2_X1 U13539 ( .A1(n11023), .A2(n11022), .ZN(n11025) );
  INV_X1 U13540 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11470) );
  MUX2_X1 U13541 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n11470), .S(n11212), .Z(
        n11024) );
  NAND2_X1 U13542 ( .A1(n11024), .A2(n11025), .ZN(n11217) );
  OAI211_X1 U13543 ( .C1(n11025), .C2(n11024), .A(n13883), .B(n11217), .ZN(
        n11026) );
  NAND2_X1 U13544 ( .A1(n11027), .A2(n11026), .ZN(P1_U3256) );
  NAND2_X1 U13545 ( .A1(n12702), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n11028) );
  OAI21_X1 U13546 ( .B1(n11029), .B2(n12702), .A(n11028), .ZN(P3_U3520) );
  NAND2_X1 U13547 ( .A1(n14657), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11031) );
  NOR2_X1 U13548 ( .A1(n11034), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n14637) );
  INV_X1 U13549 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11030) );
  MUX2_X1 U13550 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n11030), .S(n14643), .Z(
        n14638) );
  OAI21_X1 U13551 ( .B1(n14639), .B2(n14637), .A(n14638), .ZN(n14641) );
  OAI21_X1 U13552 ( .B1(n14643), .B2(P2_REG2_REG_12__SCAN_IN), .A(n14641), 
        .ZN(n14654) );
  INV_X1 U13553 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11460) );
  MUX2_X1 U13554 ( .A(n11460), .B(P2_REG2_REG_13__SCAN_IN), .S(n14657), .Z(
        n14653) );
  NAND2_X1 U13555 ( .A1(n11031), .A2(n14655), .ZN(n12225) );
  XNOR2_X1 U13556 ( .A(n12226), .B(n12225), .ZN(n11032) );
  NOR2_X1 U13557 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n11032), .ZN(n12227) );
  AOI21_X1 U13558 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n11032), .A(n12227), 
        .ZN(n11044) );
  INV_X1 U13559 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n14381) );
  INV_X1 U13560 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n14388) );
  AOI21_X1 U13561 ( .B1(n11034), .B2(P2_REG1_REG_11__SCAN_IN), .A(n11033), 
        .ZN(n14636) );
  MUX2_X1 U13562 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n14388), .S(n14643), .Z(
        n14635) );
  MUX2_X1 U13563 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n14381), .S(n14657), .Z(
        n14650) );
  NAND2_X1 U13564 ( .A1(n14651), .A2(n14650), .ZN(n14649) );
  OAI21_X1 U13565 ( .B1(n14381), .B2(n11036), .A(n14649), .ZN(n11038) );
  XNOR2_X1 U13566 ( .A(n12239), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n11037) );
  NAND2_X1 U13567 ( .A1(n11037), .A2(n11038), .ZN(n12237) );
  OAI211_X1 U13568 ( .C1(n11038), .C2(n11037), .A(n14688), .B(n12237), .ZN(
        n11043) );
  NOR2_X1 U13569 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11039), .ZN(n11041) );
  NOR2_X1 U13570 ( .A1(n14620), .A2(n12239), .ZN(n11040) );
  AOI211_X1 U13571 ( .C1(n14684), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n11041), 
        .B(n11040), .ZN(n11042) );
  OAI211_X1 U13572 ( .C1(n11044), .C2(n14652), .A(n11043), .B(n11042), .ZN(
        P2_U3228) );
  NAND2_X1 U13573 ( .A1(n12702), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n11045) );
  OAI21_X1 U13574 ( .B1(n12494), .B2(n12702), .A(n11045), .ZN(P3_U3521) );
  OAI21_X1 U13575 ( .B1(n11048), .B2(n11047), .A(n11046), .ZN(n11051) );
  OAI22_X1 U13576 ( .A1(n11050), .A2(n13624), .B1(n11049), .B2(n13633), .ZN(
        n11847) );
  AOI21_X1 U13577 ( .B1(n11051), .B2(n14526), .A(n11847), .ZN(n11277) );
  AOI21_X1 U13578 ( .B1(n11052), .B2(n11851), .A(n14119), .ZN(n11053) );
  AND2_X1 U13579 ( .A1(n11053), .A2(n11241), .ZN(n11279) );
  INV_X1 U13580 ( .A(n11851), .ZN(n11054) );
  NOR2_X1 U13581 ( .A1(n14482), .A2(n11054), .ZN(n11057) );
  OAI22_X1 U13582 ( .A1(n14080), .A2(n11055), .B1(n11849), .B2(n14477), .ZN(
        n11056) );
  AOI211_X1 U13583 ( .C1(n11279), .C2(n14485), .A(n11057), .B(n11056), .ZN(
        n11062) );
  OAI21_X1 U13584 ( .B1(n11060), .B2(n11059), .A(n11058), .ZN(n11280) );
  NAND2_X1 U13585 ( .A1(n11280), .A2(n14092), .ZN(n11061) );
  OAI211_X1 U13586 ( .C1(n11277), .C2(n14479), .A(n11062), .B(n11061), .ZN(
        P1_U3284) );
  INV_X1 U13587 ( .A(n11063), .ZN(n11065) );
  OAI22_X1 U13588 ( .A1(n12543), .A2(P3_U3151), .B1(SI_22_), .B2(n12303), .ZN(
        n11064) );
  AOI21_X1 U13589 ( .B1(n11065), .B2(n14270), .A(n11064), .ZN(P3_U3273) );
  INV_X1 U13590 ( .A(n11066), .ZN(n11069) );
  INV_X1 U13591 ( .A(n11067), .ZN(n11068) );
  OAI22_X1 U13592 ( .A1(n12125), .A2(n11071), .B1(n14520), .B2(n12092), .ZN(
        n11075) );
  OAI22_X1 U13593 ( .A1(n11071), .A2(n12092), .B1(n14520), .B2(n12090), .ZN(
        n11072) );
  XOR2_X1 U13594 ( .A(n12265), .B(n11072), .Z(n11117) );
  INV_X1 U13595 ( .A(n11117), .ZN(n11073) );
  AOI22_X1 U13596 ( .A1(n12282), .A2(n11990), .B1(n13770), .B2(n12275), .ZN(
        n11077) );
  XOR2_X1 U13597 ( .A(n12265), .B(n11077), .Z(n11425) );
  OAI22_X1 U13598 ( .A1(n6627), .A2(n12092), .B1(n11078), .B2(n12125), .ZN(
        n11426) );
  XNOR2_X1 U13599 ( .A(n11425), .B(n11426), .ZN(n11079) );
  XNOR2_X1 U13600 ( .A(n6605), .B(n11079), .ZN(n11084) );
  AOI22_X1 U13601 ( .A1(n13771), .A2(n13913), .B1(n13717), .B2(n13769), .ZN(
        n11987) );
  NAND2_X1 U13602 ( .A1(n6468), .A2(n11990), .ZN(n11081) );
  OAI211_X1 U13603 ( .C1(n11987), .C2(n13739), .A(n11081), .B(n11080), .ZN(
        n11082) );
  AOI21_X1 U13604 ( .B1(n11994), .B2(n13742), .A(n11082), .ZN(n11083) );
  OAI21_X1 U13605 ( .B1(n11084), .B2(n13731), .A(n11083), .ZN(P1_U3227) );
  AOI211_X1 U13606 ( .C1(n14430), .C2(n11087), .A(n11086), .B(n11085), .ZN(
        n11092) );
  INV_X1 U13607 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n11088) );
  OAI22_X1 U13608 ( .A1(n14232), .A2(n11565), .B1(n14549), .B2(n11088), .ZN(
        n11089) );
  INV_X1 U13609 ( .A(n11089), .ZN(n11090) );
  OAI21_X1 U13610 ( .B1(n11092), .B2(n14547), .A(n11090), .ZN(P1_U3483) );
  AOI22_X1 U13611 ( .A1(n14163), .A2(n11552), .B1(n14558), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n11091) );
  OAI21_X1 U13612 ( .B1(n11092), .B2(n14558), .A(n11091), .ZN(P1_U3536) );
  XNOR2_X1 U13613 ( .A(n14710), .B(n12199), .ZN(n11093) );
  NAND2_X1 U13614 ( .A1(n13301), .A2(n6477), .ZN(n11094) );
  NAND2_X1 U13615 ( .A1(n11093), .A2(n11094), .ZN(n11163) );
  INV_X1 U13616 ( .A(n11093), .ZN(n11096) );
  INV_X1 U13617 ( .A(n11094), .ZN(n11095) );
  NAND2_X1 U13618 ( .A1(n11096), .A2(n11095), .ZN(n11097) );
  NAND2_X1 U13619 ( .A1(n11163), .A2(n11097), .ZN(n11106) );
  NAND2_X1 U13620 ( .A1(n11099), .A2(n11098), .ZN(n11101) );
  INV_X1 U13621 ( .A(n11164), .ZN(n11104) );
  AOI21_X1 U13622 ( .B1(n11106), .B2(n11105), .A(n11104), .ZN(n11113) );
  INV_X1 U13623 ( .A(n14704), .ZN(n11110) );
  NAND2_X1 U13624 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n14616) );
  OAI22_X1 U13625 ( .A1(n11108), .A2(n13254), .B1(n11107), .B2(n13256), .ZN(
        n14702) );
  NAND2_X1 U13626 ( .A1(n13257), .A2(n14702), .ZN(n11109) );
  OAI211_X1 U13627 ( .C1(n13259), .C2(n11110), .A(n14616), .B(n11109), .ZN(
        n11111) );
  AOI21_X1 U13628 ( .B1(n14710), .B2(n13262), .A(n11111), .ZN(n11112) );
  OAI21_X1 U13629 ( .B1(n11113), .B2(n13267), .A(n11112), .ZN(P2_U3203) );
  AOI211_X1 U13630 ( .C1(n11117), .C2(n11116), .A(n13731), .B(n11115), .ZN(
        n11118) );
  INV_X1 U13631 ( .A(n11118), .ZN(n11122) );
  NAND2_X1 U13632 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n12142) );
  OAI21_X1 U13633 ( .B1(n13739), .B2(n14518), .A(n12142), .ZN(n11119) );
  AOI21_X1 U13634 ( .B1(n6468), .B2(n11120), .A(n11119), .ZN(n11121) );
  OAI211_X1 U13635 ( .C1(n14417), .C2(n11123), .A(n11122), .B(n11121), .ZN(
        P1_U3230) );
  XNOR2_X1 U13636 ( .A(n11124), .B(n11132), .ZN(n14781) );
  AOI21_X1 U13637 ( .B1(n11125), .B2(n11129), .A(n11505), .ZN(n11127) );
  NAND2_X1 U13638 ( .A1(n11127), .A2(n11126), .ZN(n14782) );
  AOI22_X1 U13639 ( .A1(n14706), .A2(n11129), .B1(n14705), .B2(n11128), .ZN(
        n11130) );
  OAI21_X1 U13640 ( .B1(n14714), .B2(n14782), .A(n11130), .ZN(n11138) );
  NAND3_X1 U13641 ( .A1(n10996), .A2(n11132), .A3(n11131), .ZN(n11133) );
  NAND2_X1 U13642 ( .A1(n10831), .A2(n11133), .ZN(n11134) );
  NAND2_X1 U13643 ( .A1(n11134), .A2(n14725), .ZN(n11136) );
  NAND2_X1 U13644 ( .A1(n11136), .A2(n11135), .ZN(n14785) );
  MUX2_X1 U13645 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n14785), .S(n14733), .Z(
        n11137) );
  AOI211_X1 U13646 ( .C1(n13426), .C2(n14781), .A(n11138), .B(n11137), .ZN(
        n11139) );
  INV_X1 U13647 ( .A(n11139), .ZN(P2_U3260) );
  INV_X1 U13648 ( .A(n11234), .ZN(n11147) );
  OAI211_X1 U13649 ( .C1(n11142), .C2(n11141), .A(n11140), .B(n12670), .ZN(
        n11146) );
  NOR2_X1 U13650 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11143), .ZN(n14932) );
  OAI22_X1 U13651 ( .A1(n15018), .A2(n12676), .B1(n11388), .B2(n12665), .ZN(
        n11144) );
  AOI211_X1 U13652 ( .C1(n12648), .C2(n11233), .A(n14932), .B(n11144), .ZN(
        n11145) );
  OAI211_X1 U13653 ( .C1(n11147), .C2(n11500), .A(n11146), .B(n11145), .ZN(
        P3_U3153) );
  INV_X1 U13654 ( .A(n11148), .ZN(n11185) );
  OAI222_X1 U13655 ( .A1(n11150), .A2(P1_U3086), .B1(n14251), .B2(n11185), 
        .C1(n11149), .C2(n14245), .ZN(P1_U3335) );
  AOI21_X1 U13656 ( .B1(n11157), .B2(n11151), .A(n6601), .ZN(n14800) );
  OAI211_X1 U13657 ( .C1(n11152), .C2(n14797), .A(n14711), .B(n11440), .ZN(
        n14795) );
  AOI22_X1 U13658 ( .A1(n14706), .A2(n11154), .B1(n14705), .B2(n11153), .ZN(
        n11155) );
  OAI21_X1 U13659 ( .B1(n14795), .B2(n14714), .A(n11155), .ZN(n11161) );
  XOR2_X1 U13660 ( .A(n11156), .B(n11157), .Z(n11159) );
  OAI21_X1 U13661 ( .B1(n11159), .B2(n13462), .A(n11158), .ZN(n14799) );
  MUX2_X1 U13662 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n14799), .S(n14733), .Z(
        n11160) );
  AOI211_X1 U13663 ( .C1(n14800), .C2(n13426), .A(n11161), .B(n11160), .ZN(
        n11162) );
  INV_X1 U13664 ( .A(n11162), .ZN(P2_U3257) );
  XNOR2_X1 U13665 ( .A(n14813), .B(n12199), .ZN(n11365) );
  NAND2_X1 U13666 ( .A1(n13300), .A2(n12193), .ZN(n11364) );
  XNOR2_X1 U13667 ( .A(n11365), .B(n11364), .ZN(n11366) );
  XNOR2_X1 U13668 ( .A(n11367), .B(n11366), .ZN(n11172) );
  INV_X1 U13669 ( .A(n11328), .ZN(n11169) );
  NAND2_X1 U13670 ( .A1(n13299), .A2(n13172), .ZN(n11166) );
  NAND2_X1 U13671 ( .A1(n13301), .A2(n13171), .ZN(n11165) );
  NAND2_X1 U13672 ( .A1(n11166), .A2(n11165), .ZN(n11325) );
  NOR2_X1 U13673 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11167), .ZN(n14622) );
  AOI21_X1 U13674 ( .B1(n13257), .B2(n11325), .A(n14622), .ZN(n11168) );
  OAI21_X1 U13675 ( .B1(n11169), .B2(n13259), .A(n11168), .ZN(n11170) );
  AOI21_X1 U13676 ( .B1(n14813), .B2(n13262), .A(n11170), .ZN(n11171) );
  OAI21_X1 U13677 ( .B1(n11172), .B2(n13267), .A(n11171), .ZN(P2_U3189) );
  XNOR2_X1 U13678 ( .A(n11173), .B(n9474), .ZN(n11175) );
  AOI21_X1 U13679 ( .B1(n11175), .B2(n14725), .A(n11174), .ZN(n14754) );
  XNOR2_X1 U13680 ( .A(n9474), .B(n11176), .ZN(n14751) );
  INV_X1 U13681 ( .A(n11177), .ZN(n11179) );
  AOI21_X1 U13682 ( .B1(n14746), .B2(n11180), .A(n11505), .ZN(n11178) );
  NAND2_X1 U13683 ( .A1(n11179), .A2(n11178), .ZN(n14753) );
  AOI22_X1 U13684 ( .A1(n14736), .A2(P2_REG2_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(n14705), .ZN(n11182) );
  NAND2_X1 U13685 ( .A1(n14706), .A2(n11180), .ZN(n11181) );
  OAI211_X1 U13686 ( .C1(n14714), .C2(n14753), .A(n11182), .B(n11181), .ZN(
        n11183) );
  AOI21_X1 U13687 ( .B1(n14751), .B2(n13426), .A(n11183), .ZN(n11184) );
  OAI21_X1 U13688 ( .B1(n14736), .B2(n14754), .A(n11184), .ZN(P2_U3264) );
  OAI222_X1 U13689 ( .A1(n13591), .A2(n6950), .B1(P2_U3088), .B2(n8681), .C1(
        n13589), .C2(n11185), .ZN(P2_U3307) );
  NOR2_X1 U13690 ( .A1(n14092), .A2(n14071), .ZN(n11192) );
  OAI22_X1 U13691 ( .A1(n14479), .A2(n11187), .B1(n11186), .B2(n14477), .ZN(
        n11190) );
  AOI21_X1 U13692 ( .B1(n13956), .B2(n14482), .A(n11188), .ZN(n11189) );
  AOI211_X1 U13693 ( .C1(n14479), .C2(P1_REG2_REG_0__SCAN_IN), .A(n11190), .B(
        n11189), .ZN(n11191) );
  OAI21_X1 U13694 ( .B1(n11193), .B2(n11192), .A(n11191), .ZN(P1_U3293) );
  INV_X1 U13695 ( .A(n14541), .ZN(n14532) );
  OAI21_X1 U13696 ( .B1(n11195), .B2(n11200), .A(n11194), .ZN(n14487) );
  AOI211_X1 U13697 ( .C1(n14475), .C2(n11197), .A(n14119), .B(n11196), .ZN(
        n14484) );
  NAND2_X1 U13698 ( .A1(n13767), .A2(n13717), .ZN(n11199) );
  NAND2_X1 U13699 ( .A1(n13769), .A2(n13913), .ZN(n11198) );
  NAND2_X1 U13700 ( .A1(n11199), .A2(n11198), .ZN(n11596) );
  XNOR2_X1 U13701 ( .A(n11201), .B(n11200), .ZN(n11202) );
  NOR2_X1 U13702 ( .A1(n11202), .A2(n14534), .ZN(n11203) );
  AOI211_X1 U13703 ( .C1(n14546), .C2(n14487), .A(n11596), .B(n11203), .ZN(
        n14490) );
  INV_X1 U13704 ( .A(n14490), .ZN(n11204) );
  AOI211_X1 U13705 ( .C1(n14532), .C2(n14487), .A(n14484), .B(n11204), .ZN(
        n11209) );
  AOI22_X1 U13706 ( .A1(n14163), .A2(n14475), .B1(n14558), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n11205) );
  OAI21_X1 U13707 ( .B1(n11209), .B2(n14558), .A(n11205), .ZN(P1_U3535) );
  INV_X1 U13708 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n11206) );
  NOR2_X1 U13709 ( .A1(n14549), .A2(n11206), .ZN(n11207) );
  AOI21_X1 U13710 ( .B1(n9158), .B2(n14475), .A(n11207), .ZN(n11208) );
  OAI21_X1 U13711 ( .B1(n11209), .B2(n14547), .A(n11208), .ZN(P1_U3480) );
  MUX2_X1 U13712 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n11210), .S(n11695), .Z(
        n11214) );
  OAI21_X1 U13713 ( .B1(n11214), .B2(n11213), .A(n11694), .ZN(n11224) );
  NAND2_X1 U13714 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14400)
         );
  INV_X1 U13715 ( .A(n14400), .ZN(n11215) );
  AOI21_X1 U13716 ( .B1(n13827), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n11215), 
        .ZN(n11222) );
  MUX2_X1 U13717 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n11216), .S(n11695), .Z(
        n11220) );
  OAI21_X1 U13718 ( .B1(n11218), .B2(n11470), .A(n11217), .ZN(n11219) );
  NAND2_X1 U13719 ( .A1(n11220), .A2(n11219), .ZN(n11703) );
  OAI211_X1 U13720 ( .C1(n11220), .C2(n11219), .A(n13883), .B(n11703), .ZN(
        n11221) );
  OAI211_X1 U13721 ( .C1(n13806), .C2(n11704), .A(n11222), .B(n11221), .ZN(
        n11223) );
  AOI21_X1 U13722 ( .B1(n14462), .B2(n11224), .A(n11223), .ZN(n11225) );
  INV_X1 U13723 ( .A(n11225), .ZN(P1_U3257) );
  XNOR2_X1 U13724 ( .A(n11227), .B(n11226), .ZN(n11232) );
  OAI21_X1 U13725 ( .B1(n11229), .B2(n12504), .A(n11228), .ZN(n15107) );
  OAI22_X1 U13726 ( .A1(n11388), .A2(n14339), .B1(n15018), .B2(n14341), .ZN(
        n11230) );
  AOI21_X1 U13727 ( .B1(n15107), .B2(n15070), .A(n11230), .ZN(n11231) );
  OAI21_X1 U13728 ( .B1(n11232), .B2(n15045), .A(n11231), .ZN(n15105) );
  INV_X1 U13729 ( .A(n15105), .ZN(n11238) );
  INV_X1 U13730 ( .A(n12852), .ZN(n15078) );
  AND2_X1 U13731 ( .A1(n11233), .A2(n15071), .ZN(n15106) );
  AOI22_X1 U13732 ( .A1(n15036), .A2(n15106), .B1(n15077), .B2(n11234), .ZN(
        n11235) );
  OAI21_X1 U13733 ( .B1(n11642), .B2(n15080), .A(n11235), .ZN(n11236) );
  AOI21_X1 U13734 ( .B1(n15107), .B2(n15078), .A(n11236), .ZN(n11237) );
  OAI21_X1 U13735 ( .B1(n11238), .B2(n15082), .A(n11237), .ZN(P3_U3226) );
  XNOR2_X1 U13736 ( .A(n11239), .B(n11246), .ZN(n11342) );
  NAND2_X1 U13737 ( .A1(n13766), .A2(n13913), .ZN(n11337) );
  OAI21_X1 U13738 ( .B1(n14477), .B2(n11881), .A(n11337), .ZN(n11240) );
  MUX2_X1 U13739 ( .A(n11240), .B(P1_REG2_REG_10__SCAN_IN), .S(n14491), .Z(
        n11244) );
  AOI211_X1 U13740 ( .C1(n11883), .C2(n11241), .A(n14119), .B(n11298), .ZN(
        n11339) );
  INV_X1 U13741 ( .A(n11339), .ZN(n11242) );
  OR2_X1 U13742 ( .A1(n12007), .A2(n13633), .ZN(n11338) );
  AOI21_X1 U13743 ( .B1(n11242), .B2(n11338), .A(n14085), .ZN(n11243) );
  AOI211_X1 U13744 ( .C1(n14082), .C2(n11883), .A(n11244), .B(n11243), .ZN(
        n11249) );
  OAI21_X1 U13745 ( .B1(n11247), .B2(n11246), .A(n11245), .ZN(n11340) );
  NAND2_X1 U13746 ( .A1(n11340), .A2(n14092), .ZN(n11248) );
  OAI211_X1 U13747 ( .C1(n11342), .C2(n14042), .A(n11249), .B(n11248), .ZN(
        P1_U3283) );
  OAI222_X1 U13748 ( .A1(n11251), .A2(P1_U3086), .B1(n14251), .B2(n11266), 
        .C1(n11250), .C2(n14245), .ZN(P1_U3334) );
  XNOR2_X1 U13749 ( .A(n11253), .B(n11252), .ZN(n15104) );
  INV_X1 U13750 ( .A(n15104), .ZN(n11265) );
  OAI211_X1 U13751 ( .C1(n11255), .C2(n12507), .A(n11254), .B(n15060), .ZN(
        n11259) );
  OAI22_X1 U13752 ( .A1(n15029), .A2(n14341), .B1(n11354), .B2(n14339), .ZN(
        n11256) );
  INV_X1 U13753 ( .A(n11256), .ZN(n11258) );
  NAND2_X1 U13754 ( .A1(n15104), .A2(n15070), .ZN(n11257) );
  NAND3_X1 U13755 ( .A1(n11259), .A2(n11258), .A3(n11257), .ZN(n15102) );
  MUX2_X1 U13756 ( .A(n15102), .B(P3_REG2_REG_6__SCAN_IN), .S(n15082), .Z(
        n11260) );
  INV_X1 U13757 ( .A(n11260), .ZN(n11264) );
  AND2_X1 U13758 ( .A1(n11261), .A2(n15071), .ZN(n15103) );
  AOI22_X1 U13759 ( .A1(n15036), .A2(n15103), .B1(n15077), .B2(n11262), .ZN(
        n11263) );
  OAI211_X1 U13760 ( .C1(n11265), .C2(n12852), .A(n11264), .B(n11263), .ZN(
        P3_U3227) );
  OAI222_X1 U13761 ( .A1(n13591), .A2(n11268), .B1(P2_U3088), .B2(n11267), 
        .C1(n13589), .C2(n11266), .ZN(P2_U3306) );
  INV_X1 U13762 ( .A(n11269), .ZN(n11358) );
  OAI211_X1 U13763 ( .C1(n11272), .C2(n11271), .A(n11270), .B(n12670), .ZN(
        n11276) );
  NOR2_X1 U13764 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11273), .ZN(n14949) );
  OAI22_X1 U13765 ( .A1(n11354), .A2(n12676), .B1(n12387), .B2(n12665), .ZN(
        n11274) );
  AOI211_X1 U13766 ( .C1(n12648), .C2(n11360), .A(n14949), .B(n11274), .ZN(
        n11275) );
  OAI211_X1 U13767 ( .C1(n11358), .C2(n11500), .A(n11276), .B(n11275), .ZN(
        P3_U3161) );
  INV_X1 U13768 ( .A(n11277), .ZN(n11278) );
  AOI211_X1 U13769 ( .C1(n14430), .C2(n11280), .A(n11279), .B(n11278), .ZN(
        n11285) );
  AOI22_X1 U13770 ( .A1(n14163), .A2(n11851), .B1(n14558), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n11281) );
  OAI21_X1 U13771 ( .B1(n11285), .B2(n14558), .A(n11281), .ZN(P1_U3537) );
  INV_X1 U13772 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n11282) );
  NOR2_X1 U13773 ( .A1(n14549), .A2(n11282), .ZN(n11283) );
  AOI21_X1 U13774 ( .B1(n9158), .B2(n11851), .A(n11283), .ZN(n11284) );
  OAI21_X1 U13775 ( .B1(n11285), .B2(n14547), .A(n11284), .ZN(P1_U3486) );
  NAND2_X1 U13776 ( .A1(n11286), .A2(n14270), .ZN(n11287) );
  OAI211_X1 U13777 ( .C1(n11288), .C2(n12303), .A(n11287), .B(n12546), .ZN(
        P3_U3272) );
  XNOR2_X1 U13778 ( .A(n11289), .B(n11295), .ZN(n11290) );
  NAND2_X1 U13779 ( .A1(n11290), .A2(n14526), .ZN(n11293) );
  NAND2_X1 U13780 ( .A1(n13765), .A2(n13913), .ZN(n11291) );
  OAI21_X1 U13781 ( .B1(n12016), .B2(n13633), .A(n11291), .ZN(n14412) );
  INV_X1 U13782 ( .A(n14412), .ZN(n11292) );
  NAND2_X1 U13783 ( .A1(n11293), .A2(n11292), .ZN(n14427) );
  INV_X1 U13784 ( .A(n14427), .ZN(n11304) );
  OAI21_X1 U13785 ( .B1(n11296), .B2(n11295), .A(n11294), .ZN(n14429) );
  INV_X1 U13786 ( .A(n11415), .ZN(n11297) );
  OAI211_X1 U13787 ( .C1(n14426), .C2(n11298), .A(n11297), .B(n14493), .ZN(
        n14425) );
  OAI22_X1 U13788 ( .A1(n14080), .A2(n11299), .B1(n14416), .B2(n14477), .ZN(
        n11300) );
  AOI21_X1 U13789 ( .B1(n14413), .B2(n14082), .A(n11300), .ZN(n11301) );
  OAI21_X1 U13790 ( .B1(n14425), .B2(n14085), .A(n11301), .ZN(n11302) );
  AOI21_X1 U13791 ( .B1(n14429), .B2(n14092), .A(n11302), .ZN(n11303) );
  OAI21_X1 U13792 ( .B1(n11304), .B2(n14491), .A(n11303), .ZN(P1_U3282) );
  XNOR2_X1 U13793 ( .A(n11306), .B(n11305), .ZN(n14826) );
  NAND2_X1 U13794 ( .A1(n14826), .A2(n14801), .ZN(n11315) );
  NAND3_X1 U13795 ( .A1(n11324), .A2(n11308), .A3(n11307), .ZN(n11309) );
  NAND2_X1 U13796 ( .A1(n11310), .A2(n11309), .ZN(n11313) );
  NAND2_X1 U13797 ( .A1(n13298), .A2(n13172), .ZN(n11312) );
  NAND2_X1 U13798 ( .A1(n13300), .A2(n13171), .ZN(n11311) );
  NAND2_X1 U13799 ( .A1(n11312), .A2(n11311), .ZN(n11378) );
  AOI21_X1 U13800 ( .B1(n11313), .B2(n14725), .A(n11378), .ZN(n11314) );
  INV_X1 U13801 ( .A(n12193), .ZN(n11440) );
  OAI21_X1 U13802 ( .B1(n11327), .B2(n14823), .A(n11440), .ZN(n11316) );
  OR2_X1 U13803 ( .A1(n11316), .A2(n11441), .ZN(n14821) );
  AOI22_X1 U13804 ( .A1(n14736), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n11376), 
        .B2(n14705), .ZN(n11318) );
  NAND2_X1 U13805 ( .A1(n11382), .A2(n14706), .ZN(n11317) );
  OAI211_X1 U13806 ( .C1(n14821), .C2(n14714), .A(n11318), .B(n11317), .ZN(
        n11319) );
  AOI21_X1 U13807 ( .B1(n14826), .B2(n11320), .A(n11319), .ZN(n11321) );
  OAI21_X1 U13808 ( .B1(n14828), .B2(n14736), .A(n11321), .ZN(P2_U3254) );
  NAND2_X1 U13809 ( .A1(n11322), .A2(n11332), .ZN(n11323) );
  NAND2_X1 U13810 ( .A1(n11324), .A2(n11323), .ZN(n11326) );
  AOI21_X1 U13811 ( .B1(n11326), .B2(n14725), .A(n11325), .ZN(n14816) );
  AOI211_X1 U13812 ( .C1(n14813), .C2(n14712), .A(n11505), .B(n11327), .ZN(
        n14812) );
  INV_X1 U13813 ( .A(n14813), .ZN(n11330) );
  AOI22_X1 U13814 ( .A1(n14736), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n11328), 
        .B2(n14705), .ZN(n11329) );
  OAI21_X1 U13815 ( .B1(n11330), .B2(n13453), .A(n11329), .ZN(n11335) );
  OAI21_X1 U13816 ( .B1(n11333), .B2(n11332), .A(n11331), .ZN(n14818) );
  NOR2_X1 U13817 ( .A1(n14818), .A2(n14715), .ZN(n11334) );
  AOI211_X1 U13818 ( .C1(n13473), .C2(n14812), .A(n11335), .B(n11334), .ZN(
        n11336) );
  OAI21_X1 U13819 ( .B1(n14736), .B2(n14816), .A(n11336), .ZN(P2_U3255) );
  NAND2_X1 U13820 ( .A1(n11338), .A2(n11337), .ZN(n11879) );
  AOI211_X1 U13821 ( .C1(n11340), .C2(n14430), .A(n11339), .B(n11879), .ZN(
        n11341) );
  OAI21_X1 U13822 ( .B1(n14534), .B2(n11342), .A(n11341), .ZN(n11348) );
  OAI22_X1 U13823 ( .A1(n11346), .A2(n14186), .B1(n14560), .B2(n10547), .ZN(
        n11343) );
  AOI21_X1 U13824 ( .B1(n11348), .B2(n14560), .A(n11343), .ZN(n11344) );
  INV_X1 U13825 ( .A(n11344), .ZN(P1_U3538) );
  INV_X1 U13826 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n11345) );
  OAI22_X1 U13827 ( .A1(n11346), .A2(n14232), .B1(n14549), .B2(n11345), .ZN(
        n11347) );
  AOI21_X1 U13828 ( .B1(n11348), .B2(n14549), .A(n11347), .ZN(n11349) );
  INV_X1 U13829 ( .A(n11349), .ZN(P1_U3489) );
  OR2_X1 U13830 ( .A1(n11350), .A2(n12503), .ZN(n11351) );
  NAND2_X1 U13831 ( .A1(n11352), .A2(n11351), .ZN(n15111) );
  INV_X1 U13832 ( .A(n15111), .ZN(n11363) );
  XOR2_X1 U13833 ( .A(n12503), .B(n11353), .Z(n11357) );
  OAI22_X1 U13834 ( .A1(n12387), .A2(n14339), .B1(n11354), .B2(n14341), .ZN(
        n11355) );
  AOI21_X1 U13835 ( .B1(n15111), .B2(n15070), .A(n11355), .ZN(n11356) );
  OAI21_X1 U13836 ( .B1(n11357), .B2(n15045), .A(n11356), .ZN(n15109) );
  NAND2_X1 U13837 ( .A1(n15109), .A2(n15080), .ZN(n11362) );
  OAI22_X1 U13838 ( .A1(n15080), .A2(n11648), .B1(n11358), .B2(n15009), .ZN(
        n11359) );
  AOI21_X1 U13839 ( .B1(n15004), .B2(n11360), .A(n11359), .ZN(n11361) );
  OAI211_X1 U13840 ( .C1(n11363), .C2(n12852), .A(n11362), .B(n11361), .ZN(
        P3_U3225) );
  XNOR2_X1 U13841 ( .A(n11382), .B(n12199), .ZN(n11368) );
  NAND2_X1 U13842 ( .A1(n13299), .A2(n12193), .ZN(n11369) );
  NAND2_X1 U13843 ( .A1(n11368), .A2(n11369), .ZN(n11394) );
  INV_X1 U13844 ( .A(n11368), .ZN(n11371) );
  INV_X1 U13845 ( .A(n11369), .ZN(n11370) );
  NAND2_X1 U13846 ( .A1(n11371), .A2(n11370), .ZN(n11372) );
  NAND2_X1 U13847 ( .A1(n11394), .A2(n11372), .ZN(n11374) );
  INV_X1 U13848 ( .A(n11395), .ZN(n11373) );
  AOI21_X1 U13849 ( .B1(n11375), .B2(n11374), .A(n11373), .ZN(n11384) );
  INV_X1 U13850 ( .A(n11376), .ZN(n11380) );
  AOI21_X1 U13851 ( .B1(n13257), .B2(n11378), .A(n11377), .ZN(n11379) );
  OAI21_X1 U13852 ( .B1(n11380), .B2(n13259), .A(n11379), .ZN(n11381) );
  AOI21_X1 U13853 ( .B1(n11382), .B2(n13262), .A(n11381), .ZN(n11383) );
  OAI21_X1 U13854 ( .B1(n11384), .B2(n13267), .A(n11383), .ZN(P2_U3208) );
  AOI21_X1 U13855 ( .B1(n11387), .B2(n11386), .A(n11385), .ZN(n11393) );
  AND2_X1 U13856 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n14968) );
  OAI22_X1 U13857 ( .A1(n11388), .A2(n12676), .B1(n14342), .B2(n12665), .ZN(
        n11389) );
  AOI211_X1 U13858 ( .C1(n12648), .C2(n15003), .A(n14968), .B(n11389), .ZN(
        n11392) );
  NAND2_X1 U13859 ( .A1(n12678), .A2(n11390), .ZN(n11391) );
  OAI211_X1 U13860 ( .C1(n11393), .C2(n12650), .A(n11392), .B(n11391), .ZN(
        P3_U3171) );
  NAND2_X1 U13861 ( .A1(n11395), .A2(n11394), .ZN(n11503) );
  XNOR2_X1 U13862 ( .A(n11443), .B(n12199), .ZN(n11396) );
  NAND2_X1 U13863 ( .A1(n13298), .A2(n6477), .ZN(n11397) );
  AND2_X1 U13864 ( .A1(n11396), .A2(n11397), .ZN(n11502) );
  INV_X1 U13865 ( .A(n11502), .ZN(n11400) );
  INV_X1 U13866 ( .A(n11396), .ZN(n11399) );
  INV_X1 U13867 ( .A(n11397), .ZN(n11398) );
  NAND2_X1 U13868 ( .A1(n11399), .A2(n11398), .ZN(n11501) );
  NAND2_X1 U13869 ( .A1(n11400), .A2(n11501), .ZN(n11401) );
  XNOR2_X1 U13870 ( .A(n11503), .B(n11401), .ZN(n11407) );
  INV_X1 U13871 ( .A(n11442), .ZN(n11404) );
  OAI22_X1 U13872 ( .A1(n11402), .A2(n13254), .B1(n7107), .B2(n13256), .ZN(
        n11436) );
  AOI22_X1 U13873 ( .A1(n13257), .A2(n11436), .B1(P2_REG3_REG_12__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11403) );
  OAI21_X1 U13874 ( .B1(n11404), .B2(n13259), .A(n11403), .ZN(n11405) );
  AOI21_X1 U13875 ( .B1(n11443), .B2(n13262), .A(n11405), .ZN(n11406) );
  OAI21_X1 U13876 ( .B1(n11407), .B2(n13267), .A(n11406), .ZN(P2_U3196) );
  OAI21_X1 U13877 ( .B1(n11409), .B2(n7347), .A(n11408), .ZN(n11576) );
  XNOR2_X1 U13878 ( .A(n11410), .B(n11411), .ZN(n11412) );
  AOI22_X1 U13879 ( .A1(n13764), .A2(n13913), .B1(n13717), .B2(n13762), .ZN(
        n13647) );
  OAI21_X1 U13880 ( .B1(n11412), .B2(n14534), .A(n13647), .ZN(n11413) );
  AOI21_X1 U13881 ( .B1(n14546), .B2(n11576), .A(n11413), .ZN(n11578) );
  INV_X1 U13882 ( .A(n11414), .ZN(n14486) );
  OAI211_X1 U13883 ( .C1(n11415), .C2(n13652), .A(n14493), .B(n11472), .ZN(
        n11577) );
  OAI22_X1 U13884 ( .A1(n14080), .A2(n11416), .B1(n13645), .B2(n14477), .ZN(
        n11417) );
  AOI21_X1 U13885 ( .B1(n11418), .B2(n14082), .A(n11417), .ZN(n11419) );
  OAI21_X1 U13886 ( .B1(n11577), .B2(n14085), .A(n11419), .ZN(n11420) );
  AOI21_X1 U13887 ( .B1(n11576), .B2(n14486), .A(n11420), .ZN(n11421) );
  OAI21_X1 U13888 ( .B1(n11578), .B2(n14491), .A(n11421), .ZN(P1_U3281) );
  NAND2_X1 U13889 ( .A1(n14411), .A2(n14536), .ZN(n11422) );
  OAI211_X1 U13890 ( .C1(n14417), .C2(n11424), .A(n11423), .B(n11422), .ZN(
        n11433) );
  INV_X1 U13891 ( .A(n11426), .ZN(n11427) );
  NAND2_X1 U13892 ( .A1(n14537), .A2(n12282), .ZN(n11429) );
  NAND2_X1 U13893 ( .A1(n13769), .A2(n12275), .ZN(n11428) );
  NAND2_X1 U13894 ( .A1(n11429), .A2(n11428), .ZN(n11430) );
  XNOR2_X1 U13895 ( .A(n11430), .B(n12265), .ZN(n11536) );
  AOI22_X1 U13896 ( .A1(n14537), .A2(n12285), .B1(n12284), .B2(n13769), .ZN(
        n11541) );
  XNOR2_X1 U13897 ( .A(n11536), .B(n11541), .ZN(n11537) );
  XNOR2_X1 U13898 ( .A(n11538), .B(n11537), .ZN(n11431) );
  NOR2_X1 U13899 ( .A1(n11431), .A2(n13731), .ZN(n11432) );
  AOI211_X1 U13900 ( .C1(n14537), .C2(n6468), .A(n11433), .B(n11432), .ZN(
        n11434) );
  INV_X1 U13901 ( .A(n11434), .ZN(P1_U3239) );
  XNOR2_X1 U13902 ( .A(n11435), .B(n11438), .ZN(n11437) );
  AOI21_X1 U13903 ( .B1(n11437), .B2(n14725), .A(n11436), .ZN(n14384) );
  XOR2_X1 U13904 ( .A(n11439), .B(n11438), .Z(n14382) );
  INV_X1 U13905 ( .A(n14382), .ZN(n11447) );
  OAI211_X1 U13906 ( .C1(n11441), .C2(n14385), .A(n11440), .B(n11456), .ZN(
        n14383) );
  AOI22_X1 U13907 ( .A1(n14736), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n11442), 
        .B2(n14705), .ZN(n11445) );
  NAND2_X1 U13908 ( .A1(n11443), .A2(n14706), .ZN(n11444) );
  OAI211_X1 U13909 ( .C1(n14383), .C2(n14714), .A(n11445), .B(n11444), .ZN(
        n11446) );
  AOI21_X1 U13910 ( .B1(n11447), .B2(n13426), .A(n11446), .ZN(n11448) );
  OAI21_X1 U13911 ( .B1(n14736), .B2(n14384), .A(n11448), .ZN(P2_U3253) );
  XNOR2_X1 U13912 ( .A(n11449), .B(n11454), .ZN(n11450) );
  NAND2_X1 U13913 ( .A1(n11450), .A2(n14725), .ZN(n11453) );
  NAND2_X1 U13914 ( .A1(n13296), .A2(n13172), .ZN(n11452) );
  NAND2_X1 U13915 ( .A1(n13298), .A2(n13171), .ZN(n11451) );
  AND2_X1 U13916 ( .A1(n11452), .A2(n11451), .ZN(n11513) );
  NAND2_X1 U13917 ( .A1(n11453), .A2(n11513), .ZN(n14378) );
  INV_X1 U13918 ( .A(n14378), .ZN(n11465) );
  XOR2_X1 U13919 ( .A(n11455), .B(n11454), .Z(n14380) );
  INV_X1 U13920 ( .A(n11456), .ZN(n11458) );
  INV_X1 U13921 ( .A(n11504), .ZN(n14377) );
  OAI211_X1 U13922 ( .C1(n11458), .C2(n14377), .A(n11440), .B(n11760), .ZN(
        n14376) );
  INV_X1 U13923 ( .A(n11515), .ZN(n11459) );
  OAI22_X1 U13924 ( .A1(n14733), .A2(n11460), .B1(n11459), .B2(n14724), .ZN(
        n11461) );
  AOI21_X1 U13925 ( .B1(n11504), .B2(n14706), .A(n11461), .ZN(n11462) );
  OAI21_X1 U13926 ( .B1(n14376), .B2(n14714), .A(n11462), .ZN(n11463) );
  AOI21_X1 U13927 ( .B1(n14380), .B2(n13426), .A(n11463), .ZN(n11464) );
  OAI21_X1 U13928 ( .B1(n14736), .B2(n11465), .A(n11464), .ZN(P2_U3252) );
  INV_X1 U13929 ( .A(n11466), .ZN(n11467) );
  OAI222_X1 U13930 ( .A1(n7977), .A2(P3_U3151), .B1(n13138), .B2(n11467), .C1(
        n6810), .C2(n12303), .ZN(P3_U3271) );
  OAI21_X1 U13931 ( .B1(n11469), .B2(n11474), .A(n11468), .ZN(n11486) );
  INV_X1 U13932 ( .A(n11486), .ZN(n11482) );
  OAI22_X1 U13933 ( .A1(n14080), .A2(n11470), .B1(n13695), .B2(n14477), .ZN(
        n11471) );
  AOI21_X1 U13934 ( .B1(n12024), .B2(n14082), .A(n11471), .ZN(n11481) );
  AOI21_X1 U13935 ( .B1(n11472), .B2(n12024), .A(n14119), .ZN(n11473) );
  NAND2_X1 U13936 ( .A1(n11473), .A2(n11519), .ZN(n11483) );
  XNOR2_X1 U13937 ( .A(n11475), .B(n11474), .ZN(n11476) );
  NAND2_X1 U13938 ( .A1(n11476), .A2(n14526), .ZN(n11484) );
  NAND2_X1 U13939 ( .A1(n13761), .A2(n13717), .ZN(n11478) );
  NAND2_X1 U13940 ( .A1(n13763), .A2(n13913), .ZN(n11477) );
  AND2_X1 U13941 ( .A1(n11478), .A2(n11477), .ZN(n13697) );
  OAI211_X1 U13942 ( .C1(n14023), .C2(n11483), .A(n11484), .B(n13697), .ZN(
        n11479) );
  NAND2_X1 U13943 ( .A1(n11479), .A2(n14080), .ZN(n11480) );
  OAI211_X1 U13944 ( .C1(n11482), .C2(n14073), .A(n11481), .B(n11480), .ZN(
        P1_U3280) );
  NAND3_X1 U13945 ( .A1(n11484), .A2(n13697), .A3(n11483), .ZN(n11485) );
  AOI21_X1 U13946 ( .B1(n14430), .B2(n11486), .A(n11485), .ZN(n11491) );
  INV_X1 U13947 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n11487) );
  OAI22_X1 U13948 ( .A1(n13702), .A2(n14232), .B1(n14549), .B2(n11487), .ZN(
        n11488) );
  INV_X1 U13949 ( .A(n11488), .ZN(n11489) );
  OAI21_X1 U13950 ( .B1(n11491), .B2(n14547), .A(n11489), .ZN(P1_U3498) );
  AOI22_X1 U13951 ( .A1(n12024), .A2(n14163), .B1(n14558), .B2(
        P1_REG1_REG_13__SCAN_IN), .ZN(n11490) );
  OAI21_X1 U13952 ( .B1(n11491), .B2(n14558), .A(n11490), .ZN(P1_U3541) );
  INV_X1 U13953 ( .A(n11492), .ZN(n11591) );
  OAI211_X1 U13954 ( .C1(n11495), .C2(n11494), .A(n11493), .B(n12670), .ZN(
        n11499) );
  NOR2_X1 U13955 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11496), .ZN(n14979) );
  OAI22_X1 U13956 ( .A1(n11825), .A2(n12665), .B1(n12681), .B2(n15114), .ZN(
        n11497) );
  AOI211_X1 U13957 ( .C1(n12663), .C2(n12695), .A(n14979), .B(n11497), .ZN(
        n11498) );
  OAI211_X1 U13958 ( .C1(n11591), .C2(n11500), .A(n11499), .B(n11498), .ZN(
        P3_U3157) );
  XNOR2_X1 U13959 ( .A(n11504), .B(n12209), .ZN(n11506) );
  AND2_X1 U13960 ( .A1(n13297), .A2(n11505), .ZN(n11507) );
  NAND2_X1 U13961 ( .A1(n11506), .A2(n11507), .ZN(n11721) );
  INV_X1 U13962 ( .A(n11506), .ZN(n11509) );
  INV_X1 U13963 ( .A(n11507), .ZN(n11508) );
  NAND2_X1 U13964 ( .A1(n11509), .A2(n11508), .ZN(n11510) );
  AND2_X1 U13965 ( .A1(n11721), .A2(n11510), .ZN(n11511) );
  OAI211_X1 U13966 ( .C1(n11512), .C2(n11511), .A(n11722), .B(n13241), .ZN(
        n11517) );
  OAI22_X1 U13967 ( .A1(n13272), .A2(n11513), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8386), .ZN(n11514) );
  AOI21_X1 U13968 ( .B1(n11515), .B2(n13274), .A(n11514), .ZN(n11516) );
  OAI211_X1 U13969 ( .C1(n14377), .C2(n13278), .A(n11517), .B(n11516), .ZN(
        P2_U3206) );
  OAI21_X1 U13970 ( .B1(n6593), .B2(n8899), .A(n11518), .ZN(n14422) );
  AOI21_X1 U13971 ( .B1(n14419), .B2(n11519), .A(n14119), .ZN(n11521) );
  NAND2_X1 U13972 ( .A1(n11521), .A2(n11743), .ZN(n14420) );
  INV_X1 U13973 ( .A(n14420), .ZN(n11529) );
  INV_X1 U13974 ( .A(n14419), .ZN(n11527) );
  NAND2_X1 U13975 ( .A1(n13762), .A2(n13913), .ZN(n11522) );
  OAI21_X1 U13976 ( .B1(n11523), .B2(n13633), .A(n11522), .ZN(n14418) );
  INV_X1 U13977 ( .A(n14418), .ZN(n11524) );
  OAI22_X1 U13978 ( .A1(n14479), .A2(n11524), .B1(n14402), .B2(n14477), .ZN(
        n11525) );
  AOI21_X1 U13979 ( .B1(n14479), .B2(P1_REG2_REG_14__SCAN_IN), .A(n11525), 
        .ZN(n11526) );
  OAI21_X1 U13980 ( .B1(n11527), .B2(n14482), .A(n11526), .ZN(n11528) );
  AOI21_X1 U13981 ( .B1(n11529), .B2(n14485), .A(n11528), .ZN(n11532) );
  XNOR2_X1 U13982 ( .A(n11530), .B(n8899), .ZN(n14424) );
  NAND2_X1 U13983 ( .A1(n14424), .A2(n14071), .ZN(n11531) );
  OAI211_X1 U13984 ( .C1(n14422), .C2(n14073), .A(n11532), .B(n11531), .ZN(
        P1_U3279) );
  AOI222_X1 U13985 ( .A1(n11534), .A2(n12220), .B1(n11533), .B2(
        P2_STATE_REG_SCAN_IN), .C1(P1_DATAO_REG_22__SCAN_IN), .C2(n13593), 
        .ZN(n11535) );
  INV_X1 U13986 ( .A(n11535), .ZN(P2_U3305) );
  INV_X1 U13987 ( .A(n11536), .ZN(n11540) );
  NOR2_X1 U13988 ( .A1(n11542), .A2(n12125), .ZN(n11543) );
  AOI21_X1 U13989 ( .B1(n14475), .B2(n12275), .A(n11543), .ZN(n11545) );
  AOI22_X1 U13990 ( .A1(n14475), .A2(n12282), .B1(n12285), .B2(n13768), .ZN(
        n11544) );
  XNOR2_X1 U13991 ( .A(n11544), .B(n12265), .ZN(n11546) );
  XOR2_X1 U13992 ( .A(n11545), .B(n11546), .Z(n11600) );
  INV_X1 U13993 ( .A(n11545), .ZN(n11548) );
  INV_X1 U13994 ( .A(n11546), .ZN(n11547) );
  NAND2_X1 U13995 ( .A1(n11552), .A2(n12282), .ZN(n11550) );
  NAND2_X1 U13996 ( .A1(n13767), .A2(n12285), .ZN(n11549) );
  NAND2_X1 U13997 ( .A1(n11550), .A2(n11549), .ZN(n11551) );
  XNOR2_X1 U13998 ( .A(n11551), .B(n12265), .ZN(n11556) );
  NAND2_X1 U13999 ( .A1(n11552), .A2(n12285), .ZN(n11554) );
  NAND2_X1 U14000 ( .A1(n12284), .A2(n13767), .ZN(n11553) );
  NAND2_X1 U14001 ( .A1(n11554), .A2(n11553), .ZN(n11555) );
  NOR2_X1 U14002 ( .A1(n11556), .A2(n11555), .ZN(n11835) );
  AOI21_X1 U14003 ( .B1(n11556), .B2(n11555), .A(n11835), .ZN(n11557) );
  OAI21_X1 U14004 ( .B1(n6606), .B2(n11557), .A(n11836), .ZN(n11558) );
  NAND2_X1 U14005 ( .A1(n11558), .A2(n14409), .ZN(n11564) );
  NOR2_X1 U14006 ( .A1(n14417), .A2(n11559), .ZN(n11560) );
  AOI211_X1 U14007 ( .C1(n14411), .C2(n11562), .A(n11561), .B(n11560), .ZN(
        n11563) );
  OAI211_X1 U14008 ( .C1(n11565), .C2(n13745), .A(n11564), .B(n11563), .ZN(
        P1_U3221) );
  INV_X1 U14009 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n11571) );
  XNOR2_X1 U14010 ( .A(n11566), .B(n12511), .ZN(n15002) );
  INV_X1 U14011 ( .A(n12511), .ZN(n11568) );
  OAI211_X1 U14012 ( .C1(n6602), .C2(n11568), .A(n15060), .B(n11567), .ZN(
        n11570) );
  AOI22_X1 U14013 ( .A1(n12694), .A2(n15063), .B1(n15062), .B2(n12696), .ZN(
        n11569) );
  NAND2_X1 U14014 ( .A1(n11570), .A2(n11569), .ZN(n15001) );
  AOI21_X1 U14015 ( .B1(n15002), .B2(n15100), .A(n15001), .ZN(n11573) );
  MUX2_X1 U14016 ( .A(n11571), .B(n11573), .S(n15120), .Z(n11572) );
  OAI21_X1 U14017 ( .B1(n13121), .B2(n6844), .A(n11572), .ZN(P3_U3417) );
  INV_X1 U14018 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n11574) );
  MUX2_X1 U14019 ( .A(n11574), .B(n11573), .S(n15131), .Z(n11575) );
  OAI21_X1 U14020 ( .B1(n13063), .B2(n6844), .A(n11575), .ZN(P3_U3468) );
  INV_X1 U14021 ( .A(n11576), .ZN(n11579) );
  OAI211_X1 U14022 ( .C1(n11579), .C2(n14541), .A(n11578), .B(n11577), .ZN(
        n11584) );
  OAI22_X1 U14023 ( .A1(n13652), .A2(n14186), .B1(n14560), .B2(n8864), .ZN(
        n11580) );
  AOI21_X1 U14024 ( .B1(n11584), .B2(n14560), .A(n11580), .ZN(n11581) );
  INV_X1 U14025 ( .A(n11581), .ZN(P1_U3540) );
  INV_X1 U14026 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n11582) );
  OAI22_X1 U14027 ( .A1(n13652), .A2(n14232), .B1(n14549), .B2(n11582), .ZN(
        n11583) );
  AOI21_X1 U14028 ( .B1(n11584), .B2(n14549), .A(n11583), .ZN(n11585) );
  INV_X1 U14029 ( .A(n11585), .ZN(P1_U3495) );
  XNOR2_X1 U14030 ( .A(n11586), .B(n12505), .ZN(n15117) );
  OAI211_X1 U14031 ( .C1(n11588), .C2(n12505), .A(n11587), .B(n15060), .ZN(
        n11590) );
  AOI22_X1 U14032 ( .A1(n15062), .A2(n12695), .B1(n12693), .B2(n15063), .ZN(
        n11589) );
  OAI211_X1 U14033 ( .C1(n15117), .C2(n11829), .A(n11590), .B(n11589), .ZN(
        n15119) );
  NAND2_X1 U14034 ( .A1(n15119), .A2(n15080), .ZN(n11595) );
  OAI22_X1 U14035 ( .A1(n15080), .A2(n11658), .B1(n11591), .B2(n15009), .ZN(
        n11592) );
  AOI21_X1 U14036 ( .B1(n15004), .B2(n11593), .A(n11592), .ZN(n11594) );
  OAI211_X1 U14037 ( .C1(n15117), .C2(n12852), .A(n11595), .B(n11594), .ZN(
        P3_U3223) );
  NAND2_X1 U14038 ( .A1(n14411), .A2(n11596), .ZN(n11597) );
  OAI211_X1 U14039 ( .C1(n14417), .C2(n14476), .A(n11598), .B(n11597), .ZN(
        n11603) );
  XNOR2_X1 U14040 ( .A(n11599), .B(n11600), .ZN(n11601) );
  NOR2_X1 U14041 ( .A1(n11601), .A2(n13731), .ZN(n11602) );
  AOI211_X1 U14042 ( .C1(n14475), .C2(n6468), .A(n11603), .B(n11602), .ZN(
        n11604) );
  INV_X1 U14043 ( .A(n11604), .ZN(P1_U3213) );
  NOR2_X1 U14044 ( .A1(n11668), .A2(n11606), .ZN(n11607) );
  AOI22_X1 U14045 ( .A1(n11670), .A2(P3_REG2_REG_4__SCAN_IN), .B1(n11627), 
        .B2(n14878), .ZN(n14871) );
  AOI21_X1 U14046 ( .B1(P3_REG2_REG_4__SCAN_IN), .B2(n14878), .A(n14870), .ZN(
        n11608) );
  NOR2_X1 U14047 ( .A1(n11672), .A2(n11608), .ZN(n11609) );
  AOI22_X1 U14048 ( .A1(n11674), .A2(P3_REG2_REG_6__SCAN_IN), .B1(n11610), 
        .B2(n14913), .ZN(n14905) );
  NOR2_X1 U14049 ( .A1(n11612), .A2(n11613), .ZN(n11614) );
  AOI22_X1 U14050 ( .A1(n11677), .A2(P3_REG2_REG_8__SCAN_IN), .B1(n11648), 
        .B2(n14947), .ZN(n14940) );
  NOR2_X1 U14051 ( .A1(n11615), .A2(n11616), .ZN(n11617) );
  NOR2_X1 U14052 ( .A1(n11652), .A2(n14958), .ZN(n14957) );
  NAND2_X1 U14053 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n11665), .ZN(n11618) );
  OAI21_X1 U14054 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n11665), .A(n11618), 
        .ZN(n14989) );
  AOI21_X1 U14055 ( .B1(n7512), .B2(n11619), .A(n11799), .ZN(n11689) );
  INV_X1 U14056 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n11620) );
  MUX2_X1 U14057 ( .A(n11621), .B(n11620), .S(n12776), .Z(n11622) );
  NAND2_X1 U14058 ( .A1(n11622), .A2(n11668), .ZN(n11625) );
  INV_X1 U14059 ( .A(n11622), .ZN(n11623) );
  NAND2_X1 U14060 ( .A1(n11623), .A2(n14861), .ZN(n11624) );
  NAND2_X1 U14061 ( .A1(n11625), .A2(n11624), .ZN(n14856) );
  INV_X1 U14062 ( .A(n11625), .ZN(n14873) );
  INV_X1 U14063 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n11626) );
  MUX2_X1 U14064 ( .A(n11627), .B(n11626), .S(n12776), .Z(n11628) );
  NAND2_X1 U14065 ( .A1(n11628), .A2(n11670), .ZN(n14891) );
  INV_X1 U14066 ( .A(n11628), .ZN(n11629) );
  NAND2_X1 U14067 ( .A1(n11629), .A2(n14878), .ZN(n11630) );
  AND2_X1 U14068 ( .A1(n14891), .A2(n11630), .ZN(n14872) );
  OAI21_X1 U14069 ( .B1(n14874), .B2(n14873), .A(n14872), .ZN(n14892) );
  INV_X1 U14070 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n11631) );
  MUX2_X1 U14071 ( .A(n11632), .B(n11631), .S(n12776), .Z(n11633) );
  NAND2_X1 U14072 ( .A1(n11633), .A2(n11672), .ZN(n11636) );
  INV_X1 U14073 ( .A(n11633), .ZN(n11634) );
  NAND2_X1 U14074 ( .A1(n11634), .A2(n14895), .ZN(n11635) );
  NAND2_X1 U14075 ( .A1(n11636), .A2(n11635), .ZN(n14890) );
  INV_X1 U14076 ( .A(n11636), .ZN(n14908) );
  INV_X1 U14077 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n11637) );
  MUX2_X1 U14078 ( .A(n11610), .B(n11637), .S(n6473), .Z(n11638) );
  NAND2_X1 U14079 ( .A1(n11638), .A2(n11674), .ZN(n14926) );
  INV_X1 U14080 ( .A(n11638), .ZN(n11639) );
  NAND2_X1 U14081 ( .A1(n11639), .A2(n14913), .ZN(n11640) );
  AND2_X1 U14082 ( .A1(n14926), .A2(n11640), .ZN(n14907) );
  OAI21_X1 U14083 ( .B1(n14909), .B2(n14908), .A(n14907), .ZN(n14927) );
  INV_X1 U14084 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n11641) );
  MUX2_X1 U14085 ( .A(n11642), .B(n11641), .S(n12776), .Z(n11643) );
  NAND2_X1 U14086 ( .A1(n11643), .A2(n11612), .ZN(n11646) );
  INV_X1 U14087 ( .A(n11643), .ZN(n11644) );
  NAND2_X1 U14088 ( .A1(n11644), .A2(n14930), .ZN(n11645) );
  NAND2_X1 U14089 ( .A1(n11646), .A2(n11645), .ZN(n14925) );
  INV_X1 U14090 ( .A(n11646), .ZN(n14942) );
  INV_X1 U14091 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n11647) );
  MUX2_X1 U14092 ( .A(n11648), .B(n11647), .S(n6473), .Z(n11649) );
  NAND2_X1 U14093 ( .A1(n11649), .A2(n11677), .ZN(n14960) );
  INV_X1 U14094 ( .A(n11649), .ZN(n11650) );
  NAND2_X1 U14095 ( .A1(n11650), .A2(n14947), .ZN(n11651) );
  AND2_X1 U14096 ( .A1(n14960), .A2(n11651), .ZN(n14941) );
  OAI21_X1 U14097 ( .B1(n14943), .B2(n14942), .A(n14941), .ZN(n14961) );
  MUX2_X1 U14098 ( .A(n11652), .B(n11574), .S(n12776), .Z(n11653) );
  NAND2_X1 U14099 ( .A1(n11653), .A2(n11615), .ZN(n11656) );
  INV_X1 U14100 ( .A(n11653), .ZN(n11654) );
  NAND2_X1 U14101 ( .A1(n11654), .A2(n14965), .ZN(n11655) );
  NAND2_X1 U14102 ( .A1(n11656), .A2(n11655), .ZN(n14959) );
  INV_X1 U14103 ( .A(n11656), .ZN(n14983) );
  INV_X1 U14104 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n11657) );
  MUX2_X1 U14105 ( .A(n11658), .B(n11657), .S(n6473), .Z(n11659) );
  NAND2_X1 U14106 ( .A1(n11659), .A2(n14995), .ZN(n11662) );
  INV_X1 U14107 ( .A(n11659), .ZN(n11660) );
  NAND2_X1 U14108 ( .A1(n11660), .A2(n11665), .ZN(n11661) );
  AND2_X1 U14109 ( .A1(n11662), .A2(n11661), .ZN(n14982) );
  OAI21_X1 U14110 ( .B1(n14984), .B2(n14983), .A(n14982), .ZN(n14987) );
  NAND2_X1 U14111 ( .A1(n14987), .A2(n11662), .ZN(n11664) );
  MUX2_X1 U14112 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n6473), .Z(n11810) );
  XNOR2_X1 U14113 ( .A(n11810), .B(n11811), .ZN(n11663) );
  NAND2_X1 U14114 ( .A1(n11664), .A2(n11663), .ZN(n11815) );
  OAI21_X1 U14115 ( .B1(n11664), .B2(n11663), .A(n11815), .ZN(n11687) );
  NAND2_X1 U14116 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n11665), .ZN(n11680) );
  AOI22_X1 U14117 ( .A1(n14995), .A2(n11657), .B1(P3_REG1_REG_10__SCAN_IN), 
        .B2(n11665), .ZN(n14978) );
  AOI22_X1 U14118 ( .A1(n11677), .A2(n11647), .B1(P3_REG1_REG_8__SCAN_IN), 
        .B2(n14947), .ZN(n14951) );
  AOI22_X1 U14119 ( .A1(n11674), .A2(n11637), .B1(P3_REG1_REG_6__SCAN_IN), 
        .B2(n14913), .ZN(n14917) );
  AOI22_X1 U14120 ( .A1(n11670), .A2(n11626), .B1(P3_REG1_REG_4__SCAN_IN), 
        .B2(n14878), .ZN(n14882) );
  NAND2_X1 U14121 ( .A1(n14861), .A2(n11667), .ZN(n11669) );
  XNOR2_X1 U14122 ( .A(n11668), .B(n11667), .ZN(n14865) );
  NAND2_X1 U14123 ( .A1(P3_REG1_REG_3__SCAN_IN), .A2(n14865), .ZN(n14864) );
  NAND2_X1 U14124 ( .A1(n11669), .A2(n14864), .ZN(n14883) );
  NAND2_X1 U14125 ( .A1(n14882), .A2(n14883), .ZN(n14881) );
  NAND2_X1 U14126 ( .A1(n14895), .A2(n11671), .ZN(n11673) );
  NAND2_X1 U14127 ( .A1(P3_REG1_REG_5__SCAN_IN), .A2(n14899), .ZN(n14898) );
  NAND2_X1 U14128 ( .A1(n11673), .A2(n14898), .ZN(n14918) );
  NAND2_X1 U14129 ( .A1(n14917), .A2(n14918), .ZN(n14916) );
  NAND2_X1 U14130 ( .A1(n14930), .A2(n11675), .ZN(n11676) );
  XNOR2_X1 U14131 ( .A(n11612), .B(n11675), .ZN(n14934) );
  NAND2_X1 U14132 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n14934), .ZN(n14933) );
  NAND2_X1 U14133 ( .A1(n14951), .A2(n14952), .ZN(n14950) );
  NAND2_X1 U14134 ( .A1(n14965), .A2(n11678), .ZN(n11679) );
  NAND2_X1 U14135 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n14971), .ZN(n14970) );
  NAND2_X1 U14136 ( .A1(n11679), .A2(n14970), .ZN(n14977) );
  XNOR2_X1 U14137 ( .A(n11811), .B(n11802), .ZN(n11681) );
  NAND2_X1 U14138 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n11681), .ZN(n11804) );
  OAI21_X1 U14139 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n11681), .A(n11804), 
        .ZN(n11682) );
  NAND2_X1 U14140 ( .A1(n11682), .A2(n6467), .ZN(n11685) );
  NOR2_X1 U14141 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11683), .ZN(n11781) );
  AOI21_X1 U14142 ( .B1(n14969), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n11781), 
        .ZN(n11684) );
  OAI211_X1 U14143 ( .C1(n14966), .C2(n11803), .A(n11685), .B(n11684), .ZN(
        n11686) );
  AOI21_X1 U14144 ( .B1(n11687), .B2(n14962), .A(n11686), .ZN(n11688) );
  OAI21_X1 U14145 ( .B1(n11689), .B2(n14991), .A(n11688), .ZN(P3_U3193) );
  INV_X1 U14146 ( .A(n11690), .ZN(n11692) );
  OAI222_X1 U14147 ( .A1(P3_U3151), .A2(n11693), .B1(n13138), .B2(n11692), 
        .C1(n11691), .C2(n12303), .ZN(P3_U3270) );
  NAND2_X1 U14148 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n13656)
         );
  OAI21_X1 U14149 ( .B1(n14473), .B2(n9717), .A(n13656), .ZN(n11702) );
  NAND2_X1 U14150 ( .A1(n11697), .A2(n11696), .ZN(n11698) );
  NAND2_X1 U14151 ( .A1(n14461), .A2(n14460), .ZN(n14459) );
  NAND2_X1 U14152 ( .A1(n11698), .A2(n14459), .ZN(n11700) );
  XNOR2_X1 U14153 ( .A(n13847), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n11699) );
  NOR2_X1 U14154 ( .A1(n11699), .A2(n11700), .ZN(n13846) );
  AOI211_X1 U14155 ( .C1(n11700), .C2(n11699), .A(n13846), .B(n13880), .ZN(
        n11701) );
  AOI211_X1 U14156 ( .C1(n14465), .C2(n13847), .A(n11702), .B(n11701), .ZN(
        n11710) );
  OAI21_X1 U14157 ( .B1(n11216), .B2(n11704), .A(n11703), .ZN(n11705) );
  NOR2_X1 U14158 ( .A1(n14464), .A2(n11705), .ZN(n11706) );
  XNOR2_X1 U14159 ( .A(n14464), .B(n11705), .ZN(n14458) );
  NOR2_X1 U14160 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14458), .ZN(n14457) );
  NOR2_X1 U14161 ( .A1(n11706), .A2(n14457), .ZN(n11708) );
  XNOR2_X1 U14162 ( .A(n13847), .B(n11864), .ZN(n11707) );
  NAND2_X1 U14163 ( .A1(n11707), .A2(n11708), .ZN(n13839) );
  OAI211_X1 U14164 ( .C1(n11708), .C2(n11707), .A(n13883), .B(n13839), .ZN(
        n11709) );
  NAND2_X1 U14165 ( .A1(n11710), .A2(n11709), .ZN(P1_U3259) );
  XNOR2_X1 U14166 ( .A(n6469), .B(n11713), .ZN(n11712) );
  AOI22_X1 U14167 ( .A1(n13294), .A2(n13172), .B1(n13296), .B2(n13171), .ZN(
        n13271) );
  OAI21_X1 U14168 ( .B1(n11712), .B2(n13462), .A(n13271), .ZN(n11773) );
  INV_X1 U14169 ( .A(n11773), .ZN(n11720) );
  XNOR2_X1 U14170 ( .A(n11714), .B(n11713), .ZN(n11775) );
  INV_X1 U14171 ( .A(n12161), .ZN(n13279) );
  INV_X1 U14172 ( .A(n11715), .ZN(n11759) );
  OAI211_X1 U14173 ( .C1(n13279), .C2(n11759), .A(n6491), .B(n11440), .ZN(
        n11772) );
  AOI22_X1 U14174 ( .A1(n14736), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n13275), 
        .B2(n14705), .ZN(n11717) );
  NAND2_X1 U14175 ( .A1(n12161), .A2(n14706), .ZN(n11716) );
  OAI211_X1 U14176 ( .C1(n11772), .C2(n14714), .A(n11717), .B(n11716), .ZN(
        n11718) );
  AOI21_X1 U14177 ( .B1(n11775), .B2(n13426), .A(n11718), .ZN(n11719) );
  OAI21_X1 U14178 ( .B1(n11720), .B2(n14736), .A(n11719), .ZN(P2_U3250) );
  XNOR2_X1 U14179 ( .A(n13557), .B(n12199), .ZN(n12158) );
  NAND2_X1 U14180 ( .A1(n13296), .A2(n11505), .ZN(n12157) );
  XNOR2_X1 U14181 ( .A(n12158), .B(n12157), .ZN(n11726) );
  INV_X1 U14182 ( .A(n11726), .ZN(n11723) );
  INV_X1 U14183 ( .A(n12160), .ZN(n11724) );
  AOI21_X1 U14184 ( .B1(n11726), .B2(n11725), .A(n11724), .ZN(n11733) );
  INV_X1 U14185 ( .A(n11761), .ZN(n11730) );
  NAND2_X1 U14186 ( .A1(n13295), .A2(n13172), .ZN(n11728) );
  NAND2_X1 U14187 ( .A1(n13297), .A2(n13171), .ZN(n11727) );
  NAND2_X1 U14188 ( .A1(n11728), .A2(n11727), .ZN(n11757) );
  AOI22_X1 U14189 ( .A1(n13257), .A2(n11757), .B1(P2_REG3_REG_14__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11729) );
  OAI21_X1 U14190 ( .B1(n11730), .B2(n13259), .A(n11729), .ZN(n11731) );
  AOI21_X1 U14191 ( .B1(n13557), .B2(n13262), .A(n11731), .ZN(n11732) );
  OAI21_X1 U14192 ( .B1(n11733), .B2(n13267), .A(n11732), .ZN(P2_U3187) );
  OAI21_X1 U14193 ( .B1(n11735), .B2(n8912), .A(n11734), .ZN(n11790) );
  XNOR2_X1 U14194 ( .A(n11736), .B(n8912), .ZN(n11793) );
  NAND2_X1 U14195 ( .A1(n11793), .A2(n14092), .ZN(n11747) );
  NAND2_X1 U14196 ( .A1(n13759), .A2(n13717), .ZN(n11738) );
  NAND2_X1 U14197 ( .A1(n13761), .A2(n13913), .ZN(n11737) );
  AND2_X1 U14198 ( .A1(n11738), .A2(n11737), .ZN(n13738) );
  INV_X1 U14199 ( .A(n13738), .ZN(n11740) );
  INV_X1 U14200 ( .A(n11739), .ZN(n13741) );
  AOI22_X1 U14201 ( .A1(n14080), .A2(n11740), .B1(n13741), .B2(n14034), .ZN(
        n11741) );
  OAI21_X1 U14202 ( .B1(n11742), .B2(n14080), .A(n11741), .ZN(n11745) );
  INV_X1 U14203 ( .A(n12041), .ZN(n13746) );
  OAI211_X1 U14204 ( .C1(n13746), .C2(n11520), .A(n11854), .B(n14493), .ZN(
        n11789) );
  NOR2_X1 U14205 ( .A1(n11789), .A2(n14085), .ZN(n11744) );
  AOI211_X1 U14206 ( .C1(n14082), .C2(n12041), .A(n11745), .B(n11744), .ZN(
        n11746) );
  OAI211_X1 U14207 ( .C1(n11790), .C2(n14042), .A(n11747), .B(n11746), .ZN(
        P1_U3278) );
  INV_X1 U14208 ( .A(n11752), .ZN(n11750) );
  NAND2_X1 U14209 ( .A1(n13593), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n11748) );
  OAI211_X1 U14210 ( .C1(n11750), .C2(n13596), .A(n11749), .B(n11748), .ZN(
        P2_U3304) );
  NAND2_X1 U14211 ( .A1(n11752), .A2(n11751), .ZN(n11754) );
  OAI211_X1 U14212 ( .C1(n11755), .C2(n14245), .A(n11754), .B(n11753), .ZN(
        P1_U3332) );
  XNOR2_X1 U14213 ( .A(n11756), .B(n11763), .ZN(n11758) );
  AOI21_X1 U14214 ( .B1(n11758), .B2(n14725), .A(n11757), .ZN(n13559) );
  AOI211_X1 U14215 ( .C1(n13557), .C2(n11760), .A(n11505), .B(n11759), .ZN(
        n13556) );
  AOI22_X1 U14216 ( .A1(n14736), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n11761), 
        .B2(n14705), .ZN(n11762) );
  OAI21_X1 U14217 ( .B1(n6886), .B2(n13453), .A(n11762), .ZN(n11766) );
  XNOR2_X1 U14218 ( .A(n11764), .B(n11763), .ZN(n13560) );
  NOR2_X1 U14219 ( .A1(n13560), .A2(n14715), .ZN(n11765) );
  AOI211_X1 U14220 ( .C1(n13556), .C2(n13473), .A(n11766), .B(n11765), .ZN(
        n11767) );
  OAI21_X1 U14221 ( .B1(n14736), .B2(n13559), .A(n11767), .ZN(P2_U3251) );
  INV_X1 U14222 ( .A(n11768), .ZN(n11769) );
  OAI222_X1 U14223 ( .A1(P3_U3151), .A2(n11771), .B1(n12303), .B2(n11770), 
        .C1(n13138), .C2(n11769), .ZN(P3_U3269) );
  OAI21_X1 U14224 ( .B1(n13279), .B2(n14822), .A(n11772), .ZN(n11774) );
  AOI211_X1 U14225 ( .C1(n11775), .C2(n14809), .A(n11774), .B(n11773), .ZN(
        n11778) );
  NAND2_X1 U14226 ( .A1(n14829), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n11776) );
  OAI21_X1 U14227 ( .B1(n11778), .B2(n14829), .A(n11776), .ZN(P2_U3475) );
  NAND2_X1 U14228 ( .A1(n14850), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n11777) );
  OAI21_X1 U14229 ( .B1(n11778), .B2(n14850), .A(n11777), .ZN(P2_U3514) );
  NAND2_X1 U14230 ( .A1(n7387), .A2(n11779), .ZN(n11780) );
  XNOR2_X1 U14231 ( .A(n11780), .B(n12693), .ZN(n11787) );
  AOI21_X1 U14232 ( .B1(n12694), .B2(n12663), .A(n11781), .ZN(n11785) );
  NAND2_X1 U14233 ( .A1(n12678), .A2(n14335), .ZN(n11784) );
  NAND2_X1 U14234 ( .A1(n12648), .A2(n14334), .ZN(n11783) );
  NAND2_X1 U14235 ( .A1(n12692), .A2(n12674), .ZN(n11782) );
  NAND4_X1 U14236 ( .A1(n11785), .A2(n11784), .A3(n11783), .A4(n11782), .ZN(
        n11786) );
  AOI21_X1 U14237 ( .B1(n11787), .B2(n12670), .A(n11786), .ZN(n11788) );
  INV_X1 U14238 ( .A(n11788), .ZN(P3_U3176) );
  OAI211_X1 U14239 ( .C1(n13746), .C2(n14528), .A(n11789), .B(n13738), .ZN(
        n11792) );
  NOR2_X1 U14240 ( .A1(n11790), .A2(n14534), .ZN(n11791) );
  AOI211_X1 U14241 ( .C1(n11793), .C2(n14430), .A(n11792), .B(n11791), .ZN(
        n11796) );
  NAND2_X1 U14242 ( .A1(n14547), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n11794) );
  OAI21_X1 U14243 ( .B1(n11796), .B2(n14547), .A(n11794), .ZN(P1_U3504) );
  NAND2_X1 U14244 ( .A1(n14558), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n11795) );
  OAI21_X1 U14245 ( .B1(n11796), .B2(n14558), .A(n11795), .ZN(P1_U3543) );
  NOR2_X1 U14246 ( .A1(n11811), .A2(n11797), .ZN(n11798) );
  AOI22_X1 U14247 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n12706), .B1(n12708), 
        .B2(n7696), .ZN(n11800) );
  AOI21_X1 U14248 ( .B1(n11801), .B2(n11800), .A(n12703), .ZN(n11822) );
  INV_X1 U14249 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14363) );
  AOI22_X1 U14250 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n12708), .B1(n12706), 
        .B2(n14363), .ZN(n11807) );
  NAND2_X1 U14251 ( .A1(n11803), .A2(n11802), .ZN(n11805) );
  NAND2_X1 U14252 ( .A1(n11805), .A2(n11804), .ZN(n11806) );
  OAI21_X1 U14253 ( .B1(n11807), .B2(n11806), .A(n12705), .ZN(n11820) );
  INV_X1 U14254 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11808) );
  NOR2_X1 U14255 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11808), .ZN(n11899) );
  AOI21_X1 U14256 ( .B1(n14969), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n11899), 
        .ZN(n11809) );
  OAI21_X1 U14257 ( .B1(n14966), .B2(n12708), .A(n11809), .ZN(n11819) );
  INV_X1 U14258 ( .A(n11810), .ZN(n11812) );
  NAND2_X1 U14259 ( .A1(n11812), .A2(n11811), .ZN(n11814) );
  MUX2_X1 U14260 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12776), .Z(n12709) );
  XNOR2_X1 U14261 ( .A(n12709), .B(n12706), .ZN(n11813) );
  NAND3_X1 U14262 ( .A1(n11815), .A2(n11814), .A3(n11813), .ZN(n12712) );
  INV_X1 U14263 ( .A(n12712), .ZN(n11817) );
  AOI21_X1 U14264 ( .B1(n11815), .B2(n11814), .A(n11813), .ZN(n11816) );
  NOR3_X1 U14265 ( .A1(n11817), .A2(n11816), .A3(n14985), .ZN(n11818) );
  AOI211_X1 U14266 ( .C1(n6467), .C2(n11820), .A(n11819), .B(n11818), .ZN(
        n11821) );
  OAI21_X1 U14267 ( .B1(n11822), .B2(n14991), .A(n11821), .ZN(P3_U3194) );
  XNOR2_X1 U14268 ( .A(n11823), .B(n12514), .ZN(n11824) );
  OAI222_X1 U14269 ( .A1(n14339), .A2(n14328), .B1(n14341), .B2(n11825), .C1(
        n11824), .C2(n15045), .ZN(n14360) );
  INV_X1 U14270 ( .A(n14360), .ZN(n11833) );
  OAI21_X1 U14271 ( .B1(n11828), .B2(n11827), .A(n11826), .ZN(n14362) );
  NAND2_X1 U14272 ( .A1(n11829), .A2(n15054), .ZN(n15019) );
  NAND2_X1 U14273 ( .A1(n15080), .A2(n15019), .ZN(n12960) );
  AOI22_X1 U14274 ( .A1(n15082), .A2(P3_REG2_REG_12__SCAN_IN), .B1(n15077), 
        .B2(n11898), .ZN(n11830) );
  OAI21_X1 U14275 ( .B1(n13007), .B2(n14359), .A(n11830), .ZN(n11831) );
  AOI21_X1 U14276 ( .B1(n14362), .B2(n14346), .A(n11831), .ZN(n11832) );
  OAI21_X1 U14277 ( .B1(n11833), .B2(n15082), .A(n11832), .ZN(P3_U3221) );
  AOI22_X1 U14278 ( .A1(n11851), .A2(n12282), .B1(n12275), .B2(n13766), .ZN(
        n11834) );
  XOR2_X1 U14279 ( .A(n12265), .B(n11834), .Z(n11845) );
  AOI22_X1 U14280 ( .A1(n11851), .A2(n12285), .B1(n12284), .B2(n13766), .ZN(
        n11838) );
  NAND2_X1 U14281 ( .A1(n11837), .A2(n11838), .ZN(n11876) );
  INV_X1 U14282 ( .A(n11838), .ZN(n11839) );
  NAND2_X1 U14283 ( .A1(n11840), .A2(n11839), .ZN(n11841) );
  INV_X1 U14284 ( .A(n11845), .ZN(n11843) );
  INV_X1 U14285 ( .A(n11877), .ZN(n11844) );
  AOI21_X1 U14286 ( .B1(n11845), .B2(n11842), .A(n11844), .ZN(n11853) );
  INV_X1 U14287 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n11846) );
  NOR2_X1 U14288 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11846), .ZN(n13826) );
  AOI21_X1 U14289 ( .B1(n14411), .B2(n11847), .A(n13826), .ZN(n11848) );
  OAI21_X1 U14290 ( .B1(n14417), .B2(n11849), .A(n11848), .ZN(n11850) );
  AOI21_X1 U14291 ( .B1(n11851), .B2(n6468), .A(n11850), .ZN(n11852) );
  OAI21_X1 U14292 ( .B1(n11853), .B2(n13731), .A(n11852), .ZN(P1_U3231) );
  AOI211_X1 U14293 ( .C1(n14189), .C2(n11854), .A(n14119), .B(n11924), .ZN(
        n14188) );
  OAI21_X1 U14294 ( .B1(n6589), .B2(n11856), .A(n11855), .ZN(n11858) );
  AOI22_X1 U14295 ( .A1(n13760), .A2(n13913), .B1(n13717), .B2(n13758), .ZN(
        n13657) );
  INV_X1 U14296 ( .A(n13657), .ZN(n11857) );
  AOI21_X1 U14297 ( .B1(n11858), .B2(n14526), .A(n11857), .ZN(n14191) );
  INV_X1 U14298 ( .A(n14191), .ZN(n11859) );
  AOI21_X1 U14299 ( .B1(n14188), .B2(n11860), .A(n11859), .ZN(n11868) );
  OAI21_X1 U14300 ( .B1(n11863), .B2(n11862), .A(n11861), .ZN(n14187) );
  NOR2_X1 U14301 ( .A1(n12049), .A2(n14482), .ZN(n11866) );
  OAI22_X1 U14302 ( .A1(n14080), .A2(n11864), .B1(n13655), .B2(n14477), .ZN(
        n11865) );
  AOI211_X1 U14303 ( .C1(n14187), .C2(n14092), .A(n11866), .B(n11865), .ZN(
        n11867) );
  OAI21_X1 U14304 ( .B1(n11868), .B2(n14479), .A(n11867), .ZN(P1_U3277) );
  NAND2_X1 U14305 ( .A1(n11883), .A2(n12282), .ZN(n11870) );
  NAND2_X1 U14306 ( .A1(n13765), .A2(n12275), .ZN(n11869) );
  NAND2_X1 U14307 ( .A1(n11870), .A2(n11869), .ZN(n11871) );
  XNOR2_X1 U14308 ( .A(n11871), .B(n12265), .ZN(n11875) );
  NAND2_X1 U14309 ( .A1(n11883), .A2(n12285), .ZN(n11873) );
  NAND2_X1 U14310 ( .A1(n12284), .A2(n13765), .ZN(n11872) );
  NAND2_X1 U14311 ( .A1(n11873), .A2(n11872), .ZN(n11874) );
  NOR2_X1 U14312 ( .A1(n11875), .A2(n11874), .ZN(n12005) );
  AND2_X1 U14313 ( .A1(n11875), .A2(n11874), .ZN(n14405) );
  NOR2_X1 U14314 ( .A1(n12005), .A2(n14405), .ZN(n11878) );
  XOR2_X1 U14315 ( .A(n11878), .B(n12004), .Z(n11885) );
  AOI22_X1 U14316 ( .A1(n14411), .A2(n11879), .B1(P1_REG3_REG_10__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11880) );
  OAI21_X1 U14317 ( .B1(n11881), .B2(n14417), .A(n11880), .ZN(n11882) );
  AOI21_X1 U14318 ( .B1(n11883), .B2(n6468), .A(n11882), .ZN(n11884) );
  OAI21_X1 U14319 ( .B1(n11885), .B2(n13731), .A(n11884), .ZN(P1_U3217) );
  INV_X1 U14320 ( .A(n11886), .ZN(n11888) );
  OAI222_X1 U14321 ( .A1(P3_U3151), .A2(n6473), .B1(n13138), .B2(n11888), .C1(
        n11887), .C2(n12303), .ZN(P3_U3268) );
  INV_X1 U14322 ( .A(n11889), .ZN(n13200) );
  XNOR2_X1 U14323 ( .A(n11890), .B(n11892), .ZN(n11891) );
  AOI22_X1 U14324 ( .A1(n13293), .A2(n13172), .B1(n13171), .B2(n13295), .ZN(
        n13198) );
  OAI21_X1 U14325 ( .B1(n11891), .B2(n13462), .A(n13198), .ZN(n13551) );
  AOI21_X1 U14326 ( .B1(n13200), .B2(n14705), .A(n13551), .ZN(n11897) );
  AOI211_X1 U14327 ( .C1(n13553), .C2(n6491), .A(n11505), .B(n11963), .ZN(
        n13552) );
  INV_X1 U14328 ( .A(n13553), .ZN(n13203) );
  INV_X1 U14329 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n12231) );
  OAI22_X1 U14330 ( .A1(n13203), .A2(n13453), .B1(n12231), .B2(n14733), .ZN(
        n11895) );
  XNOR2_X1 U14331 ( .A(n11893), .B(n11892), .ZN(n13555) );
  NOR2_X1 U14332 ( .A1(n13555), .A2(n14715), .ZN(n11894) );
  AOI211_X1 U14333 ( .C1(n13552), .C2(n13473), .A(n11895), .B(n11894), .ZN(
        n11896) );
  OAI21_X1 U14334 ( .B1(n14736), .B2(n11897), .A(n11896), .ZN(P2_U3249) );
  NAND2_X1 U14335 ( .A1(n12678), .A2(n11898), .ZN(n11901) );
  AOI21_X1 U14336 ( .B1(n12663), .B2(n12693), .A(n11899), .ZN(n11900) );
  OAI211_X1 U14337 ( .C1(n14328), .C2(n12665), .A(n11901), .B(n11900), .ZN(
        n11907) );
  XNOR2_X1 U14338 ( .A(n11902), .B(n12692), .ZN(n11903) );
  XNOR2_X1 U14339 ( .A(n11904), .B(n11903), .ZN(n11905) );
  NOR2_X1 U14340 ( .A1(n11905), .A2(n12650), .ZN(n11906) );
  AOI211_X1 U14341 ( .C1(n12648), .C2(n11908), .A(n11907), .B(n11906), .ZN(
        n11909) );
  INV_X1 U14342 ( .A(n11909), .ZN(P3_U3164) );
  XOR2_X1 U14343 ( .A(n12517), .B(n11910), .Z(n14355) );
  INV_X1 U14344 ( .A(n12690), .ZN(n13000) );
  XNOR2_X1 U14345 ( .A(n11911), .B(n12517), .ZN(n11912) );
  OAI222_X1 U14346 ( .A1(n14339), .A2(n13000), .B1(n14341), .B2(n14340), .C1(
        n11912), .C2(n15045), .ZN(n14357) );
  NAND2_X1 U14347 ( .A1(n14357), .A2(n15080), .ZN(n11918) );
  INV_X1 U14348 ( .A(n14353), .ZN(n11916) );
  INV_X1 U14349 ( .A(n11913), .ZN(n11914) );
  OAI22_X1 U14350 ( .A1(n15080), .A2(n7722), .B1(n11914), .B2(n15009), .ZN(
        n11915) );
  AOI21_X1 U14351 ( .B1(n11916), .B2(n15004), .A(n11915), .ZN(n11917) );
  OAI211_X1 U14352 ( .C1(n12960), .C2(n14355), .A(n11918), .B(n11917), .ZN(
        P3_U3220) );
  INV_X1 U14353 ( .A(n11922), .ZN(n11919) );
  XNOR2_X1 U14354 ( .A(n11920), .B(n11919), .ZN(n14181) );
  XOR2_X1 U14355 ( .A(n11922), .B(n11921), .Z(n14183) );
  NAND2_X1 U14356 ( .A1(n14183), .A2(n14092), .ZN(n11930) );
  INV_X1 U14357 ( .A(n14077), .ZN(n11923) );
  OAI211_X1 U14358 ( .C1(n14233), .C2(n11924), .A(n11923), .B(n14493), .ZN(
        n14179) );
  INV_X1 U14359 ( .A(n14179), .ZN(n11928) );
  OAI22_X1 U14360 ( .A1(n13625), .A2(n13633), .B1(n12048), .B2(n13624), .ZN(
        n13666) );
  INV_X1 U14361 ( .A(n13666), .ZN(n14180) );
  OAI22_X1 U14362 ( .A1(n14479), .A2(n14180), .B1(n13668), .B2(n14477), .ZN(
        n11925) );
  AOI21_X1 U14363 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n14479), .A(n11925), 
        .ZN(n11926) );
  OAI21_X1 U14364 ( .B1(n14233), .B2(n14482), .A(n11926), .ZN(n11927) );
  AOI21_X1 U14365 ( .B1(n11928), .B2(n14485), .A(n11927), .ZN(n11929) );
  OAI211_X1 U14366 ( .C1(n14181), .C2(n14042), .A(n11930), .B(n11929), .ZN(
        P1_U3276) );
  OAI211_X1 U14367 ( .C1(n11933), .C2(n11932), .A(n11931), .B(n12670), .ZN(
        n11938) );
  NOR2_X1 U14368 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11934), .ZN(n12732) );
  AOI21_X1 U14369 ( .B1(n12663), .B2(n12691), .A(n12732), .ZN(n11935) );
  OAI21_X1 U14370 ( .B1(n14329), .B2(n12665), .A(n11935), .ZN(n11936) );
  AOI21_X1 U14371 ( .B1(n14331), .B2(n12678), .A(n11936), .ZN(n11937) );
  OAI211_X1 U14372 ( .C1(n12681), .C2(n14330), .A(n11938), .B(n11937), .ZN(
        P3_U3155) );
  INV_X1 U14373 ( .A(n11939), .ZN(n11944) );
  OAI222_X1 U14374 ( .A1(n11941), .A2(P1_U3086), .B1(n14251), .B2(n11944), 
        .C1(n11940), .C2(n14245), .ZN(P1_U3331) );
  INV_X1 U14375 ( .A(n11942), .ZN(n11945) );
  OAI222_X1 U14376 ( .A1(n11945), .A2(P2_U3088), .B1(n13589), .B2(n11944), 
        .C1(n11943), .C2(n13591), .ZN(P2_U3303) );
  INV_X1 U14377 ( .A(n11946), .ZN(n13247) );
  XNOR2_X1 U14378 ( .A(n11947), .B(n6985), .ZN(n11948) );
  NAND2_X1 U14379 ( .A1(n11948), .A2(n14725), .ZN(n11950) );
  AND2_X1 U14380 ( .A1(n13293), .A2(n13171), .ZN(n11949) );
  AOI21_X1 U14381 ( .B1(n13291), .B2(n13172), .A(n11949), .ZN(n13245) );
  NAND2_X1 U14382 ( .A1(n11950), .A2(n13245), .ZN(n13544) );
  AOI21_X1 U14383 ( .B1(n13247), .B2(n14705), .A(n13544), .ZN(n11958) );
  NAND2_X1 U14384 ( .A1(n11952), .A2(n11951), .ZN(n11953) );
  NAND2_X1 U14385 ( .A1(n7397), .A2(n11953), .ZN(n13540) );
  OAI21_X1 U14386 ( .B1(n11964), .B2(n13543), .A(n11440), .ZN(n11954) );
  OR2_X1 U14387 ( .A1(n13465), .A2(n11954), .ZN(n13541) );
  AOI22_X1 U14388 ( .A1(n12171), .A2(n14706), .B1(n14736), .B2(
        P2_REG2_REG_18__SCAN_IN), .ZN(n11955) );
  OAI21_X1 U14389 ( .B1(n13541), .B2(n14714), .A(n11955), .ZN(n11956) );
  AOI21_X1 U14390 ( .B1(n13540), .B2(n13426), .A(n11956), .ZN(n11957) );
  OAI21_X1 U14391 ( .B1(n11958), .B2(n14736), .A(n11957), .ZN(P2_U3247) );
  XOR2_X1 U14392 ( .A(n11959), .B(n11968), .Z(n11962) );
  NAND2_X1 U14393 ( .A1(n13292), .A2(n13172), .ZN(n11961) );
  NAND2_X1 U14394 ( .A1(n13294), .A2(n13171), .ZN(n11960) );
  NAND2_X1 U14395 ( .A1(n11961), .A2(n11960), .ZN(n13209) );
  AOI21_X1 U14396 ( .B1(n11962), .B2(n14725), .A(n13209), .ZN(n13549) );
  INV_X1 U14397 ( .A(n11963), .ZN(n11965) );
  AOI211_X1 U14398 ( .C1(n13547), .C2(n11965), .A(n11505), .B(n11964), .ZN(
        n13546) );
  INV_X1 U14399 ( .A(n11966), .ZN(n13213) );
  AOI22_X1 U14400 ( .A1(n14736), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n13213), 
        .B2(n14705), .ZN(n11967) );
  OAI21_X1 U14401 ( .B1(n13216), .B2(n13453), .A(n11967), .ZN(n11973) );
  OR2_X1 U14402 ( .A1(n11969), .A2(n11968), .ZN(n11970) );
  NAND2_X1 U14403 ( .A1(n11971), .A2(n11970), .ZN(n13550) );
  NOR2_X1 U14404 ( .A1(n13550), .A2(n14715), .ZN(n11972) );
  AOI211_X1 U14405 ( .C1(n13546), .C2(n13473), .A(n11973), .B(n11972), .ZN(
        n11974) );
  OAI21_X1 U14406 ( .B1(n14736), .B2(n13549), .A(n11974), .ZN(P2_U3248) );
  INV_X1 U14407 ( .A(n11975), .ZN(n11979) );
  OAI222_X1 U14408 ( .A1(n13591), .A2(n11977), .B1(n13589), .B2(n11979), .C1(
        n11976), .C2(P2_U3088), .ZN(P2_U3302) );
  OAI222_X1 U14409 ( .A1(P1_U3086), .A2(n11980), .B1(n14251), .B2(n11979), 
        .C1(n11978), .C2(n14245), .ZN(P1_U3330) );
  XNOR2_X1 U14410 ( .A(n11982), .B(n11981), .ZN(n11989) );
  NAND2_X1 U14411 ( .A1(n11984), .A2(n11983), .ZN(n11985) );
  NAND2_X1 U14412 ( .A1(n11986), .A2(n11985), .ZN(n14531) );
  NAND2_X1 U14413 ( .A1(n14531), .A2(n14546), .ZN(n11988) );
  OAI211_X1 U14414 ( .C1(n14534), .C2(n11989), .A(n11988), .B(n11987), .ZN(
        n14529) );
  MUX2_X1 U14415 ( .A(n14529), .B(P1_REG2_REG_5__SCAN_IN), .S(n14491), .Z(
        n12000) );
  AOI21_X1 U14416 ( .B1(n11991), .B2(n11990), .A(n14119), .ZN(n11993) );
  NAND2_X1 U14417 ( .A1(n11993), .A2(n11992), .ZN(n14527) );
  NAND2_X1 U14418 ( .A1(n14531), .A2(n14486), .ZN(n11998) );
  INV_X1 U14419 ( .A(n11994), .ZN(n11995) );
  OAI22_X1 U14420 ( .A1(n14482), .A2(n6627), .B1(n14477), .B2(n11995), .ZN(
        n11996) );
  INV_X1 U14421 ( .A(n11996), .ZN(n11997) );
  OAI211_X1 U14422 ( .C1(n14085), .C2(n14527), .A(n11998), .B(n11997), .ZN(
        n11999) );
  OR2_X1 U14423 ( .A1(n12000), .A2(n11999), .ZN(P1_U3288) );
  NAND2_X1 U14424 ( .A1(n13751), .A2(n13913), .ZN(n12002) );
  NAND2_X1 U14425 ( .A1(n13749), .A2(n13717), .ZN(n12001) );
  NAND2_X1 U14426 ( .A1(n12002), .A2(n12001), .ZN(n13968) );
  AOI22_X1 U14427 ( .A1(n14411), .A2(n13968), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12003) );
  OAI21_X1 U14428 ( .B1(n13969), .B2(n14417), .A(n12003), .ZN(n12138) );
  OAI22_X1 U14429 ( .A1(n14426), .A2(n12090), .B1(n12007), .B2(n12092), .ZN(
        n12008) );
  XNOR2_X1 U14430 ( .A(n12008), .B(n12265), .ZN(n12013) );
  OR2_X1 U14431 ( .A1(n14426), .A2(n12092), .ZN(n12010) );
  NAND2_X1 U14432 ( .A1(n13764), .A2(n12284), .ZN(n12009) );
  NAND2_X1 U14433 ( .A1(n12010), .A2(n12009), .ZN(n12012) );
  XNOR2_X1 U14434 ( .A(n12013), .B(n12012), .ZN(n14404) );
  NOR2_X1 U14435 ( .A1(n14404), .A2(n14405), .ZN(n12011) );
  OR2_X1 U14436 ( .A1(n12013), .A2(n12012), .ZN(n12014) );
  OAI22_X1 U14437 ( .A1(n13652), .A2(n12090), .B1(n12016), .B2(n12092), .ZN(
        n12015) );
  XNOR2_X1 U14438 ( .A(n12015), .B(n12265), .ZN(n12019) );
  OAI22_X1 U14439 ( .A1(n13652), .A2(n12092), .B1(n12016), .B2(n12125), .ZN(
        n12018) );
  XNOR2_X1 U14440 ( .A(n12019), .B(n12018), .ZN(n13641) );
  NAND2_X1 U14441 ( .A1(n12019), .A2(n12018), .ZN(n12020) );
  OAI22_X1 U14442 ( .A1(n13702), .A2(n12090), .B1(n12022), .B2(n12092), .ZN(
        n12021) );
  XNOR2_X1 U14443 ( .A(n12021), .B(n12265), .ZN(n12031) );
  NOR2_X1 U14444 ( .A1(n12022), .A2(n12125), .ZN(n12023) );
  AOI21_X1 U14445 ( .B1(n12024), .B2(n12285), .A(n12023), .ZN(n12032) );
  XNOR2_X1 U14446 ( .A(n12031), .B(n12032), .ZN(n13694) );
  NAND2_X1 U14447 ( .A1(n14419), .A2(n12282), .ZN(n12026) );
  NAND2_X1 U14448 ( .A1(n13761), .A2(n12275), .ZN(n12025) );
  NAND2_X1 U14449 ( .A1(n12026), .A2(n12025), .ZN(n12028) );
  XNOR2_X1 U14450 ( .A(n12028), .B(n12027), .ZN(n12036) );
  NOR2_X1 U14451 ( .A1(n12125), .A2(n12029), .ZN(n12030) );
  AOI21_X1 U14452 ( .B1(n14419), .B2(n12275), .A(n12030), .ZN(n12035) );
  XNOR2_X1 U14453 ( .A(n12036), .B(n12035), .ZN(n14394) );
  INV_X1 U14454 ( .A(n12031), .ZN(n12033) );
  NOR2_X1 U14455 ( .A1(n12033), .A2(n12032), .ZN(n14395) );
  NOR2_X1 U14456 ( .A1(n14394), .A2(n14395), .ZN(n12034) );
  NAND2_X1 U14457 ( .A1(n14393), .A2(n12034), .ZN(n14397) );
  NAND2_X1 U14458 ( .A1(n12036), .A2(n12035), .ZN(n12037) );
  NAND2_X1 U14459 ( .A1(n14397), .A2(n12037), .ZN(n12044) );
  NAND2_X1 U14460 ( .A1(n12041), .A2(n12282), .ZN(n12039) );
  NAND2_X1 U14461 ( .A1(n13760), .A2(n12285), .ZN(n12038) );
  NAND2_X1 U14462 ( .A1(n12039), .A2(n12038), .ZN(n12040) );
  XNOR2_X1 U14463 ( .A(n12040), .B(n12265), .ZN(n12042) );
  XNOR2_X1 U14464 ( .A(n12044), .B(n12042), .ZN(n13734) );
  AOI22_X1 U14465 ( .A1(n12041), .A2(n12285), .B1(n12284), .B2(n13760), .ZN(
        n13735) );
  INV_X1 U14466 ( .A(n12042), .ZN(n12043) );
  NAND2_X1 U14467 ( .A1(n12044), .A2(n12043), .ZN(n12045) );
  NAND2_X1 U14468 ( .A1(n13733), .A2(n12045), .ZN(n13653) );
  OR2_X1 U14469 ( .A1(n12049), .A2(n12092), .ZN(n12047) );
  NAND2_X1 U14470 ( .A1(n13759), .A2(n12284), .ZN(n12046) );
  NAND2_X1 U14471 ( .A1(n12047), .A2(n12046), .ZN(n12052) );
  OAI22_X1 U14472 ( .A1(n12049), .A2(n12090), .B1(n12048), .B2(n12092), .ZN(
        n12050) );
  XNOR2_X1 U14473 ( .A(n12050), .B(n12265), .ZN(n12051) );
  XOR2_X1 U14474 ( .A(n12052), .B(n12051), .Z(n13654) );
  INV_X1 U14475 ( .A(n12051), .ZN(n12054) );
  INV_X1 U14476 ( .A(n12052), .ZN(n12053) );
  NAND2_X1 U14477 ( .A1(n12054), .A2(n12053), .ZN(n12055) );
  NAND2_X1 U14478 ( .A1(n13670), .A2(n12282), .ZN(n12058) );
  NAND2_X1 U14479 ( .A1(n13758), .A2(n12275), .ZN(n12057) );
  NAND2_X1 U14480 ( .A1(n12058), .A2(n12057), .ZN(n12059) );
  XNOR2_X1 U14481 ( .A(n12059), .B(n12265), .ZN(n13663) );
  NAND2_X1 U14482 ( .A1(n13670), .A2(n12285), .ZN(n12061) );
  NAND2_X1 U14483 ( .A1(n12284), .A2(n13758), .ZN(n12060) );
  NAND2_X1 U14484 ( .A1(n12061), .A2(n12060), .ZN(n13662) );
  NAND2_X1 U14485 ( .A1(n13663), .A2(n13662), .ZN(n12062) );
  OAI22_X1 U14486 ( .A1(n14228), .A2(n12090), .B1(n13625), .B2(n12092), .ZN(
        n12063) );
  XNOR2_X1 U14487 ( .A(n12063), .B(n12265), .ZN(n12071) );
  OAI22_X1 U14488 ( .A1(n14228), .A2(n12092), .B1(n13625), .B2(n12125), .ZN(
        n12070) );
  XNOR2_X1 U14489 ( .A(n12071), .B(n12070), .ZN(n13715) );
  NAND2_X1 U14490 ( .A1(n12069), .A2(n12282), .ZN(n12065) );
  NAND2_X1 U14491 ( .A1(n13756), .A2(n12285), .ZN(n12064) );
  NAND2_X1 U14492 ( .A1(n12065), .A2(n12064), .ZN(n12067) );
  XNOR2_X1 U14493 ( .A(n12067), .B(n12027), .ZN(n12072) );
  AND2_X1 U14494 ( .A1(n13756), .A2(n12284), .ZN(n12068) );
  AOI21_X1 U14495 ( .B1(n12069), .B2(n12275), .A(n12068), .ZN(n12073) );
  XNOR2_X1 U14496 ( .A(n12072), .B(n12073), .ZN(n13620) );
  NOR2_X1 U14497 ( .A1(n12071), .A2(n12070), .ZN(n13621) );
  INV_X1 U14498 ( .A(n12072), .ZN(n12075) );
  INV_X1 U14499 ( .A(n12073), .ZN(n12074) );
  AND2_X1 U14500 ( .A1(n13755), .A2(n12284), .ZN(n12076) );
  AOI21_X1 U14501 ( .B1(n14222), .B2(n12285), .A(n12076), .ZN(n12079) );
  AOI22_X1 U14502 ( .A1(n14222), .A2(n12282), .B1(n12275), .B2(n13755), .ZN(
        n12077) );
  XNOR2_X1 U14503 ( .A(n12077), .B(n12265), .ZN(n12078) );
  XOR2_X1 U14504 ( .A(n12079), .B(n12078), .Z(n13685) );
  INV_X1 U14505 ( .A(n12078), .ZN(n12081) );
  INV_X1 U14506 ( .A(n12079), .ZN(n12080) );
  NAND2_X1 U14507 ( .A1(n12081), .A2(n12080), .ZN(n12082) );
  NAND2_X1 U14508 ( .A1(n14155), .A2(n12282), .ZN(n12085) );
  NAND2_X1 U14509 ( .A1(n13754), .A2(n12275), .ZN(n12084) );
  NAND2_X1 U14510 ( .A1(n12085), .A2(n12084), .ZN(n12086) );
  XNOR2_X1 U14511 ( .A(n12086), .B(n12027), .ZN(n12089) );
  AND2_X1 U14512 ( .A1(n13754), .A2(n12284), .ZN(n12087) );
  AOI21_X1 U14513 ( .B1(n14155), .B2(n12285), .A(n12087), .ZN(n12088) );
  NAND2_X1 U14514 ( .A1(n12089), .A2(n12088), .ZN(n13703) );
  OAI21_X1 U14515 ( .B1(n12089), .B2(n12088), .A(n13703), .ZN(n13632) );
  OAI22_X1 U14516 ( .A1(n14218), .A2(n12090), .B1(n13634), .B2(n12092), .ZN(
        n12091) );
  XNOR2_X1 U14517 ( .A(n12091), .B(n12027), .ZN(n12095) );
  OR2_X1 U14518 ( .A1(n14218), .A2(n12092), .ZN(n12094) );
  NAND2_X1 U14519 ( .A1(n13753), .A2(n12284), .ZN(n12093) );
  AND2_X1 U14520 ( .A1(n12094), .A2(n12093), .ZN(n12096) );
  NAND2_X1 U14521 ( .A1(n12095), .A2(n12096), .ZN(n13615) );
  INV_X1 U14522 ( .A(n12095), .ZN(n12098) );
  INV_X1 U14523 ( .A(n12096), .ZN(n12097) );
  NAND2_X1 U14524 ( .A1(n12098), .A2(n12097), .ZN(n12099) );
  NAND2_X1 U14525 ( .A1(n14142), .A2(n12282), .ZN(n12101) );
  NAND2_X1 U14526 ( .A1(n13752), .A2(n12285), .ZN(n12100) );
  NAND2_X1 U14527 ( .A1(n12101), .A2(n12100), .ZN(n12102) );
  XNOR2_X1 U14528 ( .A(n12102), .B(n12027), .ZN(n12105) );
  NOR2_X1 U14529 ( .A1(n12103), .A2(n12125), .ZN(n12104) );
  AOI21_X1 U14530 ( .B1(n14142), .B2(n12285), .A(n12104), .ZN(n12106) );
  NAND2_X1 U14531 ( .A1(n12105), .A2(n12106), .ZN(n13677) );
  INV_X1 U14532 ( .A(n12105), .ZN(n12108) );
  INV_X1 U14533 ( .A(n12106), .ZN(n12107) );
  NAND2_X1 U14534 ( .A1(n12108), .A2(n12107), .ZN(n12109) );
  NAND2_X1 U14535 ( .A1(n14212), .A2(n12282), .ZN(n12111) );
  NAND2_X1 U14536 ( .A1(n13751), .A2(n12275), .ZN(n12110) );
  NAND2_X1 U14537 ( .A1(n12111), .A2(n12110), .ZN(n12112) );
  XNOR2_X1 U14538 ( .A(n12112), .B(n12027), .ZN(n12115) );
  NOR2_X1 U14539 ( .A1(n12113), .A2(n12125), .ZN(n12114) );
  AOI21_X1 U14540 ( .B1(n14212), .B2(n12275), .A(n12114), .ZN(n12116) );
  NAND2_X1 U14541 ( .A1(n12115), .A2(n12116), .ZN(n12136) );
  INV_X1 U14542 ( .A(n12115), .ZN(n12118) );
  INV_X1 U14543 ( .A(n12116), .ZN(n12117) );
  NAND2_X1 U14544 ( .A1(n12118), .A2(n12117), .ZN(n12119) );
  AND2_X1 U14545 ( .A1(n12136), .A2(n12119), .ZN(n12121) );
  AND2_X1 U14546 ( .A1(n13613), .A2(n12121), .ZN(n12120) );
  INV_X1 U14547 ( .A(n12121), .ZN(n13676) );
  OR2_X1 U14548 ( .A1(n13676), .A2(n13677), .ZN(n12133) );
  AND2_X1 U14549 ( .A1(n12136), .A2(n12133), .ZN(n12259) );
  NAND2_X1 U14550 ( .A1(n12262), .A2(n12259), .ZN(n12132) );
  NAND2_X1 U14551 ( .A1(n14208), .A2(n12282), .ZN(n12123) );
  NAND2_X1 U14552 ( .A1(n13750), .A2(n12275), .ZN(n12122) );
  NAND2_X1 U14553 ( .A1(n12123), .A2(n12122), .ZN(n12124) );
  XNOR2_X1 U14554 ( .A(n12124), .B(n12027), .ZN(n12128) );
  NOR2_X1 U14555 ( .A1(n12126), .A2(n12125), .ZN(n12127) );
  AOI21_X1 U14556 ( .B1(n14208), .B2(n12275), .A(n12127), .ZN(n12129) );
  NAND2_X1 U14557 ( .A1(n12128), .A2(n12129), .ZN(n12258) );
  INV_X1 U14558 ( .A(n12128), .ZN(n12131) );
  INV_X1 U14559 ( .A(n12129), .ZN(n12130) );
  NAND2_X1 U14560 ( .A1(n12131), .A2(n12130), .ZN(n12260) );
  AND2_X1 U14561 ( .A1(n12258), .A2(n12260), .ZN(n12134) );
  NAND2_X1 U14562 ( .A1(n12132), .A2(n12134), .ZN(n12137) );
  INV_X1 U14563 ( .A(n12134), .ZN(n12135) );
  XOR2_X1 U14564 ( .A(n12140), .B(n12139), .Z(n12149) );
  NAND2_X1 U14565 ( .A1(n13827), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n12141) );
  OAI211_X1 U14566 ( .C1(n13806), .C2(n12143), .A(n12142), .B(n12141), .ZN(
        n12148) );
  AOI211_X1 U14567 ( .C1(n12146), .C2(n12145), .A(n12144), .B(n13880), .ZN(
        n12147) );
  AOI211_X1 U14568 ( .C1(n13883), .C2(n12149), .A(n12148), .B(n12147), .ZN(
        n12156) );
  NAND2_X1 U14569 ( .A1(n14256), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n13783) );
  INV_X1 U14570 ( .A(n12150), .ZN(n12151) );
  MUX2_X1 U14571 ( .A(n13783), .B(n12151), .S(n14248), .Z(n12155) );
  NAND2_X1 U14572 ( .A1(n12153), .A2(n12152), .ZN(n12154) );
  OAI211_X1 U14573 ( .C1(n12155), .C2(n6483), .A(n13775), .B(n12154), .ZN(
        n13804) );
  NAND2_X1 U14574 ( .A1(n12156), .A2(n13804), .ZN(P1_U3247) );
  NAND2_X1 U14575 ( .A1(n12158), .A2(n12157), .ZN(n12159) );
  NAND2_X1 U14576 ( .A1(n12160), .A2(n12159), .ZN(n12162) );
  XOR2_X1 U14577 ( .A(n12209), .B(n12161), .Z(n12163) );
  NAND2_X1 U14578 ( .A1(n13295), .A2(n11505), .ZN(n13268) );
  INV_X1 U14579 ( .A(n12162), .ZN(n12165) );
  INV_X1 U14580 ( .A(n12163), .ZN(n12164) );
  NOR2_X2 U14581 ( .A1(n13266), .A2(n7373), .ZN(n13195) );
  XNOR2_X1 U14582 ( .A(n13553), .B(n12209), .ZN(n12166) );
  NAND2_X1 U14583 ( .A1(n13294), .A2(n11505), .ZN(n12167) );
  XNOR2_X1 U14584 ( .A(n12166), .B(n12167), .ZN(n13194) );
  INV_X1 U14585 ( .A(n12166), .ZN(n12168) );
  NAND2_X1 U14586 ( .A1(n12168), .A2(n12167), .ZN(n13204) );
  XNOR2_X1 U14587 ( .A(n13547), .B(n12199), .ZN(n12170) );
  NAND2_X1 U14588 ( .A1(n13293), .A2(n11505), .ZN(n12169) );
  XNOR2_X1 U14589 ( .A(n12170), .B(n12169), .ZN(n13205) );
  XNOR2_X1 U14590 ( .A(n12171), .B(n12199), .ZN(n12173) );
  NAND2_X1 U14591 ( .A1(n13292), .A2(n11505), .ZN(n12172) );
  NOR2_X1 U14592 ( .A1(n12173), .A2(n12172), .ZN(n12174) );
  AOI21_X1 U14593 ( .B1(n12173), .B2(n12172), .A(n12174), .ZN(n13243) );
  INV_X1 U14594 ( .A(n12174), .ZN(n12175) );
  NAND2_X1 U14595 ( .A1(n13242), .A2(n12175), .ZN(n13169) );
  NAND2_X1 U14596 ( .A1(n13291), .A2(n11505), .ZN(n12177) );
  XNOR2_X1 U14597 ( .A(n13537), .B(n12209), .ZN(n12176) );
  XOR2_X1 U14598 ( .A(n12177), .B(n12176), .Z(n13170) );
  INV_X1 U14599 ( .A(n12176), .ZN(n12178) );
  XNOR2_X1 U14600 ( .A(n13531), .B(n12199), .ZN(n12180) );
  NAND2_X1 U14601 ( .A1(n13290), .A2(n11505), .ZN(n12179) );
  NOR2_X1 U14602 ( .A1(n12180), .A2(n12179), .ZN(n13224) );
  NAND2_X1 U14603 ( .A1(n13289), .A2(n11505), .ZN(n12182) );
  XNOR2_X1 U14604 ( .A(n13526), .B(n12209), .ZN(n12181) );
  XOR2_X1 U14605 ( .A(n12182), .B(n12181), .Z(n13178) );
  XNOR2_X1 U14606 ( .A(n13518), .B(n12209), .ZN(n12184) );
  NOR2_X1 U14607 ( .A1(n13180), .A2(n11440), .ZN(n13232) );
  AOI21_X2 U14608 ( .B1(n13233), .B2(n13232), .A(n7388), .ZN(n12188) );
  XNOR2_X1 U14609 ( .A(n13514), .B(n12209), .ZN(n12186) );
  NOR2_X1 U14610 ( .A1(n13234), .A2(n11440), .ZN(n13153) );
  INV_X1 U14611 ( .A(n12186), .ZN(n12187) );
  NOR2_X1 U14612 ( .A1(n12188), .A2(n12187), .ZN(n12189) );
  XNOR2_X1 U14613 ( .A(n13507), .B(n12209), .ZN(n12190) );
  NOR2_X1 U14614 ( .A1(n13187), .A2(n11440), .ZN(n12191) );
  XNOR2_X1 U14615 ( .A(n12190), .B(n12191), .ZN(n13218) );
  NAND2_X1 U14616 ( .A1(n12190), .A2(n12191), .ZN(n12192) );
  OAI21_X2 U14617 ( .B1(n13217), .B2(n13218), .A(n12192), .ZN(n13185) );
  XNOR2_X1 U14618 ( .A(n13382), .B(n12209), .ZN(n12194) );
  NOR2_X1 U14619 ( .A1(n13255), .A2(n11440), .ZN(n12195) );
  XNOR2_X1 U14620 ( .A(n12194), .B(n12195), .ZN(n13186) );
  NAND2_X1 U14621 ( .A1(n13185), .A2(n13186), .ZN(n12198) );
  INV_X1 U14622 ( .A(n12194), .ZN(n12196) );
  NAND2_X1 U14623 ( .A1(n12196), .A2(n12195), .ZN(n12197) );
  NAND2_X1 U14624 ( .A1(n12198), .A2(n12197), .ZN(n13250) );
  INV_X1 U14625 ( .A(n13250), .ZN(n12203) );
  XNOR2_X1 U14626 ( .A(n13497), .B(n12199), .ZN(n12201) );
  NAND2_X1 U14627 ( .A1(n13284), .A2(n11505), .ZN(n12200) );
  NAND2_X1 U14628 ( .A1(n12201), .A2(n12200), .ZN(n12204) );
  OAI21_X1 U14629 ( .B1(n12201), .B2(n12200), .A(n12204), .ZN(n13253) );
  INV_X1 U14630 ( .A(n13253), .ZN(n12202) );
  NAND2_X1 U14631 ( .A1(n13283), .A2(n11505), .ZN(n12206) );
  XNOR2_X1 U14632 ( .A(n13492), .B(n12209), .ZN(n12205) );
  XOR2_X1 U14633 ( .A(n12206), .B(n12205), .Z(n13144) );
  INV_X1 U14634 ( .A(n12205), .ZN(n12207) );
  NAND2_X1 U14635 ( .A1(n13282), .A2(n11505), .ZN(n12208) );
  XOR2_X1 U14636 ( .A(n12209), .B(n12208), .Z(n12210) );
  XNOR2_X1 U14637 ( .A(n13341), .B(n12210), .ZN(n12211) );
  INV_X1 U14638 ( .A(n12212), .ZN(n13342) );
  NAND2_X1 U14639 ( .A1(n13283), .A2(n13171), .ZN(n12213) );
  OAI21_X1 U14640 ( .B1(n12214), .B2(n13256), .A(n12213), .ZN(n13335) );
  AOI22_X1 U14641 ( .A1(n13257), .A2(n13335), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12215) );
  OAI21_X1 U14642 ( .B1(n13342), .B2(n13259), .A(n12215), .ZN(n12216) );
  AOI21_X1 U14643 ( .B1(n13487), .B2(n13262), .A(n12216), .ZN(n12217) );
  INV_X1 U14644 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n12218) );
  NAND3_X1 U14645 ( .A1(n12218), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n12223) );
  NAND2_X1 U14646 ( .A1(n12219), .A2(n12220), .ZN(n12222) );
  NAND2_X1 U14647 ( .A1(n13593), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n12221) );
  OAI211_X1 U14648 ( .C1(n7128), .C2(n12223), .A(n12222), .B(n12221), .ZN(
        P2_U3296) );
  INV_X1 U14649 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n12232) );
  NOR2_X1 U14650 ( .A1(n12245), .A2(n12232), .ZN(n12224) );
  AOI21_X1 U14651 ( .B1(n12232), .B2(n12245), .A(n12224), .ZN(n14694) );
  XNOR2_X1 U14652 ( .A(n12236), .B(n12231), .ZN(n14675) );
  NOR2_X1 U14653 ( .A1(n12226), .A2(n12225), .ZN(n12228) );
  NOR2_X1 U14654 ( .A1(n12228), .A2(n12227), .ZN(n12229) );
  NAND2_X1 U14655 ( .A1(n14662), .A2(n12229), .ZN(n12230) );
  XOR2_X1 U14656 ( .A(n14662), .B(n12229), .Z(n14664) );
  NAND2_X1 U14657 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n14664), .ZN(n14663) );
  NAND2_X1 U14658 ( .A1(n12230), .A2(n14663), .ZN(n14676) );
  NAND2_X1 U14659 ( .A1(n14675), .A2(n14676), .ZN(n14674) );
  OAI21_X1 U14660 ( .B1(n14671), .B2(n12231), .A(n14674), .ZN(n14693) );
  NAND2_X1 U14661 ( .A1(n14694), .A2(n14693), .ZN(n14691) );
  OAI21_X1 U14662 ( .B1(n12245), .B2(n12232), .A(n14691), .ZN(n12233) );
  NOR2_X1 U14663 ( .A1(n13318), .A2(n12233), .ZN(n12234) );
  XNOR2_X1 U14664 ( .A(n13318), .B(n12233), .ZN(n13312) );
  NOR2_X1 U14665 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n13312), .ZN(n13311) );
  NOR2_X1 U14666 ( .A1(n12234), .A2(n13311), .ZN(n12235) );
  XOR2_X1 U14667 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n12235), .Z(n12252) );
  INV_X1 U14668 ( .A(n12252), .ZN(n12250) );
  INV_X1 U14669 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n12244) );
  XNOR2_X1 U14670 ( .A(n12245), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n14690) );
  INV_X1 U14671 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n12243) );
  XOR2_X1 U14672 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n12236), .Z(n14678) );
  INV_X1 U14673 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n12238) );
  NAND2_X1 U14674 ( .A1(n14662), .A2(n12240), .ZN(n12242) );
  XNOR2_X1 U14675 ( .A(n12241), .B(n12240), .ZN(n14666) );
  NAND2_X1 U14676 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n14666), .ZN(n14665) );
  NAND2_X1 U14677 ( .A1(n12242), .A2(n14665), .ZN(n14679) );
  NAND2_X1 U14678 ( .A1(n14690), .A2(n14689), .ZN(n14687) );
  OAI21_X1 U14679 ( .B1(n12245), .B2(n12244), .A(n14687), .ZN(n12247) );
  INV_X1 U14680 ( .A(n12247), .ZN(n12246) );
  XNOR2_X1 U14681 ( .A(n13318), .B(n12246), .ZN(n13317) );
  NAND2_X1 U14682 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n13317), .ZN(n13316) );
  NAND2_X1 U14683 ( .A1(n13318), .A2(n12247), .ZN(n12248) );
  NOR2_X1 U14684 ( .A1(n12251), .A2(n14595), .ZN(n12249) );
  AOI211_X1 U14685 ( .C1(n12250), .C2(n14692), .A(n14685), .B(n12249), .ZN(
        n12254) );
  AOI22_X1 U14686 ( .A1(n12252), .A2(n14692), .B1(n14688), .B2(n12251), .ZN(
        n12253) );
  MUX2_X1 U14687 ( .A(n12254), .B(n12253), .S(n14720), .Z(n12255) );
  NAND2_X1 U14688 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13174)
         );
  OAI211_X1 U14689 ( .C1(n12256), .C2(n14647), .A(n12255), .B(n13174), .ZN(
        P2_U3233) );
  INV_X1 U14690 ( .A(n12257), .ZN(n13580) );
  OAI222_X1 U14691 ( .A1(P1_U3086), .A2(n6474), .B1(n14251), .B2(n13580), .C1(
        n12301), .C2(n14245), .ZN(P1_U3325) );
  AND2_X1 U14692 ( .A1(n12259), .A2(n12258), .ZN(n12261) );
  NAND2_X1 U14693 ( .A1(n14117), .A2(n12282), .ZN(n12264) );
  NAND2_X1 U14694 ( .A1(n13749), .A2(n12285), .ZN(n12263) );
  NAND2_X1 U14695 ( .A1(n12264), .A2(n12263), .ZN(n12266) );
  XNOR2_X1 U14696 ( .A(n12266), .B(n12265), .ZN(n12270) );
  NAND2_X1 U14697 ( .A1(n14117), .A2(n12285), .ZN(n12268) );
  NAND2_X1 U14698 ( .A1(n12284), .A2(n13749), .ZN(n12267) );
  NAND2_X1 U14699 ( .A1(n12268), .A2(n12267), .ZN(n12269) );
  NOR2_X1 U14700 ( .A1(n12270), .A2(n12269), .ZN(n12271) );
  AOI21_X1 U14701 ( .B1(n12270), .B2(n12269), .A(n12271), .ZN(n13724) );
  NAND2_X1 U14702 ( .A1(n14203), .A2(n12282), .ZN(n12273) );
  NAND2_X1 U14703 ( .A1(n13748), .A2(n12275), .ZN(n12272) );
  NAND2_X1 U14704 ( .A1(n12273), .A2(n12272), .ZN(n12274) );
  XNOR2_X1 U14705 ( .A(n12274), .B(n12265), .ZN(n12279) );
  NAND2_X1 U14706 ( .A1(n14203), .A2(n12275), .ZN(n12277) );
  NAND2_X1 U14707 ( .A1(n12284), .A2(n13748), .ZN(n12276) );
  NAND2_X1 U14708 ( .A1(n12277), .A2(n12276), .ZN(n12278) );
  NOR2_X1 U14709 ( .A1(n12279), .A2(n12278), .ZN(n12280) );
  AOI21_X1 U14710 ( .B1(n12279), .B2(n12278), .A(n12280), .ZN(n13601) );
  INV_X1 U14711 ( .A(n12280), .ZN(n12281) );
  NAND2_X1 U14712 ( .A1(n13600), .A2(n12281), .ZN(n12289) );
  AOI22_X1 U14713 ( .A1(n13926), .A2(n12282), .B1(n12285), .B2(n13914), .ZN(
        n12283) );
  XNOR2_X1 U14714 ( .A(n12283), .B(n12265), .ZN(n12287) );
  AOI22_X1 U14715 ( .A1(n13926), .A2(n12285), .B1(n12284), .B2(n13914), .ZN(
        n12286) );
  XNOR2_X1 U14716 ( .A(n12287), .B(n12286), .ZN(n12288) );
  XNOR2_X1 U14717 ( .A(n12289), .B(n12288), .ZN(n12295) );
  NOR2_X1 U14718 ( .A1(n14417), .A2(n13924), .ZN(n12293) );
  OAI22_X1 U14719 ( .A1(n13739), .A2(n12291), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12290), .ZN(n12292) );
  AOI211_X1 U14720 ( .C1(n13926), .C2(n6468), .A(n12293), .B(n12292), .ZN(
        n12294) );
  OAI21_X1 U14721 ( .B1(n12295), .B2(n13731), .A(n12294), .ZN(P1_U3220) );
  INV_X1 U14722 ( .A(n12296), .ZN(n13586) );
  OAI222_X1 U14723 ( .A1(n6483), .A2(P1_U3086), .B1(n14251), .B2(n13586), .C1(
        n12297), .C2(n14245), .ZN(P1_U3327) );
  INV_X1 U14724 ( .A(n12298), .ZN(n12299) );
  INV_X1 U14725 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13582) );
  INV_X1 U14726 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13578) );
  NAND2_X1 U14727 ( .A1(n13578), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12307) );
  NAND2_X1 U14728 ( .A1(n12301), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12302) );
  NAND2_X1 U14729 ( .A1(n12307), .A2(n12302), .ZN(n12308) );
  XNOR2_X1 U14730 ( .A(n12309), .B(n12308), .ZN(n12323) );
  INV_X1 U14731 ( .A(n12323), .ZN(n12304) );
  INV_X1 U14732 ( .A(SI_30_), .ZN(n12324) );
  OAI222_X1 U14733 ( .A1(P3_U3151), .A2(n7475), .B1(n13138), .B2(n12304), .C1(
        n12324), .C2(n12303), .ZN(P3_U3265) );
  INV_X1 U14734 ( .A(n12305), .ZN(n12306) );
  OAI21_X1 U14735 ( .B1(n12309), .B2(n12308), .A(n12307), .ZN(n12311) );
  XNOR2_X1 U14736 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n12310) );
  XNOR2_X1 U14737 ( .A(n12311), .B(n12310), .ZN(n13127) );
  INV_X1 U14738 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n12313) );
  OR2_X1 U14739 ( .A1(n12314), .A2(n12313), .ZN(n12320) );
  NAND2_X1 U14740 ( .A1(n12315), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12319) );
  INV_X1 U14741 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n12316) );
  OR2_X1 U14742 ( .A1(n12317), .A2(n12316), .ZN(n12318) );
  NAND4_X1 U14743 ( .A1(n12321), .A2(n12320), .A3(n12319), .A4(n12318), .ZN(
        n12835) );
  INV_X1 U14744 ( .A(n12835), .ZN(n12327) );
  NAND2_X1 U14745 ( .A1(n12323), .A2(n12322), .ZN(n12326) );
  OR2_X1 U14746 ( .A1(n9431), .A2(n12324), .ZN(n12325) );
  OAI21_X1 U14747 ( .B1(n12494), .B2(n12327), .A(n13068), .ZN(n12328) );
  NOR2_X1 U14748 ( .A1(n13066), .A2(n12835), .ZN(n12529) );
  INV_X1 U14749 ( .A(n13066), .ZN(n12329) );
  NOR2_X1 U14750 ( .A1(n13068), .A2(n12494), .ZN(n12493) );
  NAND2_X1 U14751 ( .A1(n12329), .A2(n12493), .ZN(n12330) );
  NAND2_X1 U14752 ( .A1(n12331), .A2(n12330), .ZN(n12332) );
  INV_X1 U14753 ( .A(n12336), .ZN(n12540) );
  NAND2_X1 U14754 ( .A1(n12339), .A2(n12337), .ZN(n12338) );
  NAND2_X1 U14755 ( .A1(n12338), .A2(n12488), .ZN(n12341) );
  NAND3_X1 U14756 ( .A1(n12345), .A2(n12339), .A3(n12543), .ZN(n12340) );
  NAND2_X1 U14757 ( .A1(n12341), .A2(n12340), .ZN(n12344) );
  NAND2_X1 U14758 ( .A1(n15067), .A2(n12342), .ZN(n12343) );
  NAND3_X1 U14759 ( .A1(n12344), .A2(n12343), .A3(n12348), .ZN(n12349) );
  NAND3_X1 U14760 ( .A1(n12349), .A2(n15044), .A3(n12345), .ZN(n12347) );
  NAND3_X1 U14761 ( .A1(n12347), .A2(n12352), .A3(n12346), .ZN(n12357) );
  NAND3_X1 U14762 ( .A1(n12349), .A2(n15044), .A3(n12348), .ZN(n12355) );
  AND2_X1 U14763 ( .A1(n12351), .A2(n12350), .ZN(n12354) );
  INV_X1 U14764 ( .A(n12352), .ZN(n12353) );
  AOI21_X1 U14765 ( .B1(n12355), .B2(n12354), .A(n12353), .ZN(n12356) );
  MUX2_X1 U14766 ( .A(n12357), .B(n12356), .S(n12496), .Z(n12360) );
  NAND3_X1 U14767 ( .A1(n12701), .A2(n12358), .A3(n12488), .ZN(n12359) );
  NAND3_X1 U14768 ( .A1(n12360), .A2(n15025), .A3(n12359), .ZN(n12363) );
  OR2_X1 U14769 ( .A1(n12361), .A2(n12496), .ZN(n12362) );
  NAND3_X1 U14770 ( .A1(n12363), .A2(n15015), .A3(n12362), .ZN(n12367) );
  NAND2_X1 U14771 ( .A1(n12377), .A2(n12364), .ZN(n12365) );
  NAND2_X1 U14772 ( .A1(n12365), .A2(n12488), .ZN(n12366) );
  NAND2_X1 U14773 ( .A1(n12367), .A2(n12366), .ZN(n12372) );
  NAND3_X1 U14774 ( .A1(n12700), .A2(n12496), .A3(n15034), .ZN(n12368) );
  NAND2_X1 U14775 ( .A1(n12372), .A2(n12368), .ZN(n12370) );
  NAND3_X1 U14776 ( .A1(n12370), .A2(n12371), .A3(n12369), .ZN(n12375) );
  NAND2_X1 U14777 ( .A1(n12372), .A2(n12371), .ZN(n12373) );
  NAND2_X1 U14778 ( .A1(n12373), .A2(n12488), .ZN(n12374) );
  NAND3_X1 U14779 ( .A1(n12375), .A2(n12374), .A3(n12504), .ZN(n12380) );
  NAND3_X1 U14780 ( .A1(n12697), .A2(n12376), .A3(n12488), .ZN(n12379) );
  NOR2_X1 U14781 ( .A1(n12377), .A2(n12488), .ZN(n12378) );
  AOI21_X1 U14782 ( .B1(n12380), .B2(n12379), .A(n12378), .ZN(n12386) );
  OAI21_X1 U14783 ( .B1(n12381), .B2(n12488), .A(n12503), .ZN(n12385) );
  MUX2_X1 U14784 ( .A(n12383), .B(n12382), .S(n12488), .Z(n12384) );
  OAI211_X1 U14785 ( .C1(n12386), .C2(n12385), .A(n12511), .B(n12384), .ZN(
        n12391) );
  NAND2_X1 U14786 ( .A1(n12387), .A2(n15003), .ZN(n12389) );
  NAND2_X1 U14787 ( .A1(n12695), .A2(n6844), .ZN(n12388) );
  MUX2_X1 U14788 ( .A(n12389), .B(n12388), .S(n12488), .Z(n12390) );
  NAND3_X1 U14789 ( .A1(n12391), .A2(n7237), .A3(n12390), .ZN(n12393) );
  NAND3_X1 U14790 ( .A1(n12694), .A2(n12496), .A3(n15114), .ZN(n12392) );
  NAND2_X1 U14791 ( .A1(n12393), .A2(n12392), .ZN(n12394) );
  NAND2_X1 U14792 ( .A1(n12394), .A2(n14337), .ZN(n12401) );
  INV_X1 U14793 ( .A(n12395), .ZN(n12396) );
  NAND2_X1 U14794 ( .A1(n14337), .A2(n12396), .ZN(n12398) );
  NAND3_X1 U14795 ( .A1(n12398), .A2(n12406), .A3(n12397), .ZN(n12399) );
  NAND2_X1 U14796 ( .A1(n12399), .A2(n12488), .ZN(n12400) );
  NAND2_X1 U14797 ( .A1(n12401), .A2(n12400), .ZN(n12405) );
  AOI21_X1 U14798 ( .B1(n12404), .B2(n12402), .A(n12488), .ZN(n12403) );
  AOI21_X1 U14799 ( .B1(n12405), .B2(n12404), .A(n12403), .ZN(n12411) );
  OAI21_X1 U14800 ( .B1(n12406), .B2(n12488), .A(n12517), .ZN(n12410) );
  INV_X1 U14801 ( .A(n14325), .ZN(n12518) );
  MUX2_X1 U14802 ( .A(n12408), .B(n12407), .S(n12496), .Z(n12409) );
  OAI211_X1 U14803 ( .C1(n12411), .C2(n12410), .A(n12518), .B(n12409), .ZN(
        n12415) );
  MUX2_X1 U14804 ( .A(n12413), .B(n12412), .S(n12496), .Z(n12414) );
  NAND2_X1 U14805 ( .A1(n12415), .A2(n12414), .ZN(n12416) );
  NAND2_X1 U14806 ( .A1(n12416), .A2(n13003), .ZN(n12421) );
  NAND2_X1 U14807 ( .A1(n12424), .A2(n12417), .ZN(n12418) );
  NAND2_X1 U14808 ( .A1(n12418), .A2(n12488), .ZN(n12420) );
  INV_X1 U14809 ( .A(n12423), .ZN(n12419) );
  AOI21_X1 U14810 ( .B1(n12421), .B2(n12420), .A(n12419), .ZN(n12426) );
  AOI21_X1 U14811 ( .B1(n12423), .B2(n12422), .A(n12488), .ZN(n12425) );
  OAI22_X1 U14812 ( .A1(n12426), .A2(n12425), .B1(n12424), .B2(n12488), .ZN(
        n12432) );
  INV_X1 U14813 ( .A(n12433), .ZN(n12431) );
  AND2_X1 U14814 ( .A1(n12428), .A2(n12496), .ZN(n12429) );
  OAI211_X1 U14815 ( .C1(n12431), .C2(n12430), .A(n12438), .B(n12429), .ZN(
        n12435) );
  AOI22_X1 U14816 ( .A1(n12432), .A2(n12980), .B1(n6866), .B2(n12435), .ZN(
        n12437) );
  NAND3_X1 U14817 ( .A1(n12439), .A2(n12433), .A3(n12488), .ZN(n12434) );
  NAND2_X1 U14818 ( .A1(n12435), .A2(n12434), .ZN(n12436) );
  OAI21_X1 U14819 ( .B1(n12437), .B2(n12970), .A(n12436), .ZN(n12441) );
  INV_X1 U14820 ( .A(n12937), .ZN(n12941) );
  MUX2_X1 U14821 ( .A(n12439), .B(n12438), .S(n12488), .Z(n12440) );
  NAND3_X1 U14822 ( .A1(n12441), .A2(n12941), .A3(n12440), .ZN(n12445) );
  MUX2_X1 U14823 ( .A(n12443), .B(n12442), .S(n12496), .Z(n12444) );
  AOI21_X1 U14824 ( .B1(n12445), .B2(n12444), .A(n12933), .ZN(n12450) );
  MUX2_X1 U14825 ( .A(n12447), .B(n12446), .S(n12496), .Z(n12448) );
  INV_X1 U14826 ( .A(n12448), .ZN(n12449) );
  OAI21_X1 U14827 ( .B1(n12450), .B2(n12449), .A(n12912), .ZN(n12454) );
  MUX2_X1 U14828 ( .A(n12452), .B(n12451), .S(n12496), .Z(n12453) );
  NAND3_X1 U14829 ( .A1(n12454), .A2(n12897), .A3(n12453), .ZN(n12456) );
  NAND3_X1 U14830 ( .A1(n13024), .A2(n12915), .A3(n12496), .ZN(n12455) );
  NAND2_X1 U14831 ( .A1(n12456), .A2(n12455), .ZN(n12458) );
  NAND3_X1 U14832 ( .A1(n12458), .A2(n12457), .A3(n12873), .ZN(n12466) );
  OR2_X1 U14833 ( .A1(n12592), .A2(n12885), .ZN(n12460) );
  MUX2_X1 U14834 ( .A(n12460), .B(n12459), .S(n12496), .Z(n12465) );
  XNOR2_X1 U14835 ( .A(n12461), .B(n12496), .ZN(n12462) );
  OR3_X1 U14836 ( .A1(n12868), .A2(n12463), .A3(n12462), .ZN(n12464) );
  NAND4_X1 U14837 ( .A1(n12525), .A2(n12466), .A3(n12465), .A4(n12464), .ZN(
        n12476) );
  AND2_X1 U14838 ( .A1(n12476), .A2(n7384), .ZN(n12468) );
  INV_X1 U14839 ( .A(n12481), .ZN(n12471) );
  NAND3_X1 U14840 ( .A1(n12476), .A2(n12526), .A3(n12475), .ZN(n12478) );
  NAND2_X1 U14841 ( .A1(n12478), .A2(n12477), .ZN(n12480) );
  NAND2_X1 U14842 ( .A1(n12480), .A2(n12479), .ZN(n12482) );
  NAND2_X1 U14843 ( .A1(n12482), .A2(n12481), .ZN(n12483) );
  MUX2_X1 U14844 ( .A(n12484), .B(n12483), .S(n12488), .Z(n12486) );
  XNOR2_X1 U14845 ( .A(n13068), .B(n12494), .ZN(n12530) );
  INV_X1 U14846 ( .A(n12487), .ZN(n12489) );
  NOR2_X1 U14847 ( .A1(n12489), .A2(n12488), .ZN(n12490) );
  INV_X1 U14848 ( .A(n12493), .ZN(n12497) );
  INV_X1 U14849 ( .A(n12912), .ZN(n12916) );
  NAND4_X1 U14850 ( .A1(n12504), .A2(n15044), .A3(n15015), .A4(n12503), .ZN(
        n12506) );
  NOR2_X1 U14851 ( .A1(n12506), .A2(n12505), .ZN(n12513) );
  NOR2_X1 U14852 ( .A1(n12507), .A2(n15068), .ZN(n12510) );
  AND4_X1 U14853 ( .A1(n12510), .A2(n15025), .A3(n12509), .A4(n12508), .ZN(
        n12512) );
  NAND4_X1 U14854 ( .A1(n12513), .A2(n12512), .A3(n14337), .A4(n12511), .ZN(
        n12515) );
  NOR2_X1 U14855 ( .A1(n12515), .A2(n12514), .ZN(n12516) );
  NAND4_X1 U14856 ( .A1(n13003), .A2(n12518), .A3(n12517), .A4(n12516), .ZN(
        n12519) );
  NOR2_X1 U14857 ( .A1(n12986), .A2(n12519), .ZN(n12520) );
  NAND3_X1 U14858 ( .A1(n12964), .A2(n12980), .A3(n12520), .ZN(n12521) );
  OR3_X1 U14859 ( .A1(n12937), .A2(n12951), .A3(n12521), .ZN(n12522) );
  OR4_X1 U14860 ( .A1(n12901), .A2(n12933), .A3(n12916), .A4(n12522), .ZN(
        n12523) );
  NOR2_X1 U14861 ( .A1(n12887), .A2(n12523), .ZN(n12524) );
  INV_X1 U14862 ( .A(n12530), .ZN(n12531) );
  XNOR2_X1 U14863 ( .A(n12532), .B(n12818), .ZN(n12533) );
  OAI22_X1 U14864 ( .A1(n12536), .A2(n12542), .B1(n12534), .B2(n12533), .ZN(
        n12535) );
  NAND2_X1 U14865 ( .A1(n12538), .A2(n12537), .ZN(n12539) );
  NOR4_X1 U14866 ( .A1(n14341), .A2(n12542), .A3(n13139), .A4(n12541), .ZN(
        n12545) );
  OAI21_X1 U14867 ( .B1(n12546), .B2(n12543), .A(P3_B_REG_SCAN_IN), .ZN(n12544) );
  OAI22_X1 U14868 ( .A1(n12547), .A2(n12546), .B1(n12545), .B2(n12544), .ZN(
        P3_U3296) );
  NOR2_X1 U14869 ( .A1(n15009), .A2(n12548), .ZN(n12836) );
  NOR2_X1 U14870 ( .A1(n12549), .A2(n13007), .ZN(n12550) );
  AOI211_X1 U14871 ( .C1(n15082), .C2(P3_REG2_REG_29__SCAN_IN), .A(n12836), 
        .B(n12550), .ZN(n12553) );
  OR2_X1 U14872 ( .A1(n12551), .A2(n12960), .ZN(n12552) );
  OAI211_X1 U14873 ( .C1(n12554), .C2(n15082), .A(n12553), .B(n12552), .ZN(
        P3_U3204) );
  AOI22_X1 U14874 ( .A1(n12870), .A2(n12663), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12559) );
  OAI21_X1 U14875 ( .B1(n12560), .B2(n12665), .A(n12559), .ZN(n12562) );
  NOR2_X1 U14876 ( .A1(n13080), .A2(n12681), .ZN(n12561) );
  AOI211_X1 U14877 ( .C1(n12849), .C2(n12678), .A(n12562), .B(n12561), .ZN(
        n12563) );
  NAND2_X1 U14878 ( .A1(n12564), .A2(n12563), .ZN(P3_U3154) );
  INV_X1 U14879 ( .A(n12566), .ZN(n12567) );
  NAND2_X1 U14880 ( .A1(n12565), .A2(n12567), .ZN(n12624) );
  OAI21_X1 U14881 ( .B1(n12565), .B2(n12567), .A(n12624), .ZN(n12568) );
  NOR2_X1 U14882 ( .A1(n12568), .A2(n12685), .ZN(n12627) );
  AOI21_X1 U14883 ( .B1(n12685), .B2(n12568), .A(n12627), .ZN(n12573) );
  NAND2_X1 U14884 ( .A1(n12678), .A2(n12905), .ZN(n12570) );
  AOI22_X1 U14885 ( .A1(n12663), .A2(n12927), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12569) );
  OAI211_X1 U14886 ( .C1(n12601), .C2(n12665), .A(n12570), .B(n12569), .ZN(
        n12571) );
  AOI21_X1 U14887 ( .B1(n13024), .B2(n12648), .A(n12571), .ZN(n12572) );
  OAI21_X1 U14888 ( .B1(n12573), .B2(n12650), .A(n12572), .ZN(P3_U3156) );
  XNOR2_X1 U14889 ( .A(n12574), .B(n12966), .ZN(n12575) );
  XNOR2_X1 U14890 ( .A(n12576), .B(n12575), .ZN(n12581) );
  NAND2_X1 U14891 ( .A1(n12952), .A2(n12663), .ZN(n12577) );
  NAND2_X1 U14892 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12817)
         );
  OAI211_X1 U14893 ( .C1(n12955), .C2(n12665), .A(n12577), .B(n12817), .ZN(
        n12579) );
  NOR2_X1 U14894 ( .A1(n13105), .A2(n12681), .ZN(n12578) );
  AOI211_X1 U14895 ( .C1(n12956), .C2(n12678), .A(n12579), .B(n12578), .ZN(
        n12580) );
  OAI21_X1 U14896 ( .B1(n12581), .B2(n12650), .A(n12580), .ZN(P3_U3159) );
  INV_X1 U14897 ( .A(n12582), .ZN(n12583) );
  AOI21_X1 U14898 ( .B1(n12585), .B2(n12584), .A(n12583), .ZN(n12591) );
  AOI22_X1 U14899 ( .A1(n12926), .A2(n12663), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12587) );
  NAND2_X1 U14900 ( .A1(n12678), .A2(n12929), .ZN(n12586) );
  OAI211_X1 U14901 ( .C1(n12588), .C2(n12665), .A(n12587), .B(n12586), .ZN(
        n12589) );
  AOI21_X1 U14902 ( .B1(n13033), .B2(n12648), .A(n12589), .ZN(n12590) );
  OAI21_X1 U14903 ( .B1(n12591), .B2(n12650), .A(n12590), .ZN(P3_U3163) );
  INV_X1 U14904 ( .A(n12593), .ZN(n12628) );
  INV_X1 U14905 ( .A(n12594), .ZN(n12596) );
  NOR3_X1 U14906 ( .A1(n12628), .A2(n12596), .A3(n12595), .ZN(n12599) );
  INV_X1 U14907 ( .A(n12597), .ZN(n12598) );
  OAI21_X1 U14908 ( .B1(n12599), .B2(n12598), .A(n12670), .ZN(n12604) );
  AOI22_X1 U14909 ( .A1(n12870), .A2(n12674), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12600) );
  OAI21_X1 U14910 ( .B1(n12601), .B2(n12676), .A(n12600), .ZN(n12602) );
  AOI21_X1 U14911 ( .B1(n12875), .B2(n12678), .A(n12602), .ZN(n12603) );
  OAI211_X1 U14912 ( .C1(n13084), .C2(n12681), .A(n12604), .B(n12603), .ZN(
        P3_U3165) );
  INV_X1 U14913 ( .A(n12614), .ZN(n12605) );
  AOI21_X1 U14914 ( .B1(n12607), .B2(n12606), .A(n12605), .ZN(n12612) );
  AOI22_X1 U14915 ( .A1(n12688), .A2(n12674), .B1(P3_REG3_REG_16__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12609) );
  NAND2_X1 U14916 ( .A1(n12678), .A2(n12993), .ZN(n12608) );
  OAI211_X1 U14917 ( .C1(n14329), .C2(n12676), .A(n12609), .B(n12608), .ZN(
        n12610) );
  AOI21_X1 U14918 ( .B1(n12992), .B2(n12648), .A(n12610), .ZN(n12611) );
  OAI21_X1 U14919 ( .B1(n12612), .B2(n12650), .A(n12611), .ZN(P3_U3166) );
  NAND2_X1 U14920 ( .A1(n12614), .A2(n12613), .ZN(n12616) );
  AOI21_X1 U14921 ( .B1(n12616), .B2(n12615), .A(n12650), .ZN(n12618) );
  NAND2_X1 U14922 ( .A1(n12618), .A2(n12617), .ZN(n12622) );
  NAND2_X1 U14923 ( .A1(n12689), .A2(n12663), .ZN(n12619) );
  NAND2_X1 U14924 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n14313)
         );
  OAI211_X1 U14925 ( .C1(n12978), .C2(n12665), .A(n12619), .B(n14313), .ZN(
        n12620) );
  AOI21_X1 U14926 ( .B1(n12981), .B2(n12678), .A(n12620), .ZN(n12621) );
  OAI211_X1 U14927 ( .C1(n13113), .C2(n12681), .A(n12622), .B(n12621), .ZN(
        P3_U3168) );
  INV_X1 U14928 ( .A(n13020), .ZN(n12894) );
  INV_X1 U14929 ( .A(n12623), .ZN(n12626) );
  INV_X1 U14930 ( .A(n12624), .ZN(n12625) );
  NOR3_X1 U14931 ( .A1(n12627), .A2(n12626), .A3(n12625), .ZN(n12629) );
  OAI21_X1 U14932 ( .B1(n12629), .B2(n12628), .A(n12670), .ZN(n12634) );
  NOR2_X1 U14933 ( .A1(n12676), .A2(n12915), .ZN(n12632) );
  OAI22_X1 U14934 ( .A1(n12885), .A2(n12665), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12630), .ZN(n12631) );
  AOI211_X1 U14935 ( .C1(n12892), .C2(n12678), .A(n12632), .B(n12631), .ZN(
        n12633) );
  OAI211_X1 U14936 ( .C1(n12894), .C2(n12681), .A(n12634), .B(n12633), .ZN(
        P3_U3169) );
  XNOR2_X1 U14937 ( .A(n12636), .B(n12635), .ZN(n12641) );
  AOI22_X1 U14938 ( .A1(n12686), .A2(n12674), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12638) );
  NAND2_X1 U14939 ( .A1(n12678), .A2(n12944), .ZN(n12637) );
  OAI211_X1 U14940 ( .C1(n12966), .C2(n12676), .A(n12638), .B(n12637), .ZN(
        n12639) );
  AOI21_X1 U14941 ( .B1(n12943), .B2(n12648), .A(n12639), .ZN(n12640) );
  OAI21_X1 U14942 ( .B1(n12641), .B2(n12650), .A(n12640), .ZN(P3_U3173) );
  INV_X1 U14943 ( .A(n12642), .ZN(n12643) );
  AOI21_X1 U14944 ( .B1(n12927), .B2(n12644), .A(n12643), .ZN(n12651) );
  AOI22_X1 U14945 ( .A1(n12686), .A2(n12663), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12646) );
  NAND2_X1 U14946 ( .A1(n12678), .A2(n12919), .ZN(n12645) );
  OAI211_X1 U14947 ( .C1(n12915), .C2(n12665), .A(n12646), .B(n12645), .ZN(
        n12647) );
  AOI21_X1 U14948 ( .B1(n12918), .B2(n12648), .A(n12647), .ZN(n12649) );
  OAI21_X1 U14949 ( .B1(n12651), .B2(n12650), .A(n12649), .ZN(P3_U3175) );
  OAI211_X1 U14950 ( .C1(n12654), .C2(n12653), .A(n12652), .B(n12670), .ZN(
        n12658) );
  NAND2_X1 U14951 ( .A1(n12688), .A2(n12663), .ZN(n12655) );
  NAND2_X1 U14952 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12792)
         );
  OAI211_X1 U14953 ( .C1(n12966), .C2(n12665), .A(n12655), .B(n12792), .ZN(
        n12656) );
  AOI21_X1 U14954 ( .B1(n12971), .B2(n12678), .A(n12656), .ZN(n12657) );
  OAI211_X1 U14955 ( .C1(n13109), .C2(n12681), .A(n12658), .B(n12657), .ZN(
        P3_U3178) );
  OAI21_X1 U14956 ( .B1(n12661), .B2(n12660), .A(n12659), .ZN(n12662) );
  NAND2_X1 U14957 ( .A1(n12662), .A2(n12670), .ZN(n12669) );
  AOI22_X1 U14958 ( .A1(n12684), .A2(n12663), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12664) );
  OAI21_X1 U14959 ( .B1(n12666), .B2(n12665), .A(n12664), .ZN(n12667) );
  AOI21_X1 U14960 ( .B1(n12860), .B2(n12678), .A(n12667), .ZN(n12668) );
  OAI211_X1 U14961 ( .C1(n12862), .C2(n12681), .A(n12669), .B(n12668), .ZN(
        P3_U3180) );
  OAI211_X1 U14962 ( .C1(n12673), .C2(n12672), .A(n12671), .B(n12670), .ZN(
        n12680) );
  NOR2_X1 U14963 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n7750), .ZN(n12765) );
  AOI21_X1 U14964 ( .B1(n12689), .B2(n12674), .A(n12765), .ZN(n12675) );
  OAI21_X1 U14965 ( .B1(n13000), .B2(n12676), .A(n12675), .ZN(n12677) );
  AOI21_X1 U14966 ( .B1(n13005), .B2(n12678), .A(n12677), .ZN(n12679) );
  OAI211_X1 U14967 ( .C1(n13122), .C2(n12681), .A(n12680), .B(n12679), .ZN(
        P3_U3181) );
  MUX2_X1 U14968 ( .A(n12835), .B(P3_DATAO_REG_31__SCAN_IN), .S(n12702), .Z(
        P3_U3522) );
  MUX2_X1 U14969 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12682), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14970 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12683), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14971 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n12870), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U14972 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12684), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14973 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n6647), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U14974 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n12685), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U14975 ( .A(n12927), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12702), .Z(
        P3_U3513) );
  MUX2_X1 U14976 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12686), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14977 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12926), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14978 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n12687), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U14979 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12952), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14980 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12688), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14981 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12689), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14982 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n7255), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U14983 ( .A(n12690), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12702), .Z(
        P3_U3505) );
  MUX2_X1 U14984 ( .A(n12691), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12702), .Z(
        P3_U3504) );
  MUX2_X1 U14985 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12692), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14986 ( .A(n12693), .B(P3_DATAO_REG_11__SCAN_IN), .S(n12702), .Z(
        P3_U3502) );
  MUX2_X1 U14987 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12694), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14988 ( .A(n12695), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12702), .Z(
        P3_U3500) );
  MUX2_X1 U14989 ( .A(n12696), .B(P3_DATAO_REG_8__SCAN_IN), .S(n12702), .Z(
        P3_U3499) );
  MUX2_X1 U14990 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12697), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14991 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12698), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14992 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12699), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14993 ( .A(n12700), .B(P3_DATAO_REG_4__SCAN_IN), .S(n12702), .Z(
        P3_U3495) );
  MUX2_X1 U14994 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12701), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14995 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n15064), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14996 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n10406), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U14997 ( .A(n10404), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12702), .Z(
        P3_U3491) );
  AOI21_X1 U14998 ( .B1(n7722), .B2(n12704), .A(n6521), .ZN(n12721) );
  INV_X1 U14999 ( .A(n12727), .ZN(n12736) );
  XNOR2_X1 U15000 ( .A(n12736), .B(n12726), .ZN(n12707) );
  NAND2_X1 U15001 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n12707), .ZN(n12728) );
  OAI21_X1 U15002 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n12707), .A(n12728), 
        .ZN(n12719) );
  NAND2_X1 U15003 ( .A1(n12709), .A2(n12708), .ZN(n12711) );
  MUX2_X1 U15004 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n6473), .Z(n12735) );
  XNOR2_X1 U15005 ( .A(n12735), .B(n12736), .ZN(n12710) );
  NAND3_X1 U15006 ( .A1(n12712), .A2(n12711), .A3(n12710), .ZN(n12743) );
  INV_X1 U15007 ( .A(n12743), .ZN(n12714) );
  AOI21_X1 U15008 ( .B1(n12712), .B2(n12711), .A(n12710), .ZN(n12713) );
  OAI21_X1 U15009 ( .B1(n12714), .B2(n12713), .A(n14962), .ZN(n12717) );
  AOI21_X1 U15010 ( .B1(n14969), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n12715), 
        .ZN(n12716) );
  OAI211_X1 U15011 ( .C1(n14966), .C2(n12727), .A(n12717), .B(n12716), .ZN(
        n12718) );
  AOI21_X1 U15012 ( .B1(n6467), .B2(n12719), .A(n12718), .ZN(n12720) );
  OAI21_X1 U15013 ( .B1(n12721), .B2(n14991), .A(n12720), .ZN(P3_U3195) );
  NOR2_X1 U15014 ( .A1(n12736), .A2(n12722), .ZN(n12723) );
  NAND2_X1 U15015 ( .A1(n12734), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12758) );
  OR2_X1 U15016 ( .A1(n12734), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12724) );
  NAND2_X1 U15017 ( .A1(n12758), .A2(n12724), .ZN(n12738) );
  AOI21_X1 U15018 ( .B1(n12725), .B2(n12738), .A(n12751), .ZN(n12750) );
  NAND2_X1 U15019 ( .A1(n12727), .A2(n12726), .ZN(n12729) );
  NAND2_X1 U15020 ( .A1(n12729), .A2(n12728), .ZN(n12731) );
  NAND2_X1 U15021 ( .A1(n12734), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12757) );
  OR2_X1 U15022 ( .A1(n12734), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12730) );
  AND2_X1 U15023 ( .A1(n12757), .A2(n12730), .ZN(n12739) );
  NAND2_X1 U15024 ( .A1(n12739), .A2(n12731), .ZN(n12755) );
  OAI21_X1 U15025 ( .B1(n12731), .B2(n12739), .A(n12755), .ZN(n12748) );
  AOI21_X1 U15026 ( .B1(n14969), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n12732), 
        .ZN(n12733) );
  OAI21_X1 U15027 ( .B1(n14966), .B2(n12734), .A(n12733), .ZN(n12747) );
  INV_X1 U15028 ( .A(n12735), .ZN(n12737) );
  NAND2_X1 U15029 ( .A1(n12737), .A2(n12736), .ZN(n12742) );
  INV_X1 U15030 ( .A(n12738), .ZN(n12740) );
  MUX2_X1 U15031 ( .A(n12740), .B(n12739), .S(n12776), .Z(n12741) );
  NAND3_X1 U15032 ( .A1(n12743), .A2(n12742), .A3(n12741), .ZN(n12760) );
  INV_X1 U15033 ( .A(n12760), .ZN(n12745) );
  AOI21_X1 U15034 ( .B1(n12743), .B2(n12742), .A(n12741), .ZN(n12744) );
  NOR3_X1 U15035 ( .A1(n12745), .A2(n12744), .A3(n14985), .ZN(n12746) );
  AOI211_X1 U15036 ( .C1(n6467), .C2(n12748), .A(n12747), .B(n12746), .ZN(
        n12749) );
  OAI21_X1 U15037 ( .B1(n12750), .B2(n14991), .A(n12749), .ZN(P3_U3196) );
  INV_X1 U15038 ( .A(n12751), .ZN(n12752) );
  AOI21_X1 U15039 ( .B1(n12754), .B2(n12753), .A(n12783), .ZN(n12771) );
  NAND2_X1 U15040 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n12756), .ZN(n12796) );
  OAI21_X1 U15041 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n12756), .A(n12796), 
        .ZN(n12769) );
  MUX2_X1 U15042 ( .A(n12758), .B(n12757), .S(n6473), .Z(n12759) );
  NAND2_X1 U15043 ( .A1(n12760), .A2(n12759), .ZN(n12772) );
  XNOR2_X1 U15044 ( .A(n12772), .B(n12795), .ZN(n12762) );
  MUX2_X1 U15045 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12776), .Z(n12761) );
  AOI21_X1 U15046 ( .B1(n12762), .B2(n12761), .A(n12773), .ZN(n12767) );
  NOR2_X1 U15047 ( .A1(n15000), .A2(n12763), .ZN(n12764) );
  AOI211_X1 U15048 ( .C1(n14996), .C2(n12774), .A(n12765), .B(n12764), .ZN(
        n12766) );
  OAI21_X1 U15049 ( .B1(n12767), .B2(n14985), .A(n12766), .ZN(n12768) );
  AOI21_X1 U15050 ( .B1(n6467), .B2(n12769), .A(n12768), .ZN(n12770) );
  OAI21_X1 U15051 ( .B1(n12771), .B2(n14991), .A(n12770), .ZN(P3_U3197) );
  MUX2_X1 U15052 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12776), .Z(n12780) );
  MUX2_X1 U15053 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12776), .Z(n12778) );
  INV_X1 U15054 ( .A(n12772), .ZN(n12775) );
  AOI21_X1 U15055 ( .B1(n12775), .B2(n12774), .A(n12773), .ZN(n14294) );
  INV_X1 U15056 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13057) );
  MUX2_X1 U15057 ( .A(n12784), .B(n13057), .S(n6473), .Z(n12777) );
  NOR2_X1 U15058 ( .A1(n12777), .A2(n14289), .ZN(n14290) );
  NAND2_X1 U15059 ( .A1(n12777), .A2(n14289), .ZN(n14291) );
  OAI21_X1 U15060 ( .B1(n14294), .B2(n14290), .A(n14291), .ZN(n14317) );
  XNOR2_X1 U15061 ( .A(n12778), .B(n12798), .ZN(n14318) );
  NOR2_X1 U15062 ( .A1(n14317), .A2(n14318), .ZN(n14316) );
  XNOR2_X1 U15063 ( .A(n12825), .B(n12824), .ZN(n12779) );
  NOR2_X1 U15064 ( .A1(n12779), .A2(n12780), .ZN(n12823) );
  AOI21_X1 U15065 ( .B1(n12780), .B2(n12779), .A(n12823), .ZN(n12809) );
  AND2_X1 U15066 ( .A1(n12795), .A2(n12781), .ZN(n12782) );
  AOI22_X1 U15067 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n14289), .B1(n12793), 
        .B2(n12784), .ZN(n14301) );
  XOR2_X1 U15068 ( .A(n12798), .B(n12785), .Z(n14308) );
  INV_X1 U15069 ( .A(n14307), .ZN(n12790) );
  OR2_X1 U15070 ( .A1(n12785), .A2(n14312), .ZN(n12789) );
  OR2_X1 U15071 ( .A1(n12824), .A2(n12786), .ZN(n12810) );
  NAND2_X1 U15072 ( .A1(n12824), .A2(n12786), .ZN(n12787) );
  NAND2_X1 U15073 ( .A1(n12810), .A2(n12787), .ZN(n12788) );
  AND3_X1 U15074 ( .A1(n12790), .A2(n12789), .A3(n12788), .ZN(n12791) );
  OAI21_X1 U15075 ( .B1(n12811), .B2(n12791), .A(n14300), .ZN(n12808) );
  OAI21_X1 U15076 ( .B1(n15000), .B2(n9779), .A(n12792), .ZN(n12806) );
  AOI22_X1 U15077 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12793), .B1(n14289), 
        .B2(n13057), .ZN(n14297) );
  NAND2_X1 U15078 ( .A1(n12795), .A2(n12794), .ZN(n12797) );
  NAND2_X1 U15079 ( .A1(n12797), .A2(n12796), .ZN(n14296) );
  NAND2_X1 U15080 ( .A1(n14297), .A2(n14296), .ZN(n14295) );
  NAND2_X1 U15081 ( .A1(n12799), .A2(n12798), .ZN(n12801) );
  XNOR2_X1 U15082 ( .A(n12799), .B(n14312), .ZN(n14311) );
  NAND2_X1 U15083 ( .A1(P3_REG1_REG_17__SCAN_IN), .A2(n14311), .ZN(n14310) );
  INV_X1 U15084 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13049) );
  XNOR2_X1 U15085 ( .A(n12824), .B(n13049), .ZN(n12800) );
  INV_X1 U15086 ( .A(n12813), .ZN(n12804) );
  NAND3_X1 U15087 ( .A1(n12801), .A2(n14310), .A3(n12800), .ZN(n12803) );
  INV_X1 U15088 ( .A(n6467), .ZN(n12802) );
  AOI21_X1 U15089 ( .B1(n12804), .B2(n12803), .A(n12802), .ZN(n12805) );
  AOI211_X1 U15090 ( .C1(n14996), .C2(n12824), .A(n12806), .B(n12805), .ZN(
        n12807) );
  OAI211_X1 U15091 ( .C1(n12809), .C2(n14985), .A(n12808), .B(n12807), .ZN(
        P3_U3200) );
  XNOR2_X1 U15092 ( .A(n12818), .B(n12812), .ZN(n12819) );
  AOI21_X1 U15093 ( .B1(P3_REG1_REG_18__SCAN_IN), .B2(n12814), .A(n12813), 
        .ZN(n12815) );
  XNOR2_X1 U15094 ( .A(n12818), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12822) );
  XNOR2_X1 U15095 ( .A(n12815), .B(n12822), .ZN(n12831) );
  NAND2_X1 U15096 ( .A1(n14969), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12816) );
  OAI211_X1 U15097 ( .C1(n14966), .C2(n12818), .A(n12817), .B(n12816), .ZN(
        n12830) );
  INV_X1 U15098 ( .A(n12819), .ZN(n12821) );
  MUX2_X1 U15099 ( .A(n12822), .B(n12821), .S(n12820), .Z(n12827) );
  AOI21_X1 U15100 ( .B1(n12825), .B2(n12824), .A(n12823), .ZN(n12826) );
  XOR2_X1 U15101 ( .A(n12827), .B(n12826), .Z(n12828) );
  NOR2_X1 U15102 ( .A1(n12828), .A2(n14985), .ZN(n12829) );
  NAND2_X1 U15103 ( .A1(n15082), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12837) );
  INV_X1 U15104 ( .A(n12833), .ZN(n12834) );
  AND2_X1 U15105 ( .A1(n12835), .A2(n12834), .ZN(n13064) );
  OAI21_X1 U15106 ( .B1(n13064), .B2(n12836), .A(n15080), .ZN(n12838) );
  OAI211_X1 U15107 ( .C1(n13066), .C2(n13007), .A(n12837), .B(n12838), .ZN(
        P3_U3202) );
  INV_X1 U15108 ( .A(n13068), .ZN(n12840) );
  NAND2_X1 U15109 ( .A1(n15082), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n12839) );
  OAI211_X1 U15110 ( .C1(n12840), .C2(n13007), .A(n12839), .B(n12838), .ZN(
        P3_U3203) );
  INV_X1 U15111 ( .A(n12841), .ZN(n12842) );
  OAI22_X1 U15112 ( .A1(n15080), .A2(n12843), .B1(n12842), .B2(n15009), .ZN(
        n12846) );
  NOR2_X1 U15113 ( .A1(n12844), .A2(n12960), .ZN(n12845) );
  AOI211_X1 U15114 ( .C1(n15004), .C2(n7997), .A(n12846), .B(n12845), .ZN(
        n12847) );
  OAI21_X1 U15115 ( .B1(n12848), .B2(n15082), .A(n12847), .ZN(P3_U3205) );
  INV_X1 U15116 ( .A(n12849), .ZN(n12850) );
  OAI22_X1 U15117 ( .A1(n15080), .A2(n12851), .B1(n12850), .B2(n15009), .ZN(
        n12855) );
  NOR2_X1 U15118 ( .A1(n12853), .A2(n12852), .ZN(n12854) );
  AOI211_X1 U15119 ( .C1(n15004), .C2(n12856), .A(n12855), .B(n12854), .ZN(
        n12857) );
  OAI21_X1 U15120 ( .B1(n12858), .B2(n15082), .A(n12857), .ZN(P3_U3206) );
  INV_X1 U15121 ( .A(n12859), .ZN(n12866) );
  AOI22_X1 U15122 ( .A1(n15082), .A2(P3_REG2_REG_26__SCAN_IN), .B1(n12860), 
        .B2(n15077), .ZN(n12861) );
  OAI21_X1 U15123 ( .B1(n12862), .B2(n13007), .A(n12861), .ZN(n12863) );
  AOI21_X1 U15124 ( .B1(n12864), .B2(n15078), .A(n12863), .ZN(n12865) );
  OAI21_X1 U15125 ( .B1(n12866), .B2(n15082), .A(n12865), .ZN(P3_U3207) );
  OAI211_X1 U15126 ( .C1(n12869), .C2(n12868), .A(n12867), .B(n15060), .ZN(
        n12872) );
  AOI22_X1 U15127 ( .A1(n15062), .A2(n6647), .B1(n12870), .B2(n15063), .ZN(
        n12871) );
  NAND2_X1 U15128 ( .A1(n12872), .A2(n12871), .ZN(n13016) );
  INV_X1 U15129 ( .A(n13016), .ZN(n12879) );
  XNOR2_X1 U15130 ( .A(n12874), .B(n12873), .ZN(n13017) );
  AOI22_X1 U15131 ( .A1(n15082), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n15077), 
        .B2(n12875), .ZN(n12876) );
  OAI21_X1 U15132 ( .B1(n13084), .B2(n13007), .A(n12876), .ZN(n12877) );
  AOI21_X1 U15133 ( .B1(n13017), .B2(n14346), .A(n12877), .ZN(n12878) );
  OAI21_X1 U15134 ( .B1(n12879), .B2(n15082), .A(n12878), .ZN(P3_U3208) );
  NAND2_X1 U15135 ( .A1(n12880), .A2(n12881), .ZN(n12882) );
  NAND2_X1 U15136 ( .A1(n12882), .A2(n12887), .ZN(n12884) );
  NAND2_X1 U15137 ( .A1(n12884), .A2(n12883), .ZN(n13021) );
  OAI22_X1 U15138 ( .A1(n12885), .A2(n14339), .B1(n12915), .B2(n14341), .ZN(
        n12891) );
  OAI211_X1 U15139 ( .C1(n12888), .C2(n12887), .A(n12886), .B(n15060), .ZN(
        n12889) );
  INV_X1 U15140 ( .A(n12889), .ZN(n12890) );
  AOI211_X1 U15141 ( .C1(n15070), .C2(n13021), .A(n12891), .B(n12890), .ZN(
        n13023) );
  AOI22_X1 U15142 ( .A1(n15082), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n15077), 
        .B2(n12892), .ZN(n12893) );
  OAI21_X1 U15143 ( .B1(n12894), .B2(n13007), .A(n12893), .ZN(n12895) );
  AOI21_X1 U15144 ( .B1(n13021), .B2(n15078), .A(n12895), .ZN(n12896) );
  OAI21_X1 U15145 ( .B1(n13023), .B2(n15082), .A(n12896), .ZN(P3_U3209) );
  OR2_X1 U15146 ( .A1(n12898), .A2(n12897), .ZN(n12899) );
  AND2_X1 U15147 ( .A1(n12880), .A2(n12899), .ZN(n13026) );
  INV_X1 U15148 ( .A(n13026), .ZN(n12911) );
  OAI211_X1 U15149 ( .C1(n12902), .C2(n12901), .A(n12900), .B(n15060), .ZN(
        n12904) );
  AOI22_X1 U15150 ( .A1(n6647), .A2(n15063), .B1(n15062), .B2(n12927), .ZN(
        n12903) );
  NAND2_X1 U15151 ( .A1(n12904), .A2(n12903), .ZN(n13025) );
  NAND2_X1 U15152 ( .A1(n13025), .A2(n15080), .ZN(n12910) );
  INV_X1 U15153 ( .A(n12905), .ZN(n12906) );
  OAI22_X1 U15154 ( .A1(n15080), .A2(n12907), .B1(n12906), .B2(n15009), .ZN(
        n12908) );
  AOI21_X1 U15155 ( .B1(n13024), .B2(n15004), .A(n12908), .ZN(n12909) );
  OAI211_X1 U15156 ( .C1(n12911), .C2(n12960), .A(n12910), .B(n12909), .ZN(
        P3_U3210) );
  XNOR2_X1 U15157 ( .A(n12913), .B(n12912), .ZN(n12914) );
  OAI222_X1 U15158 ( .A1(n14341), .A2(n12940), .B1(n14339), .B2(n12915), .C1(
        n15045), .C2(n12914), .ZN(n13029) );
  INV_X1 U15159 ( .A(n13029), .ZN(n12923) );
  XNOR2_X1 U15160 ( .A(n12917), .B(n12916), .ZN(n13030) );
  INV_X1 U15161 ( .A(n12918), .ZN(n13093) );
  AOI22_X1 U15162 ( .A1(n15082), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n15077), 
        .B2(n12919), .ZN(n12920) );
  OAI21_X1 U15163 ( .B1(n13093), .B2(n13007), .A(n12920), .ZN(n12921) );
  AOI21_X1 U15164 ( .B1(n13030), .B2(n14346), .A(n12921), .ZN(n12922) );
  OAI21_X1 U15165 ( .B1(n12923), .B2(n15082), .A(n12922), .ZN(P3_U3211) );
  OAI21_X1 U15166 ( .B1(n12925), .B2(n12933), .A(n12924), .ZN(n12928) );
  AOI222_X1 U15167 ( .A1(n15060), .A2(n12928), .B1(n12927), .B2(n15063), .C1(
        n12926), .C2(n15062), .ZN(n13034) );
  INV_X1 U15168 ( .A(n12929), .ZN(n12930) );
  OAI22_X1 U15169 ( .A1(n15080), .A2(n12931), .B1(n12930), .B2(n15009), .ZN(
        n12932) );
  AOI21_X1 U15170 ( .B1(n13033), .B2(n15004), .A(n12932), .ZN(n12936) );
  XNOR2_X1 U15171 ( .A(n12934), .B(n12933), .ZN(n13036) );
  NAND2_X1 U15172 ( .A1(n13036), .A2(n14346), .ZN(n12935) );
  OAI211_X1 U15173 ( .C1(n13034), .C2(n15082), .A(n12936), .B(n12935), .ZN(
        P3_U3212) );
  XNOR2_X1 U15174 ( .A(n12938), .B(n12937), .ZN(n12939) );
  OAI222_X1 U15175 ( .A1(n14339), .A2(n12940), .B1(n14341), .B2(n12966), .C1(
        n12939), .C2(n15045), .ZN(n13039) );
  INV_X1 U15176 ( .A(n13039), .ZN(n12948) );
  XNOR2_X1 U15177 ( .A(n12942), .B(n12941), .ZN(n13040) );
  INV_X1 U15178 ( .A(n12943), .ZN(n13101) );
  AOI22_X1 U15179 ( .A1(n15082), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n15077), 
        .B2(n12944), .ZN(n12945) );
  OAI21_X1 U15180 ( .B1(n13101), .B2(n13007), .A(n12945), .ZN(n12946) );
  AOI21_X1 U15181 ( .B1(n13040), .B2(n14346), .A(n12946), .ZN(n12947) );
  OAI21_X1 U15182 ( .B1(n12948), .B2(n15082), .A(n12947), .ZN(P3_U3213) );
  XNOR2_X1 U15183 ( .A(n12949), .B(n12951), .ZN(n13044) );
  INV_X1 U15184 ( .A(n13044), .ZN(n12961) );
  OAI211_X1 U15185 ( .C1(n6561), .C2(n12951), .A(n12950), .B(n15060), .ZN(
        n12954) );
  NAND2_X1 U15186 ( .A1(n12952), .A2(n15062), .ZN(n12953) );
  OAI211_X1 U15187 ( .C1(n12955), .C2(n14339), .A(n12954), .B(n12953), .ZN(
        n13043) );
  AOI22_X1 U15188 ( .A1(n15082), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15077), 
        .B2(n12956), .ZN(n12957) );
  OAI21_X1 U15189 ( .B1(n13105), .B2(n13007), .A(n12957), .ZN(n12958) );
  AOI21_X1 U15190 ( .B1(n13043), .B2(n15080), .A(n12958), .ZN(n12959) );
  OAI21_X1 U15191 ( .B1(n12961), .B2(n12960), .A(n12959), .ZN(P3_U3214) );
  AOI21_X1 U15192 ( .B1(n12964), .B2(n12963), .A(n12962), .ZN(n12965) );
  OAI222_X1 U15193 ( .A1(n14339), .A2(n12966), .B1(n14341), .B2(n12989), .C1(
        n15045), .C2(n12965), .ZN(n13047) );
  INV_X1 U15194 ( .A(n13047), .ZN(n12975) );
  INV_X1 U15195 ( .A(n12967), .ZN(n12968) );
  AOI21_X1 U15196 ( .B1(n12970), .B2(n12969), .A(n12968), .ZN(n13048) );
  AOI22_X1 U15197 ( .A1(n15082), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n15077), 
        .B2(n12971), .ZN(n12972) );
  OAI21_X1 U15198 ( .B1(n13109), .B2(n13007), .A(n12972), .ZN(n12973) );
  AOI21_X1 U15199 ( .B1(n13048), .B2(n14346), .A(n12973), .ZN(n12974) );
  OAI21_X1 U15200 ( .B1(n12975), .B2(n15082), .A(n12974), .ZN(P3_U3215) );
  XNOR2_X1 U15201 ( .A(n12976), .B(n12980), .ZN(n12977) );
  OAI222_X1 U15202 ( .A1(n14339), .A2(n12978), .B1(n14341), .B2(n13001), .C1(
        n12977), .C2(n15045), .ZN(n13051) );
  INV_X1 U15203 ( .A(n13051), .ZN(n12985) );
  XNOR2_X1 U15204 ( .A(n12979), .B(n12980), .ZN(n13052) );
  AOI22_X1 U15205 ( .A1(n15082), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15077), 
        .B2(n12981), .ZN(n12982) );
  OAI21_X1 U15206 ( .B1(n13113), .B2(n13007), .A(n12982), .ZN(n12983) );
  AOI21_X1 U15207 ( .B1(n13052), .B2(n14346), .A(n12983), .ZN(n12984) );
  OAI21_X1 U15208 ( .B1(n12985), .B2(n15082), .A(n12984), .ZN(P3_U3216) );
  XNOR2_X1 U15209 ( .A(n12987), .B(n12986), .ZN(n12988) );
  OAI222_X1 U15210 ( .A1(n14339), .A2(n12989), .B1(n14341), .B2(n14329), .C1(
        n12988), .C2(n15045), .ZN(n13055) );
  INV_X1 U15211 ( .A(n13055), .ZN(n12997) );
  XNOR2_X1 U15212 ( .A(n12991), .B(n12990), .ZN(n13056) );
  INV_X1 U15213 ( .A(n12992), .ZN(n13117) );
  AOI22_X1 U15214 ( .A1(n15082), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15077), 
        .B2(n12993), .ZN(n12994) );
  OAI21_X1 U15215 ( .B1(n13117), .B2(n13007), .A(n12994), .ZN(n12995) );
  AOI21_X1 U15216 ( .B1(n13056), .B2(n14346), .A(n12995), .ZN(n12996) );
  OAI21_X1 U15217 ( .B1(n12997), .B2(n15082), .A(n12996), .ZN(P3_U3217) );
  XNOR2_X1 U15218 ( .A(n12998), .B(n13003), .ZN(n12999) );
  OAI222_X1 U15219 ( .A1(n14339), .A2(n13001), .B1(n14341), .B2(n13000), .C1(
        n12999), .C2(n15045), .ZN(n13059) );
  INV_X1 U15220 ( .A(n13059), .ZN(n13010) );
  OAI21_X1 U15221 ( .B1(n13004), .B2(n13003), .A(n13002), .ZN(n13060) );
  AOI22_X1 U15222 ( .A1(n15082), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15077), 
        .B2(n13005), .ZN(n13006) );
  OAI21_X1 U15223 ( .B1(n13122), .B2(n13007), .A(n13006), .ZN(n13008) );
  AOI21_X1 U15224 ( .B1(n13060), .B2(n14346), .A(n13008), .ZN(n13009) );
  OAI21_X1 U15225 ( .B1(n13010), .B2(n15082), .A(n13009), .ZN(P3_U3218) );
  NAND2_X1 U15226 ( .A1(n9450), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n13011) );
  NAND2_X1 U15227 ( .A1(n13064), .A2(n15131), .ZN(n13013) );
  OAI211_X1 U15228 ( .C1(n13066), .C2(n13063), .A(n13011), .B(n13013), .ZN(
        P3_U3490) );
  INV_X1 U15229 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n13015) );
  INV_X1 U15230 ( .A(n13063), .ZN(n13012) );
  NAND2_X1 U15231 ( .A1(n13068), .A2(n13012), .ZN(n13014) );
  OAI211_X1 U15232 ( .C1(n15131), .C2(n13015), .A(n13014), .B(n13013), .ZN(
        P3_U3489) );
  INV_X1 U15233 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13018) );
  AOI21_X1 U15234 ( .B1(n15100), .B2(n13017), .A(n13016), .ZN(n13081) );
  MUX2_X1 U15235 ( .A(n13018), .B(n13081), .S(n15131), .Z(n13019) );
  OAI21_X1 U15236 ( .B1(n13084), .B2(n13063), .A(n13019), .ZN(P3_U3484) );
  AOI22_X1 U15237 ( .A1(n13021), .A2(n15112), .B1(n15071), .B2(n13020), .ZN(
        n13022) );
  NAND2_X1 U15238 ( .A1(n13023), .A2(n13022), .ZN(n13085) );
  MUX2_X1 U15239 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n13085), .S(n15131), .Z(
        P3_U3483) );
  INV_X1 U15240 ( .A(n13024), .ZN(n13089) );
  INV_X1 U15241 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13027) );
  AOI21_X1 U15242 ( .B1(n13026), .B2(n15100), .A(n13025), .ZN(n13086) );
  MUX2_X1 U15243 ( .A(n13027), .B(n13086), .S(n15131), .Z(n13028) );
  OAI21_X1 U15244 ( .B1(n13089), .B2(n13063), .A(n13028), .ZN(P3_U3482) );
  INV_X1 U15245 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13031) );
  AOI21_X1 U15246 ( .B1(n15100), .B2(n13030), .A(n13029), .ZN(n13090) );
  MUX2_X1 U15247 ( .A(n13031), .B(n13090), .S(n15131), .Z(n13032) );
  OAI21_X1 U15248 ( .B1(n13093), .B2(n13063), .A(n13032), .ZN(P3_U3481) );
  INV_X1 U15249 ( .A(n13033), .ZN(n13097) );
  INV_X1 U15250 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13037) );
  INV_X1 U15251 ( .A(n13034), .ZN(n13035) );
  AOI21_X1 U15252 ( .B1(n15100), .B2(n13036), .A(n13035), .ZN(n13094) );
  MUX2_X1 U15253 ( .A(n13037), .B(n13094), .S(n15131), .Z(n13038) );
  OAI21_X1 U15254 ( .B1(n13097), .B2(n13063), .A(n13038), .ZN(P3_U3480) );
  INV_X1 U15255 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13041) );
  AOI21_X1 U15256 ( .B1(n13040), .B2(n15100), .A(n13039), .ZN(n13098) );
  MUX2_X1 U15257 ( .A(n13041), .B(n13098), .S(n15131), .Z(n13042) );
  OAI21_X1 U15258 ( .B1(n13101), .B2(n13063), .A(n13042), .ZN(P3_U3479) );
  INV_X1 U15259 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13045) );
  AOI21_X1 U15260 ( .B1(n15100), .B2(n13044), .A(n13043), .ZN(n13102) );
  MUX2_X1 U15261 ( .A(n13045), .B(n13102), .S(n15131), .Z(n13046) );
  OAI21_X1 U15262 ( .B1(n13105), .B2(n13063), .A(n13046), .ZN(P3_U3478) );
  AOI21_X1 U15263 ( .B1(n13048), .B2(n15100), .A(n13047), .ZN(n13106) );
  MUX2_X1 U15264 ( .A(n13049), .B(n13106), .S(n15131), .Z(n13050) );
  OAI21_X1 U15265 ( .B1(n13109), .B2(n13063), .A(n13050), .ZN(P3_U3477) );
  INV_X1 U15266 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13053) );
  AOI21_X1 U15267 ( .B1(n13052), .B2(n15100), .A(n13051), .ZN(n13110) );
  MUX2_X1 U15268 ( .A(n13053), .B(n13110), .S(n15131), .Z(n13054) );
  OAI21_X1 U15269 ( .B1(n13113), .B2(n13063), .A(n13054), .ZN(P3_U3476) );
  AOI21_X1 U15270 ( .B1(n13056), .B2(n15100), .A(n13055), .ZN(n13114) );
  MUX2_X1 U15271 ( .A(n13057), .B(n13114), .S(n15131), .Z(n13058) );
  OAI21_X1 U15272 ( .B1(n13117), .B2(n13063), .A(n13058), .ZN(P3_U3475) );
  INV_X1 U15273 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13061) );
  AOI21_X1 U15274 ( .B1(n15100), .B2(n13060), .A(n13059), .ZN(n13118) );
  MUX2_X1 U15275 ( .A(n13061), .B(n13118), .S(n15131), .Z(n13062) );
  OAI21_X1 U15276 ( .B1(n13122), .B2(n13063), .A(n13062), .ZN(P3_U3474) );
  NAND2_X1 U15277 ( .A1(n13064), .A2(n15120), .ZN(n13069) );
  NAND2_X1 U15278 ( .A1(n15121), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n13065) );
  OAI211_X1 U15279 ( .C1(n13066), .C2(n13121), .A(n13069), .B(n13065), .ZN(
        P3_U3458) );
  INV_X1 U15280 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n13071) );
  INV_X1 U15281 ( .A(n13121), .ZN(n13067) );
  NAND2_X1 U15282 ( .A1(n13068), .A2(n13067), .ZN(n13070) );
  OAI211_X1 U15283 ( .C1(n15120), .C2(n13071), .A(n13070), .B(n13069), .ZN(
        P3_U3457) );
  NAND2_X1 U15284 ( .A1(n13072), .A2(n15120), .ZN(n13074) );
  OR2_X1 U15285 ( .A1(n15120), .A2(n7907), .ZN(n13073) );
  OAI21_X1 U15286 ( .B1(n13075), .B2(n13121), .A(n7369), .ZN(P3_U3455) );
  INV_X1 U15287 ( .A(n13076), .ZN(n13077) );
  OAI21_X1 U15288 ( .B1(n13080), .B2(n13121), .A(n13079), .ZN(P3_U3454) );
  MUX2_X1 U15289 ( .A(n13082), .B(n13081), .S(n15120), .Z(n13083) );
  OAI21_X1 U15290 ( .B1(n13084), .B2(n13121), .A(n13083), .ZN(P3_U3452) );
  MUX2_X1 U15291 ( .A(P3_REG0_REG_24__SCAN_IN), .B(n13085), .S(n15120), .Z(
        P3_U3451) );
  MUX2_X1 U15292 ( .A(n13087), .B(n13086), .S(n15120), .Z(n13088) );
  OAI21_X1 U15293 ( .B1(n13089), .B2(n13121), .A(n13088), .ZN(P3_U3450) );
  MUX2_X1 U15294 ( .A(n13091), .B(n13090), .S(n15120), .Z(n13092) );
  OAI21_X1 U15295 ( .B1(n13093), .B2(n13121), .A(n13092), .ZN(P3_U3449) );
  MUX2_X1 U15296 ( .A(n13095), .B(n13094), .S(n15120), .Z(n13096) );
  OAI21_X1 U15297 ( .B1(n13097), .B2(n13121), .A(n13096), .ZN(P3_U3448) );
  MUX2_X1 U15298 ( .A(n13099), .B(n13098), .S(n15120), .Z(n13100) );
  OAI21_X1 U15299 ( .B1(n13101), .B2(n13121), .A(n13100), .ZN(P3_U3447) );
  MUX2_X1 U15300 ( .A(n13103), .B(n13102), .S(n15120), .Z(n13104) );
  OAI21_X1 U15301 ( .B1(n13105), .B2(n13121), .A(n13104), .ZN(P3_U3446) );
  MUX2_X1 U15302 ( .A(n13107), .B(n13106), .S(n15120), .Z(n13108) );
  OAI21_X1 U15303 ( .B1(n13109), .B2(n13121), .A(n13108), .ZN(P3_U3444) );
  MUX2_X1 U15304 ( .A(n13111), .B(n13110), .S(n15120), .Z(n13112) );
  OAI21_X1 U15305 ( .B1(n13113), .B2(n13121), .A(n13112), .ZN(P3_U3441) );
  MUX2_X1 U15306 ( .A(n13115), .B(n13114), .S(n15120), .Z(n13116) );
  OAI21_X1 U15307 ( .B1(n13117), .B2(n13121), .A(n13116), .ZN(P3_U3438) );
  MUX2_X1 U15308 ( .A(n13119), .B(n13118), .S(n15120), .Z(n13120) );
  OAI21_X1 U15309 ( .B1(n13122), .B2(n13121), .A(n13120), .ZN(P3_U3435) );
  MUX2_X1 U15310 ( .A(P3_D_REG_1__SCAN_IN), .B(n13123), .S(n13125), .Z(
        P3_U3377) );
  INV_X1 U15311 ( .A(n13124), .ZN(n13126) );
  MUX2_X1 U15312 ( .A(P3_D_REG_0__SCAN_IN), .B(n13126), .S(n13125), .Z(
        P3_U3376) );
  INV_X1 U15313 ( .A(n13127), .ZN(n13131) );
  NOR4_X1 U15314 ( .A1(n13128), .A2(P3_IR_REG_30__SCAN_IN), .A3(n7460), .A4(
        P3_U3151), .ZN(n13129) );
  AOI21_X1 U15315 ( .B1(n14268), .B2(SI_31_), .A(n13129), .ZN(n13130) );
  OAI21_X1 U15316 ( .B1(n13131), .B2(n13138), .A(n13130), .ZN(P3_U3264) );
  INV_X1 U15317 ( .A(n13132), .ZN(n13134) );
  OAI222_X1 U15318 ( .A1(n12303), .A2(n13135), .B1(n13138), .B2(n13134), .C1(
        n13133), .C2(P3_U3151), .ZN(P3_U3266) );
  INV_X1 U15319 ( .A(n13136), .ZN(n13137) );
  OAI222_X1 U15320 ( .A1(n12303), .A2(n13141), .B1(P3_U3151), .B2(n13139), 
        .C1(n13138), .C2(n13137), .ZN(P3_U3267) );
  MUX2_X1 U15321 ( .A(n13143), .B(n13142), .S(P3_STATE_REG_SCAN_IN), .Z(
        P3_U3295) );
  XNOR2_X1 U15322 ( .A(n13145), .B(n13144), .ZN(n13151) );
  INV_X1 U15323 ( .A(n13352), .ZN(n13148) );
  OAI22_X1 U15324 ( .A1(n13188), .A2(n13254), .B1(n13146), .B2(n13256), .ZN(
        n13350) );
  AOI22_X1 U15325 ( .A1(n13257), .A2(n13350), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13147) );
  OAI21_X1 U15326 ( .B1(n13148), .B2(n13259), .A(n13147), .ZN(n13149) );
  AOI21_X1 U15327 ( .B1(n13492), .B2(n13262), .A(n13149), .ZN(n13150) );
  OAI21_X1 U15328 ( .B1(n13151), .B2(n13267), .A(n13150), .ZN(P2_U3186) );
  XNOR2_X1 U15329 ( .A(n13152), .B(n13153), .ZN(n13159) );
  NOR2_X1 U15330 ( .A1(n13187), .A2(n13256), .ZN(n13154) );
  AOI21_X1 U15331 ( .B1(n13288), .B2(n13171), .A(n13154), .ZN(n13511) );
  OAI22_X1 U15332 ( .A1(n13511), .A2(n13272), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13155), .ZN(n13156) );
  AOI21_X1 U15333 ( .B1(n13403), .B2(n13274), .A(n13156), .ZN(n13158) );
  NAND2_X1 U15334 ( .A1(n13514), .A2(n13262), .ZN(n13157) );
  OAI211_X1 U15335 ( .C1(n13159), .C2(n13267), .A(n13158), .B(n13157), .ZN(
        P2_U3188) );
  AOI21_X1 U15336 ( .B1(n13160), .B2(n13161), .A(n13267), .ZN(n13163) );
  NAND2_X1 U15337 ( .A1(n13163), .A2(n13162), .ZN(n13167) );
  AOI22_X1 U15338 ( .A1(n14766), .A2(n13262), .B1(n13257), .B2(n13164), .ZN(
        n13166) );
  MUX2_X1 U15339 ( .A(n13259), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n13165) );
  NAND3_X1 U15340 ( .A1(n13167), .A2(n13166), .A3(n13165), .ZN(P2_U3190) );
  AOI21_X1 U15341 ( .B1(n13170), .B2(n13169), .A(n13168), .ZN(n13177) );
  AOI22_X1 U15342 ( .A1(n13290), .A2(n13172), .B1(n13171), .B2(n13292), .ZN(
        n13461) );
  NAND2_X1 U15343 ( .A1(n13274), .A2(n13468), .ZN(n13173) );
  OAI211_X1 U15344 ( .C1(n13461), .C2(n13272), .A(n13174), .B(n13173), .ZN(
        n13175) );
  AOI21_X1 U15345 ( .B1(n13537), .B2(n13262), .A(n13175), .ZN(n13176) );
  OAI21_X1 U15346 ( .B1(n13177), .B2(n13267), .A(n13176), .ZN(P2_U3191) );
  XNOR2_X1 U15347 ( .A(n13179), .B(n13178), .ZN(n13184) );
  OAI22_X1 U15348 ( .A1(n13180), .A2(n13256), .B1(n7119), .B2(n13254), .ZN(
        n13437) );
  AOI22_X1 U15349 ( .A1(n13437), .A2(n13257), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13181) );
  OAI21_X1 U15350 ( .B1(n13434), .B2(n13259), .A(n13181), .ZN(n13182) );
  AOI21_X1 U15351 ( .B1(n13526), .B2(n13262), .A(n13182), .ZN(n13183) );
  OAI21_X1 U15352 ( .B1(n13184), .B2(n13267), .A(n13183), .ZN(P2_U3195) );
  XNOR2_X1 U15353 ( .A(n13185), .B(n13186), .ZN(n13193) );
  INV_X1 U15354 ( .A(n13380), .ZN(n13190) );
  OAI22_X1 U15355 ( .A1(n13188), .A2(n13256), .B1(n13187), .B2(n13254), .ZN(
        n13376) );
  AOI22_X1 U15356 ( .A1(n13257), .A2(n13376), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13189) );
  OAI21_X1 U15357 ( .B1(n13190), .B2(n13259), .A(n13189), .ZN(n13191) );
  AOI21_X1 U15358 ( .B1(n13502), .B2(n13262), .A(n13191), .ZN(n13192) );
  OAI21_X1 U15359 ( .B1(n13193), .B2(n13267), .A(n13192), .ZN(P2_U3197) );
  OAI21_X1 U15360 ( .B1(n13195), .B2(n13194), .A(n13206), .ZN(n13196) );
  NAND2_X1 U15361 ( .A1(n13196), .A2(n13241), .ZN(n13202) );
  OAI22_X1 U15362 ( .A1(n13272), .A2(n13198), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13197), .ZN(n13199) );
  AOI21_X1 U15363 ( .B1(n13200), .B2(n13274), .A(n13199), .ZN(n13201) );
  OAI211_X1 U15364 ( .C1(n13203), .C2(n13278), .A(n13202), .B(n13201), .ZN(
        P2_U3198) );
  AND3_X1 U15365 ( .A1(n13206), .A2(n13205), .A3(n13204), .ZN(n13207) );
  OAI21_X1 U15366 ( .B1(n13208), .B2(n13207), .A(n13241), .ZN(n13215) );
  INV_X1 U15367 ( .A(n13209), .ZN(n13211) );
  OAI22_X1 U15368 ( .A1(n13272), .A2(n13211), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13210), .ZN(n13212) );
  AOI21_X1 U15369 ( .B1(n13213), .B2(n13274), .A(n13212), .ZN(n13214) );
  OAI211_X1 U15370 ( .C1(n13216), .C2(n13278), .A(n13215), .B(n13214), .ZN(
        P2_U3200) );
  XNOR2_X1 U15371 ( .A(n13217), .B(n13218), .ZN(n13223) );
  INV_X1 U15372 ( .A(n13394), .ZN(n13220) );
  OAI22_X1 U15373 ( .A1(n13234), .A2(n13254), .B1(n13255), .B2(n13256), .ZN(
        n13390) );
  AOI22_X1 U15374 ( .A1(n13257), .A2(n13390), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13219) );
  OAI21_X1 U15375 ( .B1(n13220), .B2(n13259), .A(n13219), .ZN(n13221) );
  AOI21_X1 U15376 ( .B1(n13507), .B2(n13262), .A(n13221), .ZN(n13222) );
  OAI21_X1 U15377 ( .B1(n13223), .B2(n13267), .A(n13222), .ZN(P2_U3201) );
  NOR2_X1 U15378 ( .A1(n13224), .A2(n6598), .ZN(n13225) );
  XNOR2_X1 U15379 ( .A(n13226), .B(n13225), .ZN(n13231) );
  INV_X1 U15380 ( .A(n13450), .ZN(n13228) );
  OAI22_X1 U15381 ( .A1(n13235), .A2(n13256), .B1(n8486), .B2(n13254), .ZN(
        n13445) );
  AOI22_X1 U15382 ( .A1(n13445), .A2(n13257), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13227) );
  OAI21_X1 U15383 ( .B1(n13228), .B2(n13259), .A(n13227), .ZN(n13229) );
  AOI21_X1 U15384 ( .B1(n13531), .B2(n13262), .A(n13229), .ZN(n13230) );
  OAI21_X1 U15385 ( .B1(n13231), .B2(n13267), .A(n13230), .ZN(P2_U3205) );
  XNOR2_X1 U15386 ( .A(n13233), .B(n13232), .ZN(n13240) );
  INV_X1 U15387 ( .A(n13420), .ZN(n13237) );
  OAI22_X1 U15388 ( .A1(n13235), .A2(n13254), .B1(n13234), .B2(n13256), .ZN(
        n13416) );
  AOI22_X1 U15389 ( .A1(n13416), .A2(n13257), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13236) );
  OAI21_X1 U15390 ( .B1(n13237), .B2(n13259), .A(n13236), .ZN(n13238) );
  AOI21_X1 U15391 ( .B1(n13518), .B2(n13262), .A(n13238), .ZN(n13239) );
  OAI21_X1 U15392 ( .B1(n13240), .B2(n13267), .A(n13239), .ZN(P2_U3207) );
  OAI211_X1 U15393 ( .C1(n13244), .C2(n13243), .A(n13242), .B(n13241), .ZN(
        n13249) );
  OAI22_X1 U15394 ( .A1(n13272), .A2(n13245), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13314), .ZN(n13246) );
  AOI21_X1 U15395 ( .B1(n13247), .B2(n13274), .A(n13246), .ZN(n13248) );
  OAI211_X1 U15396 ( .C1(n13543), .C2(n13278), .A(n13249), .B(n13248), .ZN(
        P2_U3210) );
  INV_X1 U15397 ( .A(n13251), .ZN(n13252) );
  AOI21_X1 U15398 ( .B1(n13250), .B2(n13253), .A(n13252), .ZN(n13264) );
  INV_X1 U15399 ( .A(n13366), .ZN(n13260) );
  OAI22_X1 U15400 ( .A1(n6785), .A2(n13256), .B1(n13255), .B2(n13254), .ZN(
        n13361) );
  AOI22_X1 U15401 ( .A1(n13257), .A2(n13361), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13258) );
  OAI21_X1 U15402 ( .B1(n13260), .B2(n13259), .A(n13258), .ZN(n13261) );
  AOI21_X1 U15403 ( .B1(n13497), .B2(n13262), .A(n13261), .ZN(n13263) );
  OAI21_X1 U15404 ( .B1(n13264), .B2(n13267), .A(n13263), .ZN(P2_U3212) );
  AOI211_X1 U15405 ( .C1(n13265), .C2(n13268), .A(n13267), .B(n13266), .ZN(
        n13269) );
  INV_X1 U15406 ( .A(n13269), .ZN(n13277) );
  OAI22_X1 U15407 ( .A1(n13272), .A2(n13271), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13270), .ZN(n13273) );
  AOI21_X1 U15408 ( .B1(n13275), .B2(n13274), .A(n13273), .ZN(n13276) );
  OAI211_X1 U15409 ( .C1(n13279), .C2(n13278), .A(n13277), .B(n13276), .ZN(
        P2_U3213) );
  MUX2_X1 U15410 ( .A(n13325), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13309), .Z(
        P2_U3562) );
  MUX2_X1 U15411 ( .A(n13280), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13309), .Z(
        P2_U3561) );
  MUX2_X1 U15412 ( .A(n13281), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13309), .Z(
        P2_U3560) );
  MUX2_X1 U15413 ( .A(n13282), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13309), .Z(
        P2_U3559) );
  MUX2_X1 U15414 ( .A(n13283), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13309), .Z(
        P2_U3558) );
  MUX2_X1 U15415 ( .A(n13284), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13309), .Z(
        P2_U3557) );
  MUX2_X1 U15416 ( .A(n13285), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13309), .Z(
        P2_U3556) );
  MUX2_X1 U15417 ( .A(n13286), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13309), .Z(
        P2_U3555) );
  MUX2_X1 U15418 ( .A(n13287), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13309), .Z(
        P2_U3554) );
  MUX2_X1 U15419 ( .A(n13288), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13309), .Z(
        P2_U3553) );
  MUX2_X1 U15420 ( .A(n13289), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13309), .Z(
        P2_U3552) );
  MUX2_X1 U15421 ( .A(n13290), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13309), .Z(
        P2_U3551) );
  INV_X2 U15422 ( .A(P2_U3947), .ZN(n13309) );
  MUX2_X1 U15423 ( .A(n13291), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13309), .Z(
        P2_U3550) );
  MUX2_X1 U15424 ( .A(n13292), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13309), .Z(
        P2_U3549) );
  MUX2_X1 U15425 ( .A(n13293), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13309), .Z(
        P2_U3548) );
  MUX2_X1 U15426 ( .A(n13294), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13309), .Z(
        P2_U3547) );
  MUX2_X1 U15427 ( .A(n13295), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13309), .Z(
        P2_U3546) );
  MUX2_X1 U15428 ( .A(n13296), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13309), .Z(
        P2_U3545) );
  MUX2_X1 U15429 ( .A(n13297), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13309), .Z(
        P2_U3544) );
  MUX2_X1 U15430 ( .A(n13298), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13309), .Z(
        P2_U3543) );
  MUX2_X1 U15431 ( .A(n13299), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13309), .Z(
        P2_U3542) );
  MUX2_X1 U15432 ( .A(n13300), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13309), .Z(
        P2_U3541) );
  MUX2_X1 U15433 ( .A(n13301), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13309), .Z(
        P2_U3540) );
  MUX2_X1 U15434 ( .A(n13302), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13309), .Z(
        P2_U3539) );
  MUX2_X1 U15435 ( .A(n13303), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13309), .Z(
        P2_U3538) );
  MUX2_X1 U15436 ( .A(n13304), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13309), .Z(
        P2_U3537) );
  MUX2_X1 U15437 ( .A(n13305), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13309), .Z(
        P2_U3536) );
  MUX2_X1 U15438 ( .A(n13306), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13309), .Z(
        P2_U3535) );
  MUX2_X1 U15439 ( .A(n13307), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13309), .Z(
        P2_U3534) );
  MUX2_X1 U15440 ( .A(n6995), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13309), .Z(
        P2_U3533) );
  MUX2_X1 U15441 ( .A(n13308), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13309), .Z(
        P2_U3532) );
  MUX2_X1 U15442 ( .A(n13310), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13309), .Z(
        P2_U3531) );
  AOI21_X1 U15443 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n13312), .A(n13311), 
        .ZN(n13313) );
  OR2_X1 U15444 ( .A1(n13313), .A2(n14652), .ZN(n13322) );
  NOR2_X1 U15445 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n13314), .ZN(n13315) );
  AOI21_X1 U15446 ( .B1(n14684), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n13315), 
        .ZN(n13321) );
  OAI211_X1 U15447 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n13317), .A(n14688), 
        .B(n13316), .ZN(n13320) );
  NAND2_X1 U15448 ( .A1(n14685), .A2(n13318), .ZN(n13319) );
  NAND4_X1 U15449 ( .A1(n13322), .A2(n13321), .A3(n13320), .A4(n13319), .ZN(
        P2_U3232) );
  NAND2_X1 U15450 ( .A1(n13329), .A2(n13479), .ZN(n13328) );
  XNOR2_X1 U15451 ( .A(n9634), .B(n13328), .ZN(n13323) );
  NAND2_X1 U15452 ( .A1(n13323), .A2(n11440), .ZN(n13476) );
  NAND2_X1 U15453 ( .A1(n13325), .A2(n13324), .ZN(n13477) );
  NOR2_X1 U15454 ( .A1(n14736), .A2(n13477), .ZN(n13331) );
  NOR2_X1 U15455 ( .A1(n9634), .A2(n13453), .ZN(n13326) );
  AOI211_X1 U15456 ( .C1(n14736), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13331), 
        .B(n13326), .ZN(n13327) );
  OAI21_X1 U15457 ( .B1(n13476), .B2(n14714), .A(n13327), .ZN(P2_U3234) );
  OAI211_X1 U15458 ( .C1(n13329), .C2(n13479), .A(n11440), .B(n13328), .ZN(
        n13478) );
  NOR2_X1 U15459 ( .A1(n13479), .A2(n13453), .ZN(n13330) );
  AOI211_X1 U15460 ( .C1(n14736), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13331), 
        .B(n13330), .ZN(n13332) );
  OAI21_X1 U15461 ( .B1(n14714), .B2(n13478), .A(n13332), .ZN(P2_U3235) );
  AOI211_X1 U15462 ( .C1(n13338), .C2(n13334), .A(n13462), .B(n13333), .ZN(
        n13336) );
  NOR2_X1 U15463 ( .A1(n13336), .A2(n13335), .ZN(n13489) );
  OAI21_X1 U15464 ( .B1(n13339), .B2(n13338), .A(n13337), .ZN(n13490) );
  INV_X1 U15465 ( .A(n13490), .ZN(n13347) );
  OAI211_X1 U15466 ( .C1(n13341), .C2(n6492), .A(n11440), .B(n13340), .ZN(
        n13485) );
  INV_X1 U15467 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13343) );
  OAI22_X1 U15468 ( .A1(n14733), .A2(n13343), .B1(n13342), .B2(n14724), .ZN(
        n13344) );
  AOI21_X1 U15469 ( .B1(n13487), .B2(n14706), .A(n13344), .ZN(n13345) );
  OAI21_X1 U15470 ( .B1(n13485), .B2(n14714), .A(n13345), .ZN(n13346) );
  AOI21_X1 U15471 ( .B1(n13347), .B2(n13426), .A(n13346), .ZN(n13348) );
  OAI21_X1 U15472 ( .B1(n13489), .B2(n14736), .A(n13348), .ZN(P2_U3237) );
  XNOR2_X1 U15473 ( .A(n13349), .B(n13355), .ZN(n13351) );
  AOI21_X1 U15474 ( .B1(n13351), .B2(n14725), .A(n13350), .ZN(n13494) );
  AOI211_X1 U15475 ( .C1(n13492), .C2(n13363), .A(n11505), .B(n6492), .ZN(
        n13491) );
  AOI22_X1 U15476 ( .A1(n14736), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n13352), 
        .B2(n14705), .ZN(n13353) );
  OAI21_X1 U15477 ( .B1(n6882), .B2(n13453), .A(n13353), .ZN(n13358) );
  OAI21_X1 U15478 ( .B1(n13356), .B2(n13355), .A(n13354), .ZN(n13495) );
  NOR2_X1 U15479 ( .A1(n13495), .A2(n14715), .ZN(n13357) );
  AOI211_X1 U15480 ( .C1(n13491), .C2(n13473), .A(n13358), .B(n13357), .ZN(
        n13359) );
  OAI21_X1 U15481 ( .B1(n14736), .B2(n13494), .A(n13359), .ZN(P2_U3238) );
  XNOR2_X1 U15482 ( .A(n13360), .B(n13370), .ZN(n13362) );
  AOI21_X1 U15483 ( .B1(n13362), .B2(n14725), .A(n13361), .ZN(n13499) );
  INV_X1 U15484 ( .A(n13378), .ZN(n13365) );
  INV_X1 U15485 ( .A(n13363), .ZN(n13364) );
  AOI211_X1 U15486 ( .C1(n13497), .C2(n13365), .A(n11505), .B(n13364), .ZN(
        n13496) );
  AOI22_X1 U15487 ( .A1(n14736), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n13366), 
        .B2(n14705), .ZN(n13367) );
  OAI21_X1 U15488 ( .B1(n13368), .B2(n13453), .A(n13367), .ZN(n13372) );
  XOR2_X1 U15489 ( .A(n13370), .B(n13369), .Z(n13500) );
  NOR2_X1 U15490 ( .A1(n13500), .A2(n14715), .ZN(n13371) );
  AOI211_X1 U15491 ( .C1(n13496), .C2(n13473), .A(n13372), .B(n13371), .ZN(
        n13373) );
  OAI21_X1 U15492 ( .B1(n14736), .B2(n13499), .A(n13373), .ZN(P2_U3239) );
  XNOR2_X1 U15493 ( .A(n13375), .B(n13374), .ZN(n13377) );
  AOI21_X1 U15494 ( .B1(n13377), .B2(n14725), .A(n13376), .ZN(n13504) );
  INV_X1 U15495 ( .A(n13392), .ZN(n13379) );
  AOI211_X1 U15496 ( .C1(n13502), .C2(n13379), .A(n11505), .B(n13378), .ZN(
        n13501) );
  AOI22_X1 U15497 ( .A1(n14736), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n13380), 
        .B2(n14705), .ZN(n13381) );
  OAI21_X1 U15498 ( .B1(n13382), .B2(n13453), .A(n13381), .ZN(n13387) );
  AOI21_X1 U15499 ( .B1(n13385), .B2(n13384), .A(n13383), .ZN(n13505) );
  NOR2_X1 U15500 ( .A1(n13505), .A2(n14715), .ZN(n13386) );
  AOI211_X1 U15501 ( .C1(n13501), .C2(n13473), .A(n13387), .B(n13386), .ZN(
        n13388) );
  OAI21_X1 U15502 ( .B1(n13504), .B2(n14736), .A(n13388), .ZN(P2_U3240) );
  XNOR2_X1 U15503 ( .A(n13389), .B(n13398), .ZN(n13391) );
  AOI21_X1 U15504 ( .B1(n13391), .B2(n14725), .A(n13390), .ZN(n13509) );
  INV_X1 U15505 ( .A(n13409), .ZN(n13393) );
  AOI211_X1 U15506 ( .C1(n13507), .C2(n13393), .A(n11505), .B(n13392), .ZN(
        n13506) );
  AOI22_X1 U15507 ( .A1(n14736), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n13394), 
        .B2(n14705), .ZN(n13395) );
  OAI21_X1 U15508 ( .B1(n13396), .B2(n13453), .A(n13395), .ZN(n13400) );
  XNOR2_X1 U15509 ( .A(n13397), .B(n13398), .ZN(n13510) );
  NOR2_X1 U15510 ( .A1(n13510), .A2(n14715), .ZN(n13399) );
  AOI211_X1 U15511 ( .C1(n13506), .C2(n13473), .A(n13400), .B(n13399), .ZN(
        n13401) );
  OAI21_X1 U15512 ( .B1(n13509), .B2(n14736), .A(n13401), .ZN(P2_U3241) );
  XOR2_X1 U15513 ( .A(n13402), .B(n13405), .Z(n13517) );
  INV_X1 U15514 ( .A(n13403), .ZN(n13407) );
  XOR2_X1 U15515 ( .A(n13405), .B(n13404), .Z(n13406) );
  NAND2_X1 U15516 ( .A1(n13406), .A2(n14725), .ZN(n13516) );
  OAI211_X1 U15517 ( .C1(n14724), .C2(n13407), .A(n13516), .B(n13511), .ZN(
        n13408) );
  NAND2_X1 U15518 ( .A1(n13408), .A2(n14733), .ZN(n13414) );
  AOI211_X1 U15519 ( .C1(n13514), .C2(n13418), .A(n11505), .B(n13409), .ZN(
        n13512) );
  INV_X1 U15520 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n13410) );
  OAI22_X1 U15521 ( .A1(n13411), .A2(n13453), .B1(n14733), .B2(n13410), .ZN(
        n13412) );
  AOI21_X1 U15522 ( .B1(n13512), .B2(n13473), .A(n13412), .ZN(n13413) );
  OAI211_X1 U15523 ( .C1(n13517), .C2(n14715), .A(n13414), .B(n13413), .ZN(
        P2_U3242) );
  XNOR2_X1 U15524 ( .A(n13415), .B(n13424), .ZN(n13417) );
  AOI21_X1 U15525 ( .B1(n13417), .B2(n14725), .A(n13416), .ZN(n13524) );
  AOI21_X1 U15526 ( .B1(n13518), .B2(n13431), .A(n11505), .ZN(n13419) );
  NAND2_X1 U15527 ( .A1(n13419), .A2(n13418), .ZN(n13521) );
  AOI22_X1 U15528 ( .A1(n13420), .A2(n14705), .B1(n14736), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n13422) );
  NAND2_X1 U15529 ( .A1(n13518), .A2(n14706), .ZN(n13421) );
  OAI211_X1 U15530 ( .C1(n13521), .C2(n14714), .A(n13422), .B(n13421), .ZN(
        n13423) );
  INV_X1 U15531 ( .A(n13423), .ZN(n13428) );
  NAND2_X1 U15532 ( .A1(n13425), .A2(n13424), .ZN(n13519) );
  NAND3_X1 U15533 ( .A1(n13520), .A2(n13519), .A3(n13426), .ZN(n13427) );
  OAI211_X1 U15534 ( .C1(n13524), .C2(n14736), .A(n13428), .B(n13427), .ZN(
        P2_U3243) );
  XOR2_X1 U15535 ( .A(n13429), .B(n13436), .Z(n13529) );
  NAND2_X1 U15536 ( .A1(n6885), .A2(n13526), .ZN(n13430) );
  AND3_X1 U15537 ( .A1(n13431), .A2(n13430), .A3(n11440), .ZN(n13525) );
  NAND2_X1 U15538 ( .A1(n13526), .A2(n14706), .ZN(n13433) );
  NAND2_X1 U15539 ( .A1(n14736), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n13432) );
  OAI211_X1 U15540 ( .C1(n14724), .C2(n13434), .A(n13433), .B(n13432), .ZN(
        n13440) );
  XOR2_X1 U15541 ( .A(n13436), .B(n13435), .Z(n13438) );
  AOI21_X1 U15542 ( .B1(n13438), .B2(n14725), .A(n13437), .ZN(n13528) );
  NOR2_X1 U15543 ( .A1(n13528), .A2(n14736), .ZN(n13439) );
  AOI211_X1 U15544 ( .C1(n13525), .C2(n13473), .A(n13440), .B(n13439), .ZN(
        n13441) );
  OAI21_X1 U15545 ( .B1(n14715), .B2(n13529), .A(n13441), .ZN(P2_U3244) );
  XNOR2_X1 U15546 ( .A(n13442), .B(n13443), .ZN(n13534) );
  XNOR2_X1 U15547 ( .A(n13444), .B(n13443), .ZN(n13446) );
  AOI21_X1 U15548 ( .B1(n13446), .B2(n14725), .A(n13445), .ZN(n13533) );
  INV_X1 U15549 ( .A(n13533), .ZN(n13456) );
  NAND2_X1 U15550 ( .A1(n13531), .A2(n13467), .ZN(n13447) );
  NAND2_X1 U15551 ( .A1(n13447), .A2(n11440), .ZN(n13448) );
  NOR2_X1 U15552 ( .A1(n13449), .A2(n13448), .ZN(n13530) );
  NAND2_X1 U15553 ( .A1(n13530), .A2(n13473), .ZN(n13452) );
  AOI22_X1 U15554 ( .A1(n14736), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13450), 
        .B2(n14705), .ZN(n13451) );
  OAI211_X1 U15555 ( .C1(n13454), .C2(n13453), .A(n13452), .B(n13451), .ZN(
        n13455) );
  AOI21_X1 U15556 ( .B1(n13456), .B2(n14733), .A(n13455), .ZN(n13457) );
  OAI21_X1 U15557 ( .B1(n13534), .B2(n14715), .A(n13457), .ZN(P2_U3245) );
  XNOR2_X1 U15558 ( .A(n13458), .B(n13459), .ZN(n13539) );
  XNOR2_X1 U15559 ( .A(n13460), .B(n13459), .ZN(n13463) );
  OAI21_X1 U15560 ( .B1(n13463), .B2(n13462), .A(n13461), .ZN(n13535) );
  NAND2_X1 U15561 ( .A1(n13535), .A2(n14733), .ZN(n13475) );
  OR2_X1 U15562 ( .A1(n13465), .A2(n13464), .ZN(n13466) );
  AND3_X1 U15563 ( .A1(n13467), .A2(n11440), .A3(n13466), .ZN(n13536) );
  INV_X1 U15564 ( .A(n13468), .ZN(n13471) );
  NAND2_X1 U15565 ( .A1(n13537), .A2(n14706), .ZN(n13470) );
  NAND2_X1 U15566 ( .A1(n14736), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n13469) );
  OAI211_X1 U15567 ( .C1(n14724), .C2(n13471), .A(n13470), .B(n13469), .ZN(
        n13472) );
  AOI21_X1 U15568 ( .B1(n13536), .B2(n13473), .A(n13472), .ZN(n13474) );
  OAI211_X1 U15569 ( .C1(n13539), .C2(n14715), .A(n13475), .B(n13474), .ZN(
        P2_U3246) );
  OAI211_X1 U15570 ( .C1(n9634), .C2(n14822), .A(n13476), .B(n13477), .ZN(
        n13561) );
  MUX2_X1 U15571 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13561), .S(n14853), .Z(
        P2_U3530) );
  OAI211_X1 U15572 ( .C1(n13479), .C2(n14822), .A(n13478), .B(n13477), .ZN(
        n13562) );
  MUX2_X1 U15573 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13562), .S(n14853), .Z(
        P2_U3529) );
  AOI21_X1 U15574 ( .B1(n14814), .B2(n13482), .A(n13481), .ZN(n13483) );
  INV_X1 U15575 ( .A(n13485), .ZN(n13486) );
  AOI21_X1 U15576 ( .B1(n14814), .B2(n13487), .A(n13486), .ZN(n13488) );
  OAI211_X1 U15577 ( .C1(n14817), .C2(n13490), .A(n13489), .B(n13488), .ZN(
        n13564) );
  MUX2_X1 U15578 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13564), .S(n14853), .Z(
        P2_U3527) );
  AOI21_X1 U15579 ( .B1(n14814), .B2(n13492), .A(n13491), .ZN(n13493) );
  OAI211_X1 U15580 ( .C1(n14817), .C2(n13495), .A(n13494), .B(n13493), .ZN(
        n13565) );
  MUX2_X1 U15581 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13565), .S(n14853), .Z(
        P2_U3526) );
  AOI21_X1 U15582 ( .B1(n14814), .B2(n13497), .A(n13496), .ZN(n13498) );
  OAI211_X1 U15583 ( .C1(n14817), .C2(n13500), .A(n13499), .B(n13498), .ZN(
        n13566) );
  MUX2_X1 U15584 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13566), .S(n14853), .Z(
        P2_U3525) );
  AOI21_X1 U15585 ( .B1(n14814), .B2(n13502), .A(n13501), .ZN(n13503) );
  OAI211_X1 U15586 ( .C1(n14817), .C2(n13505), .A(n13504), .B(n13503), .ZN(
        n13567) );
  MUX2_X1 U15587 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13567), .S(n14853), .Z(
        P2_U3524) );
  AOI21_X1 U15588 ( .B1(n14814), .B2(n13507), .A(n13506), .ZN(n13508) );
  OAI211_X1 U15589 ( .C1(n14817), .C2(n13510), .A(n13509), .B(n13508), .ZN(
        n13568) );
  MUX2_X1 U15590 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13568), .S(n14853), .Z(
        P2_U3523) );
  INV_X1 U15591 ( .A(n13511), .ZN(n13513) );
  AOI211_X1 U15592 ( .C1(n14814), .C2(n13514), .A(n13513), .B(n13512), .ZN(
        n13515) );
  OAI211_X1 U15593 ( .C1(n14817), .C2(n13517), .A(n13516), .B(n13515), .ZN(
        n13569) );
  MUX2_X1 U15594 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13569), .S(n14853), .Z(
        P2_U3522) );
  NAND2_X1 U15595 ( .A1(n13518), .A2(n14814), .ZN(n13523) );
  NAND3_X1 U15596 ( .A1(n13520), .A2(n13519), .A3(n14809), .ZN(n13522) );
  NAND4_X1 U15597 ( .A1(n13524), .A2(n13523), .A3(n13522), .A4(n13521), .ZN(
        n13570) );
  MUX2_X1 U15598 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13570), .S(n14853), .Z(
        P2_U3521) );
  AOI21_X1 U15599 ( .B1(n14814), .B2(n13526), .A(n13525), .ZN(n13527) );
  OAI211_X1 U15600 ( .C1(n14817), .C2(n13529), .A(n13528), .B(n13527), .ZN(
        n13571) );
  MUX2_X1 U15601 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13571), .S(n14853), .Z(
        P2_U3520) );
  AOI21_X1 U15602 ( .B1(n14814), .B2(n13531), .A(n13530), .ZN(n13532) );
  OAI211_X1 U15603 ( .C1(n14817), .C2(n13534), .A(n13533), .B(n13532), .ZN(
        n13572) );
  MUX2_X1 U15604 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13572), .S(n14853), .Z(
        P2_U3519) );
  AOI211_X1 U15605 ( .C1(n14814), .C2(n13537), .A(n13536), .B(n13535), .ZN(
        n13538) );
  OAI21_X1 U15606 ( .B1(n14817), .B2(n13539), .A(n13538), .ZN(n13573) );
  MUX2_X1 U15607 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13573), .S(n14853), .Z(
        P2_U3518) );
  NAND2_X1 U15608 ( .A1(n13540), .A2(n14809), .ZN(n13542) );
  OAI211_X1 U15609 ( .C1(n13543), .C2(n14822), .A(n13542), .B(n13541), .ZN(
        n13545) );
  MUX2_X1 U15610 ( .A(n13574), .B(P2_REG1_REG_18__SCAN_IN), .S(n14850), .Z(
        P2_U3517) );
  AOI21_X1 U15611 ( .B1(n14814), .B2(n13547), .A(n13546), .ZN(n13548) );
  OAI211_X1 U15612 ( .C1(n14817), .C2(n13550), .A(n13549), .B(n13548), .ZN(
        n13575) );
  MUX2_X1 U15613 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13575), .S(n14853), .Z(
        P2_U3516) );
  AOI211_X1 U15614 ( .C1(n14814), .C2(n13553), .A(n13552), .B(n13551), .ZN(
        n13554) );
  OAI21_X1 U15615 ( .B1(n14817), .B2(n13555), .A(n13554), .ZN(n13576) );
  MUX2_X1 U15616 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13576), .S(n14853), .Z(
        P2_U3515) );
  AOI21_X1 U15617 ( .B1(n14814), .B2(n13557), .A(n13556), .ZN(n13558) );
  OAI211_X1 U15618 ( .C1(n14817), .C2(n13560), .A(n13559), .B(n13558), .ZN(
        n13577) );
  MUX2_X1 U15619 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n13577), .S(n14853), .Z(
        P2_U3513) );
  MUX2_X1 U15620 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13561), .S(n14831), .Z(
        P2_U3498) );
  MUX2_X1 U15621 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13562), .S(n14831), .Z(
        P2_U3497) );
  MUX2_X1 U15622 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13564), .S(n14831), .Z(
        P2_U3495) );
  MUX2_X1 U15623 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13565), .S(n14831), .Z(
        P2_U3494) );
  MUX2_X1 U15624 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13566), .S(n14831), .Z(
        P2_U3493) );
  MUX2_X1 U15625 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13567), .S(n14831), .Z(
        P2_U3492) );
  MUX2_X1 U15626 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13568), .S(n14831), .Z(
        P2_U3491) );
  MUX2_X1 U15627 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13569), .S(n14831), .Z(
        P2_U3490) );
  MUX2_X1 U15628 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13570), .S(n14831), .Z(
        P2_U3489) );
  MUX2_X1 U15629 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13571), .S(n14831), .Z(
        P2_U3488) );
  MUX2_X1 U15630 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13572), .S(n14831), .Z(
        P2_U3487) );
  MUX2_X1 U15631 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13573), .S(n14831), .Z(
        P2_U3486) );
  MUX2_X1 U15632 ( .A(n13574), .B(P2_REG0_REG_18__SCAN_IN), .S(n14829), .Z(
        P2_U3484) );
  MUX2_X1 U15633 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13575), .S(n14831), .Z(
        P2_U3481) );
  MUX2_X1 U15634 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13576), .S(n14831), .Z(
        P2_U3478) );
  MUX2_X1 U15635 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n13577), .S(n14831), .Z(
        P2_U3472) );
  OAI222_X1 U15636 ( .A1(n13589), .A2(n13580), .B1(P2_U3088), .B2(n13579), 
        .C1(n13578), .C2(n13591), .ZN(P2_U3297) );
  INV_X1 U15637 ( .A(n13581), .ZN(n14243) );
  OAI222_X1 U15638 ( .A1(n13589), .A2(n14243), .B1(P2_U3088), .B2(n13583), 
        .C1(n13582), .C2(n13591), .ZN(P2_U3298) );
  AOI21_X1 U15639 ( .B1(n13593), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13584), 
        .ZN(n13585) );
  OAI21_X1 U15640 ( .B1(n13586), .B2(n13596), .A(n13585), .ZN(P2_U3299) );
  INV_X1 U15641 ( .A(n13587), .ZN(n14247) );
  OAI222_X1 U15642 ( .A1(n13591), .A2(n13590), .B1(n13589), .B2(n14247), .C1(
        P2_U3088), .C2(n13588), .ZN(P2_U3300) );
  INV_X1 U15643 ( .A(n13592), .ZN(n14250) );
  AOI22_X1 U15644 ( .A1(n13594), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n13593), .ZN(n13595) );
  OAI21_X1 U15645 ( .B1(n14250), .B2(n13596), .A(n13595), .ZN(P2_U3301) );
  INV_X1 U15646 ( .A(n13597), .ZN(n13598) );
  MUX2_X1 U15647 ( .A(n13598), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  OAI21_X1 U15648 ( .B1(n13601), .B2(n13599), .A(n13600), .ZN(n13602) );
  INV_X1 U15649 ( .A(n13602), .ZN(n13608) );
  NAND2_X1 U15650 ( .A1(n13914), .A2(n13717), .ZN(n13604) );
  NAND2_X1 U15651 ( .A1(n13749), .A2(n13913), .ZN(n13603) );
  NAND2_X1 U15652 ( .A1(n13604), .A2(n13603), .ZN(n13934) );
  AOI22_X1 U15653 ( .A1(n14411), .A2(n13934), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13605) );
  OAI21_X1 U15654 ( .B1(n13939), .B2(n14417), .A(n13605), .ZN(n13606) );
  AOI21_X1 U15655 ( .B1(n14203), .B2(n6468), .A(n13606), .ZN(n13607) );
  OAI21_X1 U15656 ( .B1(n13608), .B2(n13731), .A(n13607), .ZN(P1_U3214) );
  NAND2_X1 U15657 ( .A1(n13751), .A2(n13717), .ZN(n13609) );
  OAI21_X1 U15658 ( .B1(n13634), .B2(n13624), .A(n13609), .ZN(n14141) );
  AOI22_X1 U15659 ( .A1(n14411), .A2(n14141), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13610) );
  OAI21_X1 U15660 ( .B1(n14000), .B2(n14417), .A(n13610), .ZN(n13618) );
  NAND2_X1 U15661 ( .A1(n13611), .A2(n13613), .ZN(n13678) );
  INV_X1 U15662 ( .A(n13613), .ZN(n13614) );
  NAND3_X1 U15663 ( .A1(n13705), .A2(n13615), .A3(n13614), .ZN(n13616) );
  AOI21_X1 U15664 ( .B1(n13678), .B2(n13616), .A(n13731), .ZN(n13617) );
  AOI211_X1 U15665 ( .C1(n14142), .C2(n6468), .A(n13618), .B(n13617), .ZN(
        n13619) );
  INV_X1 U15666 ( .A(n13619), .ZN(P1_U3216) );
  OAI21_X1 U15667 ( .B1(n6514), .B2(n13621), .A(n13620), .ZN(n13623) );
  NAND3_X1 U15668 ( .A1(n13623), .A2(n14409), .A3(n13622), .ZN(n13630) );
  INV_X1 U15669 ( .A(n14066), .ZN(n13628) );
  NOR2_X1 U15670 ( .A1(n13625), .A2(n13624), .ZN(n13626) );
  AOI21_X1 U15671 ( .B1(n13755), .B2(n13717), .A(n13626), .ZN(n14165) );
  NAND2_X1 U15672 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13885)
         );
  OAI21_X1 U15673 ( .B1(n13739), .B2(n14165), .A(n13885), .ZN(n13627) );
  AOI21_X1 U15674 ( .B1(n13742), .B2(n13628), .A(n13627), .ZN(n13629) );
  OAI211_X1 U15675 ( .C1(n14167), .C2(n13745), .A(n13630), .B(n13629), .ZN(
        P1_U3219) );
  AOI21_X1 U15676 ( .B1(n13631), .B2(n13632), .A(n6490), .ZN(n13640) );
  NOR2_X1 U15677 ( .A1(n13634), .A2(n13633), .ZN(n13635) );
  AOI21_X1 U15678 ( .B1(n13755), .B2(n13913), .A(n13635), .ZN(n14033) );
  INV_X1 U15679 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n13636) );
  OAI22_X1 U15680 ( .A1(n13739), .A2(n14033), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13636), .ZN(n13638) );
  NOR2_X1 U15681 ( .A1(n14038), .A2(n13745), .ZN(n13637) );
  AOI211_X1 U15682 ( .C1(n13742), .C2(n14035), .A(n13638), .B(n13637), .ZN(
        n13639) );
  OAI21_X1 U15683 ( .B1(n13640), .B2(n13731), .A(n13639), .ZN(P1_U3223) );
  AOI21_X1 U15684 ( .B1(n13642), .B2(n13641), .A(n13731), .ZN(n13644) );
  NAND2_X1 U15685 ( .A1(n13644), .A2(n13643), .ZN(n13651) );
  INV_X1 U15686 ( .A(n13645), .ZN(n13649) );
  OAI21_X1 U15687 ( .B1(n13739), .B2(n13647), .A(n13646), .ZN(n13648) );
  AOI21_X1 U15688 ( .B1(n13742), .B2(n13649), .A(n13648), .ZN(n13650) );
  OAI211_X1 U15689 ( .C1(n13652), .C2(n13745), .A(n13651), .B(n13650), .ZN(
        P1_U3224) );
  XOR2_X1 U15690 ( .A(n13654), .B(n13653), .Z(n13661) );
  NOR2_X1 U15691 ( .A1(n14417), .A2(n13655), .ZN(n13659) );
  OAI21_X1 U15692 ( .B1(n13739), .B2(n13657), .A(n13656), .ZN(n13658) );
  AOI211_X1 U15693 ( .C1(n14189), .C2(n6468), .A(n13659), .B(n13658), .ZN(
        n13660) );
  OAI21_X1 U15694 ( .B1(n13661), .B2(n13731), .A(n13660), .ZN(P1_U3226) );
  XNOR2_X1 U15695 ( .A(n13663), .B(n13662), .ZN(n13664) );
  XNOR2_X1 U15696 ( .A(n13665), .B(n13664), .ZN(n13672) );
  NAND2_X1 U15697 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13844)
         );
  NAND2_X1 U15698 ( .A1(n14411), .A2(n13666), .ZN(n13667) );
  OAI211_X1 U15699 ( .C1(n14417), .C2(n13668), .A(n13844), .B(n13667), .ZN(
        n13669) );
  AOI21_X1 U15700 ( .B1(n13670), .B2(n6468), .A(n13669), .ZN(n13671) );
  OAI21_X1 U15701 ( .B1(n13672), .B2(n13731), .A(n13671), .ZN(P1_U3228) );
  NAND2_X1 U15702 ( .A1(n13752), .A2(n13913), .ZN(n13674) );
  NAND2_X1 U15703 ( .A1(n13750), .A2(n13717), .ZN(n13673) );
  NAND2_X1 U15704 ( .A1(n13674), .A2(n13673), .ZN(n13980) );
  AOI22_X1 U15705 ( .A1(n14411), .A2(n13980), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13675) );
  OAI21_X1 U15706 ( .B1(n13987), .B2(n14417), .A(n13675), .ZN(n13682) );
  NAND3_X1 U15707 ( .A1(n13678), .A2(n13677), .A3(n13676), .ZN(n13679) );
  AOI21_X1 U15708 ( .B1(n13680), .B2(n13679), .A(n13731), .ZN(n13681) );
  INV_X1 U15709 ( .A(n13684), .ZN(P1_U3229) );
  XNOR2_X1 U15710 ( .A(n13686), .B(n13685), .ZN(n13692) );
  NOR2_X1 U15711 ( .A1(n14417), .A2(n14055), .ZN(n13690) );
  AND2_X1 U15712 ( .A1(n13756), .A2(n13913), .ZN(n13687) );
  AOI21_X1 U15713 ( .B1(n13754), .B2(n13717), .A(n13687), .ZN(n14047) );
  OAI22_X1 U15714 ( .A1(n14047), .A2(n13739), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13688), .ZN(n13689) );
  AOI211_X1 U15715 ( .C1(n14222), .C2(n6468), .A(n13690), .B(n13689), .ZN(
        n13691) );
  OAI21_X1 U15716 ( .B1(n13692), .B2(n13731), .A(n13691), .ZN(P1_U3233) );
  OAI211_X1 U15717 ( .C1(n13694), .C2(n13693), .A(n14393), .B(n14409), .ZN(
        n13701) );
  INV_X1 U15718 ( .A(n13695), .ZN(n13699) );
  OAI21_X1 U15719 ( .B1(n13739), .B2(n13697), .A(n13696), .ZN(n13698) );
  AOI21_X1 U15720 ( .B1(n13742), .B2(n13699), .A(n13698), .ZN(n13700) );
  OAI211_X1 U15721 ( .C1(n13702), .C2(n13745), .A(n13701), .B(n13700), .ZN(
        P1_U3234) );
  NOR3_X1 U15722 ( .A1(n6490), .A2(n6732), .A3(n13704), .ZN(n13707) );
  INV_X1 U15723 ( .A(n13705), .ZN(n13706) );
  OAI21_X1 U15724 ( .B1(n13707), .B2(n13706), .A(n14409), .ZN(n13713) );
  INV_X1 U15725 ( .A(n14011), .ZN(n13711) );
  AND2_X1 U15726 ( .A1(n13752), .A2(n13717), .ZN(n13708) );
  AOI21_X1 U15727 ( .B1(n13754), .B2(n13913), .A(n13708), .ZN(n14016) );
  INV_X1 U15728 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13709) );
  OAI22_X1 U15729 ( .A1(n14016), .A2(n13739), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13709), .ZN(n13710) );
  AOI21_X1 U15730 ( .B1(n13742), .B2(n13711), .A(n13710), .ZN(n13712) );
  OAI211_X1 U15731 ( .C1(n13745), .C2(n14218), .A(n13713), .B(n13712), .ZN(
        P1_U3235) );
  AOI21_X1 U15732 ( .B1(n13715), .B2(n13714), .A(n6514), .ZN(n13721) );
  NOR2_X1 U15733 ( .A1(n14417), .A2(n14078), .ZN(n13719) );
  AND2_X1 U15734 ( .A1(n13758), .A2(n13913), .ZN(n13716) );
  AOI21_X1 U15735 ( .B1(n13756), .B2(n13717), .A(n13716), .ZN(n14173) );
  NAND2_X1 U15736 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n13858)
         );
  OAI21_X1 U15737 ( .B1(n13739), .B2(n14173), .A(n13858), .ZN(n13718) );
  AOI211_X1 U15738 ( .C1(n14083), .C2(n6468), .A(n13719), .B(n13718), .ZN(
        n13720) );
  OAI21_X1 U15739 ( .B1(n13721), .B2(n13731), .A(n13720), .ZN(P1_U3238) );
  OAI21_X1 U15740 ( .B1(n13724), .B2(n13722), .A(n13723), .ZN(n13725) );
  INV_X1 U15741 ( .A(n13725), .ZN(n13732) );
  NAND2_X1 U15742 ( .A1(n13748), .A2(n13717), .ZN(n13727) );
  NAND2_X1 U15743 ( .A1(n13750), .A2(n13913), .ZN(n13726) );
  NAND2_X1 U15744 ( .A1(n13727), .A2(n13726), .ZN(n14116) );
  AOI22_X1 U15745 ( .A1(n14411), .A2(n14116), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13728) );
  OAI21_X1 U15746 ( .B1(n13950), .B2(n14417), .A(n13728), .ZN(n13729) );
  AOI21_X1 U15747 ( .B1(n14117), .B2(n6468), .A(n13729), .ZN(n13730) );
  OAI21_X1 U15748 ( .B1(n13732), .B2(n13731), .A(n13730), .ZN(P1_U3240) );
  OAI21_X1 U15749 ( .B1(n13735), .B2(n13734), .A(n13733), .ZN(n13736) );
  NAND2_X1 U15750 ( .A1(n13736), .A2(n14409), .ZN(n13744) );
  NAND2_X1 U15751 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14471)
         );
  OAI21_X1 U15752 ( .B1(n13739), .B2(n13738), .A(n14471), .ZN(n13740) );
  AOI21_X1 U15753 ( .B1(n13742), .B2(n13741), .A(n13740), .ZN(n13743) );
  OAI211_X1 U15754 ( .C1(n13746), .C2(n13745), .A(n13744), .B(n13743), .ZN(
        P1_U3241) );
  MUX2_X1 U15755 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n13890), .S(n13775), .Z(
        P1_U3591) );
  MUX2_X1 U15756 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13910), .S(n13775), .Z(
        P1_U3590) );
  MUX2_X1 U15757 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13747), .S(n13775), .Z(
        P1_U3589) );
  MUX2_X1 U15758 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n13914), .S(n13775), .Z(
        P1_U3588) );
  MUX2_X1 U15759 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n13748), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15760 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n13749), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15761 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n13750), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15762 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n13751), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15763 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n13752), .S(n13775), .Z(
        P1_U3583) );
  MUX2_X1 U15764 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n13753), .S(n13775), .Z(
        P1_U3582) );
  MUX2_X1 U15765 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n13754), .S(n13775), .Z(
        P1_U3581) );
  MUX2_X1 U15766 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13755), .S(n13775), .Z(
        P1_U3580) );
  MUX2_X1 U15767 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n13756), .S(n13775), .Z(
        P1_U3579) );
  MUX2_X1 U15768 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n13757), .S(n13775), .Z(
        P1_U3578) );
  MUX2_X1 U15769 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n13758), .S(n13775), .Z(
        P1_U3577) );
  MUX2_X1 U15770 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n13759), .S(n13775), .Z(
        P1_U3576) );
  MUX2_X1 U15771 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n13760), .S(n13775), .Z(
        P1_U3575) );
  MUX2_X1 U15772 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13761), .S(n13775), .Z(
        P1_U3574) );
  MUX2_X1 U15773 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n13762), .S(n13775), .Z(
        P1_U3573) );
  MUX2_X1 U15774 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n13763), .S(n13775), .Z(
        P1_U3572) );
  MUX2_X1 U15775 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13764), .S(n13775), .Z(
        P1_U3571) );
  MUX2_X1 U15776 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n13765), .S(n13775), .Z(
        P1_U3570) );
  MUX2_X1 U15777 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n13766), .S(n13775), .Z(
        P1_U3569) );
  MUX2_X1 U15778 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13767), .S(n13775), .Z(
        P1_U3568) );
  MUX2_X1 U15779 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n13768), .S(n13775), .Z(
        P1_U3567) );
  MUX2_X1 U15780 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13769), .S(n13775), .Z(
        P1_U3566) );
  MUX2_X1 U15781 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13770), .S(n13775), .Z(
        P1_U3565) );
  MUX2_X1 U15782 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13771), .S(n13775), .Z(
        P1_U3564) );
  MUX2_X1 U15783 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n13772), .S(n13775), .Z(
        P1_U3563) );
  MUX2_X1 U15784 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n13773), .S(n13775), .Z(
        P1_U3562) );
  MUX2_X1 U15785 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n13774), .S(n13775), .Z(
        P1_U3561) );
  MUX2_X1 U15786 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n13776), .S(n13775), .Z(
        P1_U3560) );
  OAI22_X1 U15787 ( .A1(n14473), .A2(n9677), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13777), .ZN(n13778) );
  AOI21_X1 U15788 ( .B1(n13779), .B2(n14465), .A(n13778), .ZN(n13788) );
  AND2_X1 U15789 ( .A1(n14256), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n13781) );
  OAI211_X1 U15790 ( .C1(n13782), .C2(n13781), .A(n14462), .B(n13780), .ZN(
        n13787) );
  INV_X1 U15791 ( .A(n13783), .ZN(n13785) );
  OAI211_X1 U15792 ( .C1(n13785), .C2(n13784), .A(n13883), .B(n13795), .ZN(
        n13786) );
  NAND3_X1 U15793 ( .A1(n13788), .A2(n13787), .A3(n13786), .ZN(P1_U3244) );
  INV_X1 U15794 ( .A(n13789), .ZN(n13792) );
  OAI22_X1 U15795 ( .A1(n14473), .A2(n9678), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13790), .ZN(n13791) );
  AOI21_X1 U15796 ( .B1(n13792), .B2(n14465), .A(n13791), .ZN(n13803) );
  INV_X1 U15797 ( .A(n13793), .ZN(n13816) );
  NAND3_X1 U15798 ( .A1(n13796), .A2(n13795), .A3(n13794), .ZN(n13797) );
  NAND3_X1 U15799 ( .A1(n13883), .A2(n13816), .A3(n13797), .ZN(n13802) );
  OAI211_X1 U15800 ( .C1(n13800), .C2(n13799), .A(n14462), .B(n13798), .ZN(
        n13801) );
  NAND4_X1 U15801 ( .A1(n13804), .A2(n13803), .A3(n13802), .A4(n13801), .ZN(
        P1_U3245) );
  NOR2_X1 U15802 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n13805), .ZN(n13808) );
  NOR2_X1 U15803 ( .A1(n13806), .A2(n13812), .ZN(n13807) );
  AOI211_X1 U15804 ( .C1(n13827), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n13808), .B(
        n13807), .ZN(n13821) );
  OAI211_X1 U15805 ( .C1(n13810), .C2(n13809), .A(n14462), .B(n6765), .ZN(
        n13820) );
  INV_X1 U15806 ( .A(n13811), .ZN(n13815) );
  MUX2_X1 U15807 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n13813), .S(n13812), .Z(
        n13814) );
  NAND3_X1 U15808 ( .A1(n13816), .A2(n13815), .A3(n13814), .ZN(n13817) );
  NAND3_X1 U15809 ( .A1(n13883), .A2(n13818), .A3(n13817), .ZN(n13819) );
  NAND3_X1 U15810 ( .A1(n13821), .A2(n13820), .A3(n13819), .ZN(P1_U3246) );
  OAI21_X1 U15811 ( .B1(n13824), .B2(n13823), .A(n13822), .ZN(n13825) );
  NAND2_X1 U15812 ( .A1(n13825), .A2(n14462), .ZN(n13838) );
  AOI21_X1 U15813 ( .B1(n13827), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n13826), .ZN(
        n13837) );
  MUX2_X1 U15814 ( .A(n11055), .B(P1_REG2_REG_9__SCAN_IN), .S(n13834), .Z(
        n13830) );
  INV_X1 U15815 ( .A(n13828), .ZN(n13829) );
  NAND2_X1 U15816 ( .A1(n13830), .A2(n13829), .ZN(n13832) );
  OAI211_X1 U15817 ( .C1(n13833), .C2(n13832), .A(n13831), .B(n13883), .ZN(
        n13836) );
  NAND2_X1 U15818 ( .A1(n14465), .A2(n13834), .ZN(n13835) );
  NAND4_X1 U15819 ( .A1(n13838), .A2(n13837), .A3(n13836), .A4(n13835), .ZN(
        P1_U3252) );
  NAND2_X1 U15820 ( .A1(n13847), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n13840) );
  NAND2_X1 U15821 ( .A1(n13840), .A2(n13839), .ZN(n13843) );
  INV_X1 U15822 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n13863) );
  NOR2_X1 U15823 ( .A1(n13862), .A2(n13863), .ZN(n13841) );
  AOI21_X1 U15824 ( .B1(n13863), .B2(n13862), .A(n13841), .ZN(n13842) );
  NAND2_X1 U15825 ( .A1(n13842), .A2(n13843), .ZN(n13861) );
  OAI211_X1 U15826 ( .C1(n13843), .C2(n13842), .A(n13883), .B(n13861), .ZN(
        n13853) );
  INV_X1 U15827 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n13845) );
  OAI21_X1 U15828 ( .B1(n14473), .B2(n13845), .A(n13844), .ZN(n13851) );
  AOI21_X1 U15829 ( .B1(n13847), .B2(P1_REG1_REG_16__SCAN_IN), .A(n13846), 
        .ZN(n13849) );
  XNOR2_X1 U15830 ( .A(n13855), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n13848) );
  NOR2_X1 U15831 ( .A1(n13849), .A2(n13848), .ZN(n13854) );
  AOI211_X1 U15832 ( .C1(n13849), .C2(n13848), .A(n13854), .B(n13880), .ZN(
        n13850) );
  AOI211_X1 U15833 ( .C1(n14465), .C2(n13855), .A(n13851), .B(n13850), .ZN(
        n13852) );
  NAND2_X1 U15834 ( .A1(n13853), .A2(n13852), .ZN(P1_U3260) );
  AOI21_X1 U15835 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n13855), .A(n13854), 
        .ZN(n13869) );
  XNOR2_X1 U15836 ( .A(n13868), .B(n13869), .ZN(n13856) );
  NOR2_X1 U15837 ( .A1(n14177), .A2(n13856), .ZN(n13871) );
  AOI211_X1 U15838 ( .C1(n13856), .C2(n14177), .A(n13871), .B(n13880), .ZN(
        n13857) );
  INV_X1 U15839 ( .A(n13857), .ZN(n13867) );
  INV_X1 U15840 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n13859) );
  OAI21_X1 U15841 ( .B1(n14473), .B2(n13859), .A(n13858), .ZN(n13860) );
  AOI21_X1 U15842 ( .B1(n13875), .B2(n14465), .A(n13860), .ZN(n13866) );
  OAI21_X1 U15843 ( .B1(n13863), .B2(n13862), .A(n13861), .ZN(n13874) );
  XNOR2_X1 U15844 ( .A(n13868), .B(n13874), .ZN(n13864) );
  NAND2_X1 U15845 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n13864), .ZN(n13877) );
  OAI211_X1 U15846 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n13864), .A(n13883), 
        .B(n13877), .ZN(n13865) );
  NAND3_X1 U15847 ( .A1(n13867), .A2(n13866), .A3(n13865), .ZN(P1_U3261) );
  NOR2_X1 U15848 ( .A1(n13869), .A2(n13868), .ZN(n13870) );
  NOR2_X1 U15849 ( .A1(n13871), .A2(n13870), .ZN(n13873) );
  INV_X1 U15850 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n13872) );
  XOR2_X1 U15851 ( .A(n13873), .B(n13872), .Z(n13881) );
  NAND2_X1 U15852 ( .A1(n13875), .A2(n13874), .ZN(n13876) );
  NAND2_X1 U15853 ( .A1(n13877), .A2(n13876), .ZN(n13878) );
  XOR2_X1 U15854 ( .A(n13878), .B(P1_REG2_REG_19__SCAN_IN), .Z(n13879) );
  AOI22_X1 U15855 ( .A1(n13881), .A2(n14462), .B1(n13883), .B2(n13879), .ZN(
        n13884) );
  INV_X1 U15856 ( .A(n13879), .ZN(n13882) );
  NOR2_X1 U15857 ( .A1(n13887), .A2(n14119), .ZN(n14095) );
  NAND2_X1 U15858 ( .A1(n14095), .A2(n14485), .ZN(n13892) );
  NAND2_X1 U15859 ( .A1(n13888), .A2(P1_B_REG_SCAN_IN), .ZN(n13889) );
  AND2_X1 U15860 ( .A1(n13717), .A2(n13889), .ZN(n13909) );
  AND2_X1 U15861 ( .A1(n13890), .A2(n13909), .ZN(n14094) );
  INV_X1 U15862 ( .A(n14094), .ZN(n14098) );
  NOR2_X1 U15863 ( .A1(n14479), .A2(n14098), .ZN(n13896) );
  AOI21_X1 U15864 ( .B1(n14479), .B2(P1_REG2_REG_31__SCAN_IN), .A(n13896), 
        .ZN(n13891) );
  OAI211_X1 U15865 ( .C1(n6815), .C2(n14482), .A(n13892), .B(n13891), .ZN(
        P1_U3263) );
  NAND2_X1 U15866 ( .A1(n14198), .A2(n13907), .ZN(n13893) );
  NAND2_X1 U15867 ( .A1(n13893), .A2(n14493), .ZN(n13894) );
  OR2_X1 U15868 ( .A1(n13895), .A2(n13894), .ZN(n14099) );
  AOI21_X1 U15869 ( .B1(n14479), .B2(P1_REG2_REG_30__SCAN_IN), .A(n13896), 
        .ZN(n13898) );
  NAND2_X1 U15870 ( .A1(n14198), .A2(n14082), .ZN(n13897) );
  OAI211_X1 U15871 ( .C1(n14099), .C2(n14085), .A(n13898), .B(n13897), .ZN(
        P1_U3264) );
  NAND2_X1 U15872 ( .A1(n13900), .A2(n13899), .ZN(n13901) );
  XNOR2_X1 U15873 ( .A(n13901), .B(n13906), .ZN(n14111) );
  NOR2_X1 U15874 ( .A1(n9156), .A2(n13914), .ZN(n13903) );
  INV_X1 U15875 ( .A(n13914), .ZN(n13902) );
  OAI22_X1 U15876 ( .A1(n13904), .A2(n13903), .B1(n13902), .B2(n13926), .ZN(
        n13905) );
  XNOR2_X1 U15877 ( .A(n13906), .B(n13905), .ZN(n14109) );
  OAI21_X1 U15878 ( .B1(n14106), .B2(n13908), .A(n13907), .ZN(n14103) );
  NOR2_X1 U15879 ( .A1(n14103), .A2(n13956), .ZN(n13919) );
  NAND2_X1 U15880 ( .A1(n13910), .A2(n13909), .ZN(n14104) );
  OAI22_X1 U15881 ( .A1(n13912), .A2(n14104), .B1(n13911), .B2(n14477), .ZN(
        n13916) );
  NAND2_X1 U15882 ( .A1(n13914), .A2(n13913), .ZN(n14105) );
  NOR2_X1 U15883 ( .A1(n14491), .A2(n14105), .ZN(n13915) );
  AOI211_X1 U15884 ( .C1(n14491), .C2(P1_REG2_REG_29__SCAN_IN), .A(n13916), 
        .B(n13915), .ZN(n13917) );
  OAI21_X1 U15885 ( .B1(n14106), .B2(n14482), .A(n13917), .ZN(n13918) );
  AOI211_X1 U15886 ( .C1(n14109), .C2(n14071), .A(n13919), .B(n13918), .ZN(
        n13920) );
  OAI21_X1 U15887 ( .B1(n14111), .B2(n14073), .A(n13920), .ZN(P1_U3356) );
  INV_X1 U15888 ( .A(n13922), .ZN(n13930) );
  NAND2_X1 U15889 ( .A1(n14491), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n13923) );
  OAI21_X1 U15890 ( .B1(n14477), .B2(n13924), .A(n13923), .ZN(n13925) );
  AOI21_X1 U15891 ( .B1(n13926), .B2(n14082), .A(n13925), .ZN(n13927) );
  OAI21_X1 U15892 ( .B1(n13928), .B2(n14085), .A(n13927), .ZN(n13929) );
  AOI21_X1 U15893 ( .B1(n13930), .B2(n14092), .A(n13929), .ZN(n13931) );
  OAI21_X1 U15894 ( .B1(n13921), .B2(n14491), .A(n13931), .ZN(P1_U3265) );
  XNOR2_X1 U15895 ( .A(n13933), .B(n13932), .ZN(n13935) );
  AOI21_X1 U15896 ( .B1(n13935), .B2(n14526), .A(n13934), .ZN(n14115) );
  NAND2_X1 U15897 ( .A1(n13949), .A2(n14203), .ZN(n13937) );
  NAND3_X1 U15898 ( .A1(n13938), .A2(n14493), .A3(n13937), .ZN(n14113) );
  INV_X1 U15899 ( .A(n13939), .ZN(n13940) );
  AOI22_X1 U15900 ( .A1(n14479), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n13940), 
        .B2(n14034), .ZN(n13942) );
  NAND2_X1 U15901 ( .A1(n14203), .A2(n14082), .ZN(n13941) );
  OAI211_X1 U15902 ( .C1(n14113), .C2(n14085), .A(n13942), .B(n13941), .ZN(
        n13943) );
  AOI21_X1 U15903 ( .B1(n14112), .B2(n14092), .A(n13943), .ZN(n13944) );
  OAI21_X1 U15904 ( .B1(n14115), .B2(n14491), .A(n13944), .ZN(P1_U3266) );
  XNOR2_X1 U15905 ( .A(n13946), .B(n13945), .ZN(n14124) );
  XNOR2_X1 U15906 ( .A(n13948), .B(n13947), .ZN(n14122) );
  OAI21_X1 U15907 ( .B1(n13952), .B2(n13967), .A(n13949), .ZN(n14120) );
  INV_X1 U15908 ( .A(n14116), .ZN(n13951) );
  OAI22_X1 U15909 ( .A1(n14479), .A2(n13951), .B1(n13950), .B2(n14477), .ZN(
        n13954) );
  NOR2_X1 U15910 ( .A1(n13952), .A2(n14482), .ZN(n13953) );
  AOI211_X1 U15911 ( .C1(n14491), .C2(P1_REG2_REG_26__SCAN_IN), .A(n13954), 
        .B(n13953), .ZN(n13955) );
  OAI21_X1 U15912 ( .B1(n13956), .B2(n14120), .A(n13955), .ZN(n13957) );
  AOI21_X1 U15913 ( .B1(n14071), .B2(n14122), .A(n13957), .ZN(n13958) );
  OAI21_X1 U15914 ( .B1(n14073), .B2(n14124), .A(n13958), .ZN(P1_U3267) );
  INV_X1 U15915 ( .A(n13959), .ZN(n13961) );
  XNOR2_X1 U15916 ( .A(n13961), .B(n13960), .ZN(n14130) );
  OAI21_X1 U15917 ( .B1(n13964), .B2(n13963), .A(n13962), .ZN(n14125) );
  INV_X1 U15918 ( .A(n14125), .ZN(n13976) );
  NAND2_X1 U15919 ( .A1(n14208), .A2(n13985), .ZN(n13965) );
  NAND2_X1 U15920 ( .A1(n13965), .A2(n14493), .ZN(n13966) );
  OR2_X1 U15921 ( .A1(n13967), .A2(n13966), .ZN(n14127) );
  INV_X1 U15922 ( .A(n13968), .ZN(n14126) );
  NAND2_X1 U15923 ( .A1(n14491), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n13972) );
  INV_X1 U15924 ( .A(n13969), .ZN(n13970) );
  NAND2_X1 U15925 ( .A1(n14034), .A2(n13970), .ZN(n13971) );
  OAI211_X1 U15926 ( .C1(n14491), .C2(n14126), .A(n13972), .B(n13971), .ZN(
        n13973) );
  AOI21_X1 U15927 ( .B1(n14208), .B2(n14082), .A(n13973), .ZN(n13974) );
  OAI21_X1 U15928 ( .B1(n14127), .B2(n14085), .A(n13974), .ZN(n13975) );
  AOI21_X1 U15929 ( .B1(n13976), .B2(n14092), .A(n13975), .ZN(n13977) );
  OAI21_X1 U15930 ( .B1(n14130), .B2(n14042), .A(n13977), .ZN(P1_U3268) );
  XNOR2_X1 U15931 ( .A(n13979), .B(n13978), .ZN(n13981) );
  AOI21_X1 U15932 ( .B1(n13981), .B2(n14526), .A(n13980), .ZN(n14136) );
  NAND2_X1 U15933 ( .A1(n13982), .A2(n7070), .ZN(n13983) );
  NAND2_X1 U15934 ( .A1(n13984), .A2(n13983), .ZN(n14133) );
  AOI21_X1 U15935 ( .B1(n14212), .B2(n13999), .A(n14119), .ZN(n13986) );
  NAND2_X1 U15936 ( .A1(n13986), .A2(n13985), .ZN(n14134) );
  INV_X1 U15937 ( .A(n13987), .ZN(n13988) );
  AOI22_X1 U15938 ( .A1(n14491), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n13988), 
        .B2(n14034), .ZN(n13990) );
  NAND2_X1 U15939 ( .A1(n14212), .A2(n14082), .ZN(n13989) );
  OAI211_X1 U15940 ( .C1(n14134), .C2(n14085), .A(n13990), .B(n13989), .ZN(
        n13991) );
  AOI21_X1 U15941 ( .B1(n14133), .B2(n14092), .A(n13991), .ZN(n13992) );
  OAI21_X1 U15942 ( .B1(n14136), .B2(n14479), .A(n13992), .ZN(P1_U3269) );
  XOR2_X1 U15943 ( .A(n13993), .B(n13997), .Z(n14145) );
  INV_X1 U15944 ( .A(n13994), .ZN(n13995) );
  AOI21_X1 U15945 ( .B1(n13997), .B2(n13996), .A(n13995), .ZN(n14139) );
  NAND2_X1 U15946 ( .A1(n14139), .A2(n14092), .ZN(n14007) );
  AOI21_X1 U15947 ( .B1(n14142), .B2(n14015), .A(n14119), .ZN(n13998) );
  AND2_X1 U15948 ( .A1(n13999), .A2(n13998), .ZN(n14140) );
  NOR2_X1 U15949 ( .A1(n14477), .A2(n14000), .ZN(n14001) );
  NOR2_X1 U15950 ( .A1(n14141), .A2(n14001), .ZN(n14004) );
  NAND2_X1 U15951 ( .A1(n14142), .A2(n14082), .ZN(n14003) );
  NAND2_X1 U15952 ( .A1(n14479), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n14002) );
  OAI211_X1 U15953 ( .C1(n14491), .C2(n14004), .A(n14003), .B(n14002), .ZN(
        n14005) );
  AOI21_X1 U15954 ( .B1(n14140), .B2(n14485), .A(n14005), .ZN(n14006) );
  OAI211_X1 U15955 ( .C1(n14145), .C2(n14042), .A(n14007), .B(n14006), .ZN(
        P1_U3270) );
  OR2_X1 U15956 ( .A1(n14008), .A2(n14018), .ZN(n14009) );
  NAND2_X1 U15957 ( .A1(n14010), .A2(n14009), .ZN(n14146) );
  INV_X1 U15958 ( .A(n14146), .ZN(n14027) );
  INV_X1 U15959 ( .A(n14218), .ZN(n14014) );
  OAI22_X1 U15960 ( .A1(n14080), .A2(n14012), .B1(n14011), .B2(n14477), .ZN(
        n14013) );
  AOI21_X1 U15961 ( .B1(n14014), .B2(n14082), .A(n14013), .ZN(n14026) );
  OAI211_X1 U15962 ( .C1(n14032), .C2(n14218), .A(n14015), .B(n14493), .ZN(
        n14017) );
  AND2_X1 U15963 ( .A1(n14017), .A2(n14016), .ZN(n14148) );
  NAND2_X1 U15964 ( .A1(n14019), .A2(n14018), .ZN(n14020) );
  NAND2_X1 U15965 ( .A1(n14021), .A2(n14020), .ZN(n14022) );
  NAND2_X1 U15966 ( .A1(n14022), .A2(n14526), .ZN(n14147) );
  OAI21_X1 U15967 ( .B1(n14023), .B2(n14148), .A(n14147), .ZN(n14024) );
  NAND2_X1 U15968 ( .A1(n14024), .A2(n14080), .ZN(n14025) );
  OAI211_X1 U15969 ( .C1(n14027), .C2(n14073), .A(n14026), .B(n14025), .ZN(
        P1_U3271) );
  OAI21_X1 U15970 ( .B1(n14029), .B2(n14030), .A(n14028), .ZN(n14158) );
  XNOR2_X1 U15971 ( .A(n14031), .B(n14030), .ZN(n14152) );
  NAND2_X1 U15972 ( .A1(n14152), .A2(n14092), .ZN(n14041) );
  AOI211_X1 U15973 ( .C1(n14155), .C2(n6513), .A(n14119), .B(n14032), .ZN(
        n14153) );
  INV_X1 U15974 ( .A(n14033), .ZN(n14154) );
  AOI22_X1 U15975 ( .A1(n14080), .A2(n14154), .B1(n14035), .B2(n14034), .ZN(
        n14037) );
  NAND2_X1 U15976 ( .A1(n14479), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n14036) );
  OAI211_X1 U15977 ( .C1(n14038), .C2(n14482), .A(n14037), .B(n14036), .ZN(
        n14039) );
  AOI21_X1 U15978 ( .B1(n14153), .B2(n14485), .A(n14039), .ZN(n14040) );
  OAI211_X1 U15979 ( .C1(n14158), .C2(n14042), .A(n14041), .B(n14040), .ZN(
        P1_U3272) );
  NAND2_X1 U15980 ( .A1(n14044), .A2(n14043), .ZN(n14045) );
  NAND3_X1 U15981 ( .A1(n14046), .A2(n14526), .A3(n14045), .ZN(n14048) );
  NAND2_X1 U15982 ( .A1(n14050), .A2(n14049), .ZN(n14051) );
  NAND2_X1 U15983 ( .A1(n14052), .A2(n14051), .ZN(n14161) );
  INV_X1 U15984 ( .A(n14161), .ZN(n14059) );
  AOI21_X1 U15985 ( .B1(n14222), .B2(n14065), .A(n14119), .ZN(n14053) );
  NAND2_X1 U15986 ( .A1(n14053), .A2(n6513), .ZN(n14159) );
  NAND2_X1 U15987 ( .A1(n14491), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n14054) );
  OAI21_X1 U15988 ( .B1(n14477), .B2(n14055), .A(n14054), .ZN(n14056) );
  AOI21_X1 U15989 ( .B1(n14222), .B2(n14082), .A(n14056), .ZN(n14057) );
  OAI21_X1 U15990 ( .B1(n14159), .B2(n14085), .A(n14057), .ZN(n14058) );
  AOI21_X1 U15991 ( .B1(n14059), .B2(n14092), .A(n14058), .ZN(n14060) );
  OAI21_X1 U15992 ( .B1(n14491), .B2(n14160), .A(n14060), .ZN(P1_U3273) );
  XNOR2_X1 U15993 ( .A(n14062), .B(n14061), .ZN(n14171) );
  OAI21_X1 U15994 ( .B1(n7396), .B2(n14064), .A(n14063), .ZN(n14169) );
  OAI211_X1 U15995 ( .C1(n14167), .C2(n14075), .A(n14493), .B(n14065), .ZN(
        n14166) );
  OAI22_X1 U15996 ( .A1(n14479), .A2(n14165), .B1(n14066), .B2(n14477), .ZN(
        n14068) );
  NOR2_X1 U15997 ( .A1(n14167), .A2(n14482), .ZN(n14067) );
  AOI211_X1 U15998 ( .C1(n14491), .C2(P1_REG2_REG_19__SCAN_IN), .A(n14068), 
        .B(n14067), .ZN(n14069) );
  OAI21_X1 U15999 ( .B1(n14085), .B2(n14166), .A(n14069), .ZN(n14070) );
  AOI21_X1 U16000 ( .B1(n14169), .B2(n14071), .A(n14070), .ZN(n14072) );
  OAI21_X1 U16001 ( .B1(n14171), .B2(n14073), .A(n14072), .ZN(P1_U3274) );
  XNOR2_X1 U16002 ( .A(n14074), .B(n14088), .ZN(n14176) );
  INV_X1 U16003 ( .A(n14075), .ZN(n14076) );
  OAI211_X1 U16004 ( .C1(n14228), .C2(n14077), .A(n14076), .B(n14493), .ZN(
        n14172) );
  INV_X1 U16005 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14079) );
  OAI22_X1 U16006 ( .A1(n14080), .A2(n14079), .B1(n14078), .B2(n14477), .ZN(
        n14081) );
  AOI21_X1 U16007 ( .B1(n14083), .B2(n14082), .A(n14081), .ZN(n14084) );
  OAI21_X1 U16008 ( .B1(n14172), .B2(n14085), .A(n14084), .ZN(n14091) );
  INV_X1 U16009 ( .A(n14086), .ZN(n14089) );
  OAI211_X1 U16010 ( .C1(n14089), .C2(n14088), .A(n14087), .B(n14526), .ZN(
        n14174) );
  AOI21_X1 U16011 ( .B1(n14174), .B2(n14173), .A(n14479), .ZN(n14090) );
  AOI211_X1 U16012 ( .C1(n14176), .C2(n14092), .A(n14091), .B(n14090), .ZN(
        n14093) );
  INV_X1 U16013 ( .A(n14093), .ZN(P1_U3275) );
  NOR2_X1 U16014 ( .A1(n14095), .A2(n14094), .ZN(n14193) );
  OAI21_X1 U16015 ( .B1(n6815), .B2(n14186), .A(n14097), .ZN(P1_U3559) );
  NAND2_X1 U16016 ( .A1(n14099), .A2(n14098), .ZN(n14196) );
  MUX2_X1 U16017 ( .A(n14196), .B(P1_REG1_REG_30__SCAN_IN), .S(n14558), .Z(
        n14100) );
  INV_X1 U16018 ( .A(n14100), .ZN(n14102) );
  NAND2_X1 U16019 ( .A1(n14198), .A2(n14163), .ZN(n14101) );
  NAND2_X1 U16020 ( .A1(n14102), .A2(n14101), .ZN(P1_U3558) );
  NOR2_X1 U16021 ( .A1(n14103), .A2(n14119), .ZN(n14108) );
  OAI211_X1 U16022 ( .C1(n14106), .C2(n14528), .A(n14105), .B(n14104), .ZN(
        n14107) );
  OAI21_X1 U16023 ( .B1(n14521), .B2(n14111), .A(n14110), .ZN(n14201) );
  MUX2_X1 U16024 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14201), .S(n14560), .Z(
        P1_U3557) );
  NAND2_X1 U16025 ( .A1(n14112), .A2(n14430), .ZN(n14114) );
  AOI21_X1 U16026 ( .B1(n14117), .B2(n14538), .A(n14116), .ZN(n14118) );
  OAI21_X1 U16027 ( .B1(n14120), .B2(n14119), .A(n14118), .ZN(n14121) );
  AOI21_X1 U16028 ( .B1(n14526), .B2(n14122), .A(n14121), .ZN(n14123) );
  OAI21_X1 U16029 ( .B1(n14124), .B2(n14521), .A(n14123), .ZN(n14205) );
  MUX2_X1 U16030 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14205), .S(n14560), .Z(
        P1_U3554) );
  OR2_X1 U16031 ( .A1(n14125), .A2(n14521), .ZN(n14129) );
  AND2_X1 U16032 ( .A1(n14127), .A2(n14126), .ZN(n14128) );
  OAI211_X1 U16033 ( .C1(n14534), .C2(n14130), .A(n14129), .B(n14128), .ZN(
        n14206) );
  MUX2_X1 U16034 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14206), .S(n14560), .Z(
        n14131) );
  AOI21_X1 U16035 ( .B1(n14163), .B2(n14208), .A(n14131), .ZN(n14132) );
  INV_X1 U16036 ( .A(n14132), .ZN(P1_U3553) );
  NAND2_X1 U16037 ( .A1(n14133), .A2(n14430), .ZN(n14135) );
  NAND3_X1 U16038 ( .A1(n14136), .A2(n14135), .A3(n14134), .ZN(n14210) );
  MUX2_X1 U16039 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14210), .S(n14560), .Z(
        n14137) );
  AOI21_X1 U16040 ( .B1(n14163), .B2(n14212), .A(n14137), .ZN(n14138) );
  INV_X1 U16041 ( .A(n14138), .ZN(P1_U3552) );
  NAND2_X1 U16042 ( .A1(n14139), .A2(n14430), .ZN(n14144) );
  AOI211_X1 U16043 ( .C1(n14538), .C2(n14142), .A(n14141), .B(n14140), .ZN(
        n14143) );
  OAI211_X1 U16044 ( .C1(n14534), .C2(n14145), .A(n14144), .B(n14143), .ZN(
        n14214) );
  MUX2_X1 U16045 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14214), .S(n14560), .Z(
        P1_U3551) );
  NAND2_X1 U16046 ( .A1(n14146), .A2(n14430), .ZN(n14149) );
  NAND3_X1 U16047 ( .A1(n14149), .A2(n14148), .A3(n14147), .ZN(n14215) );
  MUX2_X1 U16048 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14215), .S(n14560), .Z(
        n14150) );
  INV_X1 U16049 ( .A(n14150), .ZN(n14151) );
  OAI21_X1 U16050 ( .B1(n14186), .B2(n14218), .A(n14151), .ZN(P1_U3550) );
  NAND2_X1 U16051 ( .A1(n14152), .A2(n14430), .ZN(n14157) );
  AOI211_X1 U16052 ( .C1(n14538), .C2(n14155), .A(n14154), .B(n14153), .ZN(
        n14156) );
  OAI211_X1 U16053 ( .C1(n14534), .C2(n14158), .A(n14157), .B(n14156), .ZN(
        n14219) );
  MUX2_X1 U16054 ( .A(n14219), .B(P1_REG1_REG_21__SCAN_IN), .S(n14558), .Z(
        P1_U3549) );
  OAI211_X1 U16055 ( .C1(n14161), .C2(n14521), .A(n14160), .B(n14159), .ZN(
        n14220) );
  MUX2_X1 U16056 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14220), .S(n14560), .Z(
        n14162) );
  AOI21_X1 U16057 ( .B1(n14163), .B2(n14222), .A(n14162), .ZN(n14164) );
  INV_X1 U16058 ( .A(n14164), .ZN(P1_U3548) );
  OAI211_X1 U16059 ( .C1(n14167), .C2(n14528), .A(n14166), .B(n14165), .ZN(
        n14168) );
  AOI21_X1 U16060 ( .B1(n14169), .B2(n14526), .A(n14168), .ZN(n14170) );
  OAI21_X1 U16061 ( .B1(n14171), .B2(n14521), .A(n14170), .ZN(n14224) );
  MUX2_X1 U16062 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14224), .S(n14560), .Z(
        P1_U3547) );
  NAND3_X1 U16063 ( .A1(n14174), .A2(n14173), .A3(n14172), .ZN(n14175) );
  AOI21_X1 U16064 ( .B1(n14176), .B2(n14430), .A(n14175), .ZN(n14225) );
  MUX2_X1 U16065 ( .A(n14177), .B(n14225), .S(n14560), .Z(n14178) );
  OAI21_X1 U16066 ( .B1(n14228), .B2(n14186), .A(n14178), .ZN(P1_U3546) );
  INV_X1 U16067 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n14184) );
  OAI211_X1 U16068 ( .C1(n14181), .C2(n14534), .A(n14180), .B(n14179), .ZN(
        n14182) );
  AOI21_X1 U16069 ( .B1(n14183), .B2(n14430), .A(n14182), .ZN(n14229) );
  MUX2_X1 U16070 ( .A(n14184), .B(n14229), .S(n14560), .Z(n14185) );
  OAI21_X1 U16071 ( .B1(n14233), .B2(n14186), .A(n14185), .ZN(P1_U3545) );
  INV_X1 U16072 ( .A(n14187), .ZN(n14192) );
  AOI21_X1 U16073 ( .B1(n14538), .B2(n14189), .A(n14188), .ZN(n14190) );
  OAI211_X1 U16074 ( .C1(n14192), .C2(n14521), .A(n14191), .B(n14190), .ZN(
        n14234) );
  MUX2_X1 U16075 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14234), .S(n14560), .Z(
        P1_U3544) );
  INV_X1 U16076 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n14194) );
  OAI21_X1 U16077 ( .B1(n6815), .B2(n14232), .A(n14195), .ZN(P1_U3527) );
  MUX2_X1 U16078 ( .A(n14196), .B(P1_REG0_REG_30__SCAN_IN), .S(n14547), .Z(
        n14197) );
  INV_X1 U16079 ( .A(n14197), .ZN(n14200) );
  NAND2_X1 U16080 ( .A1(n14198), .A2(n9158), .ZN(n14199) );
  NAND2_X1 U16081 ( .A1(n14200), .A2(n14199), .ZN(P1_U3526) );
  MUX2_X1 U16082 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14201), .S(n14549), .Z(
        P1_U3525) );
  INV_X1 U16083 ( .A(n14204), .ZN(P1_U3523) );
  MUX2_X1 U16084 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14205), .S(n14549), .Z(
        P1_U3522) );
  MUX2_X1 U16085 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14206), .S(n14549), .Z(
        n14207) );
  AOI21_X1 U16086 ( .B1(n9158), .B2(n14208), .A(n14207), .ZN(n14209) );
  INV_X1 U16087 ( .A(n14209), .ZN(P1_U3521) );
  MUX2_X1 U16088 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14210), .S(n14549), .Z(
        n14211) );
  AOI21_X1 U16089 ( .B1(n9158), .B2(n14212), .A(n14211), .ZN(n14213) );
  INV_X1 U16090 ( .A(n14213), .ZN(P1_U3520) );
  MUX2_X1 U16091 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14214), .S(n14549), .Z(
        P1_U3519) );
  MUX2_X1 U16092 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14215), .S(n14549), .Z(
        n14216) );
  INV_X1 U16093 ( .A(n14216), .ZN(n14217) );
  OAI21_X1 U16094 ( .B1(n14232), .B2(n14218), .A(n14217), .ZN(P1_U3518) );
  MUX2_X1 U16095 ( .A(n14219), .B(P1_REG0_REG_21__SCAN_IN), .S(n14547), .Z(
        P1_U3517) );
  MUX2_X1 U16096 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14220), .S(n14549), .Z(
        n14221) );
  AOI21_X1 U16097 ( .B1(n9158), .B2(n14222), .A(n14221), .ZN(n14223) );
  INV_X1 U16098 ( .A(n14223), .ZN(P1_U3516) );
  MUX2_X1 U16099 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14224), .S(n14549), .Z(
        P1_U3515) );
  INV_X1 U16100 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n14226) );
  MUX2_X1 U16101 ( .A(n14226), .B(n14225), .S(n14549), .Z(n14227) );
  OAI21_X1 U16102 ( .B1(n14228), .B2(n14232), .A(n14227), .ZN(P1_U3513) );
  INV_X1 U16103 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n14230) );
  MUX2_X1 U16104 ( .A(n14230), .B(n14229), .S(n14549), .Z(n14231) );
  OAI21_X1 U16105 ( .B1(n14233), .B2(n14232), .A(n14231), .ZN(P1_U3510) );
  MUX2_X1 U16106 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14234), .S(n14549), .Z(
        P1_U3507) );
  INV_X1 U16107 ( .A(n12219), .ZN(n14241) );
  INV_X1 U16108 ( .A(n14235), .ZN(n14237) );
  NOR4_X1 U16109 ( .A1(n14237), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), 
        .A4(n14236), .ZN(n14238) );
  AOI21_X1 U16110 ( .B1(n14239), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n14238), 
        .ZN(n14240) );
  OAI21_X1 U16111 ( .B1(n14241), .B2(n14251), .A(n14240), .ZN(P1_U3324) );
  OAI222_X1 U16112 ( .A1(P1_U3086), .A2(n14244), .B1(n14251), .B2(n14243), 
        .C1(n14242), .C2(n14245), .ZN(P1_U3326) );
  OAI222_X1 U16113 ( .A1(n14248), .A2(P1_U3086), .B1(n14251), .B2(n14247), 
        .C1(n14246), .C2(n14245), .ZN(P1_U3328) );
  OAI222_X1 U16114 ( .A1(n14252), .A2(P1_U3086), .B1(n14251), .B2(n14250), 
        .C1(n14249), .C2(n14245), .ZN(P1_U3329) );
  MUX2_X1 U16115 ( .A(n14254), .B(n14253), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  INV_X1 U16116 ( .A(n14255), .ZN(n14257) );
  MUX2_X1 U16117 ( .A(n14257), .B(n14256), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3355) );
  AOI21_X1 U16118 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14261) );
  OAI21_X1 U16119 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14261), 
        .ZN(U28) );
  OAI21_X1 U16120 ( .B1(n14264), .B2(n14263), .A(n14262), .ZN(n14265) );
  XNOR2_X1 U16121 ( .A(n14265), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  AOI22_X1 U16122 ( .A1(n14266), .A2(n14270), .B1(SI_7_), .B2(n14268), .ZN(
        n14267) );
  OAI21_X1 U16123 ( .B1(P3_U3151), .B2(n14930), .A(n14267), .ZN(P3_U3288) );
  AOI22_X1 U16124 ( .A1(n14270), .A2(n14269), .B1(SI_2_), .B2(n14268), .ZN(
        n14271) );
  OAI21_X1 U16125 ( .B1(P3_U3151), .B2(n6476), .A(n14271), .ZN(P3_U3293) );
  AOI21_X1 U16126 ( .B1(n14275), .B2(n14274), .A(n14273), .ZN(SUB_1596_U57) );
  OAI21_X1 U16127 ( .B1(n14278), .B2(n14277), .A(n14276), .ZN(SUB_1596_U55) );
  AOI21_X1 U16128 ( .B1(n14280), .B2(n14618), .A(n14279), .ZN(SUB_1596_U54) );
  AOI21_X1 U16129 ( .B1(n14283), .B2(n14282), .A(n14281), .ZN(n14284) );
  XOR2_X1 U16130 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n14284), .Z(SUB_1596_U70)
         );
  OAI21_X1 U16131 ( .B1(n14287), .B2(n14286), .A(n14285), .ZN(n14288) );
  XNOR2_X1 U16132 ( .A(n14288), .B(P2_ADDR_REG_17__SCAN_IN), .ZN(SUB_1596_U63)
         );
  AOI22_X1 U16133 ( .A1(n14996), .A2(n14289), .B1(n14969), .B2(
        P3_ADDR_REG_16__SCAN_IN), .ZN(n14306) );
  INV_X1 U16134 ( .A(n14290), .ZN(n14292) );
  NAND2_X1 U16135 ( .A1(n14292), .A2(n14291), .ZN(n14293) );
  XNOR2_X1 U16136 ( .A(n14294), .B(n14293), .ZN(n14299) );
  OAI21_X1 U16137 ( .B1(n14297), .B2(n14296), .A(n14295), .ZN(n14298) );
  AOI22_X1 U16138 ( .A1(n14299), .A2(n14962), .B1(n6467), .B2(n14298), .ZN(
        n14305) );
  NAND2_X1 U16139 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(P3_U3151), .ZN(n14304)
         );
  OAI221_X1 U16140 ( .B1(n14302), .B2(n6576), .C1(n14302), .C2(n14301), .A(
        n14300), .ZN(n14303) );
  NAND4_X1 U16141 ( .A1(n14306), .A2(n14305), .A3(n14304), .A4(n14303), .ZN(
        P3_U3198) );
  AOI21_X1 U16142 ( .B1(n14309), .B2(n14308), .A(n14307), .ZN(n14323) );
  OAI21_X1 U16143 ( .B1(n14311), .B2(P3_REG1_REG_17__SCAN_IN), .A(n14310), 
        .ZN(n14321) );
  NAND2_X1 U16144 ( .A1(n14996), .A2(n14312), .ZN(n14314) );
  OAI211_X1 U16145 ( .C1(n14315), .C2(n15000), .A(n14314), .B(n14313), .ZN(
        n14320) );
  AOI211_X1 U16146 ( .C1(n14318), .C2(n14317), .A(n14985), .B(n14316), .ZN(
        n14319) );
  AOI211_X1 U16147 ( .C1(n6467), .C2(n14321), .A(n14320), .B(n14319), .ZN(
        n14322) );
  OAI21_X1 U16148 ( .B1(n14323), .B2(n14991), .A(n14322), .ZN(P3_U3199) );
  XNOR2_X1 U16149 ( .A(n14324), .B(n14325), .ZN(n14351) );
  XNOR2_X1 U16150 ( .A(n14326), .B(n14325), .ZN(n14327) );
  OAI222_X1 U16151 ( .A1(n14339), .A2(n14329), .B1(n14341), .B2(n14328), .C1(
        n14327), .C2(n15045), .ZN(n14349) );
  AOI21_X1 U16152 ( .B1(n15019), .B2(n14351), .A(n14349), .ZN(n14333) );
  NOR2_X1 U16153 ( .A1(n14330), .A2(n15115), .ZN(n14350) );
  AOI22_X1 U16154 ( .A1(n14350), .A2(n15036), .B1(n15077), .B2(n14331), .ZN(
        n14332) );
  OAI221_X1 U16155 ( .B1(n15082), .B2(n14333), .C1(n15080), .C2(n7736), .A(
        n14332), .ZN(P3_U3219) );
  AND2_X1 U16156 ( .A1(n14334), .A2(n15071), .ZN(n14364) );
  AOI22_X1 U16157 ( .A1(n15036), .A2(n14364), .B1(n15077), .B2(n14335), .ZN(
        n14348) );
  XNOR2_X1 U16158 ( .A(n14336), .B(n14337), .ZN(n14365) );
  XNOR2_X1 U16159 ( .A(n14338), .B(n14337), .ZN(n14344) );
  OAI22_X1 U16160 ( .A1(n14342), .A2(n14341), .B1(n14340), .B2(n14339), .ZN(
        n14343) );
  AOI21_X1 U16161 ( .B1(n14344), .B2(n15060), .A(n14343), .ZN(n14367) );
  NOR2_X1 U16162 ( .A1(n14367), .A2(n15082), .ZN(n14345) );
  AOI21_X1 U16163 ( .B1(n14365), .B2(n14346), .A(n14345), .ZN(n14347) );
  OAI211_X1 U16164 ( .C1(n7512), .C2(n15080), .A(n14348), .B(n14347), .ZN(
        P3_U3222) );
  AOI211_X1 U16165 ( .C1(n15100), .C2(n14351), .A(n14350), .B(n14349), .ZN(
        n14369) );
  INV_X1 U16166 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n14352) );
  AOI22_X1 U16167 ( .A1(n15131), .A2(n14369), .B1(n14352), .B2(n9450), .ZN(
        P3_U3473) );
  OAI22_X1 U16168 ( .A1(n14355), .A2(n14354), .B1(n15115), .B2(n14353), .ZN(
        n14356) );
  NOR2_X1 U16169 ( .A1(n14357), .A2(n14356), .ZN(n14371) );
  INV_X1 U16170 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n14358) );
  AOI22_X1 U16171 ( .A1(n15131), .A2(n14371), .B1(n14358), .B2(n9450), .ZN(
        P3_U3472) );
  NOR2_X1 U16172 ( .A1(n14359), .A2(n15115), .ZN(n14361) );
  AOI211_X1 U16173 ( .C1(n15100), .C2(n14362), .A(n14361), .B(n14360), .ZN(
        n14373) );
  AOI22_X1 U16174 ( .A1(n15131), .A2(n14373), .B1(n14363), .B2(n9450), .ZN(
        P3_U3471) );
  AOI21_X1 U16175 ( .B1(n14365), .B2(n15100), .A(n14364), .ZN(n14366) );
  AND2_X1 U16176 ( .A1(n14367), .A2(n14366), .ZN(n14374) );
  INV_X1 U16177 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14368) );
  AOI22_X1 U16178 ( .A1(n15131), .A2(n14374), .B1(n14368), .B2(n9450), .ZN(
        P3_U3470) );
  INV_X1 U16179 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n14370) );
  AOI22_X1 U16180 ( .A1(n15121), .A2(n14370), .B1(n14369), .B2(n15120), .ZN(
        P3_U3432) );
  INV_X1 U16181 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14372) );
  AOI22_X1 U16182 ( .A1(n15121), .A2(n14372), .B1(n14371), .B2(n15120), .ZN(
        P3_U3429) );
  AOI22_X1 U16183 ( .A1(n15121), .A2(n7695), .B1(n14373), .B2(n15120), .ZN(
        P3_U3426) );
  INV_X1 U16184 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14375) );
  AOI22_X1 U16185 ( .A1(n15121), .A2(n14375), .B1(n14374), .B2(n15120), .ZN(
        P3_U3423) );
  OAI21_X1 U16186 ( .B1(n14377), .B2(n14822), .A(n14376), .ZN(n14379) );
  AOI211_X1 U16187 ( .C1(n14380), .C2(n14809), .A(n14379), .B(n14378), .ZN(
        n14390) );
  AOI22_X1 U16188 ( .A1(n14853), .A2(n14390), .B1(n14381), .B2(n14850), .ZN(
        P2_U3512) );
  AOI21_X1 U16189 ( .B1(n10449), .B2(n14769), .A(n14382), .ZN(n14387) );
  OAI211_X1 U16190 ( .C1(n14385), .C2(n14822), .A(n14384), .B(n14383), .ZN(
        n14386) );
  NOR2_X1 U16191 ( .A1(n14387), .A2(n14386), .ZN(n14392) );
  AOI22_X1 U16192 ( .A1(n14853), .A2(n14392), .B1(n14388), .B2(n14850), .ZN(
        P2_U3511) );
  INV_X1 U16193 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n14389) );
  AOI22_X1 U16194 ( .A1(n14831), .A2(n14390), .B1(n14389), .B2(n14829), .ZN(
        P2_U3469) );
  INV_X1 U16195 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14391) );
  AOI22_X1 U16196 ( .A1(n14831), .A2(n14392), .B1(n14391), .B2(n14829), .ZN(
        P2_U3466) );
  INV_X1 U16197 ( .A(n14393), .ZN(n14396) );
  OAI21_X1 U16198 ( .B1(n14396), .B2(n14395), .A(n14394), .ZN(n14398) );
  NAND2_X1 U16199 ( .A1(n14398), .A2(n14397), .ZN(n14399) );
  AOI222_X1 U16200 ( .A1(n6468), .A2(n14419), .B1(n14418), .B2(n14411), .C1(
        n14399), .C2(n14409), .ZN(n14401) );
  OAI211_X1 U16201 ( .C1(n14417), .C2(n14402), .A(n14401), .B(n14400), .ZN(
        P1_U3215) );
  INV_X1 U16202 ( .A(n14403), .ZN(n14406) );
  OAI21_X1 U16203 ( .B1(n14406), .B2(n14405), .A(n14404), .ZN(n14408) );
  NAND2_X1 U16204 ( .A1(n14408), .A2(n14407), .ZN(n14410) );
  AOI222_X1 U16205 ( .A1(n6468), .A2(n14413), .B1(n14412), .B2(n14411), .C1(
        n14410), .C2(n14409), .ZN(n14415) );
  OAI211_X1 U16206 ( .C1(n14417), .C2(n14416), .A(n14415), .B(n14414), .ZN(
        P1_U3236) );
  AOI21_X1 U16207 ( .B1(n14419), .B2(n14538), .A(n14418), .ZN(n14421) );
  OAI211_X1 U16208 ( .C1(n14422), .C2(n14521), .A(n14421), .B(n14420), .ZN(
        n14423) );
  AOI21_X1 U16209 ( .B1(n14526), .B2(n14424), .A(n14423), .ZN(n14432) );
  AOI22_X1 U16210 ( .A1(n14560), .A2(n14432), .B1(n11210), .B2(n14558), .ZN(
        P1_U3542) );
  OAI21_X1 U16211 ( .B1(n14426), .B2(n14528), .A(n14425), .ZN(n14428) );
  AOI211_X1 U16212 ( .C1(n14430), .C2(n14429), .A(n14428), .B(n14427), .ZN(
        n14434) );
  AOI22_X1 U16213 ( .A1(n14560), .A2(n14434), .B1(n10678), .B2(n14558), .ZN(
        P1_U3539) );
  INV_X1 U16214 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14431) );
  AOI22_X1 U16215 ( .A1(n14549), .A2(n14432), .B1(n14431), .B2(n14547), .ZN(
        P1_U3501) );
  INV_X1 U16216 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14433) );
  AOI22_X1 U16217 ( .A1(n14549), .A2(n14434), .B1(n14433), .B2(n14547), .ZN(
        P1_U3492) );
  OAI21_X1 U16218 ( .B1(n14437), .B2(n14436), .A(n14435), .ZN(n14438) );
  XNOR2_X1 U16219 ( .A(n14438), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  OAI21_X1 U16220 ( .B1(n14440), .B2(n14648), .A(n14439), .ZN(SUB_1596_U68) );
  OAI21_X1 U16221 ( .B1(n14443), .B2(n14442), .A(n14441), .ZN(n14444) );
  XNOR2_X1 U16222 ( .A(n14444), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(SUB_1596_U67)
         );
  OAI21_X1 U16223 ( .B1(n14447), .B2(n14446), .A(n14445), .ZN(n14448) );
  XNOR2_X1 U16224 ( .A(n14448), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  AOI21_X1 U16225 ( .B1(n14451), .B2(n14450), .A(n14449), .ZN(n14452) );
  XOR2_X1 U16226 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n14452), .Z(SUB_1596_U65)
         );
  AOI21_X1 U16227 ( .B1(n14455), .B2(n14454), .A(n14453), .ZN(n14456) );
  XOR2_X1 U16228 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n14456), .Z(SUB_1596_U64)
         );
  AOI21_X1 U16229 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14458), .A(n14457), 
        .ZN(n14469) );
  OAI21_X1 U16230 ( .B1(n14461), .B2(n14460), .A(n14459), .ZN(n14463) );
  NAND2_X1 U16231 ( .A1(n14463), .A2(n14462), .ZN(n14467) );
  NAND2_X1 U16232 ( .A1(n14465), .A2(n14464), .ZN(n14466) );
  OAI211_X1 U16233 ( .C1(n14469), .C2(n14468), .A(n14467), .B(n14466), .ZN(
        n14470) );
  INV_X1 U16234 ( .A(n14470), .ZN(n14472) );
  OAI211_X1 U16235 ( .C1(n14474), .C2(n14473), .A(n14472), .B(n14471), .ZN(
        P1_U3258) );
  INV_X1 U16236 ( .A(n14475), .ZN(n14481) );
  NOR2_X1 U16237 ( .A1(n14477), .A2(n14476), .ZN(n14478) );
  AOI21_X1 U16238 ( .B1(n14479), .B2(P1_REG2_REG_7__SCAN_IN), .A(n14478), .ZN(
        n14480) );
  OAI21_X1 U16239 ( .B1(n14482), .B2(n14481), .A(n14480), .ZN(n14483) );
  INV_X1 U16240 ( .A(n14483), .ZN(n14489) );
  AOI22_X1 U16241 ( .A1(n14487), .A2(n14486), .B1(n14485), .B2(n14484), .ZN(
        n14488) );
  OAI211_X1 U16242 ( .C1(n14491), .C2(n14490), .A(n14489), .B(n14488), .ZN(
        P1_U3286) );
  AND2_X1 U16243 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14492), .ZN(P1_U3294) );
  AND2_X1 U16244 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14492), .ZN(P1_U3295) );
  AND2_X1 U16245 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14492), .ZN(P1_U3296) );
  AND2_X1 U16246 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14492), .ZN(P1_U3297) );
  AND2_X1 U16247 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14492), .ZN(P1_U3298) );
  AND2_X1 U16248 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14492), .ZN(P1_U3299) );
  AND2_X1 U16249 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14492), .ZN(P1_U3300) );
  AND2_X1 U16250 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14492), .ZN(P1_U3301) );
  AND2_X1 U16251 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14492), .ZN(P1_U3302) );
  AND2_X1 U16252 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14492), .ZN(P1_U3303) );
  AND2_X1 U16253 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14492), .ZN(P1_U3304) );
  AND2_X1 U16254 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14492), .ZN(P1_U3305) );
  AND2_X1 U16255 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14492), .ZN(P1_U3306) );
  AND2_X1 U16256 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14492), .ZN(P1_U3307) );
  AND2_X1 U16257 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14492), .ZN(P1_U3308) );
  AND2_X1 U16258 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14492), .ZN(P1_U3309) );
  AND2_X1 U16259 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14492), .ZN(P1_U3310) );
  AND2_X1 U16260 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14492), .ZN(P1_U3311) );
  AND2_X1 U16261 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14492), .ZN(P1_U3312) );
  AND2_X1 U16262 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14492), .ZN(P1_U3313) );
  AND2_X1 U16263 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14492), .ZN(P1_U3314) );
  AND2_X1 U16264 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14492), .ZN(P1_U3315) );
  AND2_X1 U16265 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14492), .ZN(P1_U3316) );
  AND2_X1 U16266 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14492), .ZN(P1_U3317) );
  AND2_X1 U16267 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14492), .ZN(P1_U3318) );
  AND2_X1 U16268 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14492), .ZN(P1_U3319) );
  AND2_X1 U16269 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14492), .ZN(P1_U3320) );
  AND2_X1 U16270 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14492), .ZN(P1_U3321) );
  AND2_X1 U16271 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14492), .ZN(P1_U3322) );
  AND2_X1 U16272 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14492), .ZN(P1_U3323) );
  AOI22_X1 U16273 ( .A1(n14494), .A2(n14493), .B1(n14538), .B2(n10085), .ZN(
        n14495) );
  OAI211_X1 U16274 ( .C1(n14521), .C2(n14497), .A(n14496), .B(n14495), .ZN(
        n14498) );
  INV_X1 U16275 ( .A(n14498), .ZN(n14550) );
  INV_X1 U16276 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n14499) );
  AOI22_X1 U16277 ( .A1(n14549), .A2(n14550), .B1(n14499), .B2(n14547), .ZN(
        P1_U3462) );
  INV_X1 U16278 ( .A(n14507), .ZN(n14509) );
  INV_X1 U16279 ( .A(n14500), .ZN(n14502) );
  OAI211_X1 U16280 ( .C1(n14503), .C2(n14528), .A(n14502), .B(n14501), .ZN(
        n14504) );
  AOI21_X1 U16281 ( .B1(n14505), .B2(n14526), .A(n14504), .ZN(n14506) );
  OAI21_X1 U16282 ( .B1(n14507), .B2(n14541), .A(n14506), .ZN(n14508) );
  AOI21_X1 U16283 ( .B1(n14546), .B2(n14509), .A(n14508), .ZN(n14552) );
  AOI22_X1 U16284 ( .A1(n14549), .A2(n14552), .B1(n8711), .B2(n14547), .ZN(
        P1_U3465) );
  NAND2_X1 U16285 ( .A1(n14510), .A2(n14532), .ZN(n14513) );
  INV_X1 U16286 ( .A(n14511), .ZN(n14512) );
  OAI211_X1 U16287 ( .C1(n14514), .C2(n14528), .A(n14513), .B(n14512), .ZN(
        n14515) );
  NOR2_X1 U16288 ( .A1(n14516), .A2(n14515), .ZN(n14554) );
  INV_X1 U16289 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n14517) );
  AOI22_X1 U16290 ( .A1(n14549), .A2(n14554), .B1(n14517), .B2(n14547), .ZN(
        P1_U3468) );
  OAI211_X1 U16291 ( .C1(n14520), .C2(n14528), .A(n14519), .B(n14518), .ZN(
        n14524) );
  NOR2_X1 U16292 ( .A1(n14522), .A2(n14521), .ZN(n14523) );
  AOI211_X1 U16293 ( .C1(n14526), .C2(n14525), .A(n14524), .B(n14523), .ZN(
        n14555) );
  AOI22_X1 U16294 ( .A1(n14549), .A2(n14555), .B1(n8769), .B2(n14547), .ZN(
        P1_U3471) );
  OAI21_X1 U16295 ( .B1(n6627), .B2(n14528), .A(n14527), .ZN(n14530) );
  AOI211_X1 U16296 ( .C1(n14532), .C2(n14531), .A(n14530), .B(n14529), .ZN(
        n14557) );
  INV_X1 U16297 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n14533) );
  AOI22_X1 U16298 ( .A1(n14549), .A2(n14557), .B1(n14533), .B2(n14547), .ZN(
        P1_U3474) );
  NOR2_X1 U16299 ( .A1(n14535), .A2(n14534), .ZN(n14544) );
  INV_X1 U16300 ( .A(n14545), .ZN(n14542) );
  AOI21_X1 U16301 ( .B1(n14538), .B2(n14537), .A(n14536), .ZN(n14540) );
  OAI211_X1 U16302 ( .C1(n14542), .C2(n14541), .A(n14540), .B(n14539), .ZN(
        n14543) );
  AOI211_X1 U16303 ( .C1(n14546), .C2(n14545), .A(n14544), .B(n14543), .ZN(
        n14559) );
  INV_X1 U16304 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n14548) );
  AOI22_X1 U16305 ( .A1(n14549), .A2(n14559), .B1(n14548), .B2(n14547), .ZN(
        P1_U3477) );
  AOI22_X1 U16306 ( .A1(n14560), .A2(n14550), .B1(n10370), .B2(n14558), .ZN(
        P1_U3529) );
  AOI22_X1 U16307 ( .A1(n14560), .A2(n14552), .B1(n14551), .B2(n14558), .ZN(
        P1_U3530) );
  AOI22_X1 U16308 ( .A1(n14560), .A2(n14554), .B1(n14553), .B2(n14558), .ZN(
        P1_U3531) );
  AOI22_X1 U16309 ( .A1(n14560), .A2(n14555), .B1(n10372), .B2(n14558), .ZN(
        P1_U3532) );
  INV_X1 U16310 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n14556) );
  AOI22_X1 U16311 ( .A1(n14560), .A2(n14557), .B1(n14556), .B2(n14558), .ZN(
        P1_U3533) );
  AOI22_X1 U16312 ( .A1(n14560), .A2(n14559), .B1(n10373), .B2(n14558), .ZN(
        P1_U3534) );
  NOR2_X1 U16313 ( .A1(n14684), .A2(P2_U3947), .ZN(P2_U3087) );
  INV_X1 U16314 ( .A(n14561), .ZN(n14672) );
  OAI21_X1 U16315 ( .B1(n14672), .B2(n14562), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n14563) );
  OAI21_X1 U16316 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n14563), .ZN(n14574) );
  XOR2_X1 U16317 ( .A(n14565), .B(n14564), .Z(n14566) );
  NAND2_X1 U16318 ( .A1(n14692), .A2(n14566), .ZN(n14573) );
  NAND2_X1 U16319 ( .A1(n14568), .A2(n14567), .ZN(n14569) );
  NAND3_X1 U16320 ( .A1(n14688), .A2(n14570), .A3(n14569), .ZN(n14572) );
  NAND2_X1 U16321 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(n14684), .ZN(n14571) );
  NAND4_X1 U16322 ( .A1(n14574), .A2(n14573), .A3(n14572), .A4(n14571), .ZN(
        P2_U3216) );
  INV_X1 U16323 ( .A(n14575), .ZN(n14582) );
  AND3_X1 U16324 ( .A1(n14578), .A2(n14577), .A3(n14576), .ZN(n14579) );
  NOR3_X1 U16325 ( .A1(n14652), .A2(n14580), .A3(n14579), .ZN(n14581) );
  AOI211_X1 U16326 ( .C1(n14685), .C2(n14583), .A(n14582), .B(n14581), .ZN(
        n14588) );
  NAND2_X1 U16327 ( .A1(n14585), .A2(n14584), .ZN(n14586) );
  NAND3_X1 U16328 ( .A1(n14688), .A2(n14593), .A3(n14586), .ZN(n14587) );
  OAI211_X1 U16329 ( .C1(n14647), .C2(n14589), .A(n14588), .B(n14587), .ZN(
        P2_U3218) );
  INV_X1 U16330 ( .A(n14590), .ZN(n14598) );
  AND3_X1 U16331 ( .A1(n14593), .A2(n14592), .A3(n14591), .ZN(n14594) );
  NOR3_X1 U16332 ( .A1(n14596), .A2(n14595), .A3(n14594), .ZN(n14597) );
  AOI211_X1 U16333 ( .C1(n14685), .C2(n14599), .A(n14598), .B(n14597), .ZN(
        n14605) );
  AOI211_X1 U16334 ( .C1(n14602), .C2(n14601), .A(n14600), .B(n14652), .ZN(
        n14603) );
  INV_X1 U16335 ( .A(n14603), .ZN(n14604) );
  OAI211_X1 U16336 ( .C1(n14647), .C2(n15136), .A(n14605), .B(n14604), .ZN(
        P2_U3219) );
  INV_X1 U16337 ( .A(n14606), .ZN(n14607) );
  OAI21_X1 U16338 ( .B1(n14609), .B2(n14608), .A(n14607), .ZN(n14615) );
  OAI21_X1 U16339 ( .B1(n14612), .B2(n14611), .A(n14610), .ZN(n14613) );
  AOI222_X1 U16340 ( .A1(n14615), .A2(n14688), .B1(n14614), .B2(n14685), .C1(
        n14613), .C2(n14692), .ZN(n14617) );
  OAI211_X1 U16341 ( .C1(n14618), .C2(n14647), .A(n14617), .B(n14616), .ZN(
        P2_U3223) );
  NOR2_X1 U16342 ( .A1(n14620), .A2(n14619), .ZN(n14621) );
  AOI211_X1 U16343 ( .C1(n14684), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n14622), 
        .B(n14621), .ZN(n14632) );
  OAI211_X1 U16344 ( .C1(n14625), .C2(n14624), .A(n14623), .B(n14688), .ZN(
        n14631) );
  AOI211_X1 U16345 ( .C1(n14628), .C2(n14627), .A(n14652), .B(n14626), .ZN(
        n14629) );
  INV_X1 U16346 ( .A(n14629), .ZN(n14630) );
  NAND3_X1 U16347 ( .A1(n14632), .A2(n14631), .A3(n14630), .ZN(P2_U3224) );
  INV_X1 U16348 ( .A(n14633), .ZN(n14634) );
  OAI21_X1 U16349 ( .B1(n14636), .B2(n14635), .A(n14634), .ZN(n14644) );
  OR3_X1 U16350 ( .A1(n14639), .A2(n14638), .A3(n14637), .ZN(n14640) );
  NAND2_X1 U16351 ( .A1(n14641), .A2(n14640), .ZN(n14642) );
  AOI222_X1 U16352 ( .A1(n14644), .A2(n14688), .B1(n14643), .B2(n14685), .C1(
        n14642), .C2(n14692), .ZN(n14646) );
  NAND2_X1 U16353 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n14645)
         );
  OAI211_X1 U16354 ( .C1(n14648), .C2(n14647), .A(n14646), .B(n14645), .ZN(
        P2_U3226) );
  AOI22_X1 U16355 ( .A1(n14684), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(P2_U3088), .ZN(n14661) );
  OAI211_X1 U16356 ( .C1(n14651), .C2(n14650), .A(n14649), .B(n14688), .ZN(
        n14660) );
  AOI21_X1 U16357 ( .B1(n14654), .B2(n14653), .A(n14652), .ZN(n14656) );
  NAND2_X1 U16358 ( .A1(n14656), .A2(n14655), .ZN(n14659) );
  NAND2_X1 U16359 ( .A1(n14657), .A2(n14685), .ZN(n14658) );
  NAND4_X1 U16360 ( .A1(n14661), .A2(n14660), .A3(n14659), .A4(n14658), .ZN(
        P2_U3227) );
  AOI22_X1 U16361 ( .A1(n14684), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n14670) );
  NAND2_X1 U16362 ( .A1(n14685), .A2(n14662), .ZN(n14669) );
  OAI211_X1 U16363 ( .C1(n14664), .C2(P2_REG2_REG_15__SCAN_IN), .A(n14692), 
        .B(n14663), .ZN(n14668) );
  OAI211_X1 U16364 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n14666), .A(n14688), 
        .B(n14665), .ZN(n14667) );
  NAND4_X1 U16365 ( .A1(n14670), .A2(n14669), .A3(n14668), .A4(n14667), .ZN(
        P2_U3229) );
  OAI21_X1 U16366 ( .B1(n14672), .B2(n14671), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n14673) );
  OAI21_X1 U16367 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n14673), .ZN(n14683) );
  OAI211_X1 U16368 ( .C1(n14676), .C2(n14675), .A(n14692), .B(n14674), .ZN(
        n14682) );
  NAND2_X1 U16369 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n14684), .ZN(n14681) );
  OAI211_X1 U16370 ( .C1(n14679), .C2(n14678), .A(n14688), .B(n14677), .ZN(
        n14680) );
  NAND4_X1 U16371 ( .A1(n14683), .A2(n14682), .A3(n14681), .A4(n14680), .ZN(
        P2_U3230) );
  AOI22_X1 U16372 ( .A1(n14684), .A2(P2_ADDR_REG_17__SCAN_IN), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(P2_U3088), .ZN(n14698) );
  NAND2_X1 U16373 ( .A1(n14686), .A2(n14685), .ZN(n14697) );
  OAI211_X1 U16374 ( .C1(n14690), .C2(n14689), .A(n14688), .B(n14687), .ZN(
        n14696) );
  OAI211_X1 U16375 ( .C1(n14694), .C2(n14693), .A(n14692), .B(n14691), .ZN(
        n14695) );
  NAND4_X1 U16376 ( .A1(n14698), .A2(n14697), .A3(n14696), .A4(n14695), .ZN(
        P2_U3231) );
  NAND2_X1 U16377 ( .A1(n14700), .A2(n14699), .ZN(n14701) );
  XOR2_X1 U16378 ( .A(n14708), .B(n14701), .Z(n14703) );
  AOI21_X1 U16379 ( .B1(n14703), .B2(n14725), .A(n14702), .ZN(n14806) );
  AOI222_X1 U16380 ( .A1(n14710), .A2(n14706), .B1(P2_REG2_REG_9__SCAN_IN), 
        .B2(n14736), .C1(n14705), .C2(n14704), .ZN(n14718) );
  OAI21_X1 U16381 ( .B1(n14709), .B2(n14708), .A(n14707), .ZN(n14803) );
  AOI21_X1 U16382 ( .B1(n14711), .B2(n14710), .A(n11505), .ZN(n14713) );
  NAND2_X1 U16383 ( .A1(n14713), .A2(n14712), .ZN(n14804) );
  OAI22_X1 U16384 ( .A1(n14803), .A2(n14715), .B1(n14714), .B2(n14804), .ZN(
        n14716) );
  INV_X1 U16385 ( .A(n14716), .ZN(n14717) );
  OAI211_X1 U16386 ( .C1(n14736), .C2(n14806), .A(n14718), .B(n14717), .ZN(
        P2_U3256) );
  INV_X1 U16387 ( .A(n14749), .ZN(n14731) );
  INV_X1 U16388 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n14723) );
  AOI21_X1 U16389 ( .B1(n14720), .B2(n14745), .A(n14719), .ZN(n14722) );
  OAI22_X1 U16390 ( .A1(n14724), .A2(n14723), .B1(n14722), .B2(n14721), .ZN(
        n14730) );
  NOR2_X1 U16391 ( .A1(n14801), .A2(n14725), .ZN(n14726) );
  OR2_X1 U16392 ( .A1(n14749), .A2(n14726), .ZN(n14728) );
  AND2_X1 U16393 ( .A1(n14728), .A2(n14727), .ZN(n14748) );
  INV_X1 U16394 ( .A(n14748), .ZN(n14729) );
  AOI211_X1 U16395 ( .C1(n14732), .C2(n14731), .A(n14730), .B(n14729), .ZN(
        n14734) );
  AOI22_X1 U16396 ( .A1(n14736), .A2(n14735), .B1(n14734), .B2(n14733), .ZN(
        P2_U3265) );
  AND2_X1 U16397 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14738), .ZN(P2_U3266) );
  AND2_X1 U16398 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14738), .ZN(P2_U3267) );
  AND2_X1 U16399 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14738), .ZN(P2_U3268) );
  AND2_X1 U16400 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n14738), .ZN(P2_U3269) );
  AND2_X1 U16401 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14738), .ZN(P2_U3270) );
  AND2_X1 U16402 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14738), .ZN(P2_U3271) );
  AND2_X1 U16403 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14738), .ZN(P2_U3272) );
  AND2_X1 U16404 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14738), .ZN(P2_U3273) );
  AND2_X1 U16405 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14738), .ZN(P2_U3274) );
  AND2_X1 U16406 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14738), .ZN(P2_U3275) );
  AND2_X1 U16407 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14738), .ZN(P2_U3276) );
  AND2_X1 U16408 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14738), .ZN(P2_U3277) );
  AND2_X1 U16409 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14738), .ZN(P2_U3278) );
  AND2_X1 U16410 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14738), .ZN(P2_U3279) );
  AND2_X1 U16411 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14738), .ZN(P2_U3280) );
  AND2_X1 U16412 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14738), .ZN(P2_U3281) );
  AND2_X1 U16413 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14738), .ZN(P2_U3282) );
  AND2_X1 U16414 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14738), .ZN(P2_U3283) );
  AND2_X1 U16415 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14738), .ZN(P2_U3284) );
  AND2_X1 U16416 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14738), .ZN(P2_U3285) );
  AND2_X1 U16417 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14738), .ZN(P2_U3286) );
  AND2_X1 U16418 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14738), .ZN(P2_U3287) );
  AND2_X1 U16419 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14738), .ZN(P2_U3288) );
  AND2_X1 U16420 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14738), .ZN(P2_U3289) );
  AND2_X1 U16421 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14738), .ZN(P2_U3290) );
  AND2_X1 U16422 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14738), .ZN(P2_U3291) );
  AND2_X1 U16423 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14738), .ZN(P2_U3292) );
  AND2_X1 U16424 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14738), .ZN(P2_U3293) );
  AND2_X1 U16425 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14738), .ZN(P2_U3294) );
  AND2_X1 U16426 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14738), .ZN(P2_U3295) );
  AOI22_X1 U16427 ( .A1(n14741), .A2(n14740), .B1(n14739), .B2(n14743), .ZN(
        P2_U3416) );
  AOI21_X1 U16428 ( .B1(n14744), .B2(n14743), .A(n14742), .ZN(P2_U3417) );
  NAND2_X1 U16429 ( .A1(n14746), .A2(n14745), .ZN(n14747) );
  OAI211_X1 U16430 ( .C1(n14749), .C2(n14769), .A(n14748), .B(n14747), .ZN(
        n14832) );
  OAI22_X1 U16431 ( .A1(n14829), .A2(n14832), .B1(P2_REG0_REG_0__SCAN_IN), 
        .B2(n14831), .ZN(n14750) );
  INV_X1 U16432 ( .A(n14750), .ZN(P2_U3430) );
  INV_X1 U16433 ( .A(n14751), .ZN(n14752) );
  AOI21_X1 U16434 ( .B1(n10449), .B2(n14769), .A(n14752), .ZN(n14757) );
  OAI211_X1 U16435 ( .C1(n14755), .C2(n14822), .A(n14754), .B(n14753), .ZN(
        n14756) );
  NOR2_X1 U16436 ( .A1(n14757), .A2(n14756), .ZN(n14835) );
  AOI22_X1 U16437 ( .A1(n14831), .A2(n14835), .B1(n8190), .B2(n14829), .ZN(
        P2_U3433) );
  INV_X1 U16438 ( .A(n14769), .ZN(n14825) );
  OAI21_X1 U16439 ( .B1(n14759), .B2(n14822), .A(n14758), .ZN(n14760) );
  AOI21_X1 U16440 ( .B1(n14761), .B2(n14825), .A(n14760), .ZN(n14762) );
  AND2_X1 U16441 ( .A1(n14763), .A2(n14762), .ZN(n14837) );
  INV_X1 U16442 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n14764) );
  AOI22_X1 U16443 ( .A1(n14831), .A2(n14837), .B1(n14764), .B2(n14829), .ZN(
        P2_U3436) );
  INV_X1 U16444 ( .A(n14770), .ZN(n14772) );
  AOI21_X1 U16445 ( .B1(n14814), .B2(n14766), .A(n14765), .ZN(n14767) );
  OAI211_X1 U16446 ( .C1(n14770), .C2(n14769), .A(n14768), .B(n14767), .ZN(
        n14771) );
  AOI21_X1 U16447 ( .B1(n14801), .B2(n14772), .A(n14771), .ZN(n14839) );
  INV_X1 U16448 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n14773) );
  AOI22_X1 U16449 ( .A1(n14831), .A2(n14839), .B1(n14773), .B2(n14829), .ZN(
        P2_U3439) );
  AND2_X1 U16450 ( .A1(n14774), .A2(n14809), .ZN(n14779) );
  OAI21_X1 U16451 ( .B1(n14776), .B2(n14822), .A(n14775), .ZN(n14777) );
  NOR3_X1 U16452 ( .A1(n14779), .A2(n14778), .A3(n14777), .ZN(n14841) );
  INV_X1 U16453 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n14780) );
  AOI22_X1 U16454 ( .A1(n14831), .A2(n14841), .B1(n14780), .B2(n14829), .ZN(
        P2_U3442) );
  AND2_X1 U16455 ( .A1(n14781), .A2(n14809), .ZN(n14786) );
  OAI21_X1 U16456 ( .B1(n14783), .B2(n14822), .A(n14782), .ZN(n14784) );
  NOR3_X1 U16457 ( .A1(n14786), .A2(n14785), .A3(n14784), .ZN(n14843) );
  INV_X1 U16458 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n14787) );
  AOI22_X1 U16459 ( .A1(n14831), .A2(n14843), .B1(n14787), .B2(n14829), .ZN(
        P2_U3445) );
  AOI21_X1 U16460 ( .B1(n14814), .B2(n14789), .A(n14788), .ZN(n14790) );
  OAI211_X1 U16461 ( .C1(n14792), .C2(n14817), .A(n14791), .B(n14790), .ZN(
        n14793) );
  INV_X1 U16462 ( .A(n14793), .ZN(n14844) );
  INV_X1 U16463 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n14794) );
  AOI22_X1 U16464 ( .A1(n14831), .A2(n14844), .B1(n14794), .B2(n14829), .ZN(
        P2_U3451) );
  NAND2_X1 U16465 ( .A1(n14800), .A2(n14825), .ZN(n14796) );
  OAI211_X1 U16466 ( .C1(n14797), .C2(n14822), .A(n14796), .B(n14795), .ZN(
        n14798) );
  AOI211_X1 U16467 ( .C1(n14801), .C2(n14800), .A(n14799), .B(n14798), .ZN(
        n14846) );
  INV_X1 U16468 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n14802) );
  AOI22_X1 U16469 ( .A1(n14831), .A2(n14846), .B1(n14802), .B2(n14829), .ZN(
        P2_U3454) );
  INV_X1 U16470 ( .A(n14803), .ZN(n14810) );
  OAI21_X1 U16471 ( .B1(n14805), .B2(n14822), .A(n14804), .ZN(n14808) );
  INV_X1 U16472 ( .A(n14806), .ZN(n14807) );
  AOI211_X1 U16473 ( .C1(n14810), .C2(n14809), .A(n14808), .B(n14807), .ZN(
        n14848) );
  INV_X1 U16474 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n14811) );
  AOI22_X1 U16475 ( .A1(n14831), .A2(n14848), .B1(n14811), .B2(n14829), .ZN(
        P2_U3457) );
  AOI21_X1 U16476 ( .B1(n14814), .B2(n14813), .A(n14812), .ZN(n14815) );
  OAI211_X1 U16477 ( .C1(n14818), .C2(n14817), .A(n14816), .B(n14815), .ZN(
        n14819) );
  INV_X1 U16478 ( .A(n14819), .ZN(n14849) );
  INV_X1 U16479 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n14820) );
  AOI22_X1 U16480 ( .A1(n14831), .A2(n14849), .B1(n14820), .B2(n14829), .ZN(
        P2_U3460) );
  OAI21_X1 U16481 ( .B1(n14823), .B2(n14822), .A(n14821), .ZN(n14824) );
  AOI21_X1 U16482 ( .B1(n14826), .B2(n14825), .A(n14824), .ZN(n14827) );
  INV_X1 U16483 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n14830) );
  AOI22_X1 U16484 ( .A1(n14831), .A2(n14852), .B1(n14830), .B2(n14829), .ZN(
        P2_U3463) );
  OAI22_X1 U16485 ( .A1(n14850), .A2(n14832), .B1(P2_REG1_REG_0__SCAN_IN), 
        .B2(n14853), .ZN(n14833) );
  INV_X1 U16486 ( .A(n14833), .ZN(P2_U3499) );
  AOI22_X1 U16487 ( .A1(n14853), .A2(n14835), .B1(n14834), .B2(n14850), .ZN(
        P2_U3500) );
  AOI22_X1 U16488 ( .A1(n14853), .A2(n14837), .B1(n14836), .B2(n14850), .ZN(
        P2_U3501) );
  AOI22_X1 U16489 ( .A1(n14853), .A2(n14839), .B1(n14838), .B2(n14850), .ZN(
        P2_U3502) );
  AOI22_X1 U16490 ( .A1(n14853), .A2(n14841), .B1(n14840), .B2(n14850), .ZN(
        P2_U3503) );
  AOI22_X1 U16491 ( .A1(n14853), .A2(n14843), .B1(n14842), .B2(n14850), .ZN(
        P2_U3504) );
  AOI22_X1 U16492 ( .A1(n14853), .A2(n14844), .B1(n10256), .B2(n14850), .ZN(
        P2_U3506) );
  AOI22_X1 U16493 ( .A1(n14853), .A2(n14846), .B1(n14845), .B2(n14850), .ZN(
        P2_U3507) );
  AOI22_X1 U16494 ( .A1(n14853), .A2(n14848), .B1(n14847), .B2(n14850), .ZN(
        P2_U3508) );
  AOI22_X1 U16495 ( .A1(n14853), .A2(n14849), .B1(n10587), .B2(n14850), .ZN(
        P2_U3509) );
  AOI22_X1 U16496 ( .A1(n14853), .A2(n14852), .B1(n14851), .B2(n14850), .ZN(
        P2_U3510) );
  NOR2_X1 U16497 ( .A1(P3_U3897), .A2(n14969), .ZN(P3_U3150) );
  AOI21_X1 U16498 ( .B1(n11621), .B2(n14855), .A(n14854), .ZN(n14869) );
  AND3_X1 U16499 ( .A1(n14858), .A2(n14857), .A3(n14856), .ZN(n14859) );
  OAI21_X1 U16500 ( .B1(n14874), .B2(n14859), .A(n14962), .ZN(n14860) );
  OAI21_X1 U16501 ( .B1(n14966), .B2(n14861), .A(n14860), .ZN(n14862) );
  AOI211_X1 U16502 ( .C1(P3_ADDR_REG_3__SCAN_IN), .C2(n14969), .A(n14863), .B(
        n14862), .ZN(n14868) );
  OAI21_X1 U16503 ( .B1(P3_REG1_REG_3__SCAN_IN), .B2(n14865), .A(n14864), .ZN(
        n14866) );
  NAND2_X1 U16504 ( .A1(n6467), .A2(n14866), .ZN(n14867) );
  OAI211_X1 U16505 ( .C1(n14869), .C2(n14991), .A(n14868), .B(n14867), .ZN(
        P3_U3185) );
  AOI21_X1 U16506 ( .B1(n6615), .B2(n14871), .A(n14870), .ZN(n14887) );
  INV_X1 U16507 ( .A(n14892), .ZN(n14876) );
  NOR3_X1 U16508 ( .A1(n14874), .A2(n14873), .A3(n14872), .ZN(n14875) );
  OAI21_X1 U16509 ( .B1(n14876), .B2(n14875), .A(n14962), .ZN(n14877) );
  OAI21_X1 U16510 ( .B1(n14966), .B2(n14878), .A(n14877), .ZN(n14879) );
  AOI211_X1 U16511 ( .C1(P3_ADDR_REG_4__SCAN_IN), .C2(n14969), .A(n14880), .B(
        n14879), .ZN(n14886) );
  OAI21_X1 U16512 ( .B1(n14883), .B2(n14882), .A(n14881), .ZN(n14884) );
  NAND2_X1 U16513 ( .A1(n6467), .A2(n14884), .ZN(n14885) );
  OAI211_X1 U16514 ( .C1(n14887), .C2(n14991), .A(n14886), .B(n14885), .ZN(
        P3_U3186) );
  AOI21_X1 U16515 ( .B1(n11632), .B2(n14889), .A(n14888), .ZN(n14903) );
  AND3_X1 U16516 ( .A1(n14892), .A2(n14891), .A3(n14890), .ZN(n14893) );
  OAI21_X1 U16517 ( .B1(n14909), .B2(n14893), .A(n14962), .ZN(n14894) );
  OAI21_X1 U16518 ( .B1(n14966), .B2(n14895), .A(n14894), .ZN(n14896) );
  AOI211_X1 U16519 ( .C1(P3_ADDR_REG_5__SCAN_IN), .C2(n14969), .A(n14897), .B(
        n14896), .ZN(n14902) );
  OAI21_X1 U16520 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n14899), .A(n14898), .ZN(
        n14900) );
  NAND2_X1 U16521 ( .A1(n6467), .A2(n14900), .ZN(n14901) );
  OAI211_X1 U16522 ( .C1(n14903), .C2(n14991), .A(n14902), .B(n14901), .ZN(
        P3_U3187) );
  AOI21_X1 U16523 ( .B1(n14906), .B2(n14905), .A(n14904), .ZN(n14922) );
  INV_X1 U16524 ( .A(n14927), .ZN(n14911) );
  NOR3_X1 U16525 ( .A1(n14909), .A2(n14908), .A3(n14907), .ZN(n14910) );
  OAI21_X1 U16526 ( .B1(n14911), .B2(n14910), .A(n14962), .ZN(n14912) );
  OAI21_X1 U16527 ( .B1(n14966), .B2(n14913), .A(n14912), .ZN(n14914) );
  AOI211_X1 U16528 ( .C1(P3_ADDR_REG_6__SCAN_IN), .C2(n14969), .A(n14915), .B(
        n14914), .ZN(n14921) );
  OAI21_X1 U16529 ( .B1(n14918), .B2(n14917), .A(n14916), .ZN(n14919) );
  NAND2_X1 U16530 ( .A1(n14919), .A2(n6467), .ZN(n14920) );
  OAI211_X1 U16531 ( .C1(n14922), .C2(n14991), .A(n14921), .B(n14920), .ZN(
        P3_U3188) );
  AOI21_X1 U16532 ( .B1(n11642), .B2(n14924), .A(n14923), .ZN(n14938) );
  AND3_X1 U16533 ( .A1(n14927), .A2(n14926), .A3(n14925), .ZN(n14928) );
  OAI21_X1 U16534 ( .B1(n14943), .B2(n14928), .A(n14962), .ZN(n14929) );
  OAI21_X1 U16535 ( .B1(n14966), .B2(n14930), .A(n14929), .ZN(n14931) );
  AOI211_X1 U16536 ( .C1(P3_ADDR_REG_7__SCAN_IN), .C2(n14969), .A(n14932), .B(
        n14931), .ZN(n14937) );
  OAI21_X1 U16537 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n14934), .A(n14933), .ZN(
        n14935) );
  NAND2_X1 U16538 ( .A1(n14935), .A2(n6467), .ZN(n14936) );
  OAI211_X1 U16539 ( .C1(n14938), .C2(n14991), .A(n14937), .B(n14936), .ZN(
        P3_U3189) );
  AOI21_X1 U16540 ( .B1(n6612), .B2(n14940), .A(n14939), .ZN(n14956) );
  INV_X1 U16541 ( .A(n14961), .ZN(n14945) );
  NOR3_X1 U16542 ( .A1(n14943), .A2(n14942), .A3(n14941), .ZN(n14944) );
  OAI21_X1 U16543 ( .B1(n14945), .B2(n14944), .A(n14962), .ZN(n14946) );
  OAI21_X1 U16544 ( .B1(n14966), .B2(n14947), .A(n14946), .ZN(n14948) );
  AOI211_X1 U16545 ( .C1(P3_ADDR_REG_8__SCAN_IN), .C2(n14969), .A(n14949), .B(
        n14948), .ZN(n14955) );
  OAI21_X1 U16546 ( .B1(n14952), .B2(n14951), .A(n14950), .ZN(n14953) );
  NAND2_X1 U16547 ( .A1(n14953), .A2(n6467), .ZN(n14954) );
  OAI211_X1 U16548 ( .C1(n14956), .C2(n14991), .A(n14955), .B(n14954), .ZN(
        P3_U3190) );
  AOI21_X1 U16549 ( .B1(n11652), .B2(n14958), .A(n14957), .ZN(n14975) );
  AND3_X1 U16550 ( .A1(n14961), .A2(n14960), .A3(n14959), .ZN(n14963) );
  OAI21_X1 U16551 ( .B1(n14984), .B2(n14963), .A(n14962), .ZN(n14964) );
  OAI21_X1 U16552 ( .B1(n14966), .B2(n14965), .A(n14964), .ZN(n14967) );
  AOI211_X1 U16553 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n14969), .A(n14968), .B(
        n14967), .ZN(n14974) );
  OAI21_X1 U16554 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n14971), .A(n14970), .ZN(
        n14972) );
  NAND2_X1 U16555 ( .A1(n14972), .A2(n6467), .ZN(n14973) );
  OAI211_X1 U16556 ( .C1(n14975), .C2(n14991), .A(n14974), .B(n14973), .ZN(
        P3_U3191) );
  OAI21_X1 U16557 ( .B1(n14978), .B2(n14977), .A(n14976), .ZN(n14981) );
  AOI21_X1 U16558 ( .B1(n14981), .B2(n6467), .A(n14979), .ZN(n14998) );
  OR3_X1 U16559 ( .A1(n14984), .A2(n14983), .A3(n14982), .ZN(n14986) );
  AOI21_X1 U16560 ( .B1(n14987), .B2(n14986), .A(n14985), .ZN(n14994) );
  AOI21_X1 U16561 ( .B1(n14990), .B2(n14989), .A(n14988), .ZN(n14992) );
  NOR2_X1 U16562 ( .A1(n14992), .A2(n14991), .ZN(n14993) );
  AOI211_X1 U16563 ( .C1(n14996), .C2(n14995), .A(n14994), .B(n14993), .ZN(
        n14997) );
  OAI211_X1 U16564 ( .C1(n15000), .C2(n14999), .A(n14998), .B(n14997), .ZN(
        P3_U3192) );
  AOI21_X1 U16565 ( .B1(n15002), .B2(n15019), .A(n15001), .ZN(n15006) );
  AOI22_X1 U16566 ( .A1(n15004), .A2(n15003), .B1(P3_REG2_REG_9__SCAN_IN), 
        .B2(n15082), .ZN(n15005) );
  OAI21_X1 U16567 ( .B1(n15006), .B2(n15082), .A(n15005), .ZN(n15007) );
  INV_X1 U16568 ( .A(n15007), .ZN(n15008) );
  OAI21_X1 U16569 ( .B1(n15010), .B2(n15009), .A(n15008), .ZN(P3_U3224) );
  XNOR2_X1 U16570 ( .A(n15011), .B(n15015), .ZN(n15101) );
  INV_X1 U16571 ( .A(n15012), .ZN(n15013) );
  AOI21_X1 U16572 ( .B1(n15015), .B2(n15014), .A(n15013), .ZN(n15016) );
  OAI222_X1 U16573 ( .A1(n14339), .A2(n15018), .B1(n14341), .B2(n15017), .C1(
        n15045), .C2(n15016), .ZN(n15098) );
  AOI21_X1 U16574 ( .B1(n15101), .B2(n15019), .A(n15098), .ZN(n15023) );
  AND2_X1 U16575 ( .A1(n15020), .A2(n15071), .ZN(n15099) );
  AOI22_X1 U16576 ( .A1(n15036), .A2(n15099), .B1(n15077), .B2(n15021), .ZN(
        n15022) );
  OAI221_X1 U16577 ( .B1(n15082), .B2(n15023), .C1(n15080), .C2(n11632), .A(
        n15022), .ZN(P3_U3228) );
  OAI21_X1 U16578 ( .B1(n15026), .B2(n15025), .A(n15024), .ZN(n15096) );
  XNOR2_X1 U16579 ( .A(n15028), .B(n15027), .ZN(n15032) );
  OAI22_X1 U16580 ( .A1(n15041), .A2(n14341), .B1(n15029), .B2(n14339), .ZN(
        n15030) );
  AOI21_X1 U16581 ( .B1(n15096), .B2(n15070), .A(n15030), .ZN(n15031) );
  OAI21_X1 U16582 ( .B1(n15032), .B2(n15045), .A(n15031), .ZN(n15094) );
  AOI21_X1 U16583 ( .B1(n15033), .B2(n15096), .A(n15094), .ZN(n15038) );
  NOR2_X1 U16584 ( .A1(n15034), .A2(n15115), .ZN(n15095) );
  AOI22_X1 U16585 ( .A1(n15036), .A2(n15095), .B1(n15077), .B2(n15035), .ZN(
        n15037) );
  OAI221_X1 U16586 ( .B1(n15082), .B2(n15038), .C1(n15080), .C2(n11627), .A(
        n15037), .ZN(P3_U3229) );
  OAI21_X1 U16587 ( .B1(n15040), .B2(n15044), .A(n15039), .ZN(n15089) );
  OAI22_X1 U16588 ( .A1(n15042), .A2(n14341), .B1(n15041), .B2(n14339), .ZN(
        n15049) );
  NAND3_X1 U16589 ( .A1(n15058), .A2(n15044), .A3(n15043), .ZN(n15046) );
  AOI21_X1 U16590 ( .B1(n15047), .B2(n15046), .A(n15045), .ZN(n15048) );
  AOI211_X1 U16591 ( .C1(n15070), .C2(n15089), .A(n15049), .B(n15048), .ZN(
        n15050) );
  INV_X1 U16592 ( .A(n15050), .ZN(n15087) );
  INV_X1 U16593 ( .A(n15089), .ZN(n15055) );
  NOR2_X1 U16594 ( .A1(n15051), .A2(n15115), .ZN(n15088) );
  INV_X1 U16595 ( .A(n15088), .ZN(n15052) );
  OAI22_X1 U16596 ( .A1(n15055), .A2(n15054), .B1(n15053), .B2(n15052), .ZN(
        n15056) );
  AOI211_X1 U16597 ( .C1(P3_REG3_REG_2__SCAN_IN), .C2(n15077), .A(n15087), .B(
        n15056), .ZN(n15057) );
  AOI22_X1 U16598 ( .A1(n15082), .A2(n10331), .B1(n15057), .B2(n15080), .ZN(
        P3_U3231) );
  OAI21_X1 U16599 ( .B1(n15068), .B2(n15059), .A(n15058), .ZN(n15061) );
  NAND2_X1 U16600 ( .A1(n15061), .A2(n15060), .ZN(n15066) );
  AOI22_X1 U16601 ( .A1(n15064), .A2(n15063), .B1(n15062), .B2(n10404), .ZN(
        n15065) );
  NAND2_X1 U16602 ( .A1(n15066), .A2(n15065), .ZN(n15083) );
  INV_X1 U16603 ( .A(n15083), .ZN(n15076) );
  INV_X1 U16604 ( .A(n15067), .ZN(n15069) );
  XNOR2_X1 U16605 ( .A(n15069), .B(n15068), .ZN(n15085) );
  NAND2_X1 U16606 ( .A1(n15085), .A2(n15070), .ZN(n15075) );
  AND2_X1 U16607 ( .A1(n15072), .A2(n15071), .ZN(n15084) );
  NAND2_X1 U16608 ( .A1(n15084), .A2(n15073), .ZN(n15074) );
  AND3_X1 U16609 ( .A1(n15076), .A2(n15075), .A3(n15074), .ZN(n15081) );
  AOI22_X1 U16610 ( .A1(n15085), .A2(n15078), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15077), .ZN(n15079) );
  OAI221_X1 U16611 ( .B1(n15082), .B2(n15081), .C1(n15080), .C2(n10326), .A(
        n15079), .ZN(P3_U3232) );
  INV_X1 U16612 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15086) );
  AOI211_X1 U16613 ( .C1(n15100), .C2(n15085), .A(n15084), .B(n15083), .ZN(
        n15122) );
  AOI22_X1 U16614 ( .A1(n15121), .A2(n15086), .B1(n15122), .B2(n15120), .ZN(
        P3_U3393) );
  AOI211_X1 U16615 ( .C1(n15112), .C2(n15089), .A(n15088), .B(n15087), .ZN(
        n15123) );
  AOI22_X1 U16616 ( .A1(n15121), .A2(n7541), .B1(n15123), .B2(n15120), .ZN(
        P3_U3396) );
  INV_X1 U16617 ( .A(n15090), .ZN(n15091) );
  AOI211_X1 U16618 ( .C1(n15093), .C2(n15112), .A(n15092), .B(n15091), .ZN(
        n15124) );
  AOI22_X1 U16619 ( .A1(n15121), .A2(n7558), .B1(n15124), .B2(n15120), .ZN(
        P3_U3399) );
  INV_X1 U16620 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15097) );
  AOI211_X1 U16621 ( .C1(n15112), .C2(n15096), .A(n15095), .B(n15094), .ZN(
        n15125) );
  AOI22_X1 U16622 ( .A1(n15121), .A2(n15097), .B1(n15125), .B2(n15120), .ZN(
        P3_U3402) );
  AOI211_X1 U16623 ( .C1(n15101), .C2(n15100), .A(n15099), .B(n15098), .ZN(
        n15126) );
  AOI22_X1 U16624 ( .A1(n15121), .A2(n7589), .B1(n15126), .B2(n15120), .ZN(
        P3_U3405) );
  AOI211_X1 U16625 ( .C1(n15104), .C2(n15112), .A(n15103), .B(n15102), .ZN(
        n15127) );
  AOI22_X1 U16626 ( .A1(n15121), .A2(n7608), .B1(n15127), .B2(n15120), .ZN(
        P3_U3408) );
  AOI211_X1 U16627 ( .C1(n15112), .C2(n15107), .A(n15106), .B(n15105), .ZN(
        n15128) );
  AOI22_X1 U16628 ( .A1(n15121), .A2(n7622), .B1(n15128), .B2(n15120), .ZN(
        P3_U3411) );
  INV_X1 U16629 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15113) );
  NOR2_X1 U16630 ( .A1(n15108), .A2(n15115), .ZN(n15110) );
  AOI211_X1 U16631 ( .C1(n15112), .C2(n15111), .A(n15110), .B(n15109), .ZN(
        n15129) );
  AOI22_X1 U16632 ( .A1(n15121), .A2(n15113), .B1(n15129), .B2(n15120), .ZN(
        P3_U3414) );
  OAI22_X1 U16633 ( .A1(n15117), .A2(n15116), .B1(n15115), .B2(n15114), .ZN(
        n15118) );
  NOR2_X1 U16634 ( .A1(n15119), .A2(n15118), .ZN(n15130) );
  AOI22_X1 U16635 ( .A1(n15121), .A2(n7675), .B1(n15130), .B2(n15120), .ZN(
        P3_U3420) );
  AOI22_X1 U16636 ( .A1(n15131), .A2(n15122), .B1(n10325), .B2(n9450), .ZN(
        P3_U3460) );
  AOI22_X1 U16637 ( .A1(n15131), .A2(n15123), .B1(n10356), .B2(n9450), .ZN(
        P3_U3461) );
  AOI22_X1 U16638 ( .A1(n15131), .A2(n15124), .B1(n11620), .B2(n9450), .ZN(
        P3_U3462) );
  AOI22_X1 U16639 ( .A1(n15131), .A2(n15125), .B1(n11626), .B2(n9450), .ZN(
        P3_U3463) );
  AOI22_X1 U16640 ( .A1(n15131), .A2(n15126), .B1(n11631), .B2(n9450), .ZN(
        P3_U3464) );
  AOI22_X1 U16641 ( .A1(n15131), .A2(n15127), .B1(n11637), .B2(n9450), .ZN(
        P3_U3465) );
  AOI22_X1 U16642 ( .A1(n15131), .A2(n15128), .B1(n11641), .B2(n9450), .ZN(
        P3_U3466) );
  AOI22_X1 U16643 ( .A1(n15131), .A2(n15129), .B1(n11647), .B2(n9450), .ZN(
        P3_U3467) );
  AOI22_X1 U16644 ( .A1(n15131), .A2(n15130), .B1(n11657), .B2(n9450), .ZN(
        P3_U3469) );
  AOI21_X1 U16645 ( .B1(n15134), .B2(n15133), .A(n15132), .ZN(SUB_1596_U59) );
  OAI21_X1 U16646 ( .B1(n15137), .B2(n15136), .A(n15135), .ZN(SUB_1596_U58) );
  XOR2_X1 U16647 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15138), .Z(SUB_1596_U53) );
  OAI21_X1 U16648 ( .B1(n15141), .B2(n15140), .A(n15139), .ZN(SUB_1596_U56) );
  AOI21_X1 U16649 ( .B1(n15144), .B2(n15143), .A(n15142), .ZN(n15145) );
  XOR2_X1 U16650 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n15145), .Z(SUB_1596_U60) );
  AOI21_X1 U16651 ( .B1(n15148), .B2(n15147), .A(n15146), .ZN(SUB_1596_U5) );
  OR2_X1 U7448 ( .A1(n12337), .A2(n10898), .ZN(n12534) );
  NAND2_X1 U9061 ( .A1(n11520), .A2(n13746), .ZN(n11854) );
  CLKBUF_X1 U7221 ( .A(n7596), .Z(n6645) );
  CLKBUF_X1 U7264 ( .A(n8712), .Z(n8717) );
  CLKBUF_X3 U7297 ( .A(n8278), .Z(n9453) );
  CLKBUF_X1 U7320 ( .A(n8682), .Z(n9666) );
  CLKBUF_X1 U7666 ( .A(n7955), .Z(n12818) );
  CLKBUF_X1 U8083 ( .A(n9114), .Z(n6483) );
endmodule

