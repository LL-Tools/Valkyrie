

module b15_C_SARLock_k_64_2 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, U3445, U3446, U3447, U3448, U3213, U3212, 
        U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, 
        U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, 
        U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, 
        U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, 
        U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, 
        U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, 
        U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, 
        U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, 
        U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, 
        U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, 
        U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, 
        U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, 
        U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, 
        U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, 
        U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, 
        U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, 
        U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, 
        U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, 
        U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, 
        U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, 
        U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, 
        U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, 
        U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, 
        U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, 
        U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, 
        U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, 
        U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, 
        U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, 
        U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, 
        U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, 
        U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, 
        U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, 
        U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, 
        U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, 
        U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, 
        U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, 
        U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, 
        U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, 
        U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, 
        U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, 
        U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, 
        U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, 
        U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, 
        U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, 
        U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687;

  INV_X1 U3426 ( .A(n3499), .ZN(n5508) );
  AOI21_X1 U3427 ( .B1(n3566), .B2(n3522), .A(n3420), .ZN(n6032) );
  NAND2_X1 U3428 ( .A1(n4383), .A2(n3371), .ZN(n3541) );
  CLKBUF_X2 U3429 ( .A(n3156), .Z(n4027) );
  AND2_X1 U3430 ( .A1(n3317), .A2(n3316), .ZN(n4346) );
  CLKBUF_X2 U3431 ( .A(n3254), .Z(n4407) );
  NAND2_X1 U3432 ( .A1(n2993), .A2(n2983), .ZN(n4411) );
  NAND4_X2 U3433 ( .A1(n3170), .A2(n3169), .A3(n3168), .A4(n3167), .ZN(n4434)
         );
  AND2_X1 U3434 ( .A1(n3122), .A2(n4660), .ZN(n3282) );
  NOR2_X2 U3435 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4670) );
  CLKBUF_X1 U3436 ( .A(n4065), .Z(n2977) );
  NOR2_X1 U3437 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4065) );
  AND2_X1 U3439 ( .A1(n3121), .A2(n4660), .ZN(n2980) );
  NAND2_X1 U3440 ( .A1(n3338), .A2(n3337), .ZN(n3392) );
  NAND2_X1 U3441 ( .A1(n3563), .A2(n4407), .ZN(n4843) );
  NOR2_X1 U3442 ( .A1(n4407), .A2(n4852), .ZN(n4831) );
  INV_X2 U3443 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3114) );
  INV_X2 U3444 ( .A(n5181), .ZN(n5073) );
  AND2_X1 U34450 ( .A1(n4404), .A2(n4405), .ZN(n3587) );
  NAND2_X1 U34460 ( .A1(n4226), .A2(n4434), .ZN(n3253) );
  CLKBUF_X3 U34470 ( .A(n3568), .Z(n5521) );
  AND4_X1 U34480 ( .A1(n3155), .A2(n3154), .A3(n3153), .A4(n3152), .ZN(n3167)
         );
  INV_X1 U3449 ( .A(n5826), .ZN(n5802) );
  INV_X1 U3450 ( .A(n5889), .ZN(n5870) );
  INV_X1 U34510 ( .A(n4849), .ZN(n4325) );
  NOR2_X1 U34520 ( .A1(n3078), .A2(n3076), .ZN(n5251) );
  AND4_X1 U3454 ( .A1(n3135), .A2(n3134), .A3(n3133), .A4(n3132), .ZN(n2978)
         );
  OAI21_X2 U34550 ( .B1(n5295), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n3033), .ZN(n3034) );
  AND2_X4 U34560 ( .A1(n4341), .A2(n4657), .ZN(n3877) );
  AND2_X4 U3457 ( .A1(n4670), .A2(n4660), .ZN(n3302) );
  AND2_X4 U3458 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4660) );
  AND2_X4 U34590 ( .A1(n3115), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3121) );
  AND2_X1 U34600 ( .A1(n3026), .A2(n3027), .ZN(n4483) );
  CLKBUF_X2 U34610 ( .A(n6001), .Z(n6009) );
  XNOR2_X1 U34620 ( .A(n3393), .B(n3392), .ZN(n3568) );
  INV_X1 U34630 ( .A(n3165), .ZN(n4381) );
  INV_X2 U34640 ( .A(n3239), .ZN(n4226) );
  NAND4_X1 U34650 ( .A1(n3237), .A2(n3236), .A3(n3235), .A4(n3234), .ZN(n3254)
         );
  CLKBUF_X2 U3466 ( .A(n3877), .Z(n3971) );
  BUF_X2 U3467 ( .A(n4026), .Z(n3993) );
  CLKBUF_X2 U34680 ( .A(n3225), .Z(n3855) );
  BUF_X2 U34690 ( .A(n3841), .Z(n3893) );
  BUF_X2 U34700 ( .A(n3352), .Z(n4018) );
  BUF_X2 U34710 ( .A(n3673), .Z(n3888) );
  CLKBUF_X2 U34720 ( .A(n3300), .Z(n4039) );
  CLKBUF_X2 U34730 ( .A(n3203), .Z(n4046) );
  BUF_X2 U34740 ( .A(n3136), .Z(n4040) );
  AOI21_X1 U3475 ( .B1(n5069), .B2(n5067), .A(n5068), .ZN(n5268) );
  NOR2_X1 U3476 ( .A1(n5270), .A2(n3081), .ZN(n3078) );
  OR3_X1 U3477 ( .A1(n5270), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .A3(n5286), 
        .ZN(n5277) );
  INV_X1 U3478 ( .A(n3042), .ZN(n5680) );
  NAND2_X1 U3479 ( .A1(n3102), .A2(n3101), .ZN(n5373) );
  INV_X1 U3480 ( .A(n4822), .ZN(n3023) );
  AND2_X1 U3481 ( .A1(n3618), .A2(n2986), .ZN(n3022) );
  NAND2_X1 U3482 ( .A1(n4255), .A2(n5511), .ZN(n5737) );
  NAND2_X1 U3483 ( .A1(n3073), .A2(n4363), .ZN(n3442) );
  AND2_X2 U3484 ( .A1(n3415), .A2(n3414), .ZN(n3566) );
  AND2_X1 U3485 ( .A1(n4246), .A2(n6370), .ZN(n5484) );
  NAND2_X1 U3486 ( .A1(n3383), .A2(n3382), .ZN(n4363) );
  CLKBUF_X1 U3487 ( .A(n4357), .Z(n6143) );
  OR2_X1 U3488 ( .A1(n4120), .A2(n4119), .ZN(n4246) );
  NAND2_X1 U3489 ( .A1(n4379), .A2(n4827), .ZN(n4830) );
  NAND2_X2 U3490 ( .A1(n3560), .A2(n3559), .ZN(n4379) );
  NAND2_X1 U3491 ( .A1(n3330), .A2(n3329), .ZN(n3341) );
  NOR2_X1 U3492 ( .A1(n3258), .A2(n4232), .ZN(n3565) );
  INV_X1 U3493 ( .A(n3025), .ZN(n3024) );
  INV_X1 U3494 ( .A(n4106), .ZN(n3256) );
  NOR2_X1 U3495 ( .A1(n4344), .A2(n5028), .ZN(n4227) );
  AND2_X1 U3496 ( .A1(n3238), .A2(n4343), .ZN(n3265) );
  OAI21_X1 U3497 ( .B1(n3249), .B2(n3114), .A(n3252), .ZN(n3025) );
  OAI211_X1 U3498 ( .C1(n3193), .C2(n3192), .A(n3191), .B(n3190), .ZN(n3322)
         );
  NAND2_X1 U3499 ( .A1(n3319), .A2(n4831), .ZN(n4344) );
  AND2_X2 U3500 ( .A1(n4407), .A2(n4852), .ZN(n4849) );
  NAND2_X1 U3501 ( .A1(n4226), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4383) );
  AND2_X1 U3502 ( .A1(n4852), .A2(n4103), .ZN(n3385) );
  AND3_X2 U3503 ( .A1(n4852), .A2(STATE2_REG_0__SCAN_IN), .A3(n3239), .ZN(
        n3552) );
  OR2_X1 U3504 ( .A1(n3281), .A2(n3280), .ZN(n3405) );
  NAND2_X1 U3505 ( .A1(n3243), .A2(n3260), .ZN(n4382) );
  NAND2_X1 U3506 ( .A1(n3254), .A2(n4411), .ZN(n4218) );
  INV_X1 U3507 ( .A(n3254), .ZN(n4103) );
  NAND2_X1 U3508 ( .A1(n2994), .A2(n2978), .ZN(n3165) );
  OR2_X1 U3509 ( .A1(n3293), .A2(n3292), .ZN(n3489) );
  CLKBUF_X1 U3510 ( .A(n3260), .Z(n3261) );
  NAND2_X1 U3511 ( .A1(n3147), .A2(n3146), .ZN(n3260) );
  AND3_X1 U3512 ( .A1(n3210), .A2(n3209), .A3(n3208), .ZN(n3216) );
  AND4_X1 U3513 ( .A1(n3224), .A2(n3223), .A3(n3222), .A4(n3221), .ZN(n3236)
         );
  AND4_X1 U3514 ( .A1(n3233), .A2(n3232), .A3(n3231), .A4(n3230), .ZN(n3234)
         );
  AND4_X1 U3515 ( .A1(n3197), .A2(n3196), .A3(n3195), .A4(n3194), .ZN(n3210)
         );
  AND4_X1 U3516 ( .A1(n3207), .A2(n3206), .A3(n3205), .A4(n3204), .ZN(n3208)
         );
  AND4_X1 U3517 ( .A1(n3201), .A2(n3200), .A3(n3199), .A4(n3198), .ZN(n3209)
         );
  AND4_X1 U3518 ( .A1(n3160), .A2(n3159), .A3(n3158), .A4(n3157), .ZN(n3168)
         );
  AND4_X1 U3519 ( .A1(n3164), .A2(n3163), .A3(n3162), .A4(n3161), .ZN(n3169)
         );
  AND4_X1 U3520 ( .A1(n3126), .A2(n3125), .A3(n3124), .A4(n3123), .ZN(n3127)
         );
  AND4_X1 U3521 ( .A1(n3229), .A2(n3228), .A3(n3227), .A4(n3226), .ZN(n3235)
         );
  AND4_X1 U3522 ( .A1(n3220), .A2(n3219), .A3(n3218), .A4(n3217), .ZN(n3237)
         );
  AND4_X1 U3523 ( .A1(n3151), .A2(n3150), .A3(n3149), .A4(n3148), .ZN(n3170)
         );
  AND4_X1 U3524 ( .A1(n3140), .A2(n3139), .A3(n3138), .A4(n3137), .ZN(n3147)
         );
  INV_X2 U3525 ( .A(n6043), .ZN(n6035) );
  AND4_X1 U3526 ( .A1(n3145), .A2(n3144), .A3(n3143), .A4(n3142), .ZN(n3146)
         );
  BUF_X2 U3527 ( .A(n3141), .Z(n4021) );
  BUF_X2 U3528 ( .A(n3179), .Z(n4019) );
  BUF_X2 U3529 ( .A(n3282), .Z(n3836) );
  AND2_X2 U3530 ( .A1(n3041), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4341)
         );
  AND2_X1 U3531 ( .A1(n3116), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3122)
         );
  INV_X2 U3532 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3115) );
  NOR2_X2 U3533 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4656) );
  OAI21_X2 U3534 ( .B1(n3035), .B2(n3038), .A(n3411), .ZN(n6031) );
  AND2_X1 U3535 ( .A1(n5117), .A2(n5204), .ZN(n5192) );
  NOR2_X2 U3536 ( .A1(n5211), .A2(n5116), .ZN(n5117) );
  NOR2_X2 U3537 ( .A1(n5465), .A2(n4258), .ZN(n5695) );
  AND2_X1 U3538 ( .A1(n3121), .A2(n4660), .ZN(n2979) );
  AND2_X1 U3539 ( .A1(n3121), .A2(n4660), .ZN(n3202) );
  AND2_X1 U3540 ( .A1(n3103), .A2(n3003), .ZN(n3101) );
  NAND2_X1 U3541 ( .A1(n3166), .A2(n3165), .ZN(n3191) );
  NAND2_X1 U3542 ( .A1(n3061), .A2(n3462), .ZN(n3474) );
  INV_X1 U3543 ( .A(n3460), .ZN(n3061) );
  AOI22_X1 U3544 ( .A1(n3541), .A2(n3475), .B1(n3552), .B2(
        INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3461) );
  OR2_X1 U3545 ( .A1(n3436), .A2(n3435), .ZN(n3476) );
  NAND2_X1 U3546 ( .A1(n4121), .A2(n3058), .ZN(n4343) );
  INV_X1 U3547 ( .A(n4218), .ZN(n3058) );
  AND2_X1 U3548 ( .A1(n5085), .A2(n5154), .ZN(n3069) );
  INV_X1 U3549 ( .A(n5672), .ZN(n3081) );
  OAI21_X1 U3550 ( .B1(n3086), .B2(n3084), .A(n2999), .ZN(n3083) );
  INV_X1 U3551 ( .A(n3507), .ZN(n3084) );
  OAI21_X1 U3552 ( .B1(n3576), .B2(n3021), .A(n3019), .ZN(n3389) );
  NAND2_X1 U3553 ( .A1(n3402), .A2(n6509), .ZN(n3021) );
  AOI21_X1 U3554 ( .B1(n3020), .B2(n3402), .A(n2997), .ZN(n3019) );
  OR2_X1 U3555 ( .A1(n3389), .A2(n3388), .ZN(n3391) );
  OAI21_X1 U3556 ( .B1(n3576), .B2(STATE2_REG_0__SCAN_IN), .A(n3401), .ZN(
        n3399) );
  AND2_X2 U3557 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4657) );
  NOR2_X1 U3558 ( .A1(n4090), .A2(n3063), .ZN(n3062) );
  INV_X1 U3559 ( .A(n3065), .ZN(n3063) );
  OR2_X1 U3560 ( .A1(n2991), .A2(n5147), .ZN(n5149) );
  INV_X1 U3561 ( .A(n4086), .ZN(n4085) );
  NAND2_X1 U3562 ( .A1(n3092), .A2(n3091), .ZN(n5352) );
  AOI21_X1 U3563 ( .B1(n2982), .B2(n3095), .A(n3008), .ZN(n3091) );
  AND2_X1 U3564 ( .A1(n3094), .A2(n3093), .ZN(n2982) );
  NAND2_X1 U3565 ( .A1(n3105), .A2(n3106), .ZN(n3104) );
  INV_X1 U3566 ( .A(n5392), .ZN(n3105) );
  NAND2_X1 U3567 ( .A1(n3411), .A2(n3039), .ZN(n3038) );
  INV_X1 U3568 ( .A(n3442), .ZN(n3445) );
  NAND2_X1 U3569 ( .A1(n3060), .A2(n3059), .ZN(n3492) );
  INV_X1 U3570 ( .A(n3473), .ZN(n3059) );
  INV_X1 U3571 ( .A(n3474), .ZN(n3060) );
  OR2_X1 U3572 ( .A1(n3472), .A2(n3471), .ZN(n3485) );
  OR2_X1 U3573 ( .A1(n3455), .A2(n3454), .ZN(n3475) );
  OR2_X1 U3574 ( .A1(n3312), .A2(n3311), .ZN(n3394) );
  INV_X1 U3575 ( .A(n3394), .ZN(n3336) );
  AOI22_X1 U3576 ( .A1(n3141), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3132) );
  AOI21_X1 U3577 ( .B1(n6201), .B2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n3524), 
        .ZN(n3523) );
  AOI21_X1 U3578 ( .B1(n3248), .B2(n4411), .A(n4388), .ZN(n3190) );
  AND2_X1 U3579 ( .A1(n3066), .A2(n5160), .ZN(n3065) );
  INV_X1 U3580 ( .A(n3876), .ZN(n3066) );
  INV_X1 U3581 ( .A(n5167), .ZN(n3064) );
  AND2_X1 U3582 ( .A1(n6367), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4062) );
  AND2_X2 U3583 ( .A1(n5192), .A2(n5193), .ZN(n3785) );
  INV_X1 U3584 ( .A(n4763), .ZN(n3617) );
  INV_X1 U3585 ( .A(n2977), .ZN(n4057) );
  INV_X1 U3586 ( .A(n4374), .ZN(n3027) );
  NOR2_X1 U3587 ( .A1(n3261), .A2(n6210), .ZN(n3745) );
  INV_X1 U3588 ( .A(n3745), .ZN(n3716) );
  INV_X1 U3589 ( .A(n3079), .ZN(n3076) );
  AOI21_X1 U3590 ( .B1(n5672), .B2(n3080), .A(n3014), .ZN(n3079) );
  INV_X1 U3591 ( .A(n3513), .ZN(n3080) );
  NOR2_X1 U3592 ( .A1(n5686), .A2(n5678), .ZN(n3508) );
  NAND2_X1 U3593 ( .A1(n3047), .A2(n5194), .ZN(n3046) );
  INV_X1 U3594 ( .A(n5119), .ZN(n3047) );
  AOI21_X1 U3595 ( .B1(n3089), .B2(n3087), .A(n3000), .ZN(n3086) );
  INV_X1 U3596 ( .A(n3503), .ZN(n3087) );
  INV_X1 U3597 ( .A(n5201), .ZN(n3048) );
  INV_X1 U3598 ( .A(n5382), .ZN(n3106) );
  NAND2_X1 U3599 ( .A1(n4849), .A2(n5073), .ZN(n4208) );
  NOR2_X1 U3600 ( .A1(n3053), .A2(n3052), .ZN(n3051) );
  INV_X1 U3601 ( .A(n4760), .ZN(n3052) );
  INV_X1 U3602 ( .A(n4514), .ZN(n3050) );
  NAND2_X1 U3603 ( .A1(n4485), .A2(n3054), .ZN(n3053) );
  INV_X1 U3604 ( .A(n4398), .ZN(n3054) );
  OAI22_X1 U3605 ( .A1(n3597), .A2(n3040), .B1(n3439), .B2(n3262), .ZN(n3440)
         );
  AND2_X1 U3606 ( .A1(n3318), .A2(n4381), .ZN(n3319) );
  AND2_X1 U3607 ( .A1(n4332), .A2(n4116), .ZN(n4117) );
  INV_X1 U3608 ( .A(n4779), .ZN(n4601) );
  AOI22_X1 U3609 ( .A1(n3202), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3203), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3129) );
  AOI22_X1 U3610 ( .A1(n3156), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3130) );
  OAI21_X1 U3611 ( .B1(n6408), .B2(n4693), .A(n6395), .ZN(n4368) );
  AND2_X1 U3612 ( .A1(n6511), .A2(n4840), .ZN(n5034) );
  INV_X2 U3613 ( .A(n4060), .ZN(n4067) );
  AND2_X1 U3614 ( .A1(n3069), .A2(n3068), .ZN(n3067) );
  INV_X1 U3615 ( .A(n5144), .ZN(n3068) );
  NAND2_X1 U3616 ( .A1(n5096), .A2(n3069), .ZN(n5145) );
  NAND2_X1 U3617 ( .A1(n5096), .A2(n5154), .ZN(n5153) );
  NOR2_X1 U3618 ( .A1(n3748), .A2(n5814), .ZN(n3780) );
  NAND2_X1 U3619 ( .A1(n3005), .A2(n3718), .ZN(n5211) );
  NAND2_X1 U3620 ( .A1(n3618), .A2(n3617), .ZN(n4821) );
  NOR2_X1 U3621 ( .A1(n4922), .A2(n3611), .ZN(n3612) );
  OR3_X1 U3622 ( .A1(n3056), .A2(n3016), .A3(n5087), .ZN(n3055) );
  NOR2_X1 U3623 ( .A1(n5686), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5304)
         );
  AND2_X1 U3624 ( .A1(n5313), .A2(n3007), .ZN(n3029) );
  NOR2_X1 U3625 ( .A1(n2990), .A2(n5655), .ZN(n5176) );
  NAND2_X1 U3626 ( .A1(n5508), .A2(n3097), .ZN(n3096) );
  NAND2_X1 U3627 ( .A1(n5365), .A2(n3098), .ZN(n3097) );
  NOR2_X1 U3628 ( .A1(n5508), .A2(n3018), .ZN(n3095) );
  INV_X1 U3629 ( .A(n5375), .ZN(n3498) );
  INV_X1 U3630 ( .A(n3500), .ZN(n5507) );
  OR2_X1 U3631 ( .A1(n4908), .A2(n4907), .ZN(n4932) );
  NAND2_X1 U3632 ( .A1(n3112), .A2(n3106), .ZN(n3103) );
  AND2_X1 U3633 ( .A1(n3481), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3482)
         );
  AND2_X1 U3634 ( .A1(n6367), .A2(n4231), .ZN(n4658) );
  AND3_X1 U3635 ( .A1(n3266), .A2(n3265), .A3(n3264), .ZN(n3267) );
  NAND2_X1 U3636 ( .A1(n3391), .A2(n3390), .ZN(n3393) );
  NOR2_X1 U3637 ( .A1(n3749), .A2(n3165), .ZN(n6367) );
  INV_X1 U3638 ( .A(n4529), .ZN(n6203) );
  INV_X1 U3639 ( .A(n4869), .ZN(n6205) );
  OR2_X1 U3640 ( .A1(n3402), .A2(n3401), .ZN(n3403) );
  NAND2_X1 U3641 ( .A1(n6509), .A2(n4368), .ZN(n4779) );
  AND4_X1 U3642 ( .A1(n3214), .A2(n3213), .A3(n3212), .A4(n3211), .ZN(n3215)
         );
  NAND2_X1 U3643 ( .A1(n3877), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3211)
         );
  AND2_X1 U3644 ( .A1(n6488), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3561) );
  OR2_X1 U3645 ( .A1(n5034), .A2(n6210), .ZN(n5038) );
  INV_X1 U3646 ( .A(n5591), .ZN(n5223) );
  INV_X1 U3647 ( .A(n5242), .ZN(n5249) );
  CLKBUF_X1 U3648 ( .A(n4358), .Z(n5526) );
  AND2_X1 U3649 ( .A1(n3541), .A2(n3540), .ZN(n3543) );
  NAND2_X1 U3650 ( .A1(n3520), .A2(n3519), .ZN(n3539) );
  XNOR2_X1 U3651 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3538) );
  AND2_X1 U3652 ( .A1(n6287), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3529)
         );
  XNOR2_X1 U3653 ( .A(n4680), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3526)
         );
  BUF_X1 U3654 ( .A(n3202), .Z(n3992) );
  INV_X1 U3655 ( .A(n3401), .ZN(n3020) );
  INV_X1 U3656 ( .A(n4078), .ZN(n3347) );
  OR2_X1 U3657 ( .A1(n3248), .A2(n3262), .ZN(n4106) );
  AOI22_X1 U3658 ( .A1(n3179), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        INSTQUEUE_REG_13__6__SCAN_IN), .B2(n3877), .ZN(n3145) );
  OR2_X1 U3659 ( .A1(n5168), .A2(n5309), .ZN(n3876) );
  NOR2_X1 U3660 ( .A1(n5185), .A2(n5179), .ZN(n3072) );
  NAND2_X1 U3661 ( .A1(n3733), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3748)
         );
  NOR2_X1 U3662 ( .A1(n3639), .A2(n3635), .ZN(n3656) );
  NAND2_X1 U3663 ( .A1(n3634), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3639)
         );
  INV_X1 U3664 ( .A(n3633), .ZN(n3634) );
  NAND2_X1 U3665 ( .A1(n3567), .A2(n3760), .ZN(n3586) );
  AND2_X1 U3666 ( .A1(n3569), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3591) );
  NAND2_X1 U3667 ( .A1(n3057), .A2(n5155), .ZN(n3056) );
  INV_X1 U3668 ( .A(n5165), .ZN(n3057) );
  INV_X1 U3669 ( .A(n5357), .ZN(n3093) );
  OR2_X1 U3670 ( .A1(n3095), .A2(n3096), .ZN(n3094) );
  INV_X1 U3671 ( .A(n3492), .ZN(n3483) );
  OAI22_X1 U3672 ( .A1(n3607), .A2(n3040), .B1(n3458), .B2(n3262), .ZN(n3459)
         );
  NAND2_X1 U3673 ( .A1(n3552), .A2(n3248), .ZN(n3249) );
  AND2_X1 U3674 ( .A1(n4382), .A2(n3320), .ZN(n3241) );
  NAND2_X1 U3675 ( .A1(n3563), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3371) );
  OR2_X1 U3676 ( .A1(n3362), .A2(n3361), .ZN(n3416) );
  OR2_X1 U3677 ( .A1(n4383), .A2(n3336), .ZN(n3337) );
  INV_X1 U3678 ( .A(n3414), .ZN(n3073) );
  OR2_X1 U3679 ( .A1(n3248), .A2(n3562), .ZN(n3749) );
  NAND2_X1 U3680 ( .A1(n3352), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3213)
         );
  NAND2_X1 U3681 ( .A1(n3179), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3212) );
  AOI22_X1 U3682 ( .A1(n3202), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3301), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3175) );
  AOI22_X1 U3683 ( .A1(n3141), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3673), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3124) );
  INV_X1 U3684 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6589) );
  INV_X1 U3685 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6373) );
  AOI221_X1 U3686 ( .B1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n3523), .C1(
        n5758), .C2(n3523), .A(n3521), .ZN(n4112) );
  NOR2_X1 U3687 ( .A1(n5149), .A2(n5071), .ZN(n5055) );
  INV_X1 U3688 ( .A(n3851), .ZN(n3870) );
  AND2_X1 U3689 ( .A1(n3702), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3719)
         );
  INV_X1 U3690 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4922) );
  AND2_X1 U3691 ( .A1(n4155), .A2(n4154), .ZN(n4907) );
  INV_X1 U3692 ( .A(n6400), .ZN(n4827) );
  AND2_X1 U3693 ( .A1(n4304), .A2(n4324), .ZN(n5920) );
  NAND2_X1 U3694 ( .A1(n6011), .A2(n4303), .ZN(n4304) );
  OR2_X1 U3695 ( .A1(n4830), .A2(n4353), .ZN(n4303) );
  INV_X1 U3696 ( .A(n3760), .ZN(n4066) );
  NAND2_X1 U3697 ( .A1(n4013), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4076)
         );
  NOR2_X2 U3698 ( .A1(n5067), .A2(n5069), .ZN(n5068) );
  AND2_X1 U3699 ( .A1(n3944), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3945)
         );
  NAND2_X1 U3700 ( .A1(n3945), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3963)
         );
  AND2_X1 U3701 ( .A1(n3910), .A2(n3909), .ZN(n5160) );
  NAND3_X1 U3702 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_21__SCAN_IN), .A3(n3870), .ZN(n3873) );
  NOR2_X1 U3703 ( .A1(n3873), .A2(n6634), .ZN(n3906) );
  NOR2_X1 U3705 ( .A1(n3801), .A2(n5327), .ZN(n3802) );
  AND2_X1 U3706 ( .A1(n3785), .A2(n3072), .ZN(n5652) );
  AND2_X1 U3707 ( .A1(n3780), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3781)
         );
  NAND2_X1 U3708 ( .A1(n3781), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3801)
         );
  NAND2_X1 U3709 ( .A1(n3785), .A2(n3784), .ZN(n5187) );
  OR2_X1 U3710 ( .A1(n5804), .A2(n4057), .ZN(n3765) );
  CLKBUF_X1 U3711 ( .A(n5192), .Z(n5202) );
  AND2_X1 U3712 ( .A1(n3698), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3702)
         );
  INV_X1 U3713 ( .A(n4931), .ZN(n3028) );
  OR2_X1 U3714 ( .A1(n4931), .A2(n5002), .ZN(n5247) );
  AOI21_X1 U3715 ( .B1(n3616), .B2(n3745), .A(n3615), .ZN(n4763) );
  NOR2_X1 U3716 ( .A1(n4510), .A2(n4397), .ZN(n3026) );
  NAND2_X1 U3717 ( .A1(n3602), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3611)
         );
  NOR2_X1 U3718 ( .A1(n4980), .A2(n3592), .ZN(n3602) );
  NAND2_X1 U3719 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3592) );
  NAND2_X1 U3720 ( .A1(n3077), .A2(n3074), .ZN(n5278) );
  NOR2_X1 U3721 ( .A1(n3076), .A2(n3075), .ZN(n3074) );
  INV_X1 U3722 ( .A(n5288), .ZN(n3075) );
  OR2_X1 U3723 ( .A1(n5686), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5286)
         );
  OR2_X1 U3724 ( .A1(n5455), .A2(n4263), .ZN(n5435) );
  NOR3_X1 U3725 ( .A1(n5171), .A2(n3016), .A3(n5165), .ZN(n5156) );
  NOR2_X1 U3726 ( .A1(n5171), .A2(n5165), .ZN(n5164) );
  OR2_X1 U3727 ( .A1(n5472), .A2(n5169), .ZN(n5171) );
  NOR2_X1 U3728 ( .A1(n5700), .A2(n5711), .ZN(n4261) );
  AND2_X1 U3729 ( .A1(n5176), .A2(n4191), .ZN(n5470) );
  NAND2_X1 U3730 ( .A1(n5470), .A2(n5469), .ZN(n5472) );
  NAND2_X1 U3731 ( .A1(n5296), .A2(n4084), .ZN(n3030) );
  OR2_X1 U3732 ( .A1(n6494), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4078) );
  OAI21_X1 U3733 ( .B1(n5343), .B2(n3085), .A(n3082), .ZN(n3042) );
  NAND2_X1 U3734 ( .A1(n3089), .A2(n3507), .ZN(n3085) );
  INV_X1 U3735 ( .A(n3083), .ZN(n3082) );
  AND2_X1 U3736 ( .A1(n4183), .A2(n4182), .ZN(n5655) );
  NAND2_X1 U3737 ( .A1(n3045), .A2(n3044), .ZN(n3043) );
  INV_X1 U3738 ( .A(n3046), .ZN(n3045) );
  INV_X1 U3739 ( .A(n5188), .ZN(n3044) );
  AND2_X1 U3740 ( .A1(n4174), .A2(n4173), .ZN(n5201) );
  NOR3_X1 U3741 ( .A1(n5209), .A2(n3048), .A3(n5119), .ZN(n5198) );
  OR2_X1 U3742 ( .A1(n4348), .A2(n4242), .ZN(n4243) );
  NOR2_X1 U3743 ( .A1(n5209), .A2(n5119), .ZN(n5200) );
  OR2_X1 U3744 ( .A1(n5207), .A2(n5206), .ZN(n5209) );
  AND2_X1 U3745 ( .A1(n5514), .A2(n4163), .ZN(n5516) );
  AND2_X1 U3746 ( .A1(n5513), .A2(n5512), .ZN(n4163) );
  NAND2_X1 U3747 ( .A1(n5516), .A2(n5128), .ZN(n5207) );
  NOR2_X1 U3748 ( .A1(n4932), .A2(n4933), .ZN(n5514) );
  NAND2_X1 U3749 ( .A1(n3050), .A2(n2996), .ZN(n4908) );
  INV_X1 U3750 ( .A(n4825), .ZN(n3049) );
  NAND2_X1 U3751 ( .A1(n3050), .A2(n3051), .ZN(n4824) );
  NOR2_X1 U3752 ( .A1(n4514), .A2(n3053), .ZN(n4761) );
  NOR2_X1 U3753 ( .A1(n4975), .A2(n2998), .ZN(n6025) );
  OR2_X1 U3754 ( .A1(n4512), .A2(n4511), .ZN(n4514) );
  NOR2_X1 U3755 ( .A1(n4514), .A2(n4398), .ZN(n4486) );
  OR2_X1 U3756 ( .A1(n6056), .A2(n4316), .ZN(n4257) );
  NAND2_X1 U3757 ( .A1(n3409), .A2(n4342), .ZN(n3037) );
  NAND2_X1 U3758 ( .A1(n4127), .A2(n5073), .ZN(n4299) );
  INV_X1 U3759 ( .A(n3350), .ZN(n3100) );
  INV_X1 U3760 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4680) );
  OR3_X1 U3761 ( .A1(n4339), .A2(n4828), .A3(n4338), .ZN(n6371) );
  AND2_X1 U3762 ( .A1(n4417), .A2(n4689), .ZN(n4554) );
  AND2_X1 U3763 ( .A1(n3566), .A2(n4445), .ZN(n4737) );
  OAI21_X1 U3764 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6487), .A(n4601), 
        .ZN(n6291) );
  AOI22_X1 U3765 ( .A1(n3225), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3136), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3131) );
  AND2_X1 U3766 ( .A1(n4369), .A2(n4368), .ZN(n4491) );
  INV_X1 U3767 ( .A(n6291), .ZN(n6208) );
  NOR2_X1 U3768 ( .A1(n5790), .A2(n5647), .ZN(n5642) );
  INV_X1 U3769 ( .A(n5890), .ZN(n5876) );
  INV_X1 U3770 ( .A(n5861), .ZN(n5880) );
  OR2_X1 U3771 ( .A1(n5038), .A2(n4854), .ZN(n5826) );
  OR2_X1 U3772 ( .A1(n5038), .A2(n4850), .ZN(n5873) );
  INV_X1 U3773 ( .A(n5212), .ZN(n6519) );
  INV_X1 U3774 ( .A(n5901), .ZN(n6518) );
  NAND2_X1 U3775 ( .A1(n4387), .A2(n4386), .ZN(n5905) );
  OR3_X1 U3776 ( .A1(n4379), .A2(n6400), .A3(n4378), .ZN(n4387) );
  NAND2_X1 U3777 ( .A1(n5905), .A2(n4388), .ZN(n5901) );
  OR2_X1 U3778 ( .A1(n5097), .A2(n5096), .ZN(n5674) );
  OR2_X1 U3779 ( .A1(n5909), .A2(n4836), .ZN(n5242) );
  INV_X1 U3780 ( .A(n5909), .ZN(n5241) );
  OR2_X1 U3781 ( .A1(n4830), .A2(n6391), .ZN(n6011) );
  XNOR2_X1 U3782 ( .A(n4077), .B(n5039), .ZN(n4856) );
  OR2_X1 U3783 ( .A1(n4076), .A2(n5059), .ZN(n4077) );
  AND2_X1 U3784 ( .A1(n5067), .A2(n5146), .ZN(n5591) );
  INV_X1 U3785 ( .A(n5153), .ZN(n5152) );
  INV_X1 U3786 ( .A(n5674), .ZN(n6520) );
  OR2_X1 U3787 ( .A1(n5232), .A2(n6043), .ZN(n4095) );
  CLKBUF_X1 U3788 ( .A(n4865), .Z(n4929) );
  NOR2_X1 U3789 ( .A1(n4821), .A2(n4822), .ZN(n4867) );
  INV_X1 U3790 ( .A(n6040), .ZN(n5395) );
  INV_X1 U3791 ( .A(n6041), .ZN(n6036) );
  OR2_X1 U3792 ( .A1(n6047), .A2(n4075), .ZN(n6040) );
  OR2_X1 U3793 ( .A1(n4830), .A2(n6381), .ZN(n6041) );
  OR2_X1 U3794 ( .A1(n5077), .A2(n5076), .ZN(n5411) );
  XNOR2_X1 U3795 ( .A(n3034), .B(n4089), .ZN(n5445) );
  NOR2_X1 U3796 ( .A1(n4078), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5705) );
  NAND2_X1 U3797 ( .A1(n5343), .A2(n3503), .ZN(n3090) );
  AOI21_X1 U3798 ( .B1(n3500), .B2(n3096), .A(n3095), .ZN(n5359) );
  NAND2_X1 U3799 ( .A1(n3500), .A2(n5365), .ZN(n5506) );
  NAND2_X1 U3800 ( .A1(n3102), .A2(n3103), .ZN(n5381) );
  INV_X1 U3801 ( .A(n5705), .ZN(n6071) );
  NAND2_X1 U3802 ( .A1(n4246), .A2(n4658), .ZN(n6088) );
  AND2_X1 U3803 ( .A1(n4246), .A2(n4229), .ZN(n6100) );
  INV_X1 U3804 ( .A(n5519), .ZN(n6119) );
  INV_X1 U3805 ( .A(n6100), .ZN(n6116) );
  INV_X1 U3806 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6287) );
  NAND2_X1 U3807 ( .A1(n3271), .A2(n3270), .ZN(n3031) );
  INV_X1 U3808 ( .A(n3268), .ZN(n3271) );
  INV_X1 U3809 ( .A(n3574), .ZN(n4696) );
  INV_X1 U3810 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6125) );
  OAI21_X1 U3811 ( .B1(n4687), .B2(n6485), .A(n4779), .ZN(n6124) );
  INV_X1 U3812 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6488) );
  NAND2_X1 U3813 ( .A1(n6487), .A2(n6488), .ZN(n6494) );
  NOR2_X1 U3814 ( .A1(n5753), .A2(n4369), .ZN(n5531) );
  AND2_X1 U3815 ( .A1(n4554), .A2(n4696), .ZN(n4647) );
  NAND2_X1 U3816 ( .A1(n4453), .A2(n4696), .ZN(n5580) );
  INV_X1 U3817 ( .A(n6194), .ZN(n4815) );
  NOR2_X1 U3818 ( .A1(n5974), .A2(n4779), .ZN(n6256) );
  NOR2_X1 U3819 ( .A1(n5978), .A2(n4779), .ZN(n6262) );
  NOR2_X1 U3820 ( .A1(n5980), .A2(n4779), .ZN(n6265) );
  NOR2_X1 U3821 ( .A1(n5982), .A2(n4779), .ZN(n6270) );
  OR2_X1 U3822 ( .A1(n6253), .A2(n6252), .ZN(n6281) );
  NOR2_X1 U3823 ( .A1(n5986), .A2(n4779), .ZN(n6279) );
  INV_X1 U3824 ( .A(n5544), .ZN(n6294) );
  INV_X1 U3825 ( .A(n5552), .ZN(n6314) );
  INV_X1 U3826 ( .A(n5556), .ZN(n6322) );
  INV_X1 U3827 ( .A(n5560), .ZN(n6330) );
  INV_X1 U3828 ( .A(n6361), .ZN(n6345) );
  NOR2_X1 U3829 ( .A1(n5984), .A2(n4779), .ZN(n6350) );
  INV_X1 U3830 ( .A(n5576), .ZN(n6357) );
  OAI211_X1 U3831 ( .C1(n4633), .C2(n6487), .A(n4605), .B(n4604), .ZN(n4630)
         );
  INV_X1 U3832 ( .A(n6341), .ZN(n6354) );
  INV_X1 U3833 ( .A(n6243), .ZN(n6301) );
  INV_X1 U3834 ( .A(n6259), .ZN(n6315) );
  INV_X1 U3835 ( .A(n6262), .ZN(n6323) );
  INV_X1 U3836 ( .A(n6265), .ZN(n6331) );
  INV_X1 U3837 ( .A(n6270), .ZN(n6339) );
  AND2_X1 U3838 ( .A1(n4370), .A2(n4870), .ZN(n4606) );
  OR2_X1 U3839 ( .A1(n4602), .A2(n4529), .ZN(n4645) );
  NAND2_X1 U3840 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n4379), .ZN(n6395) );
  INV_X1 U3841 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6487) );
  NOR2_X1 U3842 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6598), .ZN(n6516) );
  OAI21_X1 U3843 ( .B1(n5343), .B2(n3088), .A(n3086), .ZN(n5323) );
  AND2_X1 U3844 ( .A1(n3064), .A2(n3065), .ZN(n2981) );
  INV_X2 U3845 ( .A(n3385), .ZN(n3262) );
  AND4_X1 U3846 ( .A1(n3175), .A2(n3177), .A3(n3176), .A4(n3171), .ZN(n2983)
         );
  OR3_X1 U3847 ( .A1(n5171), .A2(n3056), .A3(n3016), .ZN(n2984) );
  NAND2_X1 U3848 ( .A1(n3785), .A2(n3011), .ZN(n5175) );
  NAND2_X1 U3849 ( .A1(n5508), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n2985) );
  AND2_X1 U3850 ( .A1(n3617), .A2(n4866), .ZN(n2986) );
  AND2_X1 U3851 ( .A1(n3030), .A2(n3007), .ZN(n2987) );
  AND2_X1 U3852 ( .A1(n3027), .A2(n3596), .ZN(n2988) );
  AND2_X1 U3853 ( .A1(n3071), .A2(n5129), .ZN(n2989) );
  OR3_X1 U3854 ( .A1(n5209), .A2(n3048), .A3(n3043), .ZN(n2990) );
  OR2_X1 U3855 ( .A1(n5171), .A2(n3055), .ZN(n2991) );
  NAND2_X1 U3856 ( .A1(n3492), .A2(n3491), .ZN(n3499) );
  NAND2_X1 U3857 ( .A1(n5673), .A2(n5672), .ZN(n3514) );
  INV_X1 U3858 ( .A(n4510), .ZN(n3596) );
  INV_X1 U3859 ( .A(n4852), .ZN(n3563) );
  NOR2_X1 U3860 ( .A1(n5167), .A2(n3876), .ZN(n5161) );
  AND4_X1 U3861 ( .A1(n3120), .A2(n3119), .A3(n3118), .A4(n3117), .ZN(n2992)
         );
  NAND2_X1 U3862 ( .A1(n5096), .A2(n3067), .ZN(n5067) );
  AND4_X1 U3863 ( .A1(n3173), .A2(n3178), .A3(n3172), .A4(n3174), .ZN(n2993)
         );
  AND4_X1 U3864 ( .A1(n3131), .A2(n3130), .A3(n3129), .A4(n3128), .ZN(n2994)
         );
  AND2_X1 U3865 ( .A1(n3590), .A2(n3442), .ZN(n2995) );
  AND2_X1 U3866 ( .A1(n3051), .A2(n3049), .ZN(n2996) );
  INV_X1 U3867 ( .A(n5175), .ZN(n3835) );
  NOR2_X1 U3868 ( .A1(n4383), .A2(n3299), .ZN(n2997) );
  AND2_X1 U3869 ( .A1(n3426), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n2998)
         );
  NAND2_X1 U3870 ( .A1(n5686), .A2(n3506), .ZN(n2999) );
  NOR2_X1 U3871 ( .A1(n5508), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3000)
         );
  INV_X1 U3872 ( .A(n3089), .ZN(n3088) );
  AND2_X1 U3873 ( .A1(n3002), .A2(n2985), .ZN(n3089) );
  AND2_X1 U3874 ( .A1(n3090), .A2(n2985), .ZN(n3001) );
  OR2_X1 U3875 ( .A1(n5686), .A2(n5742), .ZN(n3002) );
  OR2_X1 U3876 ( .A1(n3497), .A2(n3496), .ZN(n3003) );
  NOR2_X2 U3877 ( .A1(n5909), .A2(n5028), .ZN(n3004) );
  INV_X2 U3878 ( .A(n4218), .ZN(n5181) );
  NAND2_X1 U3879 ( .A1(n4483), .A2(n4482), .ZN(n4481) );
  INV_X1 U3880 ( .A(n3262), .ZN(n6507) );
  AND2_X1 U3881 ( .A1(n3028), .A2(n2989), .ZN(n3005) );
  NOR2_X1 U3882 ( .A1(n5156), .A2(n5100), .ZN(n3006) );
  NAND2_X1 U3883 ( .A1(n5508), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3007) );
  INV_X1 U3884 ( .A(n3260), .ZN(n3575) );
  AND2_X1 U3885 ( .A1(n5686), .A2(n3501), .ZN(n3008) );
  NOR2_X1 U3886 ( .A1(n5391), .A2(n5392), .ZN(n5390) );
  NOR2_X1 U3887 ( .A1(n5390), .A2(n3112), .ZN(n3009) );
  AND2_X1 U3888 ( .A1(n4407), .A2(n4434), .ZN(n3522) );
  AND2_X1 U3889 ( .A1(n5508), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n3010)
         );
  AND2_X1 U3890 ( .A1(n3072), .A2(n5651), .ZN(n3011) );
  AND2_X1 U3891 ( .A1(n5686), .A2(n5678), .ZN(n3012) );
  XOR2_X1 U3892 ( .A(n3438), .B(n3437), .Z(n3013) );
  INV_X2 U3893 ( .A(n5508), .ZN(n5686) );
  AND2_X1 U3894 ( .A1(n5686), .A2(n5694), .ZN(n3014) );
  INV_X1 U3895 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6509) );
  NOR2_X1 U3896 ( .A1(n4931), .A2(n3070), .ZN(n3015) );
  INV_X1 U3897 ( .A(n3071), .ZN(n3070) );
  NOR2_X1 U3898 ( .A1(n5002), .A2(n5246), .ZN(n3071) );
  NAND2_X1 U3899 ( .A1(n5110), .A2(n5099), .ZN(n3016) );
  OR3_X1 U3900 ( .A1(n5209), .A2(n3048), .A3(n3046), .ZN(n3017) );
  AND2_X2 U3901 ( .A1(n3114), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4350)
         );
  AND2_X1 U3902 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3018) );
  INV_X1 U3903 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3098) );
  INV_X1 U3904 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3041) );
  NAND2_X2 U3905 ( .A1(n3031), .A2(n3315), .ZN(n3576) );
  INV_X1 U3906 ( .A(n4865), .ZN(n3655) );
  NAND2_X1 U3907 ( .A1(n3023), .A2(n3022), .ZN(n4865) );
  NAND2_X1 U3908 ( .A1(n3250), .A2(n3249), .ZN(n3331) );
  OAI21_X2 U3909 ( .B1(n3250), .B2(n3114), .A(n3024), .ZN(n3268) );
  INV_X1 U3910 ( .A(n3785), .ZN(n5184) );
  NOR2_X2 U3911 ( .A1(n4091), .A2(n5095), .ZN(n5096) );
  AND2_X2 U3912 ( .A1(n4973), .A2(n4972), .ZN(n4975) );
  AND2_X2 U3913 ( .A1(n3425), .A2(n3424), .ZN(n4973) );
  NAND2_X2 U3914 ( .A1(n3030), .A2(n3029), .ZN(n4086) );
  NOR2_X2 U3915 ( .A1(n4083), .A2(n3012), .ZN(n5296) );
  INV_X1 U3916 ( .A(n3399), .ZN(n3400) );
  NAND2_X1 U3917 ( .A1(n3268), .A2(n3269), .ZN(n3315) );
  NAND2_X1 U3918 ( .A1(n3032), .A2(n4096), .ZN(U2962) );
  NAND2_X1 U3919 ( .A1(n5445), .A2(n6036), .ZN(n3032) );
  OR2_X2 U3920 ( .A1(n5303), .A2(n4088), .ZN(n3033) );
  OAI21_X1 U3921 ( .B1(n3397), .B2(n3568), .A(n3037), .ZN(n3035) );
  AND2_X1 U3922 ( .A1(n3037), .A2(n3411), .ZN(n4315) );
  NAND2_X1 U3923 ( .A1(n3036), .A2(n3398), .ZN(n4314) );
  NAND2_X1 U3924 ( .A1(n3568), .A2(n3522), .ZN(n3036) );
  NAND2_X1 U3925 ( .A1(n3398), .A2(n3040), .ZN(n3039) );
  INV_X1 U3926 ( .A(n3522), .ZN(n3040) );
  AOI21_X2 U3927 ( .B1(n5352), .B2(n5351), .A(n3110), .ZN(n5343) );
  AOI21_X2 U3928 ( .B1(n5373), .B2(n3498), .A(n3010), .ZN(n3500) );
  OR2_X2 U3929 ( .A1(n5391), .A2(n3104), .ZN(n3102) );
  NOR2_X2 U3930 ( .A1(n4943), .A2(n3482), .ZN(n5391) );
  AND2_X1 U3931 ( .A1(n4660), .A2(n4657), .ZN(n3301) );
  AND2_X2 U3932 ( .A1(n4656), .A2(n4657), .ZN(n3136) );
  AND2_X2 U3933 ( .A1(n4350), .A2(n4657), .ZN(n3352) );
  OAI22_X2 U3934 ( .A1(n4358), .A2(STATE2_REG_0__SCAN_IN), .B1(n3384), .B2(
        n4383), .ZN(n3365) );
  NAND2_X2 U3935 ( .A1(n3366), .A2(n3351), .ZN(n4358) );
  NAND2_X1 U3936 ( .A1(n3064), .A2(n3062), .ZN(n4091) );
  NAND3_X1 U3937 ( .A1(n3442), .A2(n3590), .A3(n3522), .ZN(n3387) );
  NAND2_X1 U3938 ( .A1(n3413), .A2(n3412), .ZN(n3414) );
  NAND2_X1 U3939 ( .A1(n5270), .A2(n3513), .ZN(n5673) );
  INV_X1 U3940 ( .A(n3078), .ZN(n3077) );
  NAND2_X1 U3941 ( .A1(n3500), .A2(n2982), .ZN(n3092) );
  NAND2_X1 U3942 ( .A1(n3342), .A2(n3341), .ZN(n3099) );
  NAND2_X2 U3943 ( .A1(n3099), .A2(n3350), .ZN(n3366) );
  NAND3_X1 U3944 ( .A1(n3342), .A2(n3341), .A3(n3100), .ZN(n3351) );
  NAND2_X1 U3945 ( .A1(n3835), .A2(n3111), .ZN(n5167) );
  AND2_X1 U3946 ( .A1(n5521), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6204) );
  INV_X1 U3947 ( .A(n4481), .ZN(n3618) );
  NAND2_X1 U3948 ( .A1(n4086), .A2(n4087), .ZN(n5303) );
  AOI22_X1 U3949 ( .A1(n3673), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3352), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3142) );
  AND2_X2 U3950 ( .A1(n4341), .A2(n3122), .ZN(n3225) );
  AOI22_X1 U3951 ( .A1(n3225), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3136), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3126) );
  AND2_X1 U3952 ( .A1(n4276), .A2(n4407), .ZN(n6370) );
  XNOR2_X1 U3953 ( .A(n5068), .B(n5049), .ZN(n5259) );
  INV_X1 U3954 ( .A(n3315), .ZN(n3340) );
  XNOR2_X1 U3955 ( .A(n3460), .B(n3461), .ZN(n3607) );
  AND2_X2 U3956 ( .A1(n4350), .A2(n4670), .ZN(n3673) );
  OR2_X1 U3957 ( .A1(n3413), .A2(n3412), .ZN(n3415) );
  NAND2_X1 U3958 ( .A1(n3322), .A2(n4831), .ZN(n3255) );
  AND2_X1 U3959 ( .A1(n5312), .A2(n5168), .ZN(n3107) );
  OR2_X1 U3960 ( .A1(n3563), .A2(n4381), .ZN(n3108) );
  NOR2_X1 U3961 ( .A1(n6140), .A2(n4416), .ZN(n3109) );
  AND2_X1 U3962 ( .A1(n5686), .A2(n3502), .ZN(n3110) );
  INV_X1 U3963 ( .A(n3577), .ZN(n4060) );
  NOR2_X1 U3964 ( .A1(n3320), .A2(n6210), .ZN(n3577) );
  INV_X1 U3965 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5758) );
  INV_X1 U3966 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3496) );
  AND2_X1 U3967 ( .A1(n3834), .A2(n3833), .ZN(n3111) );
  INV_X1 U3968 ( .A(n4930), .ZN(n3654) );
  AND3_X2 U3969 ( .A1(n4834), .A2(n6007), .A3(n4833), .ZN(n5909) );
  AND2_X1 U3970 ( .A1(n3488), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3112)
         );
  AND2_X2 U3971 ( .A1(n6041), .A2(n4072), .ZN(n6047) );
  AND2_X1 U3972 ( .A1(n3459), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3113)
         );
  OR2_X1 U3973 ( .A1(n4831), .A2(n3531), .ZN(n3542) );
  INV_X1 U3974 ( .A(n3416), .ZN(n3384) );
  INV_X1 U3975 ( .A(n3561), .ZN(n3346) );
  AOI22_X1 U3976 ( .A1(n3539), .A2(n3538), .B1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n6589), .ZN(n3525) );
  INV_X1 U3977 ( .A(n3269), .ZN(n3270) );
  AND2_X1 U3978 ( .A1(n3391), .A2(n3392), .ZN(n3412) );
  NOR2_X1 U3979 ( .A1(n3525), .A2(n3526), .ZN(n3524) );
  NAND2_X1 U3980 ( .A1(n3566), .A2(n3745), .ZN(n3567) );
  AOI22_X1 U3981 ( .A1(n3541), .A2(n3476), .B1(INSTQUEUE_REG_0__4__SCAN_IN), 
        .B2(n3552), .ZN(n3443) );
  OR2_X1 U3982 ( .A1(n3328), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3329)
         );
  OR2_X1 U3983 ( .A1(n3381), .A2(n3380), .ZN(n3437) );
  NOR2_X1 U3984 ( .A1(n4012), .A2(n4011), .ZN(n4013) );
  INV_X1 U3985 ( .A(n4062), .ZN(n4036) );
  AND2_X1 U3986 ( .A1(PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n3719), .ZN(n3733)
         );
  AOI22_X1 U3987 ( .A1(n3541), .A2(n3485), .B1(INSTQUEUE_REG_0__6__SCAN_IN), 
        .B2(n3552), .ZN(n3473) );
  AND2_X1 U3988 ( .A1(n4193), .A2(n4192), .ZN(n5469) );
  NOR2_X1 U3989 ( .A1(n3490), .A2(n4383), .ZN(n3491) );
  AND2_X1 U3990 ( .A1(n3552), .A2(n3522), .ZN(n3551) );
  INV_X1 U3991 ( .A(n3963), .ZN(n3964) );
  AND2_X1 U3992 ( .A1(n4148), .A2(n4147), .ZN(n4485) );
  INV_X1 U3993 ( .A(n4090), .ZN(n3928) );
  AND2_X1 U3994 ( .A1(n3906), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3944)
         );
  INV_X1 U3995 ( .A(n5185), .ZN(n3784) );
  NAND2_X1 U3996 ( .A1(n3656), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3672)
         );
  INV_X1 U3997 ( .A(n5373), .ZN(n5374) );
  AND2_X1 U3998 ( .A1(n3440), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3441)
         );
  AND2_X1 U3999 ( .A1(n4520), .A2(n4528), .ZN(n4525) );
  NAND2_X1 U4000 ( .A1(n3370), .A2(n3369), .ZN(n6247) );
  NAND2_X1 U4001 ( .A1(n3673), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3214) );
  NAND2_X1 U4002 ( .A1(n4112), .A2(n3551), .ZN(n3560) );
  NAND2_X1 U4003 ( .A1(n3986), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4012)
         );
  AND2_X1 U4004 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n3964), .ZN(n3986)
         );
  INV_X1 U4005 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5814) );
  NOR2_X1 U4006 ( .A1(n3672), .A2(n3657), .ZN(n3698) );
  OR2_X1 U4007 ( .A1(n5034), .A2(n4913), .ZN(n5858) );
  OR3_X1 U4008 ( .A1(n5034), .A2(n4857), .A3(n6488), .ZN(n5889) );
  INV_X1 U4009 ( .A(n4658), .ZN(n4378) );
  INV_X1 U4010 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6634) );
  INV_X1 U4011 ( .A(n5210), .ZN(n3718) );
  INV_X1 U4012 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4980) );
  OR2_X1 U4013 ( .A1(n5286), .A2(n5416), .ZN(n5263) );
  AND2_X1 U4014 ( .A1(n4172), .A2(n4171), .ZN(n5119) );
  NOR2_X1 U4015 ( .A1(n4764), .A2(n3113), .ZN(n4944) );
  NOR2_X1 U4016 ( .A1(n4244), .A2(n5484), .ZN(n6056) );
  INV_X1 U4017 ( .A(n6370), .ZN(n4353) );
  OR2_X1 U4018 ( .A1(n4689), .A2(n3566), .ZN(n4869) );
  INV_X1 U4019 ( .A(n4606), .ZN(n4631) );
  OR2_X1 U4020 ( .A1(n4830), .A2(n4280), .ZN(n4292) );
  NOR2_X1 U4021 ( .A1(n5601), .A2(n5042), .ZN(n5592) );
  NOR2_X1 U4022 ( .A1(n5637), .A2(n5625), .ZN(n5609) );
  NOR2_X1 U4023 ( .A1(n6452), .A2(n5803), .ZN(n5797) );
  INV_X1 U4024 ( .A(n5887), .ZN(n5620) );
  INV_X1 U4025 ( .A(n5858), .ZN(n5875) );
  INV_X1 U4026 ( .A(n5894), .ZN(n5865) );
  INV_X1 U4027 ( .A(n5873), .ZN(n5886) );
  INV_X1 U4028 ( .A(n5905), .ZN(n6517) );
  OAI21_X1 U4029 ( .B1(n6507), .B2(n6599), .A(n5947), .ZN(n6001) );
  INV_X1 U4030 ( .A(n6011), .ZN(n6004) );
  AOI21_X1 U4031 ( .B1(n5163), .B2(n5162), .A(n2981), .ZN(n5614) );
  NAND2_X1 U4032 ( .A1(n3802), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3851)
         );
  NAND2_X1 U4033 ( .A1(n3612), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3633)
         );
  INV_X1 U4034 ( .A(n5435), .ZN(n5690) );
  NOR2_X1 U4035 ( .A1(n5731), .A2(n5737), .ZN(n5722) );
  OR2_X1 U4036 ( .A1(n5484), .A2(n5482), .ZN(n5730) );
  NAND2_X1 U4037 ( .A1(n5480), .A2(n5496), .ZN(n5511) );
  INV_X1 U4038 ( .A(n6088), .ZN(n6111) );
  INV_X1 U4039 ( .A(n6071), .ZN(n6112) );
  INV_X1 U4040 ( .A(n4257), .ZN(n6108) );
  INV_X1 U4041 ( .A(n5565), .ZN(n5573) );
  INV_X1 U4042 ( .A(n2995), .ZN(n4689) );
  INV_X1 U4043 ( .A(n6152), .ZN(n6176) );
  AND2_X1 U4044 ( .A1(n4737), .A2(n6203), .ZN(n6194) );
  NOR2_X1 U4045 ( .A1(n4869), .A2(n5521), .ZN(n4580) );
  INV_X1 U4046 ( .A(n4871), .ZN(n4903) );
  AND2_X1 U4047 ( .A1(n5521), .A2(n4696), .ZN(n4870) );
  NOR2_X1 U4048 ( .A1(n5976), .A2(n4779), .ZN(n6259) );
  INV_X1 U4049 ( .A(n5548), .ZN(n6307) );
  INV_X1 U4050 ( .A(n5564), .ZN(n6338) );
  INV_X1 U4051 ( .A(n6245), .ZN(n6295) );
  INV_X1 U4052 ( .A(n4887), .ZN(n6347) );
  INV_X1 U4053 ( .A(READY_N), .ZN(n6599) );
  INV_X1 U4054 ( .A(n6477), .ZN(n6471) );
  AND2_X1 U4055 ( .A1(n4292), .A2(n4291), .ZN(n6511) );
  INV_X1 U4056 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6638) );
  OR2_X1 U4057 ( .A1(n5034), .A2(n6487), .ZN(n5890) );
  OR2_X1 U4058 ( .A1(n5038), .A2(n4845), .ZN(n5894) );
  OR3_X1 U4059 ( .A1(n5034), .A2(n4856), .A3(n6488), .ZN(n5861) );
  AND2_X1 U4060 ( .A1(n4842), .A2(n5861), .ZN(n5899) );
  NAND2_X1 U4061 ( .A1(n5905), .A2(n3320), .ZN(n5212) );
  INV_X1 U4062 ( .A(n6519), .ZN(n5902) );
  INV_X1 U4063 ( .A(n5920), .ZN(n5945) );
  OR3_X2 U4064 ( .A1(n4830), .A2(n4829), .A3(READY_N), .ZN(n6007) );
  AND2_X1 U4065 ( .A1(n4095), .A2(n4094), .ZN(n4096) );
  OR2_X1 U4066 ( .A1(n6406), .A2(n6295), .ZN(n6043) );
  NAND2_X1 U4067 ( .A1(n4246), .A2(n4124), .ZN(n5519) );
  INV_X1 U4068 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6201) );
  AND2_X1 U4069 ( .A1(n4421), .A2(n4420), .ZN(n4637) );
  AND2_X1 U4070 ( .A1(n5540), .A2(n5539), .ZN(n5571) );
  INV_X1 U4071 ( .A(n6133), .ZN(n4546) );
  NAND2_X1 U4072 ( .A1(n4737), .A2(n4870), .ZN(n6200) );
  AND2_X1 U4073 ( .A1(n4789), .A2(n4788), .ZN(n4814) );
  NAND2_X1 U4074 ( .A1(n4580), .A2(n4696), .ZN(n4820) );
  INV_X1 U4075 ( .A(n6256), .ZN(n6308) );
  INV_X1 U4076 ( .A(n6279), .ZN(n6358) );
  NAND2_X1 U4077 ( .A1(n6205), .A2(n4870), .ZN(n6237) );
  NAND2_X1 U4078 ( .A1(n6205), .A2(n6203), .ZN(n6284) );
  AND2_X1 U4079 ( .A1(n4362), .A2(n4361), .ZN(n4505) );
  NAND2_X1 U4080 ( .A1(n3561), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6400) );
  INV_X1 U4081 ( .A(n6484), .ZN(n6480) );
  INV_X1 U4082 ( .A(n6475), .ZN(n6473) );
  AND2_X2 U4083 ( .A1(n4350), .A2(n3121), .ZN(n3156) );
  AND2_X2 U4084 ( .A1(n4656), .A2(n4670), .ZN(n3203) );
  AOI22_X1 U4085 ( .A1(n3156), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3203), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3120) );
  AND2_X2 U4086 ( .A1(n4341), .A2(n3121), .ZN(n3179) );
  AND2_X2 U4087 ( .A1(n4341), .A2(n4670), .ZN(n3841) );
  AOI22_X1 U4088 ( .A1(n3179), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3841), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3119) );
  INV_X1 U4089 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3116) );
  AND2_X2 U4090 ( .A1(n3122), .A2(n4656), .ZN(n3300) );
  AOI22_X1 U4091 ( .A1(n3282), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3300), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3118) );
  AOI22_X1 U4092 ( .A1(n3877), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3117) );
  AND2_X2 U4093 ( .A1(n3121), .A2(n4656), .ZN(n4026) );
  AOI22_X1 U4094 ( .A1(n4026), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n2979), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3125) );
  AND2_X2 U4095 ( .A1(n4350), .A2(n3122), .ZN(n3141) );
  AOI22_X1 U4096 ( .A1(n3352), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3301), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3123) );
  NAND2_X2 U4097 ( .A1(n2992), .A2(n3127), .ZN(n3239) );
  AOI22_X1 U4098 ( .A1(n3841), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3301), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3128) );
  AOI22_X1 U4099 ( .A1(n3673), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3352), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3135) );
  AOI22_X1 U4100 ( .A1(n3282), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3300), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3134) );
  AOI22_X1 U4101 ( .A1(n3179), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3877), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3133) );
  AOI22_X1 U4102 ( .A1(n3202), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3203), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3140) );
  AOI22_X1 U4103 ( .A1(n3156), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3139) );
  AOI22_X1 U4104 ( .A1(n3136), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        INSTQUEUE_REG_5__6__SCAN_IN), .B2(n3225), .ZN(n3138) );
  AOI22_X1 U4105 ( .A1(n3841), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3301), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3137) );
  AOI22_X1 U4106 ( .A1(n3282), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3300), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3144) );
  AOI22_X1 U4107 ( .A1(n3141), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3143) );
  MUX2_X1 U4108 ( .A(n3239), .B(n3165), .S(n3260), .Z(n3193) );
  NAND2_X1 U4109 ( .A1(n3673), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3151) );
  NAND2_X1 U4110 ( .A1(n3352), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3150)
         );
  NAND2_X1 U4111 ( .A1(n3300), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3149) );
  NAND2_X1 U4112 ( .A1(n3179), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3148) );
  NAND2_X1 U4113 ( .A1(n3225), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3155) );
  NAND2_X1 U4114 ( .A1(n3202), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3154)
         );
  NAND2_X1 U4115 ( .A1(n3136), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3153)
         );
  NAND2_X1 U4116 ( .A1(n3301), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3152)
         );
  NAND2_X1 U4117 ( .A1(n4026), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3160) );
  NAND2_X1 U4118 ( .A1(n3156), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3159)
         );
  NAND2_X1 U4119 ( .A1(n3841), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3158) );
  NAND2_X1 U4120 ( .A1(n3203), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3157) );
  NAND2_X1 U4121 ( .A1(n3282), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3164) );
  NAND2_X1 U4122 ( .A1(n3141), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3163) );
  NAND2_X1 U4123 ( .A1(n3877), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3162)
         );
  NAND2_X1 U4124 ( .A1(n3302), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3161) );
  AND4_X2 U4125 ( .A1(n3170), .A2(n3167), .A3(n3168), .A4(n3169), .ZN(n3243)
         );
  INV_X1 U4126 ( .A(n4382), .ZN(n3192) );
  NAND2_X1 U4127 ( .A1(n4382), .A2(n4226), .ZN(n3166) );
  NAND2_X2 U4128 ( .A1(n3575), .A2(n4434), .ZN(n3248) );
  AOI22_X1 U4129 ( .A1(n3156), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3174) );
  AOI22_X1 U4130 ( .A1(n3225), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3136), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3173) );
  AOI22_X1 U4131 ( .A1(n3179), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3203), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3172) );
  AOI22_X1 U4132 ( .A1(n3877), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3171) );
  AOI22_X1 U4133 ( .A1(n3141), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3673), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3178) );
  AOI22_X1 U4134 ( .A1(n3282), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3300), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3177) );
  AOI22_X1 U4135 ( .A1(n3352), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3841), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3176) );
  AOI22_X1 U4136 ( .A1(n3156), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3183) );
  AOI22_X1 U4137 ( .A1(n3179), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3841), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3182) );
  AOI22_X1 U4138 ( .A1(n4026), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3136), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3181) );
  AOI22_X1 U4139 ( .A1(n3282), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3180) );
  NAND4_X1 U4140 ( .A1(n3183), .A2(n3182), .A3(n3181), .A4(n3180), .ZN(n3189)
         );
  AOI22_X1 U4141 ( .A1(n3225), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3203), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3187) );
  AOI22_X1 U4142 ( .A1(n3673), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3877), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3186) );
  AOI22_X1 U4143 ( .A1(n3141), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3300), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3185) );
  AOI22_X1 U4144 ( .A1(n3352), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3301), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3184) );
  NAND4_X1 U4145 ( .A1(n3187), .A2(n3186), .A3(n3185), .A4(n3184), .ZN(n3188)
         );
  OR2_X2 U4146 ( .A1(n3189), .A2(n3188), .ZN(n3320) );
  INV_X1 U4147 ( .A(n3320), .ZN(n4388) );
  NAND2_X1 U4148 ( .A1(n3156), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3197)
         );
  NAND2_X1 U4149 ( .A1(n3136), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3196)
         );
  NAND2_X1 U4150 ( .A1(n4026), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3195) );
  NAND2_X1 U4151 ( .A1(n3225), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3194) );
  NAND2_X1 U4152 ( .A1(n3282), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3201) );
  NAND2_X1 U4153 ( .A1(n3141), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3200) );
  NAND2_X1 U4154 ( .A1(n3300), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3199) );
  NAND2_X1 U4155 ( .A1(n3302), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3198) );
  NAND2_X1 U4156 ( .A1(n2980), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3207)
         );
  NAND2_X1 U4157 ( .A1(n3841), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3206) );
  NAND2_X1 U4158 ( .A1(n3203), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3205) );
  NAND2_X1 U4159 ( .A1(n3301), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3204)
         );
  NAND2_X4 U4160 ( .A1(n3216), .A2(n3215), .ZN(n4852) );
  NAND2_X1 U4161 ( .A1(n3322), .A2(n3563), .ZN(n3246) );
  NAND2_X1 U4162 ( .A1(n3156), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3220)
         );
  NAND2_X1 U4163 ( .A1(n3673), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3219) );
  NAND2_X1 U4164 ( .A1(n3352), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3218)
         );
  NAND2_X1 U4165 ( .A1(n3841), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3217) );
  NAND2_X1 U4166 ( .A1(n3179), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3224) );
  NAND2_X1 U4167 ( .A1(n3282), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3223) );
  NAND2_X1 U4168 ( .A1(n3877), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3222)
         );
  NAND2_X1 U4169 ( .A1(n3302), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3221) );
  NAND2_X1 U4170 ( .A1(n4026), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3229) );
  NAND2_X1 U4171 ( .A1(n2980), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3228)
         );
  NAND2_X1 U4172 ( .A1(n3225), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3227) );
  NAND2_X1 U4173 ( .A1(n3136), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3226)
         );
  NAND2_X1 U4174 ( .A1(n3141), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3233) );
  NAND2_X1 U4175 ( .A1(n3300), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3232) );
  NAND2_X1 U4176 ( .A1(n3301), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3231)
         );
  NAND2_X1 U4177 ( .A1(n3203), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3230) );
  NAND3_X1 U4178 ( .A1(n4382), .A2(n3320), .A3(n4226), .ZN(n4104) );
  NAND2_X1 U4179 ( .A1(n3385), .A2(n4104), .ZN(n3238) );
  INV_X1 U4180 ( .A(n3253), .ZN(n4121) );
  INV_X1 U4181 ( .A(n3248), .ZN(n3240) );
  NAND2_X1 U4182 ( .A1(n3240), .A2(n4226), .ZN(n3242) );
  NAND2_X1 U4183 ( .A1(n3242), .A2(n3241), .ZN(n3258) );
  NAND2_X2 U4184 ( .A1(n4381), .A2(n4411), .ZN(n4232) );
  XNOR2_X1 U4185 ( .A(STATE_REG_1__SCAN_IN), .B(STATE_REG_2__SCAN_IN), .ZN(
        n4097) );
  NAND2_X1 U4186 ( .A1(n4103), .A2(n4097), .ZN(n3321) );
  NAND2_X1 U4187 ( .A1(n3321), .A2(n3243), .ZN(n3244) );
  AND2_X1 U4188 ( .A1(n3244), .A2(n4843), .ZN(n3245) );
  NAND4_X1 U4189 ( .A1(n3246), .A2(n3265), .A3(n3565), .A4(n3245), .ZN(n3247)
         );
  NAND2_X1 U4190 ( .A1(n3247), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3250) );
  MUX2_X1 U4191 ( .A(n3346), .B(n3347), .S(n6287), .Z(n3251) );
  INV_X1 U4192 ( .A(n3251), .ZN(n3252) );
  INV_X1 U4193 ( .A(n4843), .ZN(n4279) );
  NAND2_X1 U4194 ( .A1(n4279), .A2(n3253), .ZN(n4230) );
  NAND3_X1 U4195 ( .A1(n3108), .A2(n4230), .A3(n3255), .ZN(n3257) );
  NOR2_X2 U4196 ( .A1(n3257), .A2(n3256), .ZN(n4238) );
  AND2_X1 U4197 ( .A1(n3248), .A2(n3239), .ZN(n3259) );
  OAI21_X1 U4198 ( .B1(n3258), .B2(n3259), .A(n4407), .ZN(n3266) );
  NAND3_X1 U4199 ( .A1(n3262), .A2(n4103), .A3(n3261), .ZN(n3263) );
  INV_X1 U4200 ( .A(n4411), .ZN(n4380) );
  OR2_X1 U4201 ( .A1(n6494), .A2(n6509), .ZN(n6401) );
  AOI21_X1 U4202 ( .B1(n3263), .B2(n4380), .A(n6401), .ZN(n3264) );
  NAND2_X1 U4203 ( .A1(n4238), .A2(n3267), .ZN(n3269) );
  INV_X1 U4204 ( .A(n4383), .ZN(n3296) );
  AOI22_X1 U4205 ( .A1(n3855), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3275) );
  AOI22_X1 U4206 ( .A1(n3888), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3179), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3274) );
  AOI22_X1 U4207 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n2980), .B1(n4046), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3273) );
  AOI22_X1 U4208 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n3300), .B1(n4020), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3272) );
  NAND4_X1 U4209 ( .A1(n3275), .A2(n3274), .A3(n3273), .A4(n3272), .ZN(n3281)
         );
  AOI22_X1 U4210 ( .A1(n4021), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3279) );
  AOI22_X1 U4211 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n4018), .B1(n3877), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3278) );
  AOI22_X1 U4212 ( .A1(n3993), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3277) );
  INV_X1 U4213 ( .A(n3301), .ZN(n3287) );
  AOI22_X1 U4214 ( .A1(n3893), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3276) );
  NAND4_X1 U4215 ( .A1(n3279), .A2(n3278), .A3(n3277), .A4(n3276), .ZN(n3280)
         );
  INV_X1 U4216 ( .A(n3405), .ZN(n3294) );
  AOI22_X1 U4217 ( .A1(n4027), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n2980), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3286) );
  AOI22_X1 U4218 ( .A1(n3836), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3300), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3285) );
  AOI22_X1 U4219 ( .A1(n4019), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3877), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3284) );
  AOI22_X1 U4220 ( .A1(n3888), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3283) );
  NAND4_X1 U4221 ( .A1(n3286), .A2(n3285), .A3(n3284), .A4(n3283), .ZN(n3293)
         );
  AOI22_X1 U4222 ( .A1(n4018), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3893), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3291) );
  AOI22_X1 U4223 ( .A1(n3855), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3290) );
  AOI22_X1 U4224 ( .A1(n4021), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4020), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3289) );
  AOI22_X1 U4225 ( .A1(n3993), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3288) );
  NAND4_X1 U4226 ( .A1(n3291), .A2(n3290), .A3(n3289), .A4(n3288), .ZN(n3292)
         );
  XNOR2_X1 U4227 ( .A(n3294), .B(n3489), .ZN(n3295) );
  NAND2_X1 U4228 ( .A1(n3296), .A2(n3295), .ZN(n3401) );
  INV_X1 U4229 ( .A(n3552), .ZN(n3548) );
  INV_X1 U4230 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4441) );
  AOI21_X1 U4231 ( .B1(n4226), .B2(n3489), .A(n6509), .ZN(n3298) );
  NAND2_X1 U4232 ( .A1(n3563), .A2(n3405), .ZN(n3297) );
  OAI211_X1 U4233 ( .C1(n3548), .C2(n4441), .A(n3298), .B(n3297), .ZN(n3402)
         );
  INV_X1 U4234 ( .A(n3489), .ZN(n3299) );
  AOI22_X1 U4235 ( .A1(n3836), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3300), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3306) );
  AOI22_X1 U4236 ( .A1(n3855), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3993), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3305) );
  AOI22_X1 U4237 ( .A1(n3202), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3304) );
  AOI22_X1 U4238 ( .A1(n3888), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4020), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3303) );
  NAND4_X1 U4239 ( .A1(n3306), .A2(n3305), .A3(n3304), .A4(n3303), .ZN(n3312)
         );
  AOI22_X1 U4240 ( .A1(n4018), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4019), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3310) );
  AOI22_X1 U4241 ( .A1(n4021), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3309) );
  AOI22_X1 U4242 ( .A1(n3893), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3308) );
  AOI22_X1 U4243 ( .A1(n4027), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3307) );
  NAND4_X1 U4244 ( .A1(n3310), .A2(n3309), .A3(n3308), .A4(n3307), .ZN(n3311)
         );
  OR2_X1 U4245 ( .A1(n3371), .A2(n3336), .ZN(n3314) );
  NAND2_X1 U4246 ( .A1(n3552), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3313) );
  OAI211_X1 U4247 ( .C1(n4383), .C2(n3489), .A(n3314), .B(n3313), .ZN(n3388)
         );
  INV_X1 U4248 ( .A(n4104), .ZN(n3317) );
  NOR2_X1 U4249 ( .A1(n4232), .A2(n4434), .ZN(n3316) );
  AND2_X1 U4250 ( .A1(n4346), .A2(n4852), .ZN(n4275) );
  NOR2_X1 U4251 ( .A1(n4411), .A2(n4434), .ZN(n3318) );
  NAND2_X1 U4252 ( .A1(n3320), .A2(n3261), .ZN(n5028) );
  AOI21_X1 U4253 ( .B1(n4275), .B2(n3321), .A(n4227), .ZN(n3325) );
  INV_X1 U4254 ( .A(n3322), .ZN(n3324) );
  NOR2_X1 U4255 ( .A1(n3253), .A2(n4852), .ZN(n3323) );
  AND2_X2 U4256 ( .A1(n3324), .A2(n3323), .ZN(n4276) );
  NAND2_X2 U4257 ( .A1(n4276), .A2(n4103), .ZN(n4653) );
  NAND2_X1 U4258 ( .A1(n3325), .A2(n4653), .ZN(n3326) );
  NAND2_X1 U4259 ( .A1(n3326), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3333) );
  INV_X1 U4260 ( .A(n3333), .ZN(n3330) );
  XNOR2_X1 U4261 ( .A(n6287), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6140)
         );
  AND2_X1 U4262 ( .A1(n3346), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3327)
         );
  AOI21_X1 U4263 ( .B1(n3347), .B2(n6140), .A(n3327), .ZN(n3332) );
  INV_X1 U4264 ( .A(n3332), .ZN(n3328) );
  NAND2_X1 U4265 ( .A1(n3331), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3334) );
  NAND3_X1 U4266 ( .A1(n3334), .A2(n3333), .A3(n3332), .ZN(n3339) );
  NAND2_X1 U4267 ( .A1(n3341), .A2(n3339), .ZN(n3335) );
  XNOR2_X2 U4268 ( .A(n3340), .B(n3335), .ZN(n4518) );
  NAND2_X1 U4269 ( .A1(n4518), .A2(n6509), .ZN(n3338) );
  NAND2_X1 U4270 ( .A1(n3340), .A2(n3339), .ZN(n3342) );
  NAND2_X1 U4271 ( .A1(n3331), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3349) );
  AND2_X1 U4272 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3343) );
  NAND2_X1 U4273 ( .A1(n3343), .A2(n6589), .ZN(n6202) );
  INV_X1 U4274 ( .A(n3343), .ZN(n3344) );
  NAND2_X1 U4275 ( .A1(n3344), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3345) );
  NAND2_X1 U4276 ( .A1(n6202), .A2(n3345), .ZN(n4423) );
  AOI22_X1 U4277 ( .A1(n3347), .A2(n4423), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3346), .ZN(n3348) );
  NAND2_X1 U4278 ( .A1(n3349), .A2(n3348), .ZN(n3350) );
  AOI22_X1 U4279 ( .A1(n3888), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4018), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3356) );
  AOI22_X1 U4280 ( .A1(n3836), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4039), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3355) );
  AOI22_X1 U4281 ( .A1(n4019), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3354) );
  AOI22_X1 U4282 ( .A1(n4021), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4020), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3353) );
  NAND4_X1 U4283 ( .A1(n3356), .A2(n3355), .A3(n3354), .A4(n3353), .ZN(n3362)
         );
  AOI22_X1 U4284 ( .A1(n4027), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3993), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3360) );
  AOI22_X1 U4285 ( .A1(n2980), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3359) );
  AOI22_X1 U4286 ( .A1(n3855), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3358) );
  INV_X2 U4287 ( .A(n3287), .ZN(n4041) );
  AOI22_X1 U4288 ( .A1(n3893), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3357) );
  NAND4_X1 U4289 ( .A1(n3360), .A2(n3359), .A3(n3358), .A4(n3357), .ZN(n3361)
         );
  INV_X1 U4290 ( .A(n3371), .ZN(n3363) );
  AOI22_X1 U4291 ( .A1(n3363), .A2(n3416), .B1(n3552), .B2(
        INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3364) );
  XNOR2_X1 U4292 ( .A(n3365), .B(n3364), .ZN(n3413) );
  NAND2_X1 U4293 ( .A1(n3331), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3370) );
  NOR3_X1 U4294 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6589), .A3(n6373), 
        .ZN(n4742) );
  NAND2_X1 U4295 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4742), .ZN(n4734) );
  NAND2_X1 U4296 ( .A1(n6201), .A2(n4734), .ZN(n3367) );
  NAND3_X1 U4297 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4600) );
  INV_X1 U4298 ( .A(n4600), .ZN(n4367) );
  NAND2_X1 U4299 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4367), .ZN(n4509) );
  NAND2_X1 U4300 ( .A1(n3367), .A2(n4509), .ZN(n4778) );
  OAI22_X1 U4301 ( .A1(n4078), .A2(n4778), .B1(n3561), .B2(n6201), .ZN(n3368)
         );
  INV_X1 U4302 ( .A(n3368), .ZN(n3369) );
  XNOR2_X1 U4303 ( .A(n3366), .B(n6247), .ZN(n4357) );
  NAND2_X1 U4304 ( .A1(n4357), .A2(n6509), .ZN(n3383) );
  AOI22_X1 U4305 ( .A1(n3888), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3375) );
  AOI22_X1 U4306 ( .A1(n4018), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4019), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3374) );
  AOI22_X1 U4307 ( .A1(n4021), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3373) );
  AOI22_X1 U4308 ( .A1(n3971), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4020), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3372) );
  NAND4_X1 U4309 ( .A1(n3375), .A2(n3374), .A3(n3373), .A4(n3372), .ZN(n3381)
         );
  AOI22_X1 U4310 ( .A1(n3855), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4039), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3379) );
  AOI22_X1 U4311 ( .A1(n4027), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n2980), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3378) );
  AOI22_X1 U4312 ( .A1(n3893), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3377) );
  AOI22_X1 U4313 ( .A1(n3993), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3376) );
  NAND4_X1 U4314 ( .A1(n3379), .A2(n3378), .A3(n3377), .A4(n3376), .ZN(n3380)
         );
  AOI22_X1 U4315 ( .A1(n3541), .A2(n3437), .B1(n3552), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3382) );
  INV_X1 U4316 ( .A(n4363), .ZN(n4445) );
  NAND2_X1 U4317 ( .A1(n3414), .A2(n4445), .ZN(n3590) );
  NAND2_X1 U4318 ( .A1(n3394), .A2(n3405), .ZN(n3417) );
  NAND2_X1 U4319 ( .A1(n3417), .A2(n3384), .ZN(n3438) );
  NAND2_X1 U4320 ( .A1(n3013), .A2(n6507), .ZN(n3386) );
  NAND2_X1 U4321 ( .A1(n3387), .A2(n3386), .ZN(n3426) );
  INV_X1 U4322 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6106) );
  XNOR2_X1 U4323 ( .A(n3426), .B(n6106), .ZN(n4972) );
  NAND2_X1 U4324 ( .A1(n3389), .A2(n3388), .ZN(n3390) );
  OAI21_X1 U4325 ( .B1(n3405), .B2(n3394), .A(n3417), .ZN(n3396) );
  INV_X1 U4326 ( .A(n4232), .ZN(n3395) );
  OAI211_X1 U4327 ( .C1(n3396), .C2(n3262), .A(n3395), .B(n4434), .ZN(n3397)
         );
  INV_X1 U4328 ( .A(n3397), .ZN(n3398) );
  NAND2_X1 U4329 ( .A1(n3400), .A2(n3402), .ZN(n3404) );
  NAND2_X2 U4330 ( .A1(n3404), .A2(n3403), .ZN(n3574) );
  NAND2_X1 U4331 ( .A1(n3574), .A2(n3522), .ZN(n3408) );
  NAND2_X1 U4332 ( .A1(n3563), .A2(n4411), .ZN(n3418) );
  OAI21_X1 U4333 ( .B1(n3262), .B2(n3405), .A(n3418), .ZN(n3406) );
  INV_X1 U4334 ( .A(n3406), .ZN(n3407) );
  NAND2_X1 U4335 ( .A1(n3408), .A2(n3407), .ZN(n4297) );
  NAND2_X1 U4336 ( .A1(n4297), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3409)
         );
  INV_X1 U4337 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4342) );
  AND2_X1 U4338 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3410) );
  NAND2_X1 U4339 ( .A1(n4297), .A2(n3410), .ZN(n3411) );
  NAND2_X1 U4340 ( .A1(n6031), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3421)
         );
  XNOR2_X1 U4341 ( .A(n3417), .B(n3416), .ZN(n3419) );
  OAI21_X1 U4342 ( .B1(n3419), .B2(n3262), .A(n3418), .ZN(n3420) );
  NAND2_X1 U4343 ( .A1(n3421), .A2(n6032), .ZN(n3425) );
  INV_X1 U4344 ( .A(n6031), .ZN(n3423) );
  INV_X1 U4345 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3422) );
  NAND2_X1 U4346 ( .A1(n3423), .A2(n3422), .ZN(n3424) );
  AOI22_X1 U4347 ( .A1(n3888), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4018), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3430) );
  AOI22_X1 U4348 ( .A1(n3836), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4039), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3429) );
  AOI22_X1 U4349 ( .A1(n4019), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3428) );
  AOI22_X1 U4350 ( .A1(n4021), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4020), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3427) );
  NAND4_X1 U4351 ( .A1(n3430), .A2(n3429), .A3(n3428), .A4(n3427), .ZN(n3436)
         );
  AOI22_X1 U4352 ( .A1(n4027), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3993), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3434) );
  AOI22_X1 U4353 ( .A1(n2980), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3433) );
  AOI22_X1 U4354 ( .A1(n3855), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3432) );
  AOI22_X1 U4355 ( .A1(n3893), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3431) );
  NAND4_X1 U4356 ( .A1(n3434), .A2(n3433), .A3(n3432), .A4(n3431), .ZN(n3435)
         );
  XNOR2_X1 U4357 ( .A(n3442), .B(n3443), .ZN(n3597) );
  NAND2_X1 U4358 ( .A1(n3438), .A2(n3437), .ZN(n3478) );
  XOR2_X1 U4359 ( .A(n3476), .B(n3478), .Z(n3439) );
  XNOR2_X1 U4360 ( .A(n3440), .B(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6026)
         );
  NOR2_X1 U4361 ( .A1(n6025), .A2(n6026), .ZN(n6024) );
  NOR2_X1 U4362 ( .A1(n6024), .A2(n3441), .ZN(n4765) );
  INV_X1 U4363 ( .A(n3443), .ZN(n3444) );
  NAND2_X1 U4364 ( .A1(n3445), .A2(n3444), .ZN(n3460) );
  AOI22_X1 U4365 ( .A1(n4039), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4019), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3449) );
  AOI22_X1 U4366 ( .A1(n3855), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3448) );
  AOI22_X1 U4367 ( .A1(n4027), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3447) );
  AOI22_X1 U4368 ( .A1(n4018), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3446) );
  NAND4_X1 U4369 ( .A1(n3449), .A2(n3448), .A3(n3447), .A4(n3446), .ZN(n3455)
         );
  AOI22_X1 U4370 ( .A1(n3888), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3453) );
  AOI22_X1 U4371 ( .A1(n3993), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3893), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3452) );
  INV_X1 U4372 ( .A(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n6665) );
  AOI22_X1 U4373 ( .A1(n4021), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3451) );
  AOI22_X1 U4374 ( .A1(n3836), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4020), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3450) );
  NAND4_X1 U4375 ( .A1(n3453), .A2(n3452), .A3(n3451), .A4(n3450), .ZN(n3454)
         );
  INV_X1 U4376 ( .A(n3478), .ZN(n3456) );
  NAND2_X1 U4377 ( .A1(n3456), .A2(n3476), .ZN(n3457) );
  XOR2_X1 U4378 ( .A(n3475), .B(n3457), .Z(n3458) );
  XNOR2_X1 U4379 ( .A(n3459), .B(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4766)
         );
  NOR2_X1 U4380 ( .A1(n4765), .A2(n4766), .ZN(n4764) );
  INV_X1 U4381 ( .A(n3461), .ZN(n3462) );
  AOI22_X1 U4382 ( .A1(n3888), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4018), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3466) );
  AOI22_X1 U4383 ( .A1(n3836), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4039), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3465) );
  AOI22_X1 U4384 ( .A1(n4019), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3464) );
  AOI22_X1 U4385 ( .A1(n4021), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4020), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3463) );
  NAND4_X1 U4386 ( .A1(n3466), .A2(n3465), .A3(n3464), .A4(n3463), .ZN(n3472)
         );
  AOI22_X1 U4387 ( .A1(n4027), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3993), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3470) );
  AOI22_X1 U4388 ( .A1(n2980), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3469) );
  AOI22_X1 U4389 ( .A1(n3855), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3468) );
  AOI22_X1 U4390 ( .A1(n3893), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3467) );
  NAND4_X1 U4391 ( .A1(n3470), .A2(n3469), .A3(n3468), .A4(n3467), .ZN(n3471)
         );
  NAND2_X1 U4392 ( .A1(n3474), .A2(n3473), .ZN(n3616) );
  NAND2_X1 U4393 ( .A1(n3616), .A2(n3522), .ZN(n3480) );
  NAND2_X1 U4394 ( .A1(n3476), .A2(n3475), .ZN(n3477) );
  NOR2_X1 U4395 ( .A1(n3478), .A2(n3477), .ZN(n3486) );
  XNOR2_X1 U4396 ( .A(n3486), .B(n3485), .ZN(n3479) );
  OAI22_X1 U4397 ( .A1(n3483), .A2(n3480), .B1(n3479), .B2(n3262), .ZN(n3481)
         );
  XNOR2_X1 U4398 ( .A(n3481), .B(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4945)
         );
  NOR2_X1 U4399 ( .A1(n4944), .A2(n4945), .ZN(n4943) );
  AOI22_X1 U4400 ( .A1(n3541), .A2(n3489), .B1(n3552), .B2(
        INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3484) );
  XNOR2_X1 U4401 ( .A(n3492), .B(n3484), .ZN(n3619) );
  NAND2_X1 U4402 ( .A1(n3486), .A2(n3485), .ZN(n3494) );
  XOR2_X1 U4403 ( .A(n3489), .B(n3494), .Z(n3487) );
  OAI22_X1 U4404 ( .A1(n3619), .A2(n3040), .B1(n3487), .B2(n3262), .ZN(n3488)
         );
  XNOR2_X1 U4405 ( .A(n3488), .B(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n5392)
         );
  NAND2_X1 U4406 ( .A1(n6507), .A2(n3489), .ZN(n3493) );
  NAND2_X1 U4407 ( .A1(n3522), .A2(n3489), .ZN(n3490) );
  OAI21_X1 U4408 ( .B1(n3494), .B2(n3493), .A(n3499), .ZN(n3495) );
  XNOR2_X1 U4409 ( .A(n3495), .B(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5382)
         );
  INV_X1 U4410 ( .A(n3495), .ZN(n3497) );
  NOR2_X1 U4411 ( .A1(n5508), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5375)
         );
  INV_X1 U4412 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5365) );
  INV_X1 U4413 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3501) );
  NOR2_X1 U4414 ( .A1(n5686), .A2(n3501), .ZN(n5357) );
  XNOR2_X1 U4415 ( .A(n5686), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5351)
         );
  INV_X1 U4416 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3502) );
  INV_X1 U4417 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4167) );
  NAND2_X1 U4418 ( .A1(n5686), .A2(n4167), .ZN(n3503) );
  INV_X1 U4419 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5742) );
  INV_X1 U4420 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3504) );
  INV_X1 U4421 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5726) );
  NAND2_X1 U4422 ( .A1(n3504), .A2(n5726), .ZN(n3505) );
  OAI21_X1 U4423 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n3505), .A(n5508), 
        .ZN(n3507) );
  NAND3_X1 U4424 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(INSTADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n3506) );
  INV_X1 U4425 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5678) );
  NOR2_X2 U4426 ( .A1(n5680), .A2(n3508), .ZN(n4083) );
  NOR2_X1 U4427 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3509) );
  INV_X1 U4428 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5459) );
  INV_X1 U4429 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5318) );
  INV_X1 U4430 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5460) );
  NAND4_X1 U4431 ( .A1(n3509), .A2(n5459), .A3(n5318), .A4(n5460), .ZN(n3510)
         );
  NAND2_X1 U4432 ( .A1(n5508), .A2(n3510), .ZN(n3511) );
  NAND2_X1 U4433 ( .A1(n4083), .A2(n3511), .ZN(n5270) );
  NAND2_X1 U4434 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5700) );
  AND2_X1 U4435 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5297) );
  AND2_X1 U4436 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4262) );
  NAND2_X1 U4437 ( .A1(n5297), .A2(n4262), .ZN(n3512) );
  OAI21_X1 U4438 ( .B1(n5700), .B2(n3512), .A(n5686), .ZN(n3513) );
  XNOR2_X1 U4439 ( .A(n5686), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5672)
         );
  INV_X1 U4440 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5694) );
  INV_X1 U4441 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5437) );
  NOR2_X1 U4442 ( .A1(n5508), .A2(n5437), .ZN(n5288) );
  NAND2_X1 U4443 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5417) );
  NOR2_X1 U4444 ( .A1(n5278), .A2(n5417), .ZN(n5261) );
  NAND2_X1 U4445 ( .A1(n5261), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5253) );
  INV_X1 U4446 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5399) );
  INV_X1 U4447 ( .A(n3514), .ZN(n3516) );
  INV_X1 U4448 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3515) );
  INV_X1 U4449 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4210) );
  NAND2_X1 U4450 ( .A1(n3515), .A2(n4210), .ZN(n5416) );
  NOR2_X1 U4451 ( .A1(n5263), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5252)
         );
  NAND3_X1 U4452 ( .A1(n3516), .A2(n5252), .A3(n5399), .ZN(n3517) );
  OAI21_X1 U4453 ( .B1(n5253), .B2(n5399), .A(n3517), .ZN(n3518) );
  XNOR2_X1 U4454 ( .A(n3518), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4272)
         );
  XNOR2_X1 U4455 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3528) );
  NAND2_X1 U4456 ( .A1(n3529), .A2(n3528), .ZN(n3520) );
  NAND2_X1 U4457 ( .A1(n6373), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3519) );
  NOR2_X1 U4458 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6125), .ZN(n3521)
         );
  NAND2_X1 U4459 ( .A1(n4112), .A2(n3541), .ZN(n3558) );
  NAND3_X1 U4460 ( .A1(n5758), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(n3523), .ZN(n4113) );
  INV_X1 U4461 ( .A(n3551), .ZN(n3555) );
  AOI21_X1 U4462 ( .B1(n3526), .B2(n3525), .A(n3524), .ZN(n3527) );
  INV_X1 U4463 ( .A(n3527), .ZN(n4111) );
  XNOR2_X1 U4464 ( .A(n3528), .B(n3529), .ZN(n4110) );
  AOI21_X1 U4465 ( .B1(n3541), .B2(n4407), .A(n3243), .ZN(n3535) );
  AOI21_X1 U4466 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n3114), .A(n3529), 
        .ZN(n3530) );
  AOI21_X1 U4467 ( .B1(n3530), .B2(n3541), .A(n3551), .ZN(n3534) );
  AOI21_X1 U4468 ( .B1(n3530), .B2(n3253), .A(n3563), .ZN(n3532) );
  NOR2_X1 U4469 ( .A1(n3243), .A2(n4407), .ZN(n3531) );
  NOR2_X1 U4470 ( .A1(n3532), .A2(n3542), .ZN(n3533) );
  AOI211_X1 U4471 ( .C1(n3535), .C2(n4110), .A(n3534), .B(n3533), .ZN(n3537)
         );
  NOR3_X1 U4472 ( .A1(n4110), .A2(n3535), .A3(n6509), .ZN(n3536) );
  AOI211_X1 U4473 ( .C1(n4110), .C2(n3551), .A(n3537), .B(n3536), .ZN(n3547)
         );
  XNOR2_X1 U4474 ( .A(n3539), .B(n3538), .ZN(n4109) );
  INV_X1 U4475 ( .A(n4109), .ZN(n3540) );
  AOI211_X1 U4476 ( .C1(n3552), .C2(n4109), .A(n3543), .B(n3542), .ZN(n3546)
         );
  INV_X1 U4477 ( .A(n3542), .ZN(n3545) );
  INV_X1 U4478 ( .A(n3543), .ZN(n3544) );
  OAI22_X1 U4479 ( .A1(n3547), .A2(n3546), .B1(n3545), .B2(n3544), .ZN(n3550)
         );
  NAND2_X1 U4480 ( .A1(n3548), .A2(n4111), .ZN(n3549) );
  AOI22_X1 U4481 ( .A1(n3551), .A2(n4111), .B1(n3550), .B2(n3549), .ZN(n3554)
         );
  NOR2_X1 U4482 ( .A1(n3552), .A2(n4113), .ZN(n3553) );
  OAI22_X1 U4483 ( .A1(n4113), .A2(n3555), .B1(n3554), .B2(n3553), .ZN(n3556)
         );
  AOI21_X1 U4484 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6509), .A(n3556), 
        .ZN(n3557) );
  NAND2_X1 U4485 ( .A1(n3558), .A2(n3557), .ZN(n3559) );
  NAND2_X1 U4486 ( .A1(n3239), .A2(n3320), .ZN(n3562) );
  NAND2_X1 U4487 ( .A1(n3749), .A2(n3563), .ZN(n3564) );
  NAND2_X1 U4488 ( .A1(n3565), .A2(n3564), .ZN(n4334) );
  OR2_X1 U4489 ( .A1(n4334), .A2(n3253), .ZN(n6381) );
  INV_X2 U4490 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6210) );
  NAND2_X1 U4491 ( .A1(n6210), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3760) );
  NAND2_X1 U4492 ( .A1(n5521), .A2(n3745), .ZN(n3573) );
  AOI22_X1 U4493 ( .A1(n3577), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6210), .ZN(n3571) );
  INV_X1 U4494 ( .A(n5028), .ZN(n3569) );
  NAND2_X1 U4495 ( .A1(n3591), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3570) );
  AND2_X1 U4496 ( .A1(n3571), .A2(n3570), .ZN(n3572) );
  NAND2_X1 U4497 ( .A1(n3573), .A2(n3572), .ZN(n4404) );
  AOI21_X1 U4498 ( .B1(n4696), .B2(n3575), .A(n6210), .ZN(n4402) );
  AOI22_X1 U4499 ( .A1(n3577), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6210), .ZN(n3579) );
  NAND2_X1 U4500 ( .A1(n3591), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3578) );
  OAI211_X1 U4501 ( .C1(n3576), .C2(n3716), .A(n3579), .B(n3578), .ZN(n4401)
         );
  MUX2_X1 U4502 ( .A(n2977), .B(n4402), .S(n4401), .Z(n4405) );
  NAND2_X1 U4503 ( .A1(n3586), .A2(n3587), .ZN(n3585) );
  NAND2_X1 U4504 ( .A1(n3591), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3584) );
  OAI21_X1 U4505 ( .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A(n3592), .ZN(n6039) );
  NAND2_X1 U4506 ( .A1(n6039), .A2(n2977), .ZN(n3581) );
  NAND2_X1 U4507 ( .A1(n4066), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3580)
         );
  NAND2_X1 U4508 ( .A1(n3581), .A2(n3580), .ZN(n3582) );
  AOI21_X1 U4509 ( .B1(n4067), .B2(EAX_REG_2__SCAN_IN), .A(n3582), .ZN(n3583)
         );
  AND2_X1 U4510 ( .A1(n3584), .A2(n3583), .ZN(n4375) );
  NAND2_X1 U4511 ( .A1(n3585), .A2(n4375), .ZN(n3589) );
  INV_X1 U4512 ( .A(n3586), .ZN(n4376) );
  INV_X1 U4513 ( .A(n3587), .ZN(n4403) );
  NAND2_X1 U4514 ( .A1(n4376), .A2(n4403), .ZN(n3588) );
  NAND2_X1 U4515 ( .A1(n3589), .A2(n3588), .ZN(n4374) );
  INV_X1 U4516 ( .A(n3591), .ZN(n3600) );
  AOI21_X1 U4517 ( .B1(n4980), .B2(n3592), .A(n3602), .ZN(n4983) );
  OAI22_X1 U4518 ( .A1(n4983), .A2(n4057), .B1(n3760), .B2(n4980), .ZN(n3593)
         );
  AOI21_X1 U4519 ( .B1(n4067), .B2(EAX_REG_3__SCAN_IN), .A(n3593), .ZN(n3594)
         );
  OAI21_X1 U4520 ( .B1(n4680), .B2(n3600), .A(n3594), .ZN(n3595) );
  AOI21_X1 U4521 ( .B1(n2995), .B2(n3745), .A(n3595), .ZN(n4510) );
  INV_X1 U4522 ( .A(n3597), .ZN(n3606) );
  NAND2_X1 U4523 ( .A1(n6210), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3599)
         );
  NAND2_X1 U4524 ( .A1(n4067), .A2(EAX_REG_4__SCAN_IN), .ZN(n3598) );
  OAI211_X1 U4525 ( .C1(n3600), .C2(n5758), .A(n3599), .B(n3598), .ZN(n3601)
         );
  NAND2_X1 U4526 ( .A1(n3601), .A2(n4057), .ZN(n3604) );
  OAI21_X1 U4527 ( .B1(n3602), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n3611), 
        .ZN(n6030) );
  NAND2_X1 U4528 ( .A1(n6030), .A2(n2977), .ZN(n3603) );
  NAND2_X1 U4529 ( .A1(n3604), .A2(n3603), .ZN(n3605) );
  AOI21_X1 U4530 ( .B1(n3606), .B2(n3745), .A(n3605), .ZN(n4397) );
  XNOR2_X1 U4531 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .B(n3611), .ZN(n5012) );
  INV_X1 U4532 ( .A(n3607), .ZN(n3608) );
  NAND2_X1 U4533 ( .A1(n3608), .A2(n3745), .ZN(n3610) );
  AOI22_X1 U4534 ( .A1(n4067), .A2(EAX_REG_5__SCAN_IN), .B1(n4066), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3609) );
  OAI211_X1 U4535 ( .C1(n5012), .C2(n4057), .A(n3610), .B(n3609), .ZN(n4482)
         );
  OAI21_X1 U4536 ( .B1(n3612), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n3633), 
        .ZN(n6023) );
  INV_X1 U4537 ( .A(EAX_REG_6__SCAN_IN), .ZN(n5000) );
  INV_X1 U4538 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3613) );
  OAI22_X1 U4539 ( .A1(n4060), .A2(n5000), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3613), .ZN(n3614) );
  MUX2_X1 U4540 ( .A(n6023), .B(n3614), .S(n4057), .Z(n3615) );
  INV_X1 U4541 ( .A(n3619), .ZN(n3622) );
  XNOR2_X1 U4542 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .B(n3633), .ZN(n5857) );
  AOI22_X1 U4543 ( .A1(n4067), .A2(EAX_REG_7__SCAN_IN), .B1(n4066), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3620) );
  OAI21_X1 U4544 ( .B1(n5857), .B2(n4057), .A(n3620), .ZN(n3621) );
  AOI21_X1 U4545 ( .B1(n3622), .B2(n3745), .A(n3621), .ZN(n4822) );
  AOI22_X1 U4546 ( .A1(n3855), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3993), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3626) );
  AOI22_X1 U4547 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n3836), .B1(n4039), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3625) );
  AOI22_X1 U4548 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n4021), .B1(n3893), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3624) );
  AOI22_X1 U4549 ( .A1(n4046), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3623) );
  NAND4_X1 U4550 ( .A1(n3626), .A2(n3625), .A3(n3624), .A4(n3623), .ZN(n3632)
         );
  AOI22_X1 U4551 ( .A1(n3888), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4019), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3630) );
  AOI22_X1 U4552 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n4018), .B1(n3992), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3629) );
  AOI22_X1 U4553 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n4027), .B1(n4040), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3628) );
  AOI22_X1 U4554 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n3971), .B1(n4020), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3627) );
  NAND4_X1 U4555 ( .A1(n3630), .A2(n3629), .A3(n3628), .A4(n3627), .ZN(n3631)
         );
  NOR2_X1 U4556 ( .A1(n3632), .A2(n3631), .ZN(n3638) );
  INV_X1 U4557 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3635) );
  XNOR2_X1 U4558 ( .A(n3639), .B(n3635), .ZN(n5385) );
  NAND2_X1 U4559 ( .A1(n5385), .A2(n2977), .ZN(n3637) );
  AOI22_X1 U4560 ( .A1(n4067), .A2(EAX_REG_8__SCAN_IN), .B1(n4066), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3636) );
  OAI211_X1 U4561 ( .C1(n3638), .C2(n3716), .A(n3637), .B(n3636), .ZN(n4866)
         );
  XOR2_X1 U4562 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3656), .Z(n5848) );
  INV_X1 U4563 ( .A(n5848), .ZN(n5377) );
  AOI22_X1 U4564 ( .A1(n3855), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3993), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3643) );
  AOI22_X1 U4565 ( .A1(n4021), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3642) );
  AOI22_X1 U4566 ( .A1(n4027), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3893), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3641) );
  AOI22_X1 U4567 ( .A1(n4019), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3640) );
  NAND4_X1 U4568 ( .A1(n3643), .A2(n3642), .A3(n3641), .A4(n3640), .ZN(n3649)
         );
  AOI22_X1 U4569 ( .A1(n3888), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4018), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3647) );
  AOI22_X1 U4570 ( .A1(n3992), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3646) );
  AOI22_X1 U4571 ( .A1(n4039), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4020), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3645) );
  AOI22_X1 U4572 ( .A1(n4046), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3644) );
  NAND4_X1 U4573 ( .A1(n3647), .A2(n3646), .A3(n3645), .A4(n3644), .ZN(n3648)
         );
  NOR2_X1 U4574 ( .A1(n3649), .A2(n3648), .ZN(n3652) );
  NAND2_X1 U4575 ( .A1(n4067), .A2(EAX_REG_9__SCAN_IN), .ZN(n3651) );
  NAND2_X1 U4576 ( .A1(n4066), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3650)
         );
  OAI211_X1 U4577 ( .C1(n3716), .C2(n3652), .A(n3651), .B(n3650), .ZN(n3653)
         );
  AOI21_X1 U4578 ( .B1(n5377), .B2(n2977), .A(n3653), .ZN(n4930) );
  NAND2_X1 U4579 ( .A1(n3655), .A2(n3654), .ZN(n4931) );
  INV_X1 U4580 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3657) );
  XNOR2_X1 U4581 ( .A(n3672), .B(n3657), .ZN(n5368) );
  AOI22_X1 U4582 ( .A1(n3993), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3661) );
  AOI22_X1 U4583 ( .A1(n4018), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3893), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3660) );
  AOI22_X1 U4584 ( .A1(n4019), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3877), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3659) );
  AOI22_X1 U4585 ( .A1(n4021), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4020), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3658) );
  NAND4_X1 U4586 ( .A1(n3661), .A2(n3660), .A3(n3659), .A4(n3658), .ZN(n3667)
         );
  AOI22_X1 U4587 ( .A1(n3836), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4039), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3665) );
  AOI22_X1 U4588 ( .A1(n3855), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3664) );
  AOI22_X1 U4589 ( .A1(n4027), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3663) );
  AOI22_X1 U4590 ( .A1(n3888), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3662) );
  NAND4_X1 U4591 ( .A1(n3665), .A2(n3664), .A3(n3663), .A4(n3662), .ZN(n3666)
         );
  NOR2_X1 U4592 ( .A1(n3667), .A2(n3666), .ZN(n3670) );
  NAND2_X1 U4593 ( .A1(n4067), .A2(EAX_REG_10__SCAN_IN), .ZN(n3669) );
  NAND2_X1 U4594 ( .A1(n4066), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3668)
         );
  OAI211_X1 U4595 ( .C1(n3716), .C2(n3670), .A(n3669), .B(n3668), .ZN(n3671)
         );
  AOI21_X1 U4596 ( .B1(n5368), .B2(n2977), .A(n3671), .ZN(n5002) );
  XOR2_X1 U4597 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3698), .Z(n5838) );
  INV_X1 U4598 ( .A(n5838), .ZN(n6013) );
  AOI22_X1 U4599 ( .A1(n3855), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3993), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3677) );
  AOI22_X1 U4600 ( .A1(n4021), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3888), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3676) );
  AOI22_X1 U4601 ( .A1(n4027), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3675) );
  AOI22_X1 U4602 ( .A1(n4018), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3674) );
  NAND4_X1 U4603 ( .A1(n3677), .A2(n3676), .A3(n3675), .A4(n3674), .ZN(n3683)
         );
  AOI22_X1 U4604 ( .A1(n3836), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4039), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3681) );
  AOI22_X1 U4605 ( .A1(n4019), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3893), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3680) );
  AOI22_X1 U4606 ( .A1(n4040), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3679) );
  AOI22_X1 U4607 ( .A1(n3971), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4020), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3678) );
  NAND4_X1 U4608 ( .A1(n3681), .A2(n3680), .A3(n3679), .A4(n3678), .ZN(n3682)
         );
  NOR2_X1 U4609 ( .A1(n3683), .A2(n3682), .ZN(n3686) );
  NAND2_X1 U4610 ( .A1(n4067), .A2(EAX_REG_11__SCAN_IN), .ZN(n3685) );
  NAND2_X1 U4611 ( .A1(n4066), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3684)
         );
  OAI211_X1 U4612 ( .C1(n3716), .C2(n3686), .A(n3685), .B(n3684), .ZN(n3687)
         );
  AOI21_X1 U4613 ( .B1(n6013), .B2(n2977), .A(n3687), .ZN(n5246) );
  AOI22_X1 U4614 ( .A1(n3855), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3691) );
  AOI22_X1 U4615 ( .A1(n3836), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3690) );
  AOI22_X1 U4616 ( .A1(n3992), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3689) );
  AOI22_X1 U4617 ( .A1(n4018), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3688) );
  NAND4_X1 U4618 ( .A1(n3691), .A2(n3690), .A3(n3689), .A4(n3688), .ZN(n3697)
         );
  AOI22_X1 U4619 ( .A1(n4021), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4039), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3695) );
  AOI22_X1 U4620 ( .A1(n3888), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3893), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3694) );
  AOI22_X1 U4621 ( .A1(n3993), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3693) );
  AOI22_X1 U4622 ( .A1(n4019), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4020), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3692) );
  NAND4_X1 U4623 ( .A1(n3695), .A2(n3694), .A3(n3693), .A4(n3692), .ZN(n3696)
         );
  NOR2_X1 U4624 ( .A1(n3697), .A2(n3696), .ZN(n3701) );
  XNOR2_X1 U4625 ( .A(n3702), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5361)
         );
  NAND2_X1 U4626 ( .A1(n5361), .A2(n2977), .ZN(n3700) );
  AOI22_X1 U4627 ( .A1(n4067), .A2(EAX_REG_12__SCAN_IN), .B1(n4066), .B2(
        PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3699) );
  OAI211_X1 U4628 ( .C1(n3701), .C2(n3716), .A(n3700), .B(n3699), .ZN(n5129)
         );
  XOR2_X1 U4629 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .B(n3719), .Z(n5828) );
  INV_X1 U4630 ( .A(n5828), .ZN(n5353) );
  AOI22_X1 U4631 ( .A1(n3855), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3993), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3706) );
  AOI22_X1 U4632 ( .A1(n3888), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3705) );
  AOI22_X1 U4633 ( .A1(n4019), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3704) );
  AOI22_X1 U4634 ( .A1(n4039), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4020), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3703) );
  NAND4_X1 U4635 ( .A1(n3706), .A2(n3705), .A3(n3704), .A4(n3703), .ZN(n3712)
         );
  AOI22_X1 U4636 ( .A1(n4021), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3710) );
  AOI22_X1 U4637 ( .A1(n4018), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3893), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3709) );
  AOI22_X1 U4638 ( .A1(n4027), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3708) );
  AOI22_X1 U4639 ( .A1(n4046), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3707) );
  NAND4_X1 U4640 ( .A1(n3710), .A2(n3709), .A3(n3708), .A4(n3707), .ZN(n3711)
         );
  NOR2_X1 U4641 ( .A1(n3712), .A2(n3711), .ZN(n3715) );
  NAND2_X1 U4642 ( .A1(n4067), .A2(EAX_REG_13__SCAN_IN), .ZN(n3714) );
  NAND2_X1 U4643 ( .A1(n4066), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3713)
         );
  OAI211_X1 U4644 ( .C1(n3716), .C2(n3715), .A(n3714), .B(n3713), .ZN(n3717)
         );
  AOI21_X1 U4645 ( .B1(n5353), .B2(n2977), .A(n3717), .ZN(n5210) );
  INV_X1 U4646 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5120) );
  XNOR2_X1 U4647 ( .A(n3733), .B(n5120), .ZN(n5345) );
  AOI22_X1 U4648 ( .A1(n4067), .A2(EAX_REG_14__SCAN_IN), .B1(n4066), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3731) );
  AOI22_X1 U4649 ( .A1(n3855), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3723) );
  AOI22_X1 U4650 ( .A1(n3836), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4039), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3722) );
  AOI22_X1 U4651 ( .A1(n3888), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3721) );
  AOI22_X1 U4652 ( .A1(n4021), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4020), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3720) );
  NAND4_X1 U4653 ( .A1(n3723), .A2(n3722), .A3(n3721), .A4(n3720), .ZN(n3729)
         );
  AOI22_X1 U4654 ( .A1(INSTQUEUE_REG_0__6__SCAN_IN), .A2(n4018), .B1(n3893), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3727) );
  AOI22_X1 U4655 ( .A1(n4019), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3726) );
  AOI22_X1 U4656 ( .A1(n3992), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3725) );
  AOI22_X1 U4657 ( .A1(n3993), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3724) );
  NAND4_X1 U4658 ( .A1(n3727), .A2(n3726), .A3(n3725), .A4(n3724), .ZN(n3728)
         );
  OAI21_X1 U4659 ( .B1(n3729), .B2(n3728), .A(n3745), .ZN(n3730) );
  OAI211_X1 U4660 ( .C1(n5345), .C2(n4057), .A(n3731), .B(n3730), .ZN(n3732)
         );
  INV_X1 U4661 ( .A(n3732), .ZN(n5116) );
  XNOR2_X1 U4662 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n3748), .ZN(n5815)
         );
  AOI22_X1 U4663 ( .A1(n3855), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3737) );
  AOI22_X1 U4664 ( .A1(n4018), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3893), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3736) );
  AOI22_X1 U4665 ( .A1(n4021), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3877), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3735) );
  AOI22_X1 U4666 ( .A1(n4046), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3734) );
  NAND4_X1 U4667 ( .A1(n3737), .A2(n3736), .A3(n3735), .A4(n3734), .ZN(n3743)
         );
  AOI22_X1 U4668 ( .A1(n3836), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4039), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3741) );
  AOI22_X1 U4669 ( .A1(n3888), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3740) );
  AOI22_X1 U4670 ( .A1(n3993), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3739) );
  AOI22_X1 U4671 ( .A1(n4019), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4020), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3738) );
  NAND4_X1 U4672 ( .A1(n3741), .A2(n3740), .A3(n3739), .A4(n3738), .ZN(n3742)
         );
  OR2_X1 U4673 ( .A1(n3743), .A2(n3742), .ZN(n3744) );
  AOI22_X1 U4674 ( .A1(n3745), .A2(n3744), .B1(n4066), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3747) );
  NAND2_X1 U4675 ( .A1(n4067), .A2(EAX_REG_15__SCAN_IN), .ZN(n3746) );
  OAI211_X1 U4676 ( .C1(n5815), .C2(n4057), .A(n3747), .B(n3746), .ZN(n5204)
         );
  INV_X1 U4677 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5332) );
  XNOR2_X1 U4678 ( .A(n3780), .B(n5332), .ZN(n5804) );
  AOI22_X1 U4679 ( .A1(n3855), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3993), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3753) );
  AOI22_X1 U4680 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4021), .B1(n3836), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3752) );
  AOI22_X1 U4681 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n3888), .B1(n3971), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3751) );
  AOI22_X1 U4682 ( .A1(n3893), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3750) );
  NAND4_X1 U4683 ( .A1(n3753), .A2(n3752), .A3(n3751), .A4(n3750), .ZN(n3759)
         );
  AOI22_X1 U4684 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4018), .B1(n4019), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3757) );
  AOI22_X1 U4685 ( .A1(n4027), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3756) );
  AOI22_X1 U4686 ( .A1(n3992), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3755) );
  AOI22_X1 U4687 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n4039), .B1(n4020), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3754) );
  NAND4_X1 U4688 ( .A1(n3757), .A2(n3756), .A3(n3755), .A4(n3754), .ZN(n3758)
         );
  OR2_X1 U4689 ( .A1(n3759), .A2(n3758), .ZN(n3763) );
  INV_X1 U4690 ( .A(EAX_REG_16__SCAN_IN), .ZN(n3761) );
  OAI22_X1 U4691 ( .A1(n4060), .A2(n3761), .B1(n3760), .B2(n5332), .ZN(n3762)
         );
  AOI21_X1 U4692 ( .B1(n4062), .B2(n3763), .A(n3762), .ZN(n3764) );
  NAND2_X1 U4693 ( .A1(n3765), .A2(n3764), .ZN(n5193) );
  AOI22_X1 U4694 ( .A1(n4021), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4039), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3769) );
  AOI22_X1 U4695 ( .A1(n4018), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4019), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3768) );
  AOI22_X1 U4696 ( .A1(n3993), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3767) );
  AOI22_X1 U4697 ( .A1(n3893), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3766) );
  NAND4_X1 U4698 ( .A1(n3769), .A2(n3768), .A3(n3767), .A4(n3766), .ZN(n3775)
         );
  AOI22_X1 U4699 ( .A1(n3855), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3773) );
  AOI22_X1 U4700 ( .A1(n3888), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3877), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3772) );
  AOI22_X1 U4701 ( .A1(n3992), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3771) );
  AOI22_X1 U4702 ( .A1(n3836), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3770) );
  NAND4_X1 U4703 ( .A1(n3773), .A2(n3772), .A3(n3771), .A4(n3770), .ZN(n3774)
         );
  NOR2_X1 U4704 ( .A1(n3775), .A2(n3774), .ZN(n3779) );
  OAI21_X1 U4705 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6638), .A(n6210), 
        .ZN(n3776) );
  INV_X1 U4706 ( .A(n3776), .ZN(n3777) );
  AOI21_X1 U4707 ( .B1(n4067), .B2(EAX_REG_17__SCAN_IN), .A(n3777), .ZN(n3778)
         );
  OAI21_X1 U4708 ( .B1(n4036), .B2(n3779), .A(n3778), .ZN(n3783) );
  OAI21_X1 U4709 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n3781), .A(n3801), 
        .ZN(n5791) );
  OR2_X1 U4710 ( .A1(n4057), .A2(n5791), .ZN(n3782) );
  NAND2_X1 U4711 ( .A1(n3783), .A2(n3782), .ZN(n5185) );
  AOI22_X1 U4712 ( .A1(n3888), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4018), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3789) );
  AOI22_X1 U4713 ( .A1(n3836), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4039), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3788) );
  AOI22_X1 U4714 ( .A1(n4019), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4715 ( .A1(n4021), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4020), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3786) );
  NAND4_X1 U4716 ( .A1(n3789), .A2(n3788), .A3(n3787), .A4(n3786), .ZN(n3795)
         );
  AOI22_X1 U4717 ( .A1(n4027), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3993), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4718 ( .A1(n3992), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4719 ( .A1(n3855), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3791) );
  AOI22_X1 U4720 ( .A1(n3893), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3790) );
  NAND4_X1 U4721 ( .A1(n3793), .A2(n3792), .A3(n3791), .A4(n3790), .ZN(n3794)
         );
  NOR2_X1 U4722 ( .A1(n3795), .A2(n3794), .ZN(n3798) );
  INV_X1 U4723 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5327) );
  AOI21_X1 U4724 ( .B1(n5327), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3796) );
  AOI21_X1 U4725 ( .B1(n4067), .B2(EAX_REG_18__SCAN_IN), .A(n3796), .ZN(n3797)
         );
  OAI21_X1 U4726 ( .B1(n4036), .B2(n3798), .A(n3797), .ZN(n3800) );
  XNOR2_X1 U4727 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n3801), .ZN(n5783)
         );
  NAND2_X1 U4728 ( .A1(n5783), .A2(n2977), .ZN(n3799) );
  NAND2_X1 U4729 ( .A1(n3800), .A2(n3799), .ZN(n5179) );
  OR2_X1 U4730 ( .A1(n3802), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3803)
         );
  NAND2_X1 U4731 ( .A1(n3803), .A2(n3851), .ZN(n5684) );
  INV_X1 U4732 ( .A(n5684), .ZN(n3819) );
  AOI22_X1 U4733 ( .A1(n3855), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4734 ( .A1(n3836), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4039), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4735 ( .A1(n3992), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3893), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4736 ( .A1(n4021), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3804) );
  NAND4_X1 U4737 ( .A1(n3807), .A2(n3806), .A3(n3805), .A4(n3804), .ZN(n3813)
         );
  AOI22_X1 U4738 ( .A1(n3888), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4018), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3811) );
  AOI22_X1 U4739 ( .A1(n3993), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4740 ( .A1(n4019), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4020), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4741 ( .A1(n4046), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3808) );
  NAND4_X1 U4742 ( .A1(n3811), .A2(n3810), .A3(n3809), .A4(n3808), .ZN(n3812)
         );
  OR2_X1 U4743 ( .A1(n3813), .A2(n3812), .ZN(n3817) );
  INV_X1 U4744 ( .A(EAX_REG_19__SCAN_IN), .ZN(n3815) );
  NAND2_X1 U4745 ( .A1(n6210), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3814)
         );
  OAI211_X1 U4746 ( .C1(n4060), .C2(n3815), .A(n4057), .B(n3814), .ZN(n3816)
         );
  AOI21_X1 U4747 ( .B1(n4062), .B2(n3817), .A(n3816), .ZN(n3818) );
  AOI21_X1 U4748 ( .B1(n3819), .B2(n2977), .A(n3818), .ZN(n5651) );
  AOI22_X1 U4749 ( .A1(n3888), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4018), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3823) );
  AOI22_X1 U4750 ( .A1(n3836), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4039), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4751 ( .A1(n3992), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4752 ( .A1(n4019), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3820) );
  NAND4_X1 U4753 ( .A1(n3823), .A2(n3822), .A3(n3821), .A4(n3820), .ZN(n3829)
         );
  AOI22_X1 U4754 ( .A1(n4027), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3993), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4755 ( .A1(n4021), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4756 ( .A1(n3893), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3203), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4757 ( .A1(n3855), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3824) );
  NAND4_X1 U4758 ( .A1(n3827), .A2(n3826), .A3(n3825), .A4(n3824), .ZN(n3828)
         );
  NOR2_X1 U4759 ( .A1(n3829), .A2(n3828), .ZN(n3832) );
  INV_X1 U4760 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5646) );
  OAI21_X1 U4761 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5646), .A(n4057), .ZN(
        n3830) );
  AOI21_X1 U4762 ( .B1(n4067), .B2(EAX_REG_20__SCAN_IN), .A(n3830), .ZN(n3831)
         );
  OAI21_X1 U4763 ( .B1(n4036), .B2(n3832), .A(n3831), .ZN(n3834) );
  XNOR2_X1 U4764 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .B(n3851), .ZN(n5638)
         );
  NAND2_X1 U4765 ( .A1(n5638), .A2(n2977), .ZN(n3833) );
  AOI22_X1 U4766 ( .A1(n3888), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4018), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4767 ( .A1(n3836), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4039), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3839) );
  AOI22_X1 U4768 ( .A1(n4019), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3877), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3838) );
  AOI22_X1 U4769 ( .A1(n4021), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3837) );
  NAND4_X1 U4770 ( .A1(n3840), .A2(n3839), .A3(n3838), .A4(n3837), .ZN(n3847)
         );
  AOI22_X1 U4771 ( .A1(n4027), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3993), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4772 ( .A1(n3992), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4773 ( .A1(n3855), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3843) );
  AOI22_X1 U4774 ( .A1(n3893), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3842) );
  NAND4_X1 U4775 ( .A1(n3845), .A2(n3844), .A3(n3843), .A4(n3842), .ZN(n3846)
         );
  NOR2_X1 U4776 ( .A1(n3847), .A2(n3846), .ZN(n3850) );
  AOI21_X1 U4777 ( .B1(n6634), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3848) );
  AOI21_X1 U4778 ( .B1(n4067), .B2(EAX_REG_22__SCAN_IN), .A(n3848), .ZN(n3849)
         );
  OAI21_X1 U4779 ( .B1(n4036), .B2(n3850), .A(n3849), .ZN(n3854) );
  AND2_X1 U4780 ( .A1(n3873), .A2(n6634), .ZN(n3852) );
  NOR2_X1 U4781 ( .A1(n3906), .A2(n3852), .ZN(n5621) );
  NAND2_X1 U4782 ( .A1(n5621), .A2(n2977), .ZN(n3853) );
  NAND2_X1 U4783 ( .A1(n3854), .A2(n3853), .ZN(n5168) );
  AOI22_X1 U4784 ( .A1(n3888), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4019), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4785 ( .A1(n4018), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3893), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4786 ( .A1(n3855), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3857) );
  AOI22_X1 U4787 ( .A1(n3971), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3856) );
  NAND4_X1 U4788 ( .A1(n3859), .A2(n3858), .A3(n3857), .A4(n3856), .ZN(n3865)
         );
  AOI22_X1 U4789 ( .A1(n3836), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4039), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4790 ( .A1(n4027), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3862) );
  AOI22_X1 U4791 ( .A1(n3993), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3861) );
  AOI22_X1 U4792 ( .A1(n4021), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3860) );
  NAND4_X1 U4793 ( .A1(n3863), .A2(n3862), .A3(n3861), .A4(n3860), .ZN(n3864)
         );
  NOR2_X1 U4794 ( .A1(n3865), .A2(n3864), .ZN(n3869) );
  OAI21_X1 U4795 ( .B1(PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6638), .A(n6210), 
        .ZN(n3866) );
  INV_X1 U4796 ( .A(n3866), .ZN(n3867) );
  AOI21_X1 U4797 ( .B1(n4067), .B2(EAX_REG_21__SCAN_IN), .A(n3867), .ZN(n3868)
         );
  OAI21_X1 U4798 ( .B1(n4036), .B2(n3869), .A(n3868), .ZN(n3875) );
  INV_X1 U4799 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n6664) );
  NAND2_X1 U4800 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n3870), .ZN(n3871)
         );
  NAND2_X1 U4801 ( .A1(n6664), .A2(n3871), .ZN(n3872) );
  NAND2_X1 U4802 ( .A1(n3873), .A2(n3872), .ZN(n5632) );
  INV_X1 U4803 ( .A(n5632), .ZN(n5315) );
  NAND2_X1 U4804 ( .A1(n5315), .A2(n2977), .ZN(n3874) );
  NAND2_X1 U4805 ( .A1(n3875), .A2(n3874), .ZN(n5309) );
  AOI22_X1 U4806 ( .A1(n3888), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4018), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3881) );
  AOI22_X1 U4807 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n4039), .B1(n3836), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3880) );
  AOI22_X1 U4808 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4019), .B1(n3877), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3879) );
  AOI22_X1 U4809 ( .A1(n4021), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4020), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3878) );
  NAND4_X1 U4810 ( .A1(n3881), .A2(n3880), .A3(n3879), .A4(n3878), .ZN(n3887)
         );
  AOI22_X1 U4811 ( .A1(n4027), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3993), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3885) );
  AOI22_X1 U4812 ( .A1(n3992), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3884) );
  AOI22_X1 U4813 ( .A1(n3225), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3883) );
  AOI22_X1 U4814 ( .A1(n3893), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3882) );
  NAND4_X1 U4815 ( .A1(n3885), .A2(n3884), .A3(n3883), .A4(n3882), .ZN(n3886)
         );
  OR2_X1 U4816 ( .A1(n3887), .A2(n3886), .ZN(n3901) );
  AOI22_X1 U4817 ( .A1(n3888), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4018), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4818 ( .A1(n3836), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4039), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4819 ( .A1(n3179), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4820 ( .A1(n4021), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4020), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3889) );
  NAND4_X1 U4821 ( .A1(n3892), .A2(n3891), .A3(n3890), .A4(n3889), .ZN(n3899)
         );
  AOI22_X1 U4822 ( .A1(n4027), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3993), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3897) );
  AOI22_X1 U4823 ( .A1(n3992), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3896) );
  INV_X1 U4824 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n6570) );
  AOI22_X1 U4825 ( .A1(n3855), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3895) );
  AOI22_X1 U4826 ( .A1(n3893), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3894) );
  NAND4_X1 U4827 ( .A1(n3897), .A2(n3896), .A3(n3895), .A4(n3894), .ZN(n3898)
         );
  OR2_X1 U4828 ( .A1(n3899), .A2(n3898), .ZN(n3900) );
  NAND2_X1 U4829 ( .A1(n3900), .A2(n3901), .ZN(n3939) );
  OAI21_X1 U4830 ( .B1(n3901), .B2(n3900), .A(n3939), .ZN(n3905) );
  NAND2_X1 U4831 ( .A1(n6210), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3902)
         );
  NAND2_X1 U4832 ( .A1(n4057), .A2(n3902), .ZN(n3903) );
  AOI21_X1 U4833 ( .B1(n4067), .B2(EAX_REG_23__SCAN_IN), .A(n3903), .ZN(n3904)
         );
  OAI21_X1 U4834 ( .B1(n4036), .B2(n3905), .A(n3904), .ZN(n3910) );
  NOR2_X1 U4835 ( .A1(n3906), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3907)
         );
  OR2_X1 U4836 ( .A1(n3944), .A2(n3907), .ZN(n5610) );
  INV_X1 U4837 ( .A(n5610), .ZN(n3908) );
  NAND2_X1 U4838 ( .A1(n3908), .A2(n2977), .ZN(n3909) );
  AOI22_X1 U4839 ( .A1(n3855), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3914) );
  AOI22_X1 U4840 ( .A1(n3836), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4019), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3913) );
  AOI22_X1 U4841 ( .A1(n4018), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3893), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4842 ( .A1(n3203), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3911) );
  NAND4_X1 U4843 ( .A1(n3914), .A2(n3913), .A3(n3912), .A4(n3911), .ZN(n3920)
         );
  AOI22_X1 U4844 ( .A1(n4027), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3888), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3918) );
  AOI22_X1 U4845 ( .A1(n4021), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4039), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3917) );
  AOI22_X1 U4846 ( .A1(n3993), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4847 ( .A1(n3971), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4020), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3915) );
  NAND4_X1 U4848 ( .A1(n3918), .A2(n3917), .A3(n3916), .A4(n3915), .ZN(n3919)
         );
  NOR2_X1 U4849 ( .A1(n3920), .A2(n3919), .ZN(n3940) );
  NAND2_X1 U4850 ( .A1(n3940), .A2(n3939), .ZN(n3921) );
  OAI21_X1 U4851 ( .B1(n3939), .B2(n3940), .A(n3921), .ZN(n3922) );
  INV_X1 U4852 ( .A(n3922), .ZN(n3927) );
  INV_X1 U4853 ( .A(EAX_REG_24__SCAN_IN), .ZN(n3925) );
  NAND2_X1 U4854 ( .A1(n4066), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3924)
         );
  XNOR2_X1 U4855 ( .A(n3944), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5112)
         );
  NAND2_X1 U4856 ( .A1(n5112), .A2(n2977), .ZN(n3923) );
  OAI211_X1 U4857 ( .C1(n4060), .C2(n3925), .A(n3924), .B(n3923), .ZN(n3926)
         );
  AOI21_X1 U4858 ( .B1(n4062), .B2(n3927), .A(n3926), .ZN(n4090) );
  AOI22_X1 U4859 ( .A1(n3888), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4018), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3932) );
  AOI22_X1 U4860 ( .A1(n3836), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4039), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3931) );
  AOI22_X1 U4861 ( .A1(n3179), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3930) );
  AOI22_X1 U4862 ( .A1(n4021), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4020), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3929) );
  NAND4_X1 U4863 ( .A1(n3932), .A2(n3931), .A3(n3930), .A4(n3929), .ZN(n3938)
         );
  AOI22_X1 U4864 ( .A1(n4027), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3993), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3936) );
  AOI22_X1 U4865 ( .A1(n3992), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3935) );
  AOI22_X1 U4866 ( .A1(n3855), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3934) );
  AOI22_X1 U4867 ( .A1(n3893), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3933) );
  NAND4_X1 U4868 ( .A1(n3936), .A2(n3935), .A3(n3934), .A4(n3933), .ZN(n3937)
         );
  OR2_X1 U4869 ( .A1(n3938), .A2(n3937), .ZN(n3959) );
  NOR2_X1 U4870 ( .A1(n3940), .A2(n3939), .ZN(n3960) );
  XNOR2_X1 U4871 ( .A(n3959), .B(n3960), .ZN(n3943) );
  INV_X1 U4872 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5102) );
  AOI21_X1 U4873 ( .B1(n5102), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3941) );
  AOI21_X1 U4874 ( .B1(n4067), .B2(EAX_REG_25__SCAN_IN), .A(n3941), .ZN(n3942)
         );
  OAI21_X1 U4875 ( .B1(n4036), .B2(n3943), .A(n3942), .ZN(n3948) );
  OR2_X1 U4876 ( .A1(n3945), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3946)
         );
  NAND2_X1 U4877 ( .A1(n3946), .A2(n3963), .ZN(n5677) );
  INV_X1 U4878 ( .A(n5677), .ZN(n5104) );
  NAND2_X1 U4879 ( .A1(n5104), .A2(n2977), .ZN(n3947) );
  NAND2_X1 U4880 ( .A1(n3948), .A2(n3947), .ZN(n5095) );
  AOI22_X1 U4881 ( .A1(n3855), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3993), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3952) );
  AOI22_X1 U4882 ( .A1(n3888), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3893), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3951) );
  AOI22_X1 U4883 ( .A1(n4039), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3950) );
  AOI22_X1 U4884 ( .A1(n3992), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3949) );
  NAND4_X1 U4885 ( .A1(n3952), .A2(n3951), .A3(n3950), .A4(n3949), .ZN(n3958)
         );
  AOI22_X1 U4886 ( .A1(n4021), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3956) );
  AOI22_X1 U4887 ( .A1(n4027), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U4888 ( .A1(n3179), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3954) );
  AOI22_X1 U4889 ( .A1(n4018), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3953) );
  NAND4_X1 U4890 ( .A1(n3956), .A2(n3955), .A3(n3954), .A4(n3953), .ZN(n3957)
         );
  NOR2_X1 U4891 ( .A1(n3958), .A2(n3957), .ZN(n3970) );
  NAND2_X1 U4892 ( .A1(n3960), .A2(n3959), .ZN(n3969) );
  XOR2_X1 U4893 ( .A(n3970), .B(n3969), .Z(n3961) );
  NAND2_X1 U4894 ( .A1(n3961), .A2(n4062), .ZN(n3968) );
  INV_X1 U4895 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6668) );
  OAI21_X1 U4896 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6668), .A(n4057), .ZN(
        n3962) );
  AOI21_X1 U4897 ( .B1(n4067), .B2(EAX_REG_26__SCAN_IN), .A(n3962), .ZN(n3967)
         );
  NOR2_X1 U4898 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n3964), .ZN(n3965)
         );
  NOR2_X1 U4899 ( .A1(n3986), .A2(n3965), .ZN(n5597) );
  AND2_X1 U4900 ( .A1(n5597), .A2(n2977), .ZN(n3966) );
  AOI21_X1 U4901 ( .B1(n3968), .B2(n3967), .A(n3966), .ZN(n5154) );
  NOR2_X1 U4902 ( .A1(n3970), .A2(n3969), .ZN(n3991) );
  AOI22_X1 U4903 ( .A1(n3888), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4018), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3975) );
  AOI22_X1 U4904 ( .A1(n3836), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4039), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3974) );
  AOI22_X1 U4905 ( .A1(n4019), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3973) );
  AOI22_X1 U4906 ( .A1(n4021), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3972) );
  NAND4_X1 U4907 ( .A1(n3975), .A2(n3974), .A3(n3973), .A4(n3972), .ZN(n3981)
         );
  AOI22_X1 U4908 ( .A1(n4027), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3993), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3979) );
  AOI22_X1 U4909 ( .A1(n3992), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U4910 ( .A1(n3225), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U4911 ( .A1(n3893), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3976) );
  NAND4_X1 U4912 ( .A1(n3979), .A2(n3978), .A3(n3977), .A4(n3976), .ZN(n3980)
         );
  OR2_X1 U4913 ( .A1(n3981), .A2(n3980), .ZN(n3990) );
  INV_X1 U4914 ( .A(n3990), .ZN(n3982) );
  XNOR2_X1 U4915 ( .A(n3991), .B(n3982), .ZN(n3983) );
  NAND2_X1 U4916 ( .A1(n3983), .A2(n4062), .ZN(n3989) );
  NAND2_X1 U4917 ( .A1(n6210), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3984)
         );
  NAND2_X1 U4918 ( .A1(n4057), .A2(n3984), .ZN(n3985) );
  AOI21_X1 U4919 ( .B1(n4067), .B2(EAX_REG_27__SCAN_IN), .A(n3985), .ZN(n3988)
         );
  OAI21_X1 U4920 ( .B1(n3986), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n4012), 
        .ZN(n5282) );
  NOR2_X1 U4921 ( .A1(n5282), .A2(n4057), .ZN(n3987) );
  AOI21_X1 U4922 ( .B1(n3989), .B2(n3988), .A(n3987), .ZN(n5085) );
  NAND2_X1 U4923 ( .A1(n3991), .A2(n3990), .ZN(n4016) );
  AOI22_X1 U4924 ( .A1(n4018), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3997) );
  AOI22_X1 U4925 ( .A1(n4027), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3996) );
  AOI22_X1 U4926 ( .A1(n3893), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3995) );
  AOI22_X1 U4927 ( .A1(n3993), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3994) );
  NAND4_X1 U4928 ( .A1(n3997), .A2(n3996), .A3(n3995), .A4(n3994), .ZN(n4003)
         );
  AOI22_X1 U4929 ( .A1(n4021), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4039), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4001) );
  AOI22_X1 U4930 ( .A1(n3888), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4019), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4000) );
  AOI22_X1 U4931 ( .A1(n3225), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3999) );
  AOI22_X1 U4932 ( .A1(n3971), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3998) );
  NAND4_X1 U4933 ( .A1(n4001), .A2(n4000), .A3(n3999), .A4(n3998), .ZN(n4002)
         );
  NOR2_X1 U4934 ( .A1(n4003), .A2(n4002), .ZN(n4017) );
  XOR2_X1 U4935 ( .A(n4016), .B(n4017), .Z(n4004) );
  NAND2_X1 U4936 ( .A1(n4004), .A2(n4062), .ZN(n4008) );
  NAND2_X1 U4937 ( .A1(n6210), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4005)
         );
  NAND2_X1 U4938 ( .A1(n4057), .A2(n4005), .ZN(n4006) );
  AOI21_X1 U4939 ( .B1(n4067), .B2(EAX_REG_28__SCAN_IN), .A(n4006), .ZN(n4007)
         );
  NAND2_X1 U4940 ( .A1(n4008), .A2(n4007), .ZN(n4010) );
  XNOR2_X1 U4941 ( .A(n4012), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5588)
         );
  NAND2_X1 U4942 ( .A1(n5588), .A2(n2977), .ZN(n4009) );
  NAND2_X1 U4943 ( .A1(n4010), .A2(n4009), .ZN(n5144) );
  INV_X1 U4944 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4011) );
  INV_X1 U4945 ( .A(n4013), .ZN(n4014) );
  INV_X1 U4946 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5078) );
  NAND2_X1 U4947 ( .A1(n4014), .A2(n5078), .ZN(n4015) );
  NAND2_X1 U4948 ( .A1(n4076), .A2(n4015), .ZN(n5266) );
  NOR2_X1 U4949 ( .A1(n4017), .A2(n4016), .ZN(n4054) );
  AOI22_X1 U4950 ( .A1(n3888), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4018), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4025) );
  AOI22_X1 U4951 ( .A1(n3836), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4039), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4024) );
  AOI22_X1 U4952 ( .A1(n4019), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4023) );
  AOI22_X1 U4953 ( .A1(n4021), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4020), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4022) );
  NAND4_X1 U4954 ( .A1(n4025), .A2(n4024), .A3(n4023), .A4(n4022), .ZN(n4033)
         );
  AOI22_X1 U4955 ( .A1(n4027), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4026), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4031) );
  AOI22_X1 U4956 ( .A1(n3992), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4030) );
  AOI22_X1 U4957 ( .A1(n3225), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4029) );
  AOI22_X1 U4958 ( .A1(n3893), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4028) );
  NAND4_X1 U4959 ( .A1(n4031), .A2(n4030), .A3(n4029), .A4(n4028), .ZN(n4032)
         );
  OR2_X1 U4960 ( .A1(n4033), .A2(n4032), .ZN(n4053) );
  XNOR2_X1 U4961 ( .A(n4054), .B(n4053), .ZN(n4037) );
  AOI21_X1 U4962 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6210), .A(n2977), 
        .ZN(n4035) );
  NAND2_X1 U4963 ( .A1(n4067), .A2(EAX_REG_29__SCAN_IN), .ZN(n4034) );
  OAI211_X1 U4964 ( .C1(n4037), .C2(n4036), .A(n4035), .B(n4034), .ZN(n4038)
         );
  OAI21_X1 U4965 ( .B1(n4057), .B2(n5266), .A(n4038), .ZN(n5069) );
  XNOR2_X1 U4966 ( .A(n4076), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5058)
         );
  AOI22_X1 U4967 ( .A1(n3141), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3888), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4045) );
  AOI22_X1 U4968 ( .A1(n3836), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4039), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U4969 ( .A1(n3993), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U4970 ( .A1(n3893), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4042) );
  NAND4_X1 U4971 ( .A1(n4045), .A2(n4044), .A3(n4043), .A4(n4042), .ZN(n4052)
         );
  AOI22_X1 U4972 ( .A1(n3225), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4050) );
  AOI22_X1 U4973 ( .A1(n4018), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4019), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4049) );
  AOI22_X1 U4974 ( .A1(n3992), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4046), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4048) );
  AOI22_X1 U4975 ( .A1(n3971), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4047) );
  NAND4_X1 U4976 ( .A1(n4050), .A2(n4049), .A3(n4048), .A4(n4047), .ZN(n4051)
         );
  NOR2_X1 U4977 ( .A1(n4052), .A2(n4051), .ZN(n4056) );
  NAND2_X1 U4978 ( .A1(n4054), .A2(n4053), .ZN(n4055) );
  XOR2_X1 U4979 ( .A(n4056), .B(n4055), .Z(n4063) );
  INV_X1 U4980 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4059) );
  NAND2_X1 U4981 ( .A1(n6210), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4058)
         );
  OAI211_X1 U4982 ( .C1(n4060), .C2(n4059), .A(n4058), .B(n4057), .ZN(n4061)
         );
  AOI21_X1 U4983 ( .B1(n4063), .B2(n4062), .A(n4061), .ZN(n4064) );
  AOI21_X1 U4984 ( .B1(n2977), .B2(n5058), .A(n4064), .ZN(n5048) );
  NAND2_X1 U4985 ( .A1(n5068), .A2(n5048), .ZN(n4070) );
  AOI22_X1 U4986 ( .A1(n4067), .A2(EAX_REG_31__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n4066), .ZN(n4068) );
  INV_X1 U4987 ( .A(n4068), .ZN(n4069) );
  XNOR2_X2 U4988 ( .A(n4070), .B(n4069), .ZN(n5031) );
  AND2_X1 U4989 ( .A1(n6509), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4838) );
  NAND2_X1 U4990 ( .A1(n4838), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6406) );
  NOR2_X2 U4991 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6245) );
  NAND2_X1 U4992 ( .A1(n5031), .A2(n6035), .ZN(n4082) );
  AND2_X1 U4993 ( .A1(n4078), .A2(n6295), .ZN(n6512) );
  INV_X1 U4994 ( .A(n6512), .ZN(n4071) );
  NAND2_X1 U4995 ( .A1(n4071), .A2(n6509), .ZN(n4072) );
  NAND2_X1 U4996 ( .A1(n6509), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4074) );
  NAND2_X1 U4997 ( .A1(n6638), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4073) );
  NAND2_X1 U4998 ( .A1(n4074), .A2(n4073), .ZN(n6046) );
  INV_X1 U4999 ( .A(n6046), .ZN(n4075) );
  INV_X1 U5000 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5059) );
  INV_X1 U5001 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5039) );
  NAND2_X1 U5002 ( .A1(n6112), .A2(REIP_REG_31__SCAN_IN), .ZN(n4266) );
  NAND2_X1 U5003 ( .A1(n6047), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4079)
         );
  OAI211_X1 U5004 ( .C1(n6040), .C2(n4856), .A(n4266), .B(n4079), .ZN(n4080)
         );
  INV_X1 U5005 ( .A(n4080), .ZN(n4081) );
  OAI211_X1 U5006 ( .C1(n4272), .C2(n6041), .A(n4082), .B(n4081), .ZN(U2955)
         );
  NAND2_X1 U5007 ( .A1(n5686), .A2(n5318), .ZN(n4084) );
  XNOR2_X1 U5008 ( .A(n5686), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5313)
         );
  NAND2_X1 U5009 ( .A1(n4085), .A2(n5304), .ZN(n5295) );
  NAND2_X1 U5010 ( .A1(n5686), .A2(n5460), .ZN(n4087) );
  NAND3_X1 U5011 ( .A1(n5686), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4088) );
  INV_X1 U5012 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4089) );
  OAI21_X1 U5013 ( .B1(n2981), .B2(n3928), .A(n4091), .ZN(n5232) );
  INV_X1 U5014 ( .A(REIP_REG_24__SCAN_IN), .ZN(n4092) );
  NOR2_X1 U5015 ( .A1(n6071), .A2(n4092), .ZN(n5449) );
  NOR2_X1 U5016 ( .A1(n6040), .A2(n5112), .ZN(n4093) );
  AOI211_X1 U5017 ( .C1(n6047), .C2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5449), 
        .B(n4093), .ZN(n4094) );
  INV_X1 U5018 ( .A(n4097), .ZN(n4098) );
  INV_X1 U5019 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6420) );
  NAND2_X1 U5020 ( .A1(n4098), .A2(n6420), .ZN(n6413) );
  NAND2_X1 U5021 ( .A1(n4103), .A2(n6413), .ZN(n4853) );
  NAND3_X1 U5022 ( .A1(n4346), .A2(n4853), .A3(n6599), .ZN(n4099) );
  NAND3_X1 U5023 ( .A1(n4099), .A2(n4852), .A3(n5028), .ZN(n4100) );
  NAND2_X1 U5024 ( .A1(n4100), .A2(n4381), .ZN(n4101) );
  NOR2_X1 U5025 ( .A1(n4830), .A2(n4101), .ZN(n4120) );
  INV_X1 U5026 ( .A(n6367), .ZN(n4102) );
  OR3_X1 U5027 ( .A1(n4379), .A2(n4103), .A3(n4102), .ZN(n4118) );
  INV_X1 U5028 ( .A(n4276), .ZN(n4283) );
  AND2_X1 U5029 ( .A1(n3248), .A2(n4852), .ZN(n4105) );
  NAND2_X1 U5030 ( .A1(n4105), .A2(n4104), .ZN(n4235) );
  NAND2_X1 U5031 ( .A1(n4235), .A2(n4106), .ZN(n4107) );
  OR2_X1 U5032 ( .A1(n4334), .A2(n4107), .ZN(n4108) );
  NAND2_X1 U5033 ( .A1(n4283), .A2(n4108), .ZN(n4332) );
  NAND2_X1 U5034 ( .A1(n4407), .A2(n6413), .ZN(n4115) );
  NOR3_X1 U5035 ( .A1(n4111), .A2(n4110), .A3(n4109), .ZN(n4114) );
  AOI21_X1 U5036 ( .B1(n4114), .B2(n4113), .A(n4112), .ZN(n4284) );
  AND2_X1 U5037 ( .A1(n4284), .A2(n6599), .ZN(n4335) );
  NAND3_X1 U5038 ( .A1(n4115), .A2(n3165), .A3(n4335), .ZN(n4116) );
  AOI21_X1 U5039 ( .B1(n4118), .B2(n4117), .A(n6400), .ZN(n4119) );
  NOR2_X1 U5040 ( .A1(n4121), .A2(n4831), .ZN(n4122) );
  OR2_X1 U5041 ( .A1(n4334), .A2(n4122), .ZN(n4281) );
  NAND2_X1 U5042 ( .A1(n4346), .A2(n4849), .ZN(n4829) );
  NAND2_X1 U5043 ( .A1(n4227), .A2(n3239), .ZN(n4123) );
  NAND4_X1 U5044 ( .A1(n4281), .A2(n4653), .A3(n4829), .A4(n4123), .ZN(n4124)
         );
  NAND2_X1 U5045 ( .A1(n4380), .A2(n4852), .ZN(n4127) );
  MUX2_X1 U5046 ( .A(n5073), .B(n4127), .S(EBX_REG_1__SCAN_IN), .Z(n4126) );
  NAND2_X1 U5047 ( .A1(n4325), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4125)
         );
  NAND2_X1 U5048 ( .A1(n4126), .A2(n4125), .ZN(n4131) );
  NAND2_X1 U5049 ( .A1(n4127), .A2(EBX_REG_0__SCAN_IN), .ZN(n4129) );
  INV_X1 U5050 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5895) );
  NAND2_X1 U5051 ( .A1(n4218), .A2(n5895), .ZN(n4128) );
  NAND2_X1 U5052 ( .A1(n4129), .A2(n4128), .ZN(n4298) );
  XNOR2_X1 U5053 ( .A(n4131), .B(n4298), .ZN(n4847) );
  INV_X1 U5054 ( .A(n4298), .ZN(n4130) );
  NOR2_X1 U5055 ( .A1(n4131), .A2(n4130), .ZN(n4132) );
  AOI21_X1 U5056 ( .B1(n4847), .B2(n4849), .A(n4132), .ZN(n4390) );
  NAND2_X1 U5057 ( .A1(n4127), .A2(n3422), .ZN(n4134) );
  INV_X1 U5058 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4939) );
  NAND2_X1 U5059 ( .A1(n4849), .A2(n4939), .ZN(n4133) );
  NAND3_X1 U5060 ( .A1(n4134), .A2(n5073), .A3(n4133), .ZN(n4136) );
  NAND2_X1 U5061 ( .A1(n5181), .A2(n4939), .ZN(n4135) );
  NAND2_X1 U5062 ( .A1(n4136), .A2(n4135), .ZN(n4389) );
  NAND2_X1 U5063 ( .A1(n4390), .A2(n4389), .ZN(n4512) );
  INV_X1 U5064 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4981) );
  NAND2_X1 U5065 ( .A1(n4849), .A2(n4981), .ZN(n4138) );
  NAND2_X1 U5066 ( .A1(n5073), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4137)
         );
  NAND3_X1 U5067 ( .A1(n4138), .A2(n4127), .A3(n4137), .ZN(n4139) );
  OAI21_X1 U5068 ( .B1(n4208), .B2(EBX_REG_3__SCAN_IN), .A(n4139), .ZN(n4511)
         );
  INV_X1 U5069 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U5070 ( .A1(n4127), .A2(n6097), .ZN(n4141) );
  INV_X1 U5071 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4142) );
  NAND2_X1 U5072 ( .A1(n4849), .A2(n4142), .ZN(n4140) );
  NAND3_X1 U5073 ( .A1(n4141), .A2(n5073), .A3(n4140), .ZN(n4144) );
  NAND2_X1 U5074 ( .A1(n5181), .A2(n4142), .ZN(n4143) );
  AND2_X1 U5075 ( .A1(n4144), .A2(n4143), .ZN(n4398) );
  INV_X1 U5076 ( .A(n4208), .ZN(n4201) );
  INV_X1 U5077 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4924) );
  NAND2_X1 U5078 ( .A1(n4201), .A2(n4924), .ZN(n4148) );
  NAND2_X1 U5079 ( .A1(n4849), .A2(n4924), .ZN(n4146) );
  NAND2_X1 U5080 ( .A1(n5073), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4145)
         );
  NAND3_X1 U5081 ( .A1(n4146), .A2(n4127), .A3(n4145), .ZN(n4147) );
  MUX2_X1 U5082 ( .A(n5073), .B(n4127), .S(EBX_REG_6__SCAN_IN), .Z(n4150) );
  NAND2_X1 U5083 ( .A1(n4325), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4149)
         );
  NAND2_X1 U5084 ( .A1(n4150), .A2(n4149), .ZN(n4760) );
  INV_X1 U5085 ( .A(EBX_REG_7__SCAN_IN), .ZN(n6576) );
  NAND2_X1 U5086 ( .A1(n4849), .A2(n6576), .ZN(n4152) );
  NAND2_X1 U5087 ( .A1(n5073), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4151)
         );
  NAND3_X1 U5088 ( .A1(n4152), .A2(n4127), .A3(n4151), .ZN(n4153) );
  OAI21_X1 U5089 ( .B1(n4208), .B2(EBX_REG_7__SCAN_IN), .A(n4153), .ZN(n4825)
         );
  MUX2_X1 U5090 ( .A(n5073), .B(n4127), .S(EBX_REG_8__SCAN_IN), .Z(n4155) );
  NAND2_X1 U5091 ( .A1(n4325), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4154)
         );
  MUX2_X1 U5092 ( .A(n4208), .B(n5073), .S(EBX_REG_9__SCAN_IN), .Z(n4156) );
  OAI21_X1 U5093 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n4299), .A(n4156), 
        .ZN(n4933) );
  MUX2_X1 U5094 ( .A(n5073), .B(n4127), .S(EBX_REG_10__SCAN_IN), .Z(n4158) );
  NAND2_X1 U5095 ( .A1(n4325), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4157) );
  NAND2_X1 U5096 ( .A1(n4158), .A2(n4157), .ZN(n5513) );
  INV_X1 U5097 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5906) );
  NAND2_X1 U5098 ( .A1(n4201), .A2(n5906), .ZN(n4162) );
  NAND2_X1 U5099 ( .A1(n4849), .A2(n5906), .ZN(n4160) );
  NAND2_X1 U5100 ( .A1(n5073), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4159) );
  NAND3_X1 U5101 ( .A1(n4160), .A2(n4127), .A3(n4159), .ZN(n4161) );
  AND2_X1 U5102 ( .A1(n4162), .A2(n4161), .ZN(n5512) );
  MUX2_X1 U5103 ( .A(n5073), .B(n4127), .S(EBX_REG_12__SCAN_IN), .Z(n4165) );
  NAND2_X1 U5104 ( .A1(n4325), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4164) );
  NAND2_X1 U5105 ( .A1(n4165), .A2(n4164), .ZN(n5128) );
  MUX2_X1 U5106 ( .A(n4208), .B(n5073), .S(EBX_REG_13__SCAN_IN), .Z(n4166) );
  OAI21_X1 U5107 ( .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n4299), .A(n4166), 
        .ZN(n5206) );
  NAND2_X1 U5108 ( .A1(n4127), .A2(n4167), .ZN(n4169) );
  INV_X1 U5109 ( .A(EBX_REG_14__SCAN_IN), .ZN(n4170) );
  NAND2_X1 U5110 ( .A1(n4849), .A2(n4170), .ZN(n4168) );
  NAND3_X1 U5111 ( .A1(n4169), .A2(n5073), .A3(n4168), .ZN(n4172) );
  NAND2_X1 U5112 ( .A1(n5181), .A2(n4170), .ZN(n4171) );
  MUX2_X1 U5113 ( .A(n4208), .B(n5073), .S(EBX_REG_15__SCAN_IN), .Z(n4174) );
  OR2_X1 U5114 ( .A1(n4299), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4173)
         );
  INV_X1 U5115 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6557) );
  NAND2_X1 U5116 ( .A1(n4127), .A2(n6557), .ZN(n4176) );
  INV_X1 U5117 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5806) );
  NAND2_X1 U5118 ( .A1(n4849), .A2(n5806), .ZN(n4175) );
  NAND3_X1 U5119 ( .A1(n4176), .A2(n5073), .A3(n4175), .ZN(n4178) );
  NAND2_X1 U5120 ( .A1(n5181), .A2(n5806), .ZN(n4177) );
  NAND2_X1 U5121 ( .A1(n4178), .A2(n4177), .ZN(n5194) );
  MUX2_X1 U5122 ( .A(n4208), .B(n5073), .S(EBX_REG_17__SCAN_IN), .Z(n4179) );
  OAI21_X1 U5123 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n4299), .A(n4179), 
        .ZN(n5188) );
  NAND2_X1 U5124 ( .A1(n4127), .A2(n5678), .ZN(n4181) );
  INV_X1 U5125 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5664) );
  NAND2_X1 U5126 ( .A1(n4849), .A2(n5664), .ZN(n4180) );
  NAND3_X1 U5127 ( .A1(n4181), .A2(n5073), .A3(n4180), .ZN(n4183) );
  NAND2_X1 U5128 ( .A1(n5181), .A2(n5664), .ZN(n4182) );
  OR2_X1 U5129 ( .A1(n4299), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4185)
         );
  INV_X1 U5130 ( .A(EBX_REG_20__SCAN_IN), .ZN(n4188) );
  NAND2_X1 U5131 ( .A1(n4849), .A2(n4188), .ZN(n4184) );
  NAND2_X1 U5132 ( .A1(n4185), .A2(n4184), .ZN(n5177) );
  NAND2_X1 U5133 ( .A1(n4299), .A2(EBX_REG_18__SCAN_IN), .ZN(n4187) );
  NAND2_X1 U5134 ( .A1(n4325), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4186) );
  NAND2_X1 U5135 ( .A1(n4187), .A2(n4186), .ZN(n5182) );
  MUX2_X1 U5136 ( .A(n5073), .B(n5177), .S(n5182), .Z(n4190) );
  NOR2_X1 U5137 ( .A1(n5073), .A2(n4188), .ZN(n4189) );
  NOR2_X1 U5138 ( .A1(n4190), .A2(n4189), .ZN(n4191) );
  MUX2_X1 U5139 ( .A(n4208), .B(n5073), .S(EBX_REG_21__SCAN_IN), .Z(n4193) );
  OR2_X1 U5140 ( .A1(n4299), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4192)
         );
  NAND2_X1 U5141 ( .A1(n4127), .A2(n5459), .ZN(n4195) );
  INV_X1 U5142 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5172) );
  NAND2_X1 U5143 ( .A1(n4849), .A2(n5172), .ZN(n4194) );
  NAND3_X1 U5144 ( .A1(n4195), .A2(n5073), .A3(n4194), .ZN(n4197) );
  NAND2_X1 U5145 ( .A1(n5181), .A2(n5172), .ZN(n4196) );
  AND2_X1 U5146 ( .A1(n4197), .A2(n4196), .ZN(n5169) );
  MUX2_X1 U5147 ( .A(n4208), .B(n5073), .S(EBX_REG_23__SCAN_IN), .Z(n4198) );
  OAI21_X1 U5148 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n4299), .A(n4198), 
        .ZN(n5165) );
  MUX2_X1 U5149 ( .A(n5073), .B(n4127), .S(EBX_REG_24__SCAN_IN), .Z(n4200) );
  NAND2_X1 U5150 ( .A1(n4325), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4199) );
  NAND2_X1 U5151 ( .A1(n4200), .A2(n4199), .ZN(n5110) );
  INV_X1 U5152 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5106) );
  NAND2_X1 U5153 ( .A1(n4201), .A2(n5106), .ZN(n4205) );
  NAND2_X1 U5154 ( .A1(n4849), .A2(n5106), .ZN(n4203) );
  NAND2_X1 U5155 ( .A1(n5073), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4202) );
  NAND3_X1 U5156 ( .A1(n4203), .A2(n4127), .A3(n4202), .ZN(n4204) );
  AND2_X1 U5157 ( .A1(n4205), .A2(n4204), .ZN(n5099) );
  MUX2_X1 U5158 ( .A(n5073), .B(n4127), .S(EBX_REG_26__SCAN_IN), .Z(n4207) );
  NAND2_X1 U5159 ( .A1(n4325), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4206) );
  NAND2_X1 U5160 ( .A1(n4207), .A2(n4206), .ZN(n5155) );
  MUX2_X1 U5161 ( .A(n4208), .B(n5073), .S(EBX_REG_27__SCAN_IN), .Z(n4209) );
  OAI21_X1 U5162 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n4299), .A(n4209), 
        .ZN(n5087) );
  NAND2_X1 U5163 ( .A1(n4127), .A2(n4210), .ZN(n4212) );
  INV_X1 U5164 ( .A(EBX_REG_28__SCAN_IN), .ZN(n4213) );
  NAND2_X1 U5165 ( .A1(n4849), .A2(n4213), .ZN(n4211) );
  NAND3_X1 U5166 ( .A1(n4212), .A2(n5073), .A3(n4211), .ZN(n4215) );
  NAND2_X1 U5167 ( .A1(n5181), .A2(n4213), .ZN(n4214) );
  AND2_X1 U5168 ( .A1(n4215), .A2(n4214), .ZN(n5147) );
  OR2_X1 U5169 ( .A1(n4299), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4217)
         );
  INV_X1 U5170 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5143) );
  NAND2_X1 U5171 ( .A1(n4849), .A2(n5143), .ZN(n4216) );
  NAND2_X1 U5172 ( .A1(n4217), .A2(n4216), .ZN(n5071) );
  NAND2_X1 U5173 ( .A1(n5055), .A2(n4218), .ZN(n4220) );
  INV_X1 U5174 ( .A(n5149), .ZN(n5052) );
  NOR2_X1 U5175 ( .A1(n5073), .A2(EBX_REG_29__SCAN_IN), .ZN(n5072) );
  NAND2_X1 U5176 ( .A1(n5052), .A2(n5072), .ZN(n4219) );
  NAND2_X1 U5177 ( .A1(n4220), .A2(n4219), .ZN(n5077) );
  NAND2_X1 U5178 ( .A1(n4299), .A2(EBX_REG_30__SCAN_IN), .ZN(n4222) );
  NAND2_X1 U5179 ( .A1(n4325), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4221) );
  AND2_X1 U5180 ( .A1(n4222), .A2(n4221), .ZN(n5053) );
  NAND2_X1 U5181 ( .A1(n5077), .A2(n5053), .ZN(n4223) );
  INV_X1 U5182 ( .A(n5055), .ZN(n5051) );
  NAND2_X1 U5183 ( .A1(n5051), .A2(n5073), .ZN(n5054) );
  NAND2_X1 U5184 ( .A1(n4223), .A2(n5054), .ZN(n4225) );
  OAI22_X1 U5185 ( .A1(n4299), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n4325), .B2(EBX_REG_31__SCAN_IN), .ZN(n4224) );
  XNOR2_X1 U5186 ( .A(n4225), .B(n4224), .ZN(n5141) );
  INV_X1 U5187 ( .A(n5141), .ZN(n4270) );
  NAND2_X1 U5188 ( .A1(n4227), .A2(n4226), .ZN(n4228) );
  NAND2_X1 U5189 ( .A1(n4346), .A2(n6507), .ZN(n6391) );
  NAND2_X1 U5190 ( .A1(n4228), .A2(n6391), .ZN(n4229) );
  AND2_X1 U5191 ( .A1(n4230), .A2(n5181), .ZN(n4231) );
  NOR2_X1 U5192 ( .A1(n4843), .A2(n3165), .ZN(n4330) );
  OAI21_X1 U5193 ( .B1(n4330), .B2(n4299), .A(n4232), .ZN(n4236) );
  NAND2_X1 U5194 ( .A1(n5028), .A2(n3165), .ZN(n4234) );
  NAND2_X1 U5195 ( .A1(n3258), .A2(n5181), .ZN(n4233) );
  AND4_X1 U5196 ( .A1(n4236), .A2(n4235), .A3(n4234), .A4(n4233), .ZN(n4237)
         );
  NAND2_X1 U5197 ( .A1(n4238), .A2(n4237), .ZN(n4348) );
  NOR2_X1 U5198 ( .A1(n4411), .A2(n4852), .ZN(n4239) );
  NAND2_X1 U5199 ( .A1(n6367), .A2(n4239), .ZN(n4678) );
  OAI22_X1 U5200 ( .A1(n4344), .A2(n3261), .B1(n4343), .B2(n4852), .ZN(n4240)
         );
  INV_X1 U5201 ( .A(n4240), .ZN(n4241) );
  NAND2_X1 U5202 ( .A1(n4678), .A2(n4241), .ZN(n4242) );
  NAND2_X1 U5203 ( .A1(n4246), .A2(n4243), .ZN(n5479) );
  NAND2_X1 U5204 ( .A1(n6088), .A2(n5479), .ZN(n5482) );
  INV_X1 U5205 ( .A(n5730), .ZN(n6059) );
  INV_X1 U5206 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4770) );
  INV_X1 U5207 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6667) );
  OAI21_X1 U5208 ( .B1(n4342), .B2(n6667), .A(n3422), .ZN(n6091) );
  NAND3_X1 U5209 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n6091), .ZN(n4769) );
  NOR2_X1 U5210 ( .A1(n4770), .A2(n4769), .ZN(n4767) );
  NAND2_X1 U5211 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4767), .ZN(n6058)
         );
  INV_X1 U5212 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6086) );
  NOR2_X1 U5213 ( .A1(n3496), .A2(n6086), .ZN(n6075) );
  NAND3_X1 U5214 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n6075), .ZN(n4245) );
  NOR2_X1 U5215 ( .A1(n6058), .A2(n4245), .ZN(n4253) );
  INV_X1 U5216 ( .A(n4253), .ZN(n4248) );
  INV_X1 U5217 ( .A(n5479), .ZN(n4244) );
  NAND2_X1 U5218 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6094) );
  NAND2_X1 U5219 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4768) );
  NOR2_X1 U5220 ( .A1(n6094), .A2(n4768), .ZN(n4771) );
  NAND3_X1 U5221 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n4771), .ZN(n6053) );
  NOR2_X1 U5222 ( .A1(n4245), .A2(n6053), .ZN(n4254) );
  NOR2_X1 U5223 ( .A1(n5479), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4247)
         );
  NOR2_X1 U5224 ( .A1(n4246), .A2(n6112), .ZN(n4318) );
  NOR2_X1 U5225 ( .A1(n4247), .A2(n4318), .ZN(n6054) );
  OAI21_X1 U5226 ( .B1(n6056), .B2(n4254), .A(n6054), .ZN(n5497) );
  AOI21_X1 U5227 ( .B1(n6111), .B2(n4248), .A(n5497), .ZN(n5486) );
  INV_X1 U5228 ( .A(n5486), .ZN(n5728) );
  NAND3_X1 U5229 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A3(INSTADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n5483) );
  NOR2_X1 U5230 ( .A1(n4167), .A2(n5483), .ZN(n4255) );
  INV_X1 U5231 ( .A(n4255), .ZN(n5729) );
  NAND2_X1 U5232 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5731) );
  OAI21_X1 U5233 ( .B1(n5729), .B2(n5731), .A(n5730), .ZN(n4249) );
  INV_X1 U5234 ( .A(n4249), .ZN(n4250) );
  NOR2_X1 U5235 ( .A1(n5728), .A2(n4250), .ZN(n5727) );
  NAND2_X1 U5236 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4251) );
  OAI21_X1 U5237 ( .B1(n4251), .B2(n5700), .A(n5730), .ZN(n4252) );
  NAND2_X1 U5238 ( .A1(n5727), .A2(n4252), .ZN(n5476) );
  NAND2_X1 U5239 ( .A1(n6111), .A2(n4253), .ZN(n5480) );
  NOR2_X1 U5240 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5484), .ZN(n4316)
         );
  NAND2_X1 U5241 ( .A1(n4254), .A2(n6108), .ZN(n5496) );
  NAND3_X1 U5242 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n5722), .ZN(n5711) );
  INV_X1 U5243 ( .A(n4261), .ZN(n5461) );
  NAND2_X1 U5244 ( .A1(n4261), .A2(n5460), .ZN(n5473) );
  OAI21_X1 U5245 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5461), .A(n5473), 
        .ZN(n4256) );
  AOI21_X1 U5247 ( .B1(n4257), .B2(n6088), .A(n4262), .ZN(n4258) );
  AND2_X1 U5248 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5436) );
  INV_X1 U5249 ( .A(n5436), .ZN(n4259) );
  NAND2_X1 U5250 ( .A1(n5730), .A2(n4259), .ZN(n4260) );
  NAND2_X1 U5251 ( .A1(n5695), .A2(n4260), .ZN(n5431) );
  AOI21_X1 U5252 ( .B1(n5417), .B2(n5730), .A(n5431), .ZN(n5407) );
  OAI21_X1 U5253 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n6059), .A(n5407), 
        .ZN(n5404) );
  AOI21_X1 U5254 ( .B1(n5399), .B2(n5730), .A(n5404), .ZN(n4268) );
  INV_X1 U5255 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4267) );
  NAND2_X1 U5256 ( .A1(n4261), .A2(n5297), .ZN(n5455) );
  INV_X1 U5257 ( .A(n4262), .ZN(n4263) );
  NAND2_X1 U5258 ( .A1(n5690), .A2(n5436), .ZN(n5428) );
  INV_X1 U5259 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4264) );
  NOR3_X1 U5260 ( .A1(n5428), .A2(n5417), .A3(n4264), .ZN(n5400) );
  NAND3_X1 U5261 ( .A1(n5400), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n4267), .ZN(n4265) );
  OAI211_X1 U5262 ( .C1(n4268), .C2(n4267), .A(n4266), .B(n4265), .ZN(n4269)
         );
  AOI21_X1 U5263 ( .B1(n4270), .B2(n6100), .A(n4269), .ZN(n4271) );
  OAI21_X1 U5264 ( .B1(n4272), .B2(n5519), .A(n4271), .ZN(U2987) );
  AND2_X1 U5265 ( .A1(n4276), .A2(n4827), .ZN(n4273) );
  NAND2_X1 U5266 ( .A1(n4284), .A2(n4273), .ZN(n4291) );
  NAND2_X1 U5267 ( .A1(n6245), .A2(n6488), .ZN(n4913) );
  INV_X1 U5268 ( .A(n4913), .ZN(n4294) );
  INV_X1 U5269 ( .A(n4275), .ZN(n4280) );
  INV_X1 U5270 ( .A(n4292), .ZN(n5947) );
  AOI211_X1 U5271 ( .C1(MEMORYFETCH_REG_SCAN_IN), .C2(n4291), .A(n4294), .B(
        n5947), .ZN(n4274) );
  INV_X1 U5272 ( .A(n4274), .ZN(U2788) );
  INV_X1 U5273 ( .A(n4379), .ZN(n4278) );
  INV_X1 U5274 ( .A(n4831), .ZN(n4841) );
  AOI21_X1 U5275 ( .B1(n4284), .B2(n4276), .A(n4275), .ZN(n4277) );
  AOI21_X1 U5276 ( .B1(n4278), .B2(n4841), .A(n4277), .ZN(n5760) );
  NOR2_X1 U5277 ( .A1(n4279), .A2(n6507), .ZN(n4293) );
  INV_X1 U5278 ( .A(n6413), .ZN(n4324) );
  OAI21_X1 U5279 ( .B1(n4293), .B2(n4324), .A(n6599), .ZN(n6506) );
  NAND2_X1 U5280 ( .A1(n5760), .A2(n6506), .ZN(n6384) );
  AND2_X1 U5281 ( .A1(n6384), .A2(n4827), .ZN(n5767) );
  INV_X1 U5282 ( .A(MORE_REG_SCAN_IN), .ZN(n4290) );
  AND2_X1 U5283 ( .A1(n4281), .A2(n4280), .ZN(n4282) );
  OR2_X1 U5284 ( .A1(n4379), .A2(n4282), .ZN(n4287) );
  NAND2_X1 U5285 ( .A1(n4379), .A2(n4658), .ZN(n4286) );
  OR2_X1 U5286 ( .A1(n4284), .A2(n4283), .ZN(n4285) );
  AND3_X1 U5287 ( .A1(n4287), .A2(n4286), .A3(n4285), .ZN(n6382) );
  INV_X1 U5288 ( .A(n6382), .ZN(n4288) );
  NAND2_X1 U5289 ( .A1(n5767), .A2(n4288), .ZN(n4289) );
  OAI21_X1 U5290 ( .B1(n5767), .B2(n4290), .A(n4289), .ZN(U3471) );
  INV_X1 U5291 ( .A(n4293), .ZN(n4296) );
  OAI21_X1 U5292 ( .B1(n4294), .B2(READREQUEST_REG_SCAN_IN), .A(n6511), .ZN(
        n4295) );
  OAI21_X1 U5293 ( .B1(n6511), .B2(n4296), .A(n4295), .ZN(U3474) );
  XNOR2_X1 U5294 ( .A(n4297), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6042)
         );
  OAI21_X1 U5295 ( .B1(n4299), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4298), 
        .ZN(n5884) );
  OAI21_X1 U5296 ( .B1(n4318), .B2(n5484), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4300) );
  NAND2_X1 U5297 ( .A1(n6112), .A2(REIP_REG_0__SCAN_IN), .ZN(n6048) );
  OAI211_X1 U5298 ( .C1(n5884), .C2(n6116), .A(n4300), .B(n6048), .ZN(n4301)
         );
  AND2_X1 U5299 ( .A1(n5482), .A2(n6667), .ZN(n4317) );
  NOR2_X1 U5300 ( .A1(n4301), .A2(n4317), .ZN(n4302) );
  OAI21_X1 U5301 ( .B1(n6042), .B2(n5519), .A(n4302), .ZN(U3018) );
  NAND2_X1 U5302 ( .A1(n5920), .A2(n4852), .ZN(n4758) );
  NOR2_X1 U5303 ( .A1(n6488), .A2(n6210), .ZN(n4693) );
  NAND2_X1 U5304 ( .A1(n4693), .A2(n6509), .ZN(n6513) );
  INV_X2 U5305 ( .A(n6513), .ZN(n5943) );
  NOR2_X4 U5306 ( .A1(n5943), .A2(n5920), .ZN(n5934) );
  AOI22_X1 U5307 ( .A1(DATAO_REG_16__SCAN_IN), .A2(n5934), .B1(n5943), .B2(
        UWORD_REG_0__SCAN_IN), .ZN(n4305) );
  OAI21_X1 U5308 ( .B1(n3761), .B2(n4758), .A(n4305), .ZN(U2907) );
  INV_X1 U5309 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4307) );
  AOI22_X1 U5310 ( .A1(DATAO_REG_18__SCAN_IN), .A2(n5934), .B1(n5943), .B2(
        UWORD_REG_2__SCAN_IN), .ZN(n4306) );
  OAI21_X1 U5311 ( .B1(n4307), .B2(n4758), .A(n4306), .ZN(U2905) );
  INV_X1 U5312 ( .A(EAX_REG_28__SCAN_IN), .ZN(n5966) );
  AOI22_X1 U5313 ( .A1(UWORD_REG_12__SCAN_IN), .A2(n5943), .B1(n5934), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4308) );
  OAI21_X1 U5314 ( .B1(n5966), .B2(n4758), .A(n4308), .ZN(U2895) );
  INV_X1 U5315 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4310) );
  AOI22_X1 U5316 ( .A1(UWORD_REG_10__SCAN_IN), .A2(n5943), .B1(n5934), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4309) );
  OAI21_X1 U5317 ( .B1(n4310), .B2(n4758), .A(n4309), .ZN(U2897) );
  INV_X1 U5318 ( .A(EAX_REG_27__SCAN_IN), .ZN(n5963) );
  AOI22_X1 U5319 ( .A1(n5943), .A2(UWORD_REG_11__SCAN_IN), .B1(n5934), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4311) );
  OAI21_X1 U5320 ( .B1(n5963), .B2(n4758), .A(n4311), .ZN(U2896) );
  AOI22_X1 U5321 ( .A1(n5943), .A2(UWORD_REG_8__SCAN_IN), .B1(n5934), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4312) );
  OAI21_X1 U5322 ( .B1(n3925), .B2(n4758), .A(n4312), .ZN(U2899) );
  INV_X1 U5323 ( .A(EAX_REG_29__SCAN_IN), .ZN(n5969) );
  AOI22_X1 U5324 ( .A1(n5943), .A2(UWORD_REG_13__SCAN_IN), .B1(n5934), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4313) );
  OAI21_X1 U5325 ( .B1(n5969), .B2(n4758), .A(n4313), .ZN(U2894) );
  XNOR2_X1 U5326 ( .A(n4315), .B(n4314), .ZN(n4971) );
  NOR3_X1 U5327 ( .A1(n6059), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n4316), 
        .ZN(n4322) );
  XNOR2_X1 U5328 ( .A(n4847), .B(n4325), .ZN(n4406) );
  OAI21_X1 U5329 ( .B1(n4318), .B2(n4317), .A(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .ZN(n4320) );
  AND2_X1 U5330 ( .A1(n6112), .A2(REIP_REG_1__SCAN_IN), .ZN(n4966) );
  INV_X1 U5331 ( .A(n4966), .ZN(n4319) );
  OAI211_X1 U5332 ( .C1(n6116), .C2(n4406), .A(n4320), .B(n4319), .ZN(n4321)
         );
  NOR2_X1 U5333 ( .A1(n4322), .A2(n4321), .ZN(n4323) );
  OAI21_X1 U5334 ( .B1(n4971), .B2(n5519), .A(n4323), .ZN(U3017) );
  NAND2_X1 U5335 ( .A1(n6370), .A2(n4324), .ZN(n4328) );
  NAND2_X1 U5336 ( .A1(n4325), .A2(n6413), .ZN(n4326) );
  NAND2_X1 U5337 ( .A1(n4346), .A2(n4326), .ZN(n4327) );
  AOI21_X1 U5338 ( .B1(n4328), .B2(n4327), .A(READY_N), .ZN(n4329) );
  NAND2_X1 U5339 ( .A1(n4379), .A2(n4329), .ZN(n4333) );
  INV_X1 U5340 ( .A(n4330), .ZN(n4331) );
  NAND3_X1 U5341 ( .A1(n4333), .A2(n4332), .A3(n4331), .ZN(n4339) );
  NOR2_X1 U5342 ( .A1(n4334), .A2(n4841), .ZN(n4659) );
  NAND2_X1 U5343 ( .A1(n4379), .A2(n4659), .ZN(n4337) );
  INV_X1 U5344 ( .A(n4653), .ZN(n5755) );
  NAND2_X1 U5345 ( .A1(n5755), .A2(n4335), .ZN(n4336) );
  NAND2_X1 U5346 ( .A1(n4337), .A2(n4336), .ZN(n4828) );
  NOR2_X1 U5347 ( .A1(n4379), .A2(n4378), .ZN(n4338) );
  INV_X1 U5348 ( .A(n6371), .ZN(n4340) );
  NAND2_X1 U5349 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4693), .ZN(n6485) );
  INV_X1 U5350 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5766) );
  OAI22_X1 U5351 ( .A1(n4340), .A2(n6400), .B1(n6485), .B2(n5766), .ZN(n5753)
         );
  NOR2_X1 U5352 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6487), .ZN(n4369) );
  INV_X1 U5353 ( .A(n5531), .ZN(n6490) );
  OAI21_X1 U5354 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6395), .A(n6490), 
        .ZN(n6491) );
  INV_X1 U5355 ( .A(n6491), .ZN(n4356) );
  INV_X1 U5356 ( .A(n6395), .ZN(n5020) );
  NAND2_X1 U5357 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5022) );
  INV_X1 U5358 ( .A(n5022), .ZN(n4354) );
  AOI22_X1 U5359 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4267), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4342), .ZN(n5023) );
  NAND2_X1 U5360 ( .A1(n4344), .A2(n4343), .ZN(n4345) );
  NOR2_X1 U5361 ( .A1(n4346), .A2(n4345), .ZN(n4347) );
  NAND2_X1 U5362 ( .A1(n4653), .A2(n4347), .ZN(n4349) );
  NOR2_X1 U5363 ( .A1(n4349), .A2(n4348), .ZN(n4663) );
  INV_X1 U5364 ( .A(n4663), .ZN(n6368) );
  NAND2_X1 U5365 ( .A1(n4518), .A2(n6368), .ZN(n4352) );
  OAI21_X1 U5366 ( .B1(n4341), .B2(n4350), .A(n6367), .ZN(n4351) );
  OAI211_X1 U5367 ( .C1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n4353), .A(n4352), .B(n4351), .ZN(n6372) );
  INV_X1 U5368 ( .A(n6494), .ZN(n5754) );
  AOI222_X1 U5369 ( .A1(n5020), .A2(n4341), .B1(n4354), .B2(n5023), .C1(n6372), 
        .C2(n5754), .ZN(n4355) );
  OAI22_X1 U5370 ( .A1(n4356), .A2(n3041), .B1(n5531), .B2(n4355), .ZN(U3460)
         );
  INV_X1 U5371 ( .A(DATAI_6_), .ZN(n5984) );
  NAND2_X1 U5372 ( .A1(n6488), .A2(n6210), .ZN(n6508) );
  INV_X1 U5373 ( .A(n6508), .ZN(n6408) );
  INV_X1 U5374 ( .A(n6350), .ZN(n5585) );
  INV_X1 U5375 ( .A(n3576), .ZN(n6369) );
  AND2_X1 U5376 ( .A1(n6143), .A2(n6369), .ZN(n6286) );
  INV_X1 U5377 ( .A(n4518), .ZN(n5523) );
  OR2_X1 U5378 ( .A1(n5526), .A2(n5523), .ZN(n6145) );
  INV_X1 U5379 ( .A(n6145), .ZN(n4736) );
  INV_X1 U5380 ( .A(n4509), .ZN(n4359) );
  AOI21_X1 U5381 ( .B1(n6286), .B2(n4736), .A(n4359), .ZN(n4364) );
  INV_X1 U5382 ( .A(n4364), .ZN(n4360) );
  NAND2_X1 U5383 ( .A1(n4360), .A2(n6245), .ZN(n4362) );
  NAND2_X1 U5384 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n4367), .ZN(n4361) );
  NAND2_X1 U5385 ( .A1(n3566), .A2(n4363), .ZN(n4602) );
  INV_X1 U5386 ( .A(n4602), .ZN(n4370) );
  AOI21_X1 U5387 ( .B1(n4370), .B2(n5521), .A(n6043), .ZN(n4365) );
  AND2_X1 U5388 ( .A1(n6245), .A2(n6638), .ZN(n4782) );
  OAI21_X1 U5389 ( .B1(n4365), .B2(n4782), .A(n4364), .ZN(n4366) );
  OAI211_X1 U5390 ( .C1(n6245), .C2(n4367), .A(n4366), .B(n6208), .ZN(n4504)
         );
  NAND2_X1 U5391 ( .A1(n4491), .A2(n3261), .ZN(n4887) );
  NAND2_X1 U5392 ( .A1(n6035), .A2(DATAI_22_), .ZN(n6173) );
  INV_X1 U5393 ( .A(n6173), .ZN(n6348) );
  NAND2_X1 U5394 ( .A1(n5521), .A2(n3574), .ZN(n4529) );
  INV_X1 U5395 ( .A(n4645), .ZN(n4418) );
  NAND2_X1 U5396 ( .A1(n6035), .A2(DATAI_30_), .ZN(n6277) );
  INV_X1 U5397 ( .A(n6277), .ZN(n6346) );
  AOI22_X1 U5398 ( .A1(n6348), .A2(n4418), .B1(n4606), .B2(n6346), .ZN(n4371)
         );
  OAI21_X1 U5399 ( .B1(n4887), .B2(n4509), .A(n4371), .ZN(n4372) );
  AOI21_X1 U5400 ( .B1(INSTQUEUE_REG_15__6__SCAN_IN), .B2(n4504), .A(n4372), 
        .ZN(n4373) );
  OAI21_X1 U5401 ( .B1(n5585), .B2(n4505), .A(n4373), .ZN(U3146) );
  NAND3_X1 U5402 ( .A1(n4403), .A2(n4376), .A3(n4375), .ZN(n4377) );
  AND2_X1 U5403 ( .A1(n4374), .A2(n4377), .ZN(n6034) );
  INV_X1 U5404 ( .A(n6034), .ZN(n4997) );
  NAND4_X1 U5405 ( .A1(n4067), .A2(n4381), .A3(n4380), .A4(n6488), .ZN(n4385)
         );
  OR2_X1 U5406 ( .A1(n4383), .A2(n4382), .ZN(n4384) );
  NOR2_X1 U5407 ( .A1(n4385), .A2(n4384), .ZN(n4832) );
  NAND2_X1 U5408 ( .A1(n4832), .A2(n4849), .ZN(n4386) );
  OR2_X1 U5409 ( .A1(n4390), .A2(n4389), .ZN(n4391) );
  NAND2_X1 U5410 ( .A1(n4512), .A2(n4391), .ZN(n6115) );
  INV_X1 U5411 ( .A(n6115), .ZN(n4392) );
  AOI22_X1 U5412 ( .A1(n6518), .A2(n4392), .B1(n6517), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n4393) );
  OAI21_X1 U5413 ( .B1(n4997), .B2(n5902), .A(n4393), .ZN(U2857) );
  NAND2_X1 U5414 ( .A1(n4491), .A2(n4852), .ZN(n5544) );
  NAND2_X1 U5415 ( .A1(n4504), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4396)
         );
  NAND2_X1 U5416 ( .A1(n6035), .A2(DATAI_24_), .ZN(n6302) );
  INV_X1 U5417 ( .A(n6302), .ZN(n6153) );
  NAND2_X1 U5418 ( .A1(n6035), .A2(DATAI_16_), .ZN(n6156) );
  INV_X1 U5419 ( .A(DATAI_0_), .ZN(n5972) );
  NOR2_X1 U5420 ( .A1(n5972), .A2(n4779), .ZN(n6243) );
  OAI22_X1 U5421 ( .A1(n4645), .A2(n6156), .B1(n4505), .B2(n6301), .ZN(n4394)
         );
  AOI21_X1 U5422 ( .B1(n6153), .B2(n4606), .A(n4394), .ZN(n4395) );
  OAI211_X1 U5423 ( .C1(n5544), .C2(n4509), .A(n4396), .B(n4395), .ZN(U3140)
         );
  XNOR2_X1 U5424 ( .A(n2988), .B(n4397), .ZN(n6027) );
  INV_X1 U5425 ( .A(n6027), .ZN(n4837) );
  AND2_X1 U5426 ( .A1(n4514), .A2(n4398), .ZN(n4399) );
  NOR2_X1 U5427 ( .A1(n4486), .A2(n4399), .ZN(n6090) );
  AOI22_X1 U5428 ( .A1(n6518), .A2(n6090), .B1(n6517), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4400) );
  OAI21_X1 U5429 ( .B1(n4837), .B2(n5902), .A(n4400), .ZN(U2855) );
  XNOR2_X1 U5430 ( .A(n4402), .B(n4401), .ZN(n6044) );
  OAI222_X1 U5431 ( .A1(n5884), .A2(n5901), .B1(n5905), .B2(n5895), .C1(n5902), 
        .C2(n6044), .ZN(U2859) );
  INV_X1 U5432 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4846) );
  OAI21_X1 U5433 ( .B1(n4405), .B2(n4404), .A(n4403), .ZN(n4998) );
  OAI222_X1 U5434 ( .A1(n4406), .A2(n5901), .B1(n4846), .B2(n5905), .C1(n4998), 
        .C2(n5902), .ZN(U2858) );
  NAND2_X1 U5435 ( .A1(n4491), .A2(n4407), .ZN(n5548) );
  NAND2_X1 U5436 ( .A1(n4504), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4410)
         );
  NAND2_X1 U5437 ( .A1(n6035), .A2(DATAI_25_), .ZN(n6309) );
  INV_X1 U5438 ( .A(n6309), .ZN(n6157) );
  NAND2_X1 U5439 ( .A1(n6035), .A2(DATAI_17_), .ZN(n6160) );
  INV_X1 U5440 ( .A(DATAI_1_), .ZN(n5974) );
  OAI22_X1 U5441 ( .A1(n4645), .A2(n6160), .B1(n4505), .B2(n6308), .ZN(n4408)
         );
  AOI21_X1 U5442 ( .B1(n6157), .B2(n4606), .A(n4408), .ZN(n4409) );
  OAI211_X1 U5443 ( .C1(n5548), .C2(n4509), .A(n4410), .B(n4409), .ZN(U3141)
         );
  NAND2_X1 U5444 ( .A1(n4491), .A2(n4411), .ZN(n5556) );
  NAND2_X1 U5445 ( .A1(n4504), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4414)
         );
  NAND2_X1 U5446 ( .A1(n6035), .A2(DATAI_27_), .ZN(n6324) );
  INV_X1 U5447 ( .A(n6324), .ZN(n6220) );
  NAND2_X1 U5448 ( .A1(n6035), .A2(DATAI_19_), .ZN(n6223) );
  INV_X1 U5449 ( .A(DATAI_3_), .ZN(n5978) );
  OAI22_X1 U5450 ( .A1(n4645), .A2(n6223), .B1(n4505), .B2(n6323), .ZN(n4412)
         );
  AOI21_X1 U5451 ( .B1(n6220), .B2(n4606), .A(n4412), .ZN(n4413) );
  OAI211_X1 U5452 ( .C1(n5556), .C2(n4509), .A(n4414), .B(n4413), .ZN(U3143)
         );
  NAND3_X1 U5453 ( .A1(n6201), .A2(n6589), .A3(n6373), .ZN(n4551) );
  NOR2_X1 U5454 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4551), .ZN(n4640)
         );
  INV_X1 U5455 ( .A(n4640), .ZN(n4650) );
  INV_X1 U5456 ( .A(n4423), .ZN(n4415) );
  NOR2_X1 U5457 ( .A1(n4415), .A2(n6210), .ZN(n6141) );
  INV_X1 U5458 ( .A(n4778), .ZN(n4416) );
  OAI21_X1 U5459 ( .B1(n3109), .B2(n6210), .A(n4601), .ZN(n4704) );
  AOI211_X1 U5460 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4650), .A(n6141), .B(
        n4704), .ZN(n4421) );
  NOR2_X1 U5461 ( .A1(n3566), .A2(n5521), .ZN(n4417) );
  NOR3_X1 U5462 ( .A1(n4647), .A2(n4418), .A3(n6295), .ZN(n4419) );
  NAND2_X1 U5463 ( .A1(n5523), .A2(n5526), .ZN(n4575) );
  OR2_X1 U5464 ( .A1(n4575), .A2(n6143), .ZN(n4422) );
  OAI21_X1 U5465 ( .B1(n4419), .B2(n4782), .A(n4422), .ZN(n4420) );
  INV_X1 U5466 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4428) );
  INV_X1 U5467 ( .A(n6160), .ZN(n6306) );
  INV_X1 U5468 ( .A(n4422), .ZN(n4548) );
  NOR2_X1 U5469 ( .A1(n4423), .A2(n6210), .ZN(n6147) );
  AND2_X1 U5470 ( .A1(n3109), .A2(n6147), .ZN(n4424) );
  AOI21_X1 U5471 ( .B1(n4548), .B2(n6245), .A(n4424), .ZN(n4644) );
  OAI22_X1 U5472 ( .A1(n4645), .A2(n6309), .B1(n4644), .B2(n6308), .ZN(n4425)
         );
  AOI21_X1 U5473 ( .B1(n4647), .B2(n6306), .A(n4425), .ZN(n4427) );
  NAND2_X1 U5474 ( .A1(n6307), .A2(n4640), .ZN(n4426) );
  OAI211_X1 U5475 ( .C1(n4637), .C2(n4428), .A(n4427), .B(n4426), .ZN(U3021)
         );
  INV_X1 U5476 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4432) );
  NAND2_X1 U5477 ( .A1(n6035), .A2(DATAI_20_), .ZN(n6332) );
  INV_X1 U5478 ( .A(n6332), .ZN(n6266) );
  NAND2_X1 U5479 ( .A1(n6035), .A2(DATAI_28_), .ZN(n6269) );
  INV_X1 U5480 ( .A(DATAI_4_), .ZN(n5980) );
  OAI22_X1 U5481 ( .A1(n4645), .A2(n6269), .B1(n4644), .B2(n6331), .ZN(n4429)
         );
  AOI21_X1 U5482 ( .B1(n4647), .B2(n6266), .A(n4429), .ZN(n4431) );
  NAND2_X1 U5483 ( .A1(n4491), .A2(n3239), .ZN(n5560) );
  NAND2_X1 U5484 ( .A1(n6330), .A2(n4640), .ZN(n4430) );
  OAI211_X1 U5485 ( .C1(n4637), .C2(n4432), .A(n4431), .B(n4430), .ZN(U3024)
         );
  INV_X1 U5486 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4437) );
  NAND2_X1 U5487 ( .A1(n6035), .A2(DATAI_21_), .ZN(n6340) );
  INV_X1 U5488 ( .A(n6340), .ZN(n6271) );
  NAND2_X1 U5489 ( .A1(n6035), .A2(DATAI_29_), .ZN(n6274) );
  INV_X1 U5490 ( .A(DATAI_5_), .ZN(n5982) );
  OAI22_X1 U5491 ( .A1(n4645), .A2(n6274), .B1(n4644), .B2(n6339), .ZN(n4433)
         );
  AOI21_X1 U5492 ( .B1(n4647), .B2(n6271), .A(n4433), .ZN(n4436) );
  NAND2_X1 U5493 ( .A1(n4491), .A2(n4434), .ZN(n5564) );
  NAND2_X1 U5494 ( .A1(n6338), .A2(n4640), .ZN(n4435) );
  OAI211_X1 U5495 ( .C1(n4637), .C2(n4437), .A(n4436), .B(n4435), .ZN(U3025)
         );
  INV_X1 U5496 ( .A(n6156), .ZN(n6293) );
  OAI22_X1 U5497 ( .A1(n4645), .A2(n6302), .B1(n4644), .B2(n6301), .ZN(n4438)
         );
  AOI21_X1 U5498 ( .B1(n4647), .B2(n6293), .A(n4438), .ZN(n4440) );
  NAND2_X1 U5499 ( .A1(n6294), .A2(n4640), .ZN(n4439) );
  OAI211_X1 U5500 ( .C1(n4637), .C2(n4441), .A(n4440), .B(n4439), .ZN(U3020)
         );
  INV_X1 U5501 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n6655) );
  INV_X1 U5502 ( .A(n6223), .ZN(n6321) );
  OAI22_X1 U5503 ( .A1(n4645), .A2(n6324), .B1(n4644), .B2(n6323), .ZN(n4442)
         );
  AOI21_X1 U5504 ( .B1(n4647), .B2(n6321), .A(n4442), .ZN(n4444) );
  NAND2_X1 U5505 ( .A1(n6322), .A2(n4640), .ZN(n4443) );
  OAI211_X1 U5506 ( .C1(n4637), .C2(n6655), .A(n4444), .B(n4443), .ZN(U3023)
         );
  OR2_X1 U5507 ( .A1(n5521), .A2(n6638), .ZN(n4574) );
  INV_X1 U5508 ( .A(n4574), .ZN(n4446) );
  AOI21_X1 U5509 ( .B1(n4737), .B2(n4446), .A(n6295), .ZN(n4450) );
  OR2_X1 U5510 ( .A1(n5526), .A2(n4518), .ZN(n6246) );
  NOR2_X1 U5511 ( .A1(n6246), .A2(n6247), .ZN(n4699) );
  NAND3_X1 U5512 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6201), .A3(n6373), .ZN(n4701) );
  NOR2_X1 U5513 ( .A1(n6287), .A2(n4701), .ZN(n4493) );
  AOI21_X1 U5514 ( .B1(n4699), .B2(n6369), .A(n4493), .ZN(n4449) );
  INV_X1 U5515 ( .A(n4449), .ZN(n4448) );
  INV_X1 U5516 ( .A(n4701), .ZN(n4447) );
  AOI22_X1 U5517 ( .A1(n4450), .A2(n4448), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4447), .ZN(n4496) );
  AOI22_X1 U5518 ( .A1(n4450), .A2(n4449), .B1(n4701), .B2(n6295), .ZN(n4451)
         );
  NAND2_X1 U5519 ( .A1(n6208), .A2(n4451), .ZN(n4490) );
  NAND2_X1 U5520 ( .A1(n4490), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4456) );
  INV_X1 U5521 ( .A(n4737), .ZN(n4452) );
  NOR2_X1 U5522 ( .A1(n4452), .A2(n5521), .ZN(n4453) );
  NAND2_X1 U5523 ( .A1(n4453), .A2(n3574), .ZN(n6152) );
  OAI22_X1 U5524 ( .A1(n6274), .A2(n5580), .B1(n6152), .B2(n6340), .ZN(n4454)
         );
  AOI21_X1 U5525 ( .B1(n6338), .B2(n4493), .A(n4454), .ZN(n4455) );
  OAI211_X1 U5526 ( .C1(n4496), .C2(n6339), .A(n4456), .B(n4455), .ZN(U3065)
         );
  NAND2_X1 U5527 ( .A1(n4490), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4459) );
  OAI22_X1 U5528 ( .A1(n6324), .A2(n5580), .B1(n6152), .B2(n6223), .ZN(n4457)
         );
  AOI21_X1 U5529 ( .B1(n6322), .B2(n4493), .A(n4457), .ZN(n4458) );
  OAI211_X1 U5530 ( .C1(n4496), .C2(n6323), .A(n4459), .B(n4458), .ZN(U3063)
         );
  NAND2_X1 U5531 ( .A1(n4490), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4462) );
  OAI22_X1 U5532 ( .A1(n6269), .A2(n5580), .B1(n6152), .B2(n6332), .ZN(n4460)
         );
  AOI21_X1 U5533 ( .B1(n6330), .B2(n4493), .A(n4460), .ZN(n4461) );
  OAI211_X1 U5534 ( .C1(n4496), .C2(n6331), .A(n4462), .B(n4461), .ZN(U3064)
         );
  NAND2_X1 U5535 ( .A1(n4490), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4465) );
  OAI22_X1 U5536 ( .A1(n6309), .A2(n5580), .B1(n6152), .B2(n6160), .ZN(n4463)
         );
  AOI21_X1 U5537 ( .B1(n6307), .B2(n4493), .A(n4463), .ZN(n4464) );
  OAI211_X1 U5538 ( .C1(n4496), .C2(n6308), .A(n4465), .B(n4464), .ZN(U3061)
         );
  INV_X1 U5539 ( .A(DATAI_2_), .ZN(n5976) );
  NAND2_X1 U5540 ( .A1(n4490), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4468) );
  NAND2_X1 U5541 ( .A1(n4491), .A2(n3165), .ZN(n5552) );
  NAND2_X1 U5542 ( .A1(n6035), .A2(DATAI_26_), .ZN(n6316) );
  NAND2_X1 U5543 ( .A1(n6035), .A2(DATAI_18_), .ZN(n6164) );
  OAI22_X1 U5544 ( .A1(n6316), .A2(n5580), .B1(n6152), .B2(n6164), .ZN(n4466)
         );
  AOI21_X1 U5545 ( .B1(n6314), .B2(n4493), .A(n4466), .ZN(n4467) );
  OAI211_X1 U5546 ( .C1(n4496), .C2(n6315), .A(n4468), .B(n4467), .ZN(U3062)
         );
  NAND2_X1 U5547 ( .A1(n4490), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4471) );
  OAI22_X1 U5548 ( .A1(n6302), .A2(n5580), .B1(n6152), .B2(n6156), .ZN(n4469)
         );
  AOI21_X1 U5549 ( .B1(n6294), .B2(n4493), .A(n4469), .ZN(n4470) );
  OAI211_X1 U5550 ( .C1(n4496), .C2(n6301), .A(n4471), .B(n4470), .ZN(U3060)
         );
  NAND2_X1 U5551 ( .A1(n4504), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4474)
         );
  INV_X1 U5552 ( .A(n6269), .ZN(n6329) );
  OAI22_X1 U5553 ( .A1(n4645), .A2(n6332), .B1(n4505), .B2(n6331), .ZN(n4472)
         );
  AOI21_X1 U5554 ( .B1(n6329), .B2(n4606), .A(n4472), .ZN(n4473) );
  OAI211_X1 U5555 ( .C1(n5560), .C2(n4509), .A(n4474), .B(n4473), .ZN(U3144)
         );
  NAND2_X1 U5556 ( .A1(n4504), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4477)
         );
  INV_X1 U5557 ( .A(n6274), .ZN(n6337) );
  OAI22_X1 U5558 ( .A1(n4645), .A2(n6340), .B1(n4505), .B2(n6339), .ZN(n4475)
         );
  AOI21_X1 U5559 ( .B1(n6337), .B2(n4606), .A(n4475), .ZN(n4476) );
  OAI211_X1 U5560 ( .C1(n5564), .C2(n4509), .A(n4477), .B(n4476), .ZN(U3145)
         );
  NAND2_X1 U5561 ( .A1(n4490), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4480) );
  OAI22_X1 U5562 ( .A1(n6277), .A2(n5580), .B1(n6152), .B2(n6173), .ZN(n4478)
         );
  AOI21_X1 U5563 ( .B1(n6347), .B2(n4493), .A(n4478), .ZN(n4479) );
  OAI211_X1 U5564 ( .C1(n4496), .C2(n5585), .A(n4480), .B(n4479), .ZN(U3066)
         );
  OR2_X1 U5565 ( .A1(n4483), .A2(n4482), .ZN(n4484) );
  NAND2_X1 U5566 ( .A1(n4481), .A2(n4484), .ZN(n5015) );
  NOR2_X1 U5567 ( .A1(n4486), .A2(n4485), .ZN(n4487) );
  OR2_X1 U5568 ( .A1(n4761), .A2(n4487), .ZN(n4923) );
  INV_X1 U5569 ( .A(n4923), .ZN(n4488) );
  AOI22_X1 U5570 ( .A1(n4488), .A2(n6518), .B1(n6517), .B2(EBX_REG_5__SCAN_IN), 
        .ZN(n4489) );
  OAI21_X1 U5571 ( .B1(n5015), .B2(n5212), .A(n4489), .ZN(U2854) );
  INV_X1 U5572 ( .A(DATAI_7_), .ZN(n5986) );
  NAND2_X1 U5573 ( .A1(n4490), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4495) );
  NAND2_X1 U5574 ( .A1(n4491), .A2(n3320), .ZN(n5576) );
  NAND2_X1 U5575 ( .A1(n6035), .A2(DATAI_31_), .ZN(n6360) );
  NAND2_X1 U5576 ( .A1(n6035), .A2(DATAI_23_), .ZN(n6181) );
  OAI22_X1 U5577 ( .A1(n6360), .A2(n5580), .B1(n6152), .B2(n6181), .ZN(n4492)
         );
  AOI21_X1 U5578 ( .B1(n6357), .B2(n4493), .A(n4492), .ZN(n4494) );
  OAI211_X1 U5579 ( .C1(n4496), .C2(n6358), .A(n4495), .B(n4494), .ZN(U3067)
         );
  INV_X1 U5580 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4500) );
  INV_X1 U5581 ( .A(n6164), .ZN(n6313) );
  OAI22_X1 U5582 ( .A1(n4645), .A2(n6316), .B1(n4644), .B2(n6315), .ZN(n4497)
         );
  AOI21_X1 U5583 ( .B1(n4647), .B2(n6313), .A(n4497), .ZN(n4499) );
  NAND2_X1 U5584 ( .A1(n6314), .A2(n4640), .ZN(n4498) );
  OAI211_X1 U5585 ( .C1(n4637), .C2(n4500), .A(n4499), .B(n4498), .ZN(U3022)
         );
  NAND2_X1 U5586 ( .A1(n4504), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4503)
         );
  INV_X1 U5587 ( .A(n6360), .ZN(n6177) );
  OAI22_X1 U5588 ( .A1(n4645), .A2(n6181), .B1(n4505), .B2(n6358), .ZN(n4501)
         );
  AOI21_X1 U5589 ( .B1(n6177), .B2(n4606), .A(n4501), .ZN(n4502) );
  OAI211_X1 U5590 ( .C1(n5576), .C2(n4509), .A(n4503), .B(n4502), .ZN(U3147)
         );
  NAND2_X1 U5591 ( .A1(n4504), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4508)
         );
  INV_X1 U5592 ( .A(n6316), .ZN(n6161) );
  OAI22_X1 U5593 ( .A1(n4645), .A2(n6164), .B1(n4505), .B2(n6315), .ZN(n4506)
         );
  AOI21_X1 U5594 ( .B1(n6161), .B2(n4606), .A(n4506), .ZN(n4507) );
  OAI211_X1 U5595 ( .C1(n5552), .C2(n4509), .A(n4508), .B(n4507), .ZN(U3142)
         );
  AOI21_X1 U5596 ( .B1(n4510), .B2(n4374), .A(n2988), .ZN(n4994) );
  INV_X1 U5597 ( .A(n4994), .ZN(n4999) );
  NAND2_X1 U5598 ( .A1(n4512), .A2(n4511), .ZN(n4513) );
  NAND2_X1 U5599 ( .A1(n4514), .A2(n4513), .ZN(n4986) );
  INV_X1 U5600 ( .A(n4986), .ZN(n6099) );
  AOI22_X1 U5601 ( .A1(n6518), .A2(n6099), .B1(n6517), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4515) );
  OAI21_X1 U5602 ( .B1(n4999), .B2(n5902), .A(n4515), .ZN(U2856) );
  NOR2_X1 U5603 ( .A1(n4602), .A2(n4574), .ZN(n6290) );
  NAND2_X1 U5604 ( .A1(n4737), .A2(n6204), .ZN(n4733) );
  NAND2_X1 U5605 ( .A1(n4733), .A2(n4869), .ZN(n4516) );
  OAI21_X1 U5606 ( .B1(n6290), .B2(n4516), .A(n6245), .ZN(n4688) );
  INV_X1 U5607 ( .A(n6204), .ZN(n5520) );
  OAI21_X1 U5608 ( .B1(n3566), .B2(n5520), .A(n6245), .ZN(n4517) );
  NAND2_X1 U5609 ( .A1(n4688), .A2(n4517), .ZN(n4526) );
  INV_X1 U5610 ( .A(n6143), .ZN(n6241) );
  AND2_X1 U5611 ( .A1(n4518), .A2(n5526), .ZN(n4873) );
  NAND2_X1 U5612 ( .A1(n6241), .A2(n4873), .ZN(n5538) );
  OR2_X1 U5613 ( .A1(n5538), .A2(n3576), .ZN(n4520) );
  INV_X1 U5614 ( .A(n6202), .ZN(n4519) );
  NAND2_X1 U5615 ( .A1(n4519), .A2(n6201), .ZN(n4528) );
  INV_X1 U5616 ( .A(n4525), .ZN(n4521) );
  NAND2_X1 U5617 ( .A1(n4526), .A2(n4521), .ZN(n4524) );
  NAND3_X1 U5618 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6201), .A3(n6589), .ZN(n5533) );
  INV_X1 U5619 ( .A(n5533), .ZN(n4522) );
  NAND2_X1 U5620 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n4522), .ZN(n4523) );
  NAND2_X1 U5621 ( .A1(n4524), .A2(n4523), .ZN(n6133) );
  AOI22_X1 U5622 ( .A1(n4526), .A2(n4525), .B1(n5533), .B2(n6295), .ZN(n4527)
         );
  NAND2_X1 U5623 ( .A1(n6208), .A2(n4527), .ZN(n6134) );
  NAND2_X1 U5624 ( .A1(n6134), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4533) );
  INV_X1 U5625 ( .A(n4528), .ZN(n6132) );
  INV_X1 U5626 ( .A(n3566), .ZN(n4530) );
  NAND3_X1 U5627 ( .A1(n4530), .A2(n4870), .A3(n4689), .ZN(n6137) );
  NAND3_X1 U5628 ( .A1(n4530), .A2(n6203), .A3(n4689), .ZN(n6126) );
  OAI22_X1 U5629 ( .A1(n6309), .A2(n6137), .B1(n6126), .B2(n6160), .ZN(n4531)
         );
  AOI21_X1 U5630 ( .B1(n6307), .B2(n6132), .A(n4531), .ZN(n4532) );
  OAI211_X1 U5631 ( .C1(n4546), .C2(n6308), .A(n4533), .B(n4532), .ZN(U3045)
         );
  NAND2_X1 U5632 ( .A1(n6134), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4536) );
  OAI22_X1 U5633 ( .A1(n6324), .A2(n6137), .B1(n6126), .B2(n6223), .ZN(n4534)
         );
  AOI21_X1 U5634 ( .B1(n6322), .B2(n6132), .A(n4534), .ZN(n4535) );
  OAI211_X1 U5635 ( .C1(n4546), .C2(n6323), .A(n4536), .B(n4535), .ZN(U3047)
         );
  NAND2_X1 U5636 ( .A1(n6134), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4539) );
  OAI22_X1 U5637 ( .A1(n6302), .A2(n6137), .B1(n6126), .B2(n6156), .ZN(n4537)
         );
  AOI21_X1 U5638 ( .B1(n6294), .B2(n6132), .A(n4537), .ZN(n4538) );
  OAI211_X1 U5639 ( .C1(n4546), .C2(n6301), .A(n4539), .B(n4538), .ZN(U3044)
         );
  NAND2_X1 U5640 ( .A1(n6134), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4542) );
  OAI22_X1 U5641 ( .A1(n6274), .A2(n6137), .B1(n6126), .B2(n6340), .ZN(n4540)
         );
  AOI21_X1 U5642 ( .B1(n6338), .B2(n6132), .A(n4540), .ZN(n4541) );
  OAI211_X1 U5643 ( .C1(n4546), .C2(n6339), .A(n4542), .B(n4541), .ZN(U3049)
         );
  NAND2_X1 U5644 ( .A1(n6134), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4545) );
  OAI22_X1 U5645 ( .A1(n6269), .A2(n6137), .B1(n6126), .B2(n6332), .ZN(n4543)
         );
  AOI21_X1 U5646 ( .B1(n6330), .B2(n6132), .A(n4543), .ZN(n4544) );
  OAI211_X1 U5647 ( .C1(n4546), .C2(n6331), .A(n4545), .B(n4544), .ZN(U3048)
         );
  NOR2_X1 U5648 ( .A1(n6287), .A2(n4551), .ZN(n4547) );
  INV_X1 U5649 ( .A(n4547), .ZN(n4573) );
  AOI21_X1 U5650 ( .B1(n4548), .B2(n6369), .A(n4547), .ZN(n4552) );
  AOI21_X1 U5651 ( .B1(n4554), .B2(STATEBS16_REG_SCAN_IN), .A(n6295), .ZN(
        n4550) );
  AOI22_X1 U5652 ( .A1(n4552), .A2(n4550), .B1(n6295), .B2(n4551), .ZN(n4549)
         );
  NAND2_X1 U5653 ( .A1(n6208), .A2(n4549), .ZN(n4570) );
  INV_X1 U5654 ( .A(n4550), .ZN(n4553) );
  OAI22_X1 U5655 ( .A1(n4553), .A2(n4552), .B1(n6210), .B2(n4551), .ZN(n4569)
         );
  AOI22_X1 U5656 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4570), .B1(n6350), 
        .B2(n4569), .ZN(n4556) );
  NAND2_X1 U5657 ( .A1(n4554), .A2(n3574), .ZN(n5565) );
  AOI22_X1 U5658 ( .A1(n5573), .A2(n6348), .B1(n4647), .B2(n6346), .ZN(n4555)
         );
  OAI211_X1 U5659 ( .C1(n4887), .C2(n4573), .A(n4556), .B(n4555), .ZN(U3034)
         );
  AOI22_X1 U5660 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4570), .B1(n6243), 
        .B2(n4569), .ZN(n4558) );
  AOI22_X1 U5661 ( .A1(n5573), .A2(n6293), .B1(n4647), .B2(n6153), .ZN(n4557)
         );
  OAI211_X1 U5662 ( .C1(n5544), .C2(n4573), .A(n4558), .B(n4557), .ZN(U3028)
         );
  AOI22_X1 U5663 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4570), .B1(n6256), 
        .B2(n4569), .ZN(n4560) );
  AOI22_X1 U5664 ( .A1(n5573), .A2(n6306), .B1(n4647), .B2(n6157), .ZN(n4559)
         );
  OAI211_X1 U5665 ( .C1(n5548), .C2(n4573), .A(n4560), .B(n4559), .ZN(U3029)
         );
  AOI22_X1 U5666 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4570), .B1(n6262), 
        .B2(n4569), .ZN(n4562) );
  AOI22_X1 U5667 ( .A1(n5573), .A2(n6321), .B1(n4647), .B2(n6220), .ZN(n4561)
         );
  OAI211_X1 U5668 ( .C1(n5556), .C2(n4573), .A(n4562), .B(n4561), .ZN(U3031)
         );
  AOI22_X1 U5669 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4570), .B1(n6270), 
        .B2(n4569), .ZN(n4564) );
  AOI22_X1 U5670 ( .A1(n5573), .A2(n6271), .B1(n4647), .B2(n6337), .ZN(n4563)
         );
  OAI211_X1 U5671 ( .C1(n5564), .C2(n4573), .A(n4564), .B(n4563), .ZN(U3033)
         );
  AOI22_X1 U5672 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4570), .B1(n6265), 
        .B2(n4569), .ZN(n4566) );
  AOI22_X1 U5673 ( .A1(n5573), .A2(n6266), .B1(n4647), .B2(n6329), .ZN(n4565)
         );
  OAI211_X1 U5674 ( .C1(n5560), .C2(n4573), .A(n4566), .B(n4565), .ZN(U3032)
         );
  AOI22_X1 U5675 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4570), .B1(n6279), 
        .B2(n4569), .ZN(n4568) );
  INV_X1 U5676 ( .A(n6181), .ZN(n6355) );
  AOI22_X1 U5677 ( .A1(n5573), .A2(n6355), .B1(n4647), .B2(n6177), .ZN(n4567)
         );
  OAI211_X1 U5678 ( .C1(n5576), .C2(n4573), .A(n4568), .B(n4567), .ZN(U3035)
         );
  AOI22_X1 U5679 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4570), .B1(n6259), 
        .B2(n4569), .ZN(n4572) );
  AOI22_X1 U5680 ( .A1(n5573), .A2(n6313), .B1(n4647), .B2(n6161), .ZN(n4571)
         );
  OAI211_X1 U5681 ( .C1(n5552), .C2(n4573), .A(n4572), .B(n4571), .ZN(U3030)
         );
  OAI21_X1 U5682 ( .B1(n4869), .B2(n4574), .A(n6245), .ZN(n4578) );
  INV_X1 U5683 ( .A(n4575), .ZN(n4781) );
  NAND3_X1 U5684 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6589), .A3(n6373), .ZN(n4777) );
  NOR2_X1 U5685 ( .A1(n6287), .A2(n4777), .ZN(n4597) );
  AOI21_X1 U5686 ( .B1(n6286), .B2(n4781), .A(n4597), .ZN(n4579) );
  INV_X1 U5687 ( .A(n4579), .ZN(n4577) );
  AOI21_X1 U5688 ( .B1(n6295), .B2(n4777), .A(n6291), .ZN(n4576) );
  OAI21_X1 U5689 ( .B1(n4578), .B2(n4577), .A(n4576), .ZN(n4596) );
  OAI22_X1 U5690 ( .A1(n4579), .A2(n4578), .B1(n6210), .B2(n4777), .ZN(n4595)
         );
  AOI22_X1 U5691 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4596), .B1(n6350), 
        .B2(n4595), .ZN(n4582) );
  NAND2_X1 U5692 ( .A1(n4580), .A2(n3574), .ZN(n4871) );
  AOI22_X1 U5693 ( .A1(n6347), .A2(n4597), .B1(n4903), .B2(n6348), .ZN(n4581)
         );
  OAI211_X1 U5694 ( .C1(n6277), .C2(n4820), .A(n4582), .B(n4581), .ZN(U3098)
         );
  AOI22_X1 U5695 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4596), .B1(n6243), 
        .B2(n4595), .ZN(n4584) );
  AOI22_X1 U5696 ( .A1(n6294), .A2(n4597), .B1(n4903), .B2(n6293), .ZN(n4583)
         );
  OAI211_X1 U5697 ( .C1(n6302), .C2(n4820), .A(n4584), .B(n4583), .ZN(U3092)
         );
  AOI22_X1 U5698 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4596), .B1(n6256), 
        .B2(n4595), .ZN(n4586) );
  AOI22_X1 U5699 ( .A1(n6307), .A2(n4597), .B1(n4903), .B2(n6306), .ZN(n4585)
         );
  OAI211_X1 U5700 ( .C1(n6309), .C2(n4820), .A(n4586), .B(n4585), .ZN(U3093)
         );
  AOI22_X1 U5701 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4596), .B1(n6270), 
        .B2(n4595), .ZN(n4588) );
  AOI22_X1 U5702 ( .A1(n6338), .A2(n4597), .B1(n4903), .B2(n6271), .ZN(n4587)
         );
  OAI211_X1 U5703 ( .C1(n6274), .C2(n4820), .A(n4588), .B(n4587), .ZN(U3097)
         );
  AOI22_X1 U5704 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4596), .B1(n6265), 
        .B2(n4595), .ZN(n4590) );
  AOI22_X1 U5705 ( .A1(n6330), .A2(n4597), .B1(n4903), .B2(n6266), .ZN(n4589)
         );
  OAI211_X1 U5706 ( .C1(n6269), .C2(n4820), .A(n4590), .B(n4589), .ZN(U3096)
         );
  AOI22_X1 U5707 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4596), .B1(n6262), 
        .B2(n4595), .ZN(n4592) );
  AOI22_X1 U5708 ( .A1(n6322), .A2(n4597), .B1(n4903), .B2(n6321), .ZN(n4591)
         );
  OAI211_X1 U5709 ( .C1(n6324), .C2(n4820), .A(n4592), .B(n4591), .ZN(U3095)
         );
  AOI22_X1 U5710 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4596), .B1(n6259), 
        .B2(n4595), .ZN(n4594) );
  AOI22_X1 U5711 ( .A1(n6314), .A2(n4597), .B1(n4903), .B2(n6313), .ZN(n4593)
         );
  OAI211_X1 U5712 ( .C1(n6316), .C2(n4820), .A(n4594), .B(n4593), .ZN(U3094)
         );
  AOI22_X1 U5713 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4596), .B1(n6279), 
        .B2(n4595), .ZN(n4599) );
  AOI22_X1 U5714 ( .A1(n6357), .A2(n4597), .B1(n4903), .B2(n6355), .ZN(n4598)
         );
  OAI211_X1 U5715 ( .C1(n6360), .C2(n4820), .A(n4599), .B(n4598), .ZN(U3099)
         );
  NOR2_X1 U5716 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4600), .ZN(n4633)
         );
  INV_X1 U5717 ( .A(n4633), .ZN(n4629) );
  OAI21_X1 U5718 ( .B1(n6140), .B2(n6210), .A(n4601), .ZN(n6146) );
  NOR3_X1 U5719 ( .A1(n6146), .A2(n6201), .A3(n6147), .ZN(n4605) );
  OR2_X1 U5720 ( .A1(n4602), .A2(n5521), .ZN(n6244) );
  OR2_X1 U5721 ( .A1(n6244), .A2(n4696), .ZN(n6341) );
  OAI21_X1 U5722 ( .B1(n6354), .B2(n4606), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4603) );
  NAND3_X1 U5723 ( .A1(n6145), .A2(n6245), .A3(n4603), .ZN(n4604) );
  NAND2_X1 U5724 ( .A1(n4630), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4610)
         );
  NOR2_X1 U5725 ( .A1(n6145), .A2(n6295), .ZN(n6139) );
  INV_X1 U5726 ( .A(n6141), .ZN(n6239) );
  NOR2_X1 U5727 ( .A1(n6239), .A2(n6201), .ZN(n4607) );
  AOI22_X1 U5728 ( .A1(n6139), .A2(n6143), .B1(n6140), .B2(n4607), .ZN(n4636)
         );
  OAI22_X1 U5729 ( .A1(n4631), .A2(n6332), .B1(n4636), .B2(n6331), .ZN(n4608)
         );
  AOI21_X1 U5730 ( .B1(n6329), .B2(n6354), .A(n4608), .ZN(n4609) );
  OAI211_X1 U5731 ( .C1(n4629), .C2(n5560), .A(n4610), .B(n4609), .ZN(U3136)
         );
  NAND2_X1 U5732 ( .A1(n4630), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4613)
         );
  OAI22_X1 U5733 ( .A1(n4631), .A2(n6340), .B1(n4636), .B2(n6339), .ZN(n4611)
         );
  AOI21_X1 U5734 ( .B1(n6337), .B2(n6354), .A(n4611), .ZN(n4612) );
  OAI211_X1 U5735 ( .C1(n4629), .C2(n5564), .A(n4613), .B(n4612), .ZN(U3137)
         );
  NAND2_X1 U5736 ( .A1(n4630), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4616)
         );
  OAI22_X1 U5737 ( .A1(n4631), .A2(n6181), .B1(n4636), .B2(n6358), .ZN(n4614)
         );
  AOI21_X1 U5738 ( .B1(n6177), .B2(n6354), .A(n4614), .ZN(n4615) );
  OAI211_X1 U5739 ( .C1(n4629), .C2(n5576), .A(n4616), .B(n4615), .ZN(U3139)
         );
  NAND2_X1 U5740 ( .A1(n4630), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4619)
         );
  OAI22_X1 U5741 ( .A1(n4631), .A2(n6223), .B1(n4636), .B2(n6323), .ZN(n4617)
         );
  AOI21_X1 U5742 ( .B1(n6220), .B2(n6354), .A(n4617), .ZN(n4618) );
  OAI211_X1 U5743 ( .C1(n4629), .C2(n5556), .A(n4619), .B(n4618), .ZN(U3135)
         );
  NAND2_X1 U5744 ( .A1(n4630), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4622)
         );
  OAI22_X1 U5745 ( .A1(n4631), .A2(n6156), .B1(n4636), .B2(n6301), .ZN(n4620)
         );
  AOI21_X1 U5746 ( .B1(n6153), .B2(n6354), .A(n4620), .ZN(n4621) );
  OAI211_X1 U5747 ( .C1(n5544), .C2(n4629), .A(n4622), .B(n4621), .ZN(U3132)
         );
  NAND2_X1 U5748 ( .A1(n4630), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4625)
         );
  OAI22_X1 U5749 ( .A1(n4631), .A2(n6160), .B1(n4636), .B2(n6308), .ZN(n4623)
         );
  AOI21_X1 U5750 ( .B1(n6157), .B2(n6354), .A(n4623), .ZN(n4624) );
  OAI211_X1 U5751 ( .C1(n4629), .C2(n5548), .A(n4625), .B(n4624), .ZN(U3133)
         );
  NAND2_X1 U5752 ( .A1(n4630), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4628)
         );
  OAI22_X1 U5753 ( .A1(n4631), .A2(n6164), .B1(n4636), .B2(n6315), .ZN(n4626)
         );
  AOI21_X1 U5754 ( .B1(n6161), .B2(n6354), .A(n4626), .ZN(n4627) );
  OAI211_X1 U5755 ( .C1(n4629), .C2(n5552), .A(n4628), .B(n4627), .ZN(U3134)
         );
  NAND2_X1 U5756 ( .A1(n4630), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4635)
         );
  OAI22_X1 U5757 ( .A1(n4631), .A2(n6173), .B1(n6341), .B2(n6277), .ZN(n4632)
         );
  AOI21_X1 U5758 ( .B1(n6347), .B2(n4633), .A(n4632), .ZN(n4634) );
  OAI211_X1 U5759 ( .C1(n4636), .C2(n5585), .A(n4635), .B(n4634), .ZN(U3138)
         );
  INV_X1 U5760 ( .A(n4637), .ZN(n4643) );
  NAND2_X1 U5761 ( .A1(n4643), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4642) );
  INV_X1 U5762 ( .A(n4647), .ZN(n4638) );
  OAI22_X1 U5763 ( .A1(n4638), .A2(n6173), .B1(n6277), .B2(n4645), .ZN(n4639)
         );
  AOI21_X1 U5764 ( .B1(n6347), .B2(n4640), .A(n4639), .ZN(n4641) );
  OAI211_X1 U5765 ( .C1(n4644), .C2(n5585), .A(n4642), .B(n4641), .ZN(U3026)
         );
  NAND2_X1 U5766 ( .A1(n4643), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4649) );
  OAI22_X1 U5767 ( .A1(n4645), .A2(n6360), .B1(n4644), .B2(n6358), .ZN(n4646)
         );
  AOI21_X1 U5768 ( .B1(n4647), .B2(n6355), .A(n4646), .ZN(n4648) );
  OAI211_X1 U5769 ( .C1(n4650), .C2(n5576), .A(n4649), .B(n4648), .ZN(U3027)
         );
  INV_X1 U5770 ( .A(n6247), .ZN(n4651) );
  NOR2_X1 U5771 ( .A1(n3366), .A2(n4651), .ZN(n4652) );
  XNOR2_X1 U5772 ( .A(n4652), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5752)
         );
  OAI22_X1 U5773 ( .A1(n5752), .A2(n4653), .B1(n5758), .B2(n6371), .ZN(n4655)
         );
  NAND2_X1 U5774 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5766), .ZN(n4684) );
  INV_X1 U5775 ( .A(n4684), .ZN(n4654) );
  AOI22_X1 U5776 ( .A1(n4655), .A2(n6488), .B1(n4654), .B2(
        INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4686) );
  INV_X1 U5777 ( .A(n4657), .ZN(n4683) );
  XNOR2_X1 U5778 ( .A(n3115), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4666)
         );
  OR2_X1 U5779 ( .A1(n4659), .A2(n4658), .ZN(n4673) );
  INV_X1 U5780 ( .A(n4678), .ZN(n4662) );
  XNOR2_X1 U5781 ( .A(n4660), .B(n3115), .ZN(n4661) );
  MUX2_X1 U5782 ( .A(n4673), .B(n4662), .S(n4661), .Z(n4665) );
  NOR2_X1 U5783 ( .A1(n5526), .A2(n4663), .ZN(n4664) );
  AOI211_X1 U5784 ( .C1(n6370), .C2(n4666), .A(n4665), .B(n4664), .ZN(n4667)
         );
  INV_X1 U5785 ( .A(n4667), .ZN(n5025) );
  MUX2_X1 U5786 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n5025), .S(n6371), 
        .Z(n6378) );
  NAND2_X1 U5787 ( .A1(n4660), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4668) );
  NAND2_X1 U5788 ( .A1(n4668), .A2(n4680), .ZN(n4669) );
  NAND2_X1 U5789 ( .A1(n3287), .A2(n4669), .ZN(n5529) );
  MUX2_X1 U5790 ( .A(n4670), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4660), 
        .Z(n4671) );
  NOR2_X1 U5791 ( .A1(n4671), .A2(n4657), .ZN(n4672) );
  NAND2_X1 U5792 ( .A1(n4673), .A2(n4672), .ZN(n4677) );
  NAND2_X1 U5793 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4674) );
  XNOR2_X1 U5794 ( .A(n4674), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4675)
         );
  NAND2_X1 U5795 ( .A1(n6370), .A2(n4675), .ZN(n4676) );
  OAI211_X1 U5796 ( .C1(n4678), .C2(n5529), .A(n4677), .B(n4676), .ZN(n4679)
         );
  AOI21_X1 U5797 ( .B1(n6143), .B2(n6368), .A(n4679), .ZN(n5530) );
  MUX2_X1 U5798 ( .A(n4680), .B(n5530), .S(n6371), .Z(n6379) );
  INV_X1 U5799 ( .A(n6379), .ZN(n4681) );
  NAND3_X1 U5800 ( .A1(n6378), .A2(n4681), .A3(n6488), .ZN(n4682) );
  OAI211_X1 U5801 ( .C1(n4684), .C2(n4683), .A(n4682), .B(n4686), .ZN(n6386)
         );
  INV_X1 U5802 ( .A(n6386), .ZN(n4685) );
  AOI21_X1 U5803 ( .B1(n4686), .B2(n4656), .A(n4685), .ZN(n4695) );
  NOR2_X1 U5804 ( .A1(n4695), .A2(FLUSH_REG_SCAN_IN), .ZN(n4687) );
  INV_X1 U5805 ( .A(n4688), .ZN(n4691) );
  INV_X1 U5806 ( .A(n4782), .ZN(n6248) );
  AND2_X1 U5807 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6487), .ZN(n5525) );
  OAI22_X1 U5808 ( .A1(n4689), .A2(n6248), .B1(n6241), .B2(n5525), .ZN(n4690)
         );
  OAI21_X1 U5809 ( .B1(n4691), .B2(n4690), .A(n6124), .ZN(n4692) );
  OAI21_X1 U5810 ( .B1(n6124), .B2(n6201), .A(n4692), .ZN(U3462) );
  INV_X1 U5811 ( .A(n4693), .ZN(n4694) );
  NOR2_X1 U5812 ( .A1(n4695), .A2(n4694), .ZN(n6394) );
  OAI22_X1 U5813 ( .A1(n4696), .A2(n6295), .B1(n3576), .B2(n5525), .ZN(n4697)
         );
  OAI21_X1 U5814 ( .B1(n6394), .B2(n4697), .A(n6124), .ZN(n4698) );
  OAI21_X1 U5815 ( .B1(n6124), .B2(n6287), .A(n4698), .ZN(U3465) );
  NAND3_X1 U5816 ( .A1(n5580), .A2(n6245), .A3(n6126), .ZN(n4700) );
  AOI21_X1 U5817 ( .B1(n4700), .B2(n6248), .A(n4699), .ZN(n4703) );
  NOR2_X1 U5818 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4701), .ZN(n5582)
         );
  INV_X1 U5819 ( .A(n6147), .ZN(n6251) );
  OAI21_X1 U5820 ( .B1(n5582), .B2(n6487), .A(n6251), .ZN(n4702) );
  NOR3_X2 U5821 ( .A1(n4704), .A2(n4703), .A3(n4702), .ZN(n5578) );
  INV_X1 U5822 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4708) );
  NOR2_X1 U5823 ( .A1(n6246), .A2(n6295), .ZN(n6238) );
  AOI22_X1 U5824 ( .A1(n6238), .A2(n6241), .B1(n6141), .B2(n3109), .ZN(n5586)
         );
  OAI22_X1 U5825 ( .A1(n6126), .A2(n6274), .B1(n5586), .B2(n6339), .ZN(n4706)
         );
  NOR2_X1 U5826 ( .A1(n5580), .A2(n6340), .ZN(n4705) );
  AOI211_X1 U5827 ( .C1(n5582), .C2(n6338), .A(n4706), .B(n4705), .ZN(n4707)
         );
  OAI21_X1 U5828 ( .B1(n5578), .B2(n4708), .A(n4707), .ZN(U3057) );
  INV_X1 U5829 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4712) );
  OAI22_X1 U5830 ( .A1(n6126), .A2(n6269), .B1(n5586), .B2(n6331), .ZN(n4710)
         );
  NOR2_X1 U5831 ( .A1(n5580), .A2(n6332), .ZN(n4709) );
  AOI211_X1 U5832 ( .C1(n5582), .C2(n6330), .A(n4710), .B(n4709), .ZN(n4711)
         );
  OAI21_X1 U5833 ( .B1(n5578), .B2(n4712), .A(n4711), .ZN(U3056) );
  INV_X1 U5834 ( .A(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4716) );
  OAI22_X1 U5835 ( .A1(n6126), .A2(n6324), .B1(n5586), .B2(n6323), .ZN(n4714)
         );
  NOR2_X1 U5836 ( .A1(n5580), .A2(n6223), .ZN(n4713) );
  AOI211_X1 U5837 ( .C1(n5582), .C2(n6322), .A(n4714), .B(n4713), .ZN(n4715)
         );
  OAI21_X1 U5838 ( .B1(n5578), .B2(n4716), .A(n4715), .ZN(U3055) );
  INV_X1 U5839 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4720) );
  OAI22_X1 U5840 ( .A1(n6126), .A2(n6316), .B1(n5586), .B2(n6315), .ZN(n4718)
         );
  NOR2_X1 U5841 ( .A1(n5580), .A2(n6164), .ZN(n4717) );
  AOI211_X1 U5842 ( .C1(n5582), .C2(n6314), .A(n4718), .B(n4717), .ZN(n4719)
         );
  OAI21_X1 U5843 ( .B1(n5578), .B2(n4720), .A(n4719), .ZN(U3054) );
  INV_X1 U5844 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4724) );
  OAI22_X1 U5845 ( .A1(n6126), .A2(n6309), .B1(n5586), .B2(n6308), .ZN(n4722)
         );
  NOR2_X1 U5846 ( .A1(n5580), .A2(n6160), .ZN(n4721) );
  AOI211_X1 U5847 ( .C1(n5582), .C2(n6307), .A(n4722), .B(n4721), .ZN(n4723)
         );
  OAI21_X1 U5848 ( .B1(n5578), .B2(n4724), .A(n4723), .ZN(U3053) );
  INV_X1 U5849 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4728) );
  OAI22_X1 U5850 ( .A1(n6126), .A2(n6360), .B1(n5586), .B2(n6358), .ZN(n4726)
         );
  NOR2_X1 U5851 ( .A1(n5580), .A2(n6181), .ZN(n4725) );
  AOI211_X1 U5852 ( .C1(n5582), .C2(n6357), .A(n4726), .B(n4725), .ZN(n4727)
         );
  OAI21_X1 U5853 ( .B1(n5578), .B2(n4728), .A(n4727), .ZN(U3059) );
  INV_X1 U5854 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4732) );
  OAI22_X1 U5855 ( .A1(n6126), .A2(n6302), .B1(n5586), .B2(n6301), .ZN(n4730)
         );
  NOR2_X1 U5856 ( .A1(n5580), .A2(n6156), .ZN(n4729) );
  AOI211_X1 U5857 ( .C1(n5582), .C2(n6294), .A(n4730), .B(n4729), .ZN(n4731)
         );
  OAI21_X1 U5858 ( .B1(n5578), .B2(n4732), .A(n4731), .ZN(U3052) );
  NAND2_X1 U5859 ( .A1(n4733), .A2(n6245), .ZN(n4738) );
  NOR2_X1 U5860 ( .A1(n3576), .A2(n6247), .ZN(n4735) );
  INV_X1 U5861 ( .A(n4734), .ZN(n6195) );
  AOI21_X1 U5862 ( .B1(n4736), .B2(n4735), .A(n6195), .ZN(n4740) );
  INV_X1 U5863 ( .A(n4742), .ZN(n6138) );
  OAI22_X1 U5864 ( .A1(n4738), .A2(n4740), .B1(n6138), .B2(n6210), .ZN(n6196)
         );
  INV_X1 U5865 ( .A(n6196), .ZN(n4746) );
  INV_X1 U5866 ( .A(n4738), .ZN(n4739) );
  NAND2_X1 U5867 ( .A1(n4740), .A2(n4739), .ZN(n4741) );
  OAI211_X1 U5868 ( .C1(n4742), .C2(n6245), .A(n6208), .B(n4741), .ZN(n6197)
         );
  AOI22_X1 U5869 ( .A1(n6194), .A2(n6293), .B1(INSTQUEUE_REG_7__0__SCAN_IN), 
        .B2(n6197), .ZN(n4743) );
  OAI21_X1 U5870 ( .B1(n6302), .B2(n6200), .A(n4743), .ZN(n4744) );
  AOI21_X1 U5871 ( .B1(n6294), .B2(n6195), .A(n4744), .ZN(n4745) );
  OAI21_X1 U5872 ( .B1(n4746), .B2(n6301), .A(n4745), .ZN(U3076) );
  AOI22_X1 U5873 ( .A1(n5943), .A2(UWORD_REG_14__SCAN_IN), .B1(n5934), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4747) );
  OAI21_X1 U5874 ( .B1(n4059), .B2(n4758), .A(n4747), .ZN(U2893) );
  AOI22_X1 U5875 ( .A1(UWORD_REG_3__SCAN_IN), .A2(n5943), .B1(n5934), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4748) );
  OAI21_X1 U5876 ( .B1(n3815), .B2(n4758), .A(n4748), .ZN(U2904) );
  INV_X1 U5877 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4750) );
  AOI22_X1 U5878 ( .A1(n5943), .A2(UWORD_REG_5__SCAN_IN), .B1(n5934), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4749) );
  OAI21_X1 U5879 ( .B1(n4750), .B2(n4758), .A(n4749), .ZN(U2902) );
  INV_X1 U5880 ( .A(EAX_REG_23__SCAN_IN), .ZN(n6636) );
  AOI22_X1 U5881 ( .A1(n5943), .A2(UWORD_REG_7__SCAN_IN), .B1(n5934), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4751) );
  OAI21_X1 U5882 ( .B1(n6636), .B2(n4758), .A(n4751), .ZN(U2900) );
  INV_X1 U5883 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4753) );
  AOI22_X1 U5884 ( .A1(n5943), .A2(UWORD_REG_1__SCAN_IN), .B1(n5934), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4752) );
  OAI21_X1 U5885 ( .B1(n4753), .B2(n4758), .A(n4752), .ZN(U2906) );
  INV_X1 U5886 ( .A(EAX_REG_25__SCAN_IN), .ZN(n5959) );
  AOI22_X1 U5887 ( .A1(n5943), .A2(UWORD_REG_9__SCAN_IN), .B1(n5934), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4754) );
  OAI21_X1 U5888 ( .B1(n5959), .B2(n4758), .A(n4754), .ZN(U2898) );
  INV_X1 U5889 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4756) );
  AOI22_X1 U5890 ( .A1(n5943), .A2(UWORD_REG_4__SCAN_IN), .B1(n5934), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4755) );
  OAI21_X1 U5891 ( .B1(n4756), .B2(n4758), .A(n4755), .ZN(U2903) );
  INV_X1 U5892 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4759) );
  AOI22_X1 U5893 ( .A1(n5943), .A2(UWORD_REG_6__SCAN_IN), .B1(n5934), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4757) );
  OAI21_X1 U5894 ( .B1(n4759), .B2(n4758), .A(n4757), .ZN(U2901) );
  OR2_X1 U5895 ( .A1(n4761), .A2(n4760), .ZN(n4762) );
  NAND2_X1 U5896 ( .A1(n4824), .A2(n4762), .ZN(n5872) );
  XOR2_X1 U5897 ( .A(n4481), .B(n4763), .Z(n6019) );
  INV_X1 U5898 ( .A(n6019), .ZN(n5001) );
  INV_X1 U5899 ( .A(EBX_REG_6__SCAN_IN), .ZN(n5878) );
  OAI222_X1 U5900 ( .A1(n5872), .A2(n5901), .B1(n5212), .B2(n5001), .C1(n5905), 
        .C2(n5878), .ZN(U2853) );
  AOI21_X1 U5901 ( .B1(n4766), .B2(n4765), .A(n4764), .ZN(n5017) );
  INV_X1 U5902 ( .A(n4767), .ZN(n4946) );
  INV_X1 U5903 ( .A(n4768), .ZN(n6110) );
  OAI21_X1 U5904 ( .B1(n6056), .B2(n6110), .A(n6054), .ZN(n6109) );
  AOI21_X1 U5905 ( .B1(n4946), .B2(n5730), .A(n6109), .ZN(n4947) );
  AOI221_X1 U5906 ( .B1(n6088), .B2(n4770), .C1(n4769), .C2(n4770), .A(n4947), 
        .ZN(n4775) );
  NAND3_X1 U5907 ( .A1(n4771), .A2(n6108), .A3(n4770), .ZN(n4773) );
  NAND2_X1 U5908 ( .A1(n6112), .A2(REIP_REG_5__SCAN_IN), .ZN(n4772) );
  OAI211_X1 U5909 ( .C1(n4923), .C2(n6116), .A(n4773), .B(n4772), .ZN(n4774)
         );
  AOI211_X1 U5910 ( .C1(n5017), .C2(n6119), .A(n4775), .B(n4774), .ZN(n4776)
         );
  INV_X1 U5911 ( .A(n4776), .ZN(U3013) );
  NOR2_X1 U5912 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4777), .ZN(n4817)
         );
  INV_X1 U5913 ( .A(n4817), .ZN(n4802) );
  OR2_X1 U5914 ( .A1(n6140), .A2(n4778), .ZN(n6240) );
  AOI21_X1 U5915 ( .B1(n6240), .B2(STATE2_REG_2__SCAN_IN), .A(n4779), .ZN(
        n6250) );
  INV_X1 U5916 ( .A(n6250), .ZN(n4780) );
  AOI211_X1 U5917 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4802), .A(n6141), .B(
        n4780), .ZN(n4785) );
  INV_X1 U5918 ( .A(n4820), .ZN(n4804) );
  NOR3_X1 U5919 ( .A1(n4804), .A2(n6194), .A3(n6295), .ZN(n4783) );
  NAND2_X1 U5920 ( .A1(n4781), .A2(n6143), .ZN(n4786) );
  OAI21_X1 U5921 ( .B1(n4783), .B2(n4782), .A(n4786), .ZN(n4784) );
  NAND2_X1 U5922 ( .A1(n4785), .A2(n4784), .ZN(n4813) );
  NAND2_X1 U5923 ( .A1(n4813), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4792) );
  OR2_X1 U5924 ( .A1(n4786), .A2(n6295), .ZN(n4789) );
  INV_X1 U5925 ( .A(n6240), .ZN(n4787) );
  NAND2_X1 U5926 ( .A1(n6147), .A2(n4787), .ZN(n4788) );
  OAI22_X1 U5927 ( .A1(n4815), .A2(n6302), .B1(n4814), .B2(n6301), .ZN(n4790)
         );
  AOI21_X1 U5928 ( .B1(n6294), .B2(n4817), .A(n4790), .ZN(n4791) );
  OAI211_X1 U5929 ( .C1(n4820), .C2(n6156), .A(n4792), .B(n4791), .ZN(U3084)
         );
  NAND2_X1 U5930 ( .A1(n4813), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4795) );
  OAI22_X1 U5931 ( .A1(n4815), .A2(n6309), .B1(n4814), .B2(n6308), .ZN(n4793)
         );
  AOI21_X1 U5932 ( .B1(n6307), .B2(n4817), .A(n4793), .ZN(n4794) );
  OAI211_X1 U5933 ( .C1(n4820), .C2(n6160), .A(n4795), .B(n4794), .ZN(U3085)
         );
  NAND2_X1 U5934 ( .A1(n4813), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4798) );
  OAI22_X1 U5935 ( .A1(n4815), .A2(n6316), .B1(n4814), .B2(n6315), .ZN(n4796)
         );
  AOI21_X1 U5936 ( .B1(n6314), .B2(n4817), .A(n4796), .ZN(n4797) );
  OAI211_X1 U5937 ( .C1(n4820), .C2(n6164), .A(n4798), .B(n4797), .ZN(U3086)
         );
  NAND2_X1 U5938 ( .A1(n4813), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4801) );
  OAI22_X1 U5939 ( .A1(n4815), .A2(n6324), .B1(n4814), .B2(n6323), .ZN(n4799)
         );
  AOI21_X1 U5940 ( .B1(n6322), .B2(n4817), .A(n4799), .ZN(n4800) );
  OAI211_X1 U5941 ( .C1(n4820), .C2(n6223), .A(n4801), .B(n4800), .ZN(U3087)
         );
  NAND2_X1 U5942 ( .A1(n4813), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4806) );
  OAI22_X1 U5943 ( .A1(n4887), .A2(n4802), .B1(n6277), .B2(n4815), .ZN(n4803)
         );
  AOI21_X1 U5944 ( .B1(n6348), .B2(n4804), .A(n4803), .ZN(n4805) );
  OAI211_X1 U5945 ( .C1(n4814), .C2(n5585), .A(n4806), .B(n4805), .ZN(U3090)
         );
  NAND2_X1 U5946 ( .A1(n4813), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4809) );
  OAI22_X1 U5947 ( .A1(n4815), .A2(n6360), .B1(n4814), .B2(n6358), .ZN(n4807)
         );
  AOI21_X1 U5948 ( .B1(n6357), .B2(n4817), .A(n4807), .ZN(n4808) );
  OAI211_X1 U5949 ( .C1(n4820), .C2(n6181), .A(n4809), .B(n4808), .ZN(U3091)
         );
  NAND2_X1 U5950 ( .A1(n4813), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4812) );
  OAI22_X1 U5951 ( .A1(n4815), .A2(n6269), .B1(n4814), .B2(n6331), .ZN(n4810)
         );
  AOI21_X1 U5952 ( .B1(n6330), .B2(n4817), .A(n4810), .ZN(n4811) );
  OAI211_X1 U5953 ( .C1(n4820), .C2(n6332), .A(n4812), .B(n4811), .ZN(U3088)
         );
  NAND2_X1 U5954 ( .A1(n4813), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4819) );
  OAI22_X1 U5955 ( .A1(n4815), .A2(n6274), .B1(n4814), .B2(n6339), .ZN(n4816)
         );
  AOI21_X1 U5956 ( .B1(n6338), .B2(n4817), .A(n4816), .ZN(n4818) );
  OAI211_X1 U5957 ( .C1(n4820), .C2(n6340), .A(n4819), .B(n4818), .ZN(U3089)
         );
  XNOR2_X1 U5958 ( .A(n4821), .B(n4822), .ZN(n5862) );
  INV_X1 U5959 ( .A(n4908), .ZN(n4823) );
  AOI21_X1 U5960 ( .B1(n4825), .B2(n4824), .A(n4823), .ZN(n6081) );
  AOI22_X1 U5961 ( .A1(n6081), .A2(n6518), .B1(n6517), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n4826) );
  OAI21_X1 U5962 ( .B1(n5862), .B2(n5212), .A(n4826), .ZN(U2852) );
  NAND2_X1 U5963 ( .A1(n4828), .A2(n4827), .ZN(n4834) );
  NAND2_X1 U5964 ( .A1(n4832), .A2(n4831), .ZN(n4833) );
  AND2_X1 U5965 ( .A1(n3248), .A2(n3320), .ZN(n4835) );
  OR2_X2 U5966 ( .A1(n5909), .A2(n4835), .ZN(n5666) );
  INV_X1 U5967 ( .A(n4835), .ZN(n4836) );
  INV_X1 U5968 ( .A(EAX_REG_4__SCAN_IN), .ZN(n5936) );
  OAI222_X1 U5969 ( .A1(n5666), .A2(n4837), .B1(n5242), .B2(n5980), .C1(n5241), 
        .C2(n5936), .ZN(U2887) );
  INV_X1 U5970 ( .A(EAX_REG_0__SCAN_IN), .ZN(n5946) );
  OAI222_X1 U5971 ( .A1(n5666), .A2(n6044), .B1(n5242), .B2(n5972), .C1(n5241), 
        .C2(n5946), .ZN(U2891) );
  AND2_X1 U5972 ( .A1(n4838), .A2(n2977), .ZN(n6402) );
  NOR3_X1 U5973 ( .A1(n6509), .A2(n6487), .A3(n6508), .ZN(n6393) );
  OR2_X1 U5974 ( .A1(n6402), .A2(n6393), .ZN(n4839) );
  NOR2_X1 U5975 ( .A1(n6112), .A2(n4839), .ZN(n4840) );
  OR2_X1 U5976 ( .A1(n5038), .A2(n4841), .ZN(n4842) );
  NOR2_X1 U5977 ( .A1(n5038), .A2(n4843), .ZN(n5888) );
  INV_X1 U5978 ( .A(n5888), .ZN(n4958) );
  NAND2_X1 U5979 ( .A1(n6599), .A2(n6638), .ZN(n4848) );
  OR2_X1 U5980 ( .A1(n6413), .A2(n4848), .ZN(n6392) );
  INV_X1 U5981 ( .A(n4848), .ZN(n4851) );
  NOR2_X1 U5982 ( .A1(EBX_REG_31__SCAN_IN), .A2(n4851), .ZN(n4844) );
  AOI22_X1 U5983 ( .A1(n6507), .A2(n6392), .B1(n4844), .B2(n4852), .ZN(n4845)
         );
  OAI22_X1 U5984 ( .A1(n4958), .A2(n5523), .B1(n5894), .B2(n4846), .ZN(n4863)
         );
  INV_X1 U5985 ( .A(n4847), .ZN(n4855) );
  NAND3_X1 U5986 ( .A1(n4849), .A2(EBX_REG_31__SCAN_IN), .A3(n4848), .ZN(n4850) );
  NAND3_X1 U5987 ( .A1(n4853), .A2(n4852), .A3(n4851), .ZN(n4854) );
  OAI22_X1 U5988 ( .A1(n4855), .A2(n5873), .B1(n5826), .B2(REIP_REG_1__SCAN_IN), .ZN(n4862) );
  INV_X1 U5989 ( .A(n4856), .ZN(n4857) );
  NOR2_X1 U5990 ( .A1(n5889), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4861)
         );
  INV_X1 U5991 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4859) );
  NAND2_X1 U5992 ( .A1(n5034), .A2(REIP_REG_1__SCAN_IN), .ZN(n4858) );
  OAI21_X1 U5993 ( .B1(n5890), .B2(n4859), .A(n4858), .ZN(n4860) );
  NOR4_X1 U5994 ( .A1(n4863), .A2(n4862), .A3(n4861), .A4(n4860), .ZN(n4864)
         );
  OAI21_X1 U5995 ( .B1(n4998), .B2(n5899), .A(n4864), .ZN(U2826) );
  INV_X1 U5996 ( .A(EAX_REG_7__SCAN_IN), .ZN(n5930) );
  OAI222_X1 U5997 ( .A1(n5666), .A2(n5862), .B1(n5242), .B2(n5986), .C1(n5241), 
        .C2(n5930), .ZN(U2884) );
  OR2_X1 U5998 ( .A1(n4867), .A2(n4866), .ZN(n4868) );
  NAND2_X1 U5999 ( .A1(n4929), .A2(n4868), .ZN(n5383) );
  INV_X1 U6000 ( .A(DATAI_8_), .ZN(n5988) );
  INV_X1 U6001 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6550) );
  OAI222_X1 U6002 ( .A1(n5383), .A2(n5666), .B1(n5242), .B2(n5988), .C1(n5241), 
        .C2(n6550), .ZN(U2883) );
  NAND2_X1 U6003 ( .A1(n4871), .A2(n6237), .ZN(n4872) );
  AOI21_X1 U6004 ( .B1(n4872), .B2(STATEBS16_REG_SCAN_IN), .A(n6295), .ZN(
        n4876) );
  AND2_X1 U6005 ( .A1(n4873), .A2(n6143), .ZN(n6206) );
  NOR2_X1 U6006 ( .A1(n6251), .A2(n6201), .ZN(n4874) );
  AOI22_X1 U6007 ( .A1(n4876), .A2(n6206), .B1(n6140), .B2(n4874), .ZN(n4906)
         );
  NOR2_X1 U6008 ( .A1(n6141), .A2(n6146), .ZN(n5536) );
  INV_X1 U6009 ( .A(n6206), .ZN(n4875) );
  NAND3_X1 U6010 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6589), .ZN(n6211) );
  OR2_X1 U6011 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6211), .ZN(n4901)
         );
  AOI22_X1 U6012 ( .A1(n4876), .A2(n4875), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n4901), .ZN(n4877) );
  OAI211_X1 U6013 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6210), .A(n5536), .B(n4877), .ZN(n4900) );
  NAND2_X1 U6014 ( .A1(n4900), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4880)
         );
  OAI22_X1 U6015 ( .A1(n5556), .A2(n4901), .B1(n6237), .B2(n6223), .ZN(n4878)
         );
  AOI21_X1 U6016 ( .B1(n4903), .B2(n6220), .A(n4878), .ZN(n4879) );
  OAI211_X1 U6017 ( .C1(n4906), .C2(n6323), .A(n4880), .B(n4879), .ZN(U3103)
         );
  NAND2_X1 U6018 ( .A1(n4900), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4883)
         );
  OAI22_X1 U6019 ( .A1(n5544), .A2(n4901), .B1(n6237), .B2(n6156), .ZN(n4881)
         );
  AOI21_X1 U6020 ( .B1(n4903), .B2(n6153), .A(n4881), .ZN(n4882) );
  OAI211_X1 U6021 ( .C1(n4906), .C2(n6301), .A(n4883), .B(n4882), .ZN(U3100)
         );
  NAND2_X1 U6022 ( .A1(n4900), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4886)
         );
  OAI22_X1 U6023 ( .A1(n5576), .A2(n4901), .B1(n6237), .B2(n6181), .ZN(n4884)
         );
  AOI21_X1 U6024 ( .B1(n4903), .B2(n6177), .A(n4884), .ZN(n4885) );
  OAI211_X1 U6025 ( .C1(n4906), .C2(n6358), .A(n4886), .B(n4885), .ZN(U3107)
         );
  NAND2_X1 U6026 ( .A1(n4900), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4890)
         );
  OAI22_X1 U6027 ( .A1(n4887), .A2(n4901), .B1(n6237), .B2(n6173), .ZN(n4888)
         );
  AOI21_X1 U6028 ( .B1(n4903), .B2(n6346), .A(n4888), .ZN(n4889) );
  OAI211_X1 U6029 ( .C1(n4906), .C2(n5585), .A(n4890), .B(n4889), .ZN(U3106)
         );
  NAND2_X1 U6030 ( .A1(n4900), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4893)
         );
  OAI22_X1 U6031 ( .A1(n5560), .A2(n4901), .B1(n6237), .B2(n6332), .ZN(n4891)
         );
  AOI21_X1 U6032 ( .B1(n4903), .B2(n6329), .A(n4891), .ZN(n4892) );
  OAI211_X1 U6033 ( .C1(n4906), .C2(n6331), .A(n4893), .B(n4892), .ZN(U3104)
         );
  NAND2_X1 U6034 ( .A1(n4900), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4896)
         );
  OAI22_X1 U6035 ( .A1(n5552), .A2(n4901), .B1(n6237), .B2(n6164), .ZN(n4894)
         );
  AOI21_X1 U6036 ( .B1(n4903), .B2(n6161), .A(n4894), .ZN(n4895) );
  OAI211_X1 U6037 ( .C1(n4906), .C2(n6315), .A(n4896), .B(n4895), .ZN(U3102)
         );
  NAND2_X1 U6038 ( .A1(n4900), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4899)
         );
  OAI22_X1 U6039 ( .A1(n5548), .A2(n4901), .B1(n6237), .B2(n6160), .ZN(n4897)
         );
  AOI21_X1 U6040 ( .B1(n4903), .B2(n6157), .A(n4897), .ZN(n4898) );
  OAI211_X1 U6041 ( .C1(n4906), .C2(n6308), .A(n4899), .B(n4898), .ZN(U3101)
         );
  NAND2_X1 U6042 ( .A1(n4900), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4905)
         );
  OAI22_X1 U6043 ( .A1(n5564), .A2(n4901), .B1(n6237), .B2(n6340), .ZN(n4902)
         );
  AOI21_X1 U6044 ( .B1(n4903), .B2(n6337), .A(n4902), .ZN(n4904) );
  OAI211_X1 U6045 ( .C1(n4906), .C2(n6339), .A(n4905), .B(n4904), .ZN(U3105)
         );
  NAND2_X1 U6046 ( .A1(n4908), .A2(n4907), .ZN(n4909) );
  NAND2_X1 U6047 ( .A1(n4932), .A2(n4909), .ZN(n6072) );
  INV_X1 U6048 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4910) );
  OAI222_X1 U6049 ( .A1(n6072), .A2(n5901), .B1(n5905), .B2(n4910), .C1(n5212), 
        .C2(n5383), .ZN(U2851) );
  INV_X1 U6050 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6439) );
  NAND2_X1 U6051 ( .A1(REIP_REG_7__SCAN_IN), .A2(REIP_REG_6__SCAN_IN), .ZN(
        n5856) );
  NOR2_X1 U6052 ( .A1(n6439), .A2(n5856), .ZN(n5032) );
  INV_X1 U6053 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6633) );
  INV_X1 U6054 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6496) );
  INV_X1 U6055 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6431) );
  NOR3_X1 U6056 ( .A1(n6633), .A2(n6496), .A3(n6431), .ZN(n4956) );
  NAND3_X1 U6057 ( .A1(REIP_REG_5__SCAN_IN), .A2(REIP_REG_4__SCAN_IN), .A3(
        n4956), .ZN(n5033) );
  NOR2_X1 U6058 ( .A1(n5034), .A2(n5033), .ZN(n4919) );
  INV_X1 U6059 ( .A(n5034), .ZN(n5132) );
  NAND2_X1 U6060 ( .A1(n5826), .A2(n5132), .ZN(n5887) );
  AOI21_X1 U6061 ( .B1(n5032), .B2(n4919), .A(n5620), .ZN(n5847) );
  NAND3_X1 U6062 ( .A1(n5802), .A2(n4956), .A3(REIP_REG_4__SCAN_IN), .ZN(n4920) );
  INV_X1 U6063 ( .A(n4920), .ZN(n4911) );
  NAND2_X1 U6064 ( .A1(n4911), .A2(REIP_REG_5__SCAN_IN), .ZN(n5883) );
  OAI21_X1 U6065 ( .B1(n5856), .B2(n5883), .A(n6439), .ZN(n4912) );
  NAND2_X1 U6066 ( .A1(n5847), .A2(n4912), .ZN(n4918) );
  INV_X1 U6067 ( .A(n5385), .ZN(n4916) );
  OAI21_X1 U6068 ( .B1(n5890), .B2(n3635), .A(n5858), .ZN(n4915) );
  OAI22_X1 U6069 ( .A1(n4910), .A2(n5894), .B1(n5873), .B2(n6072), .ZN(n4914)
         );
  AOI211_X1 U6070 ( .C1(n5870), .C2(n4916), .A(n4915), .B(n4914), .ZN(n4917)
         );
  OAI211_X1 U6071 ( .C1(n5383), .C2(n5861), .A(n4918), .B(n4917), .ZN(U2819)
         );
  NOR2_X1 U6072 ( .A1(n5620), .A2(n4919), .ZN(n5869) );
  INV_X1 U6073 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6436) );
  NAND2_X1 U6074 ( .A1(n6436), .A2(n4920), .ZN(n4921) );
  NAND2_X1 U6075 ( .A1(n5869), .A2(n4921), .ZN(n4928) );
  OAI21_X1 U6076 ( .B1(n5890), .B2(n4922), .A(n5858), .ZN(n4926) );
  OAI22_X1 U6077 ( .A1(n4924), .A2(n5894), .B1(n5873), .B2(n4923), .ZN(n4925)
         );
  AOI211_X1 U6078 ( .C1(n5870), .C2(n5012), .A(n4926), .B(n4925), .ZN(n4927)
         );
  OAI211_X1 U6079 ( .C1(n5899), .C2(n5015), .A(n4928), .B(n4927), .ZN(U2822)
         );
  OAI21_X1 U6080 ( .B1(n3655), .B2(n3654), .A(n4931), .ZN(n5849) );
  AOI21_X1 U6081 ( .B1(n4933), .B2(n4932), .A(n5514), .ZN(n6065) );
  AOI22_X1 U6082 ( .A1(n6065), .A2(n6518), .B1(EBX_REG_9__SCAN_IN), .B2(n6517), 
        .ZN(n4934) );
  OAI21_X1 U6083 ( .B1(n5849), .B2(n5212), .A(n4934), .ZN(U2850) );
  OAI21_X1 U6084 ( .B1(n5826), .B2(REIP_REG_1__SCAN_IN), .A(n5132), .ZN(n4987)
         );
  NAND3_X1 U6085 ( .A1(n5802), .A2(REIP_REG_1__SCAN_IN), .A3(n6633), .ZN(n4938) );
  INV_X1 U6086 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n4935) );
  OAI22_X1 U6087 ( .A1(n5890), .A2(n4935), .B1(n5889), .B2(n6039), .ZN(n4936)
         );
  INV_X1 U6088 ( .A(n4936), .ZN(n4937) );
  OAI211_X1 U6089 ( .C1(n4939), .C2(n5894), .A(n4938), .B(n4937), .ZN(n4941)
         );
  OAI22_X1 U6090 ( .A1(n4958), .A2(n5526), .B1(n5873), .B2(n6115), .ZN(n4940)
         );
  AOI211_X1 U6091 ( .C1(REIP_REG_2__SCAN_IN), .C2(n4987), .A(n4941), .B(n4940), 
        .ZN(n4942) );
  OAI21_X1 U6092 ( .B1(n4997), .B2(n5899), .A(n4942), .ZN(U2825) );
  AOI21_X1 U6093 ( .B1(n4945), .B2(n4944), .A(n4943), .ZN(n6020) );
  AOI21_X1 U6094 ( .B1(n6110), .B2(n6108), .A(n6111), .ZN(n6092) );
  NOR2_X1 U6095 ( .A1(n4946), .A2(n6092), .ZN(n4949) );
  INV_X1 U6096 ( .A(n4947), .ZN(n4948) );
  MUX2_X1 U6097 ( .A(n4949), .B(n4948), .S(INSTADDRPOINTER_REG_6__SCAN_IN), 
        .Z(n4952) );
  INV_X1 U6098 ( .A(REIP_REG_6__SCAN_IN), .ZN(n4950) );
  OAI22_X1 U6099 ( .A1(n6116), .A2(n5872), .B1(n6071), .B2(n4950), .ZN(n4951)
         );
  AOI211_X1 U6100 ( .C1(n6020), .C2(n6119), .A(n4952), .B(n4951), .ZN(n4953)
         );
  INV_X1 U6101 ( .A(n4953), .ZN(U3012) );
  INV_X1 U6102 ( .A(n5899), .ZN(n4993) );
  INV_X1 U6103 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6433) );
  INV_X1 U6104 ( .A(n4956), .ZN(n4954) );
  OAI21_X1 U6105 ( .B1(n5034), .B2(n4954), .A(n5887), .ZN(n4989) );
  INV_X1 U6106 ( .A(n6030), .ZN(n4961) );
  INV_X1 U6107 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4955) );
  OAI21_X1 U6108 ( .B1(n5890), .B2(n4955), .A(n5858), .ZN(n4960) );
  NAND3_X1 U6109 ( .A1(n5802), .A2(n4956), .A3(n6433), .ZN(n4957) );
  OAI21_X1 U6110 ( .B1(n4958), .B2(n5752), .A(n4957), .ZN(n4959) );
  AOI211_X1 U6111 ( .C1(n5870), .C2(n4961), .A(n4960), .B(n4959), .ZN(n4963)
         );
  AOI22_X1 U6112 ( .A1(n5865), .A2(EBX_REG_4__SCAN_IN), .B1(n5886), .B2(n6090), 
        .ZN(n4962) );
  OAI211_X1 U6113 ( .C1(n6433), .C2(n4989), .A(n4963), .B(n4962), .ZN(n4964)
         );
  AOI21_X1 U6114 ( .B1(n6027), .B2(n4993), .A(n4964), .ZN(n4965) );
  INV_X1 U6115 ( .A(n4965), .ZN(U2823) );
  INV_X1 U6116 ( .A(n4998), .ZN(n4969) );
  AOI21_X1 U6117 ( .B1(n6047), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4966), 
        .ZN(n4967) );
  OAI21_X1 U6118 ( .B1(n6040), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4967), 
        .ZN(n4968) );
  AOI21_X1 U6119 ( .B1(n4969), .B2(n6035), .A(n4968), .ZN(n4970) );
  OAI21_X1 U6120 ( .B1(n4971), .B2(n6041), .A(n4970), .ZN(U2985) );
  NOR2_X1 U6121 ( .A1(n4972), .A2(n4973), .ZN(n4974) );
  OR2_X1 U6122 ( .A1(n4975), .A2(n4974), .ZN(n6101) );
  INV_X1 U6123 ( .A(n4983), .ZN(n4977) );
  AND2_X1 U6124 ( .A1(n6112), .A2(REIP_REG_3__SCAN_IN), .ZN(n6098) );
  AOI21_X1 U6125 ( .B1(n6047), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n6098), 
        .ZN(n4976) );
  OAI21_X1 U6126 ( .B1(n6040), .B2(n4977), .A(n4976), .ZN(n4978) );
  AOI21_X1 U6127 ( .B1(n4994), .B2(n6035), .A(n4978), .ZN(n4979) );
  OAI21_X1 U6128 ( .B1(n6041), .B2(n6101), .A(n4979), .ZN(U2983) );
  NAND2_X1 U6129 ( .A1(n5888), .A2(n6143), .ZN(n4985) );
  OAI22_X1 U6130 ( .A1(n4981), .A2(n5894), .B1(n4980), .B2(n5890), .ZN(n4982)
         );
  AOI21_X1 U6131 ( .B1(n5870), .B2(n4983), .A(n4982), .ZN(n4984) );
  OAI211_X1 U6132 ( .C1(n4986), .C2(n5873), .A(n4985), .B(n4984), .ZN(n4992)
         );
  INV_X1 U6133 ( .A(n4987), .ZN(n4988) );
  NAND2_X1 U6134 ( .A1(n4988), .A2(REIP_REG_2__SCAN_IN), .ZN(n4990) );
  AOI21_X1 U6135 ( .B1(n6431), .B2(n4990), .A(n4989), .ZN(n4991) );
  AOI211_X1 U6136 ( .C1(n4994), .C2(n4993), .A(n4992), .B(n4991), .ZN(n4995)
         );
  INV_X1 U6137 ( .A(n4995), .ZN(U2824) );
  AOI22_X1 U6138 ( .A1(n5249), .A2(DATAI_9_), .B1(EAX_REG_9__SCAN_IN), .B2(
        n5909), .ZN(n4996) );
  OAI21_X1 U6139 ( .B1(n5849), .B2(n5666), .A(n4996), .ZN(U2882) );
  INV_X1 U6140 ( .A(EAX_REG_5__SCAN_IN), .ZN(n5933) );
  OAI222_X1 U6141 ( .A1(n5015), .A2(n5666), .B1(n5242), .B2(n5982), .C1(n5241), 
        .C2(n5933), .ZN(U2886) );
  INV_X1 U6142 ( .A(EAX_REG_2__SCAN_IN), .ZN(n5940) );
  OAI222_X1 U6143 ( .A1(n4997), .A2(n5666), .B1(n5242), .B2(n5976), .C1(n5241), 
        .C2(n5940), .ZN(U2889) );
  INV_X1 U6144 ( .A(EAX_REG_1__SCAN_IN), .ZN(n5942) );
  OAI222_X1 U6145 ( .A1(n4998), .A2(n5666), .B1(n5242), .B2(n5974), .C1(n5241), 
        .C2(n5942), .ZN(U2890) );
  INV_X1 U6146 ( .A(EAX_REG_3__SCAN_IN), .ZN(n5938) );
  OAI222_X1 U6147 ( .A1(n4999), .A2(n5666), .B1(n5242), .B2(n5978), .C1(n5241), 
        .C2(n5938), .ZN(U2888) );
  OAI222_X1 U6148 ( .A1(n5242), .A2(n5984), .B1(n5666), .B2(n5001), .C1(n5000), 
        .C2(n5241), .ZN(U2885) );
  NAND2_X1 U6149 ( .A1(n4931), .A2(n5002), .ZN(n5003) );
  NAND2_X1 U6150 ( .A1(n5247), .A2(n5003), .ZN(n5372) );
  NOR3_X1 U6151 ( .A1(n5883), .A2(n6439), .A3(n5856), .ZN(n5850) );
  INV_X1 U6152 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6442) );
  XNOR2_X1 U6153 ( .A(REIP_REG_10__SCAN_IN), .B(n6442), .ZN(n5004) );
  AOI22_X1 U6154 ( .A1(REIP_REG_10__SCAN_IN), .A2(n5847), .B1(n5850), .B2(
        n5004), .ZN(n5009) );
  INV_X1 U6155 ( .A(n5368), .ZN(n5007) );
  XNOR2_X1 U6156 ( .A(n5514), .B(n5513), .ZN(n5011) );
  INV_X1 U6157 ( .A(n5011), .ZN(n6052) );
  AOI22_X1 U6158 ( .A1(n6052), .A2(n5886), .B1(n5865), .B2(EBX_REG_10__SCAN_IN), .ZN(n5005) );
  OAI211_X1 U6159 ( .C1(n5890), .C2(n3657), .A(n5005), .B(n5858), .ZN(n5006)
         );
  AOI21_X1 U6160 ( .B1(n5870), .B2(n5007), .A(n5006), .ZN(n5008) );
  OAI211_X1 U6161 ( .C1(n5861), .C2(n5372), .A(n5009), .B(n5008), .ZN(U2817)
         );
  INV_X1 U6162 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5010) );
  OAI222_X1 U6163 ( .A1(n5372), .A2(n5212), .B1(n5901), .B2(n5011), .C1(n5905), 
        .C2(n5010), .ZN(U2849) );
  INV_X1 U6164 ( .A(DATAI_10_), .ZN(n5993) );
  INV_X1 U6165 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6601) );
  OAI222_X1 U6166 ( .A1(n5372), .A2(n5666), .B1(n5242), .B2(n5993), .C1(n5241), 
        .C2(n6601), .ZN(U2881) );
  AOI22_X1 U6167 ( .A1(n6047), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .B1(n5705), 
        .B2(REIP_REG_5__SCAN_IN), .ZN(n5014) );
  NAND2_X1 U6168 ( .A1(n5395), .A2(n5012), .ZN(n5013) );
  OAI211_X1 U6169 ( .C1(n5015), .C2(n6043), .A(n5014), .B(n5013), .ZN(n5016)
         );
  AOI21_X1 U6170 ( .B1(n5017), .B2(n6036), .A(n5016), .ZN(n5018) );
  INV_X1 U6171 ( .A(n5018), .ZN(U2981) );
  INV_X1 U6172 ( .A(n4660), .ZN(n5019) );
  AOI21_X1 U6173 ( .B1(n5019), .B2(n5020), .A(n5531), .ZN(n5027) );
  NAND3_X1 U6174 ( .A1(n4660), .A2(n3115), .A3(n5020), .ZN(n5021) );
  OAI21_X1 U6175 ( .B1(n5023), .B2(n5022), .A(n5021), .ZN(n5024) );
  AOI21_X1 U6176 ( .B1(n5025), .B2(n5754), .A(n5024), .ZN(n5026) );
  OAI22_X1 U6177 ( .A1(n5027), .A2(n3115), .B1(n5531), .B2(n5026), .ZN(U3459)
         );
  NAND3_X1 U6178 ( .A1(n5031), .A2(n4388), .A3(n5241), .ZN(n5030) );
  AOI22_X1 U6179 ( .A1(n3004), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n5909), .ZN(n5029) );
  NAND2_X1 U6180 ( .A1(n5030), .A2(n5029), .ZN(U2860) );
  NAND2_X1 U6181 ( .A1(n5031), .A2(n5880), .ZN(n5047) );
  INV_X1 U6182 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6474) );
  INV_X1 U6183 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6458) );
  NAND2_X1 U6184 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5647) );
  INV_X1 U6185 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6607) );
  INV_X1 U6186 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6445) );
  NAND3_X1 U6187 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .A3(
        n5032), .ZN(n5839) );
  NOR3_X1 U6188 ( .A1(n6445), .A2(n5033), .A3(n5839), .ZN(n5133) );
  NAND2_X1 U6189 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5133), .ZN(n5825) );
  NOR2_X1 U6190 ( .A1(n6607), .A2(n5825), .ZN(n5121) );
  NAND2_X1 U6191 ( .A1(REIP_REG_14__SCAN_IN), .A2(n5121), .ZN(n5040) );
  NOR2_X1 U6192 ( .A1(n5034), .A2(n5040), .ZN(n5122) );
  NAND4_X1 U6193 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .A4(n5122), .ZN(n5648) );
  NOR3_X1 U6194 ( .A1(n6458), .A2(n5647), .A3(n5648), .ZN(n5619) );
  NAND4_X1 U6195 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5619), .ZN(n5101) );
  NAND3_X1 U6196 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n5042) );
  OAI21_X1 U6197 ( .B1(n5101), .B2(n5042), .A(n5887), .ZN(n5598) );
  INV_X1 U6198 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6470) );
  INV_X1 U6199 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6468) );
  OR2_X1 U6200 ( .A1(n6470), .A2(n6468), .ZN(n5035) );
  NAND2_X1 U6201 ( .A1(n5802), .A2(n5035), .ZN(n5036) );
  NAND2_X1 U6202 ( .A1(n5598), .A2(n5036), .ZN(n5587) );
  AOI21_X1 U6203 ( .B1(n5802), .B2(n6474), .A(n5587), .ZN(n5063) );
  OAI21_X1 U6204 ( .B1(REIP_REG_30__SCAN_IN), .B2(n5826), .A(n5063), .ZN(n5045) );
  NAND3_X1 U6205 ( .A1(n6507), .A2(EBX_REG_31__SCAN_IN), .A3(n6392), .ZN(n5037) );
  OAI22_X1 U6206 ( .A1(n5039), .A2(n5890), .B1(n5038), .B2(n5037), .ZN(n5044)
         );
  INV_X1 U6207 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6452) );
  INV_X1 U6208 ( .A(n5040), .ZN(n5801) );
  AND2_X1 U6209 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5801), .ZN(n5041) );
  NAND2_X1 U6210 ( .A1(n5802), .A2(n5041), .ZN(n5803) );
  NAND2_X1 U6211 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5797), .ZN(n5790) );
  NAND2_X1 U6212 ( .A1(REIP_REG_20__SCAN_IN), .A2(n5642), .ZN(n5637) );
  NAND2_X1 U6213 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n5625) );
  NAND2_X1 U6214 ( .A1(REIP_REG_23__SCAN_IN), .A2(n5609), .ZN(n5601) );
  NAND3_X1 U6215 ( .A1(n5592), .A2(REIP_REG_28__SCAN_IN), .A3(
        REIP_REG_27__SCAN_IN), .ZN(n5070) );
  INV_X1 U6216 ( .A(REIP_REG_30__SCAN_IN), .ZN(n5062) );
  NOR4_X1 U6217 ( .A1(n5070), .A2(REIP_REG_31__SCAN_IN), .A3(n5062), .A4(n6474), .ZN(n5043) );
  AOI211_X1 U6218 ( .C1(REIP_REG_31__SCAN_IN), .C2(n5045), .A(n5044), .B(n5043), .ZN(n5046) );
  OAI211_X1 U6219 ( .C1(n5141), .C2(n5873), .A(n5047), .B(n5046), .ZN(U2796)
         );
  INV_X1 U6220 ( .A(n5048), .ZN(n5049) );
  INV_X1 U6221 ( .A(n5259), .ZN(n5217) );
  INV_X1 U6222 ( .A(n5053), .ZN(n5050) );
  OAI211_X1 U6223 ( .C1(n5052), .C2(n5073), .A(n5051), .B(n5050), .ZN(n5057)
         );
  OAI211_X1 U6224 ( .C1(n5055), .C2(n5149), .A(n5054), .B(n5053), .ZN(n5056)
         );
  NAND2_X1 U6225 ( .A1(n5057), .A2(n5056), .ZN(n5142) );
  INV_X1 U6226 ( .A(n5058), .ZN(n5257) );
  OAI22_X1 U6227 ( .A1(n5059), .A2(n5890), .B1(n5889), .B2(n5257), .ZN(n5060)
         );
  AOI21_X1 U6228 ( .B1(EBX_REG_30__SCAN_IN), .B2(n5865), .A(n5060), .ZN(n5061)
         );
  OAI21_X1 U6229 ( .B1(n5063), .B2(n5062), .A(n5061), .ZN(n5065) );
  NOR3_X1 U6230 ( .A1(n5070), .A2(REIP_REG_30__SCAN_IN), .A3(n6474), .ZN(n5064) );
  AOI211_X1 U6231 ( .C1(n5886), .C2(n5142), .A(n5065), .B(n5064), .ZN(n5066)
         );
  OAI21_X1 U6232 ( .B1(n5217), .B2(n5861), .A(n5066), .ZN(U2797) );
  INV_X1 U6233 ( .A(n5268), .ZN(n5220) );
  INV_X1 U6234 ( .A(n5070), .ZN(n5083) );
  INV_X1 U6235 ( .A(n5071), .ZN(n5074) );
  AOI21_X1 U6236 ( .B1(n5074), .B2(n5073), .A(n5072), .ZN(n5075) );
  AND2_X1 U6237 ( .A1(n5149), .A2(n5075), .ZN(n5076) );
  OAI22_X1 U6238 ( .A1(n5078), .A2(n5890), .B1(n5889), .B2(n5266), .ZN(n5079)
         );
  AOI21_X1 U6239 ( .B1(n5865), .B2(EBX_REG_29__SCAN_IN), .A(n5079), .ZN(n5081)
         );
  NAND2_X1 U6240 ( .A1(n5587), .A2(REIP_REG_29__SCAN_IN), .ZN(n5080) );
  OAI211_X1 U6241 ( .C1(n5411), .C2(n5873), .A(n5081), .B(n5080), .ZN(n5082)
         );
  AOI21_X1 U6242 ( .B1(n5083), .B2(n6474), .A(n5082), .ZN(n5084) );
  OAI21_X1 U6243 ( .B1(n5220), .B2(n5861), .A(n5084), .ZN(U2798) );
  OAI21_X1 U6244 ( .B1(n5152), .B2(n5085), .A(n5145), .ZN(n5280) );
  INV_X1 U6245 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5086) );
  OAI22_X1 U6246 ( .A1(n5086), .A2(n5890), .B1(n6468), .B2(n5598), .ZN(n5093)
         );
  NAND2_X1 U6247 ( .A1(n2984), .A2(n5087), .ZN(n5088) );
  AND2_X1 U6248 ( .A1(n2991), .A2(n5088), .ZN(n5430) );
  INV_X1 U6249 ( .A(n5430), .ZN(n5091) );
  NOR2_X1 U6250 ( .A1(n5282), .A2(n5889), .ZN(n5089) );
  AOI21_X1 U6251 ( .B1(n5865), .B2(EBX_REG_27__SCAN_IN), .A(n5089), .ZN(n5090)
         );
  OAI21_X1 U6252 ( .B1(n5091), .B2(n5873), .A(n5090), .ZN(n5092) );
  AOI211_X1 U6253 ( .C1(n5592), .C2(n6468), .A(n5093), .B(n5092), .ZN(n5094)
         );
  OAI21_X1 U6254 ( .B1(n5280), .B2(n5861), .A(n5094), .ZN(U2800) );
  AND2_X1 U6255 ( .A1(n4091), .A2(n5095), .ZN(n5097) );
  INV_X1 U6256 ( .A(n5601), .ZN(n5098) );
  NAND2_X1 U6257 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n5600) );
  OAI211_X1 U6258 ( .C1(REIP_REG_24__SCAN_IN), .C2(REIP_REG_25__SCAN_IN), .A(
        n5098), .B(n5600), .ZN(n5109) );
  AOI21_X1 U6259 ( .B1(n5164), .B2(n5110), .A(n5099), .ZN(n5100) );
  NAND2_X1 U6260 ( .A1(n5887), .A2(n5101), .ZN(n5617) );
  INV_X1 U6261 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6465) );
  OAI22_X1 U6262 ( .A1(n5890), .A2(n5102), .B1(n5617), .B2(n6465), .ZN(n5103)
         );
  AOI21_X1 U6263 ( .B1(n5104), .B2(n5870), .A(n5103), .ZN(n5105) );
  OAI21_X1 U6264 ( .B1(n5106), .B2(n5894), .A(n5105), .ZN(n5107) );
  AOI21_X1 U6265 ( .B1(n3006), .B2(n5886), .A(n5107), .ZN(n5108) );
  OAI211_X1 U6266 ( .C1(n5674), .C2(n5861), .A(n5109), .B(n5108), .ZN(U2802)
         );
  XOR2_X1 U6267 ( .A(n5110), .B(n5164), .Z(n5450) );
  AOI22_X1 U6268 ( .A1(EBX_REG_24__SCAN_IN), .A2(n5865), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n5876), .ZN(n5111) );
  OAI21_X1 U6269 ( .B1(n4092), .B2(n5617), .A(n5111), .ZN(n5114) );
  OAI22_X1 U6270 ( .A1(n5889), .A2(n5112), .B1(REIP_REG_24__SCAN_IN), .B2(
        n5601), .ZN(n5113) );
  AOI211_X1 U6271 ( .C1(n5450), .C2(n5886), .A(n5114), .B(n5113), .ZN(n5115)
         );
  OAI21_X1 U6272 ( .B1(n5232), .B2(n5861), .A(n5115), .ZN(U2803) );
  AND2_X1 U6273 ( .A1(n5211), .A2(n5116), .ZN(n5118) );
  OR2_X1 U6274 ( .A1(n5118), .A2(n5117), .ZN(n5344) );
  AOI21_X1 U6275 ( .B1(n5119), .B2(n5209), .A(n5200), .ZN(n5492) );
  OAI21_X1 U6276 ( .B1(n5890), .B2(n5120), .A(n5858), .ZN(n5126) );
  NAND2_X1 U6277 ( .A1(n5802), .A2(n5121), .ZN(n5124) );
  INV_X1 U6278 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6449) );
  OR2_X1 U6279 ( .A1(n5620), .A2(n5122), .ZN(n5823) );
  AOI22_X1 U6280 ( .A1(EBX_REG_14__SCAN_IN), .A2(n5865), .B1(n5345), .B2(n5870), .ZN(n5123) );
  OAI221_X1 U6281 ( .B1(REIP_REG_14__SCAN_IN), .B2(n5124), .C1(n6449), .C2(
        n5823), .A(n5123), .ZN(n5125) );
  AOI211_X1 U6282 ( .C1(n5492), .C2(n5886), .A(n5126), .B(n5125), .ZN(n5127)
         );
  OAI21_X1 U6283 ( .B1(n5344), .B2(n5861), .A(n5127), .ZN(U2813) );
  OAI21_X1 U6284 ( .B1(n5516), .B2(n5128), .A(n5207), .ZN(n5495) );
  INV_X1 U6285 ( .A(n5129), .ZN(n5131) );
  INV_X1 U6286 ( .A(n3015), .ZN(n5130) );
  AOI21_X1 U6287 ( .B1(n5131), .B2(n5130), .A(n3005), .ZN(n5363) );
  NAND2_X1 U6288 ( .A1(n5363), .A2(n5880), .ZN(n5139) );
  OAI21_X1 U6289 ( .B1(n5826), .B2(n5133), .A(n5132), .ZN(n5837) );
  INV_X1 U6290 ( .A(n5133), .ZN(n5134) );
  NOR3_X1 U6291 ( .A1(n5826), .A2(REIP_REG_12__SCAN_IN), .A3(n5134), .ZN(n5834) );
  AOI21_X1 U6292 ( .B1(n5865), .B2(EBX_REG_12__SCAN_IN), .A(n5834), .ZN(n5136)
         );
  AOI21_X1 U6293 ( .B1(n5876), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n5875), 
        .ZN(n5135) );
  OAI211_X1 U6294 ( .C1(n5361), .C2(n5889), .A(n5136), .B(n5135), .ZN(n5137)
         );
  AOI21_X1 U6295 ( .B1(REIP_REG_12__SCAN_IN), .B2(n5837), .A(n5137), .ZN(n5138) );
  OAI211_X1 U6296 ( .C1(n5495), .C2(n5873), .A(n5139), .B(n5138), .ZN(U2815)
         );
  INV_X1 U6297 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5140) );
  OAI22_X1 U6298 ( .A1(n5141), .A2(n5901), .B1(n5140), .B2(n5905), .ZN(U2828)
         );
  INV_X1 U6299 ( .A(n5142), .ZN(n5402) );
  INV_X1 U6300 ( .A(EBX_REG_30__SCAN_IN), .ZN(n6560) );
  OAI222_X1 U6301 ( .A1(n5217), .A2(n5212), .B1(n5901), .B2(n5402), .C1(n5905), 
        .C2(n6560), .ZN(U2829) );
  OAI222_X1 U6302 ( .A1(n5143), .A2(n5905), .B1(n5901), .B2(n5411), .C1(n5220), 
        .C2(n5902), .ZN(U2830) );
  NAND2_X1 U6303 ( .A1(n5145), .A2(n5144), .ZN(n5146) );
  NAND2_X1 U6304 ( .A1(n2991), .A2(n5147), .ZN(n5148) );
  NAND2_X1 U6305 ( .A1(n5149), .A2(n5148), .ZN(n5589) );
  INV_X1 U6306 ( .A(n5589), .ZN(n5422) );
  AOI22_X1 U6307 ( .A1(n5422), .A2(n6518), .B1(n6517), .B2(EBX_REG_28__SCAN_IN), .ZN(n5150) );
  OAI21_X1 U6308 ( .B1(n5223), .B2(n5902), .A(n5150), .ZN(U2831) );
  AOI22_X1 U6309 ( .A1(n5430), .A2(n6518), .B1(n6517), .B2(EBX_REG_27__SCAN_IN), .ZN(n5151) );
  OAI21_X1 U6310 ( .B1(n5280), .B2(n5902), .A(n5151), .ZN(U2832) );
  OAI21_X1 U6311 ( .B1(n5154), .B2(n5096), .A(n5153), .ZN(n5603) );
  INV_X1 U6312 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5158) );
  OR2_X1 U6313 ( .A1(n5156), .A2(n5155), .ZN(n5157) );
  NAND2_X1 U6314 ( .A1(n2984), .A2(n5157), .ZN(n5602) );
  OAI222_X1 U6315 ( .A1(n5212), .A2(n5603), .B1(n5905), .B2(n5158), .C1(n5602), 
        .C2(n5901), .ZN(U2833) );
  AOI22_X1 U6316 ( .A1(n5450), .A2(n6518), .B1(EBX_REG_24__SCAN_IN), .B2(n6517), .ZN(n5159) );
  OAI21_X1 U6317 ( .B1(n5232), .B2(n5902), .A(n5159), .ZN(U2835) );
  INV_X1 U6318 ( .A(n5160), .ZN(n5163) );
  INV_X1 U6319 ( .A(n5161), .ZN(n5162) );
  INV_X1 U6320 ( .A(n5614), .ZN(n5235) );
  AOI21_X1 U6321 ( .B1(n5165), .B2(n5171), .A(n5164), .ZN(n5613) );
  AOI22_X1 U6322 ( .A1(n5613), .A2(n6518), .B1(EBX_REG_23__SCAN_IN), .B2(n6517), .ZN(n5166) );
  OAI21_X1 U6323 ( .B1(n5235), .B2(n5902), .A(n5166), .ZN(U2836) );
  OR2_X1 U6324 ( .A1(n5310), .A2(n5309), .ZN(n5312) );
  OR2_X1 U6325 ( .A1(n3107), .A2(n5161), .ZN(n5623) );
  NAND2_X1 U6326 ( .A1(n5472), .A2(n5169), .ZN(n5170) );
  NAND2_X1 U6327 ( .A1(n5171), .A2(n5170), .ZN(n5622) );
  OAI22_X1 U6328 ( .A1(n5622), .A2(n5901), .B1(n5172), .B2(n5905), .ZN(n5173)
         );
  INV_X1 U6329 ( .A(n5173), .ZN(n5174) );
  OAI21_X1 U6330 ( .B1(n5623), .B2(n5212), .A(n5174), .ZN(U2837) );
  OAI21_X1 U6331 ( .B1(n3835), .B2(n3111), .A(n5310), .ZN(n5640) );
  MUX2_X1 U6332 ( .A(n5181), .B(n5182), .S(n5176), .Z(n5178) );
  XNOR2_X1 U6333 ( .A(n5178), .B(n5177), .ZN(n5698) );
  INV_X1 U6334 ( .A(n5698), .ZN(n5639) );
  OAI222_X1 U6335 ( .A1(n5640), .A2(n5212), .B1(n5901), .B2(n5639), .C1(n5905), 
        .C2(n4188), .ZN(U2839) );
  AND2_X1 U6336 ( .A1(n5187), .A2(n5179), .ZN(n5180) );
  OR2_X1 U6337 ( .A1(n5180), .A2(n5652), .ZN(n5907) );
  XNOR2_X1 U6338 ( .A(n5182), .B(n5181), .ZN(n5654) );
  XNOR2_X1 U6339 ( .A(n2990), .B(n5654), .ZN(n5786) );
  INV_X1 U6340 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5183) );
  OAI222_X1 U6341 ( .A1(n5212), .A2(n5907), .B1(n5901), .B2(n5786), .C1(n5183), 
        .C2(n5905), .ZN(U2841) );
  NAND2_X1 U6342 ( .A1(n5184), .A2(n5185), .ZN(n5186) );
  AND2_X1 U6343 ( .A1(n5187), .A2(n5186), .ZN(n5912) );
  INV_X1 U6344 ( .A(n5912), .ZN(n5191) );
  INV_X1 U6345 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5190) );
  NAND2_X1 U6346 ( .A1(n3017), .A2(n5188), .ZN(n5189) );
  NAND2_X1 U6347 ( .A1(n2990), .A2(n5189), .ZN(n5794) );
  OAI222_X1 U6348 ( .A1(n5212), .A2(n5191), .B1(n5905), .B2(n5190), .C1(n5901), 
        .C2(n5794), .ZN(U2842) );
  OAI21_X1 U6349 ( .B1(n5202), .B2(n5193), .A(n5184), .ZN(n5336) );
  INV_X1 U6350 ( .A(n5336), .ZN(n5917) );
  OR2_X1 U6351 ( .A1(n5198), .A2(n5194), .ZN(n5195) );
  NAND2_X1 U6352 ( .A1(n3017), .A2(n5195), .ZN(n5810) );
  OAI22_X1 U6353 ( .A1(n5810), .A2(n5901), .B1(n5806), .B2(n5905), .ZN(n5196)
         );
  AOI21_X1 U6354 ( .B1(n5917), .B2(n6519), .A(n5196), .ZN(n5197) );
  INV_X1 U6355 ( .A(n5197), .ZN(U2843) );
  INV_X1 U6356 ( .A(n5198), .ZN(n5199) );
  OAI21_X1 U6357 ( .B1(n5201), .B2(n5200), .A(n5199), .ZN(n5818) );
  INV_X1 U6358 ( .A(EBX_REG_15__SCAN_IN), .ZN(n6639) );
  INV_X1 U6359 ( .A(n5202), .ZN(n5203) );
  OAI21_X1 U6360 ( .B1(n5117), .B2(n5204), .A(n5203), .ZN(n5813) );
  OAI222_X1 U6361 ( .A1(n5818), .A2(n5901), .B1(n5905), .B2(n6639), .C1(n5212), 
        .C2(n5813), .ZN(U2844) );
  AOI22_X1 U6362 ( .A1(n5492), .A2(n6518), .B1(n6517), .B2(EBX_REG_14__SCAN_IN), .ZN(n5205) );
  OAI21_X1 U6363 ( .B1(n5344), .B2(n5212), .A(n5205), .ZN(U2845) );
  NAND2_X1 U6364 ( .A1(n5207), .A2(n5206), .ZN(n5208) );
  NAND2_X1 U6365 ( .A1(n5209), .A2(n5208), .ZN(n5829) );
  INV_X1 U6366 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6621) );
  OAI21_X1 U6367 ( .B1(n3005), .B2(n3718), .A(n5211), .ZN(n5832) );
  OAI222_X1 U6368 ( .A1(n5829), .A2(n5901), .B1(n5905), .B2(n6621), .C1(n5212), 
        .C2(n5832), .ZN(U2846) );
  INV_X1 U6369 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5213) );
  INV_X1 U6370 ( .A(n5363), .ZN(n5245) );
  OAI222_X1 U6371 ( .A1(n5495), .A2(n5901), .B1(n5905), .B2(n5213), .C1(n5212), 
        .C2(n5245), .ZN(U2847) );
  NAND2_X1 U6372 ( .A1(n3243), .A2(n3320), .ZN(n5214) );
  NOR2_X2 U6373 ( .A1(n5909), .A2(n5214), .ZN(n5915) );
  AOI22_X1 U6374 ( .A1(n5915), .A2(DATAI_14_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n5909), .ZN(n5216) );
  NAND2_X1 U6375 ( .A1(n3004), .A2(DATAI_30_), .ZN(n5215) );
  OAI211_X1 U6376 ( .C1(n5217), .C2(n5666), .A(n5216), .B(n5215), .ZN(U2861)
         );
  AOI22_X1 U6377 ( .A1(n5915), .A2(DATAI_13_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n5909), .ZN(n5219) );
  NAND2_X1 U6378 ( .A1(n3004), .A2(DATAI_29_), .ZN(n5218) );
  OAI211_X1 U6379 ( .C1(n5220), .C2(n5666), .A(n5219), .B(n5218), .ZN(U2862)
         );
  AOI22_X1 U6380 ( .A1(n5915), .A2(DATAI_12_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n5909), .ZN(n5222) );
  NAND2_X1 U6381 ( .A1(n3004), .A2(DATAI_28_), .ZN(n5221) );
  OAI211_X1 U6382 ( .C1(n5223), .C2(n5666), .A(n5222), .B(n5221), .ZN(U2863)
         );
  AOI22_X1 U6383 ( .A1(n5915), .A2(DATAI_11_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n5909), .ZN(n5225) );
  NAND2_X1 U6384 ( .A1(n3004), .A2(DATAI_27_), .ZN(n5224) );
  OAI211_X1 U6385 ( .C1(n5280), .C2(n5666), .A(n5225), .B(n5224), .ZN(U2864)
         );
  AOI22_X1 U6386 ( .A1(n5915), .A2(DATAI_10_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n5909), .ZN(n5227) );
  NAND2_X1 U6387 ( .A1(n3004), .A2(DATAI_26_), .ZN(n5226) );
  OAI211_X1 U6388 ( .C1(n5603), .C2(n5666), .A(n5227), .B(n5226), .ZN(U2865)
         );
  AOI22_X1 U6389 ( .A1(n5915), .A2(DATAI_9_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n5909), .ZN(n5229) );
  NAND2_X1 U6390 ( .A1(n3004), .A2(DATAI_25_), .ZN(n5228) );
  OAI211_X1 U6391 ( .C1(n5674), .C2(n5666), .A(n5229), .B(n5228), .ZN(U2866)
         );
  AOI22_X1 U6392 ( .A1(n5915), .A2(DATAI_8_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n5909), .ZN(n5231) );
  NAND2_X1 U6393 ( .A1(n3004), .A2(DATAI_24_), .ZN(n5230) );
  OAI211_X1 U6394 ( .C1(n5232), .C2(n5666), .A(n5231), .B(n5230), .ZN(U2867)
         );
  AOI22_X1 U6395 ( .A1(n5915), .A2(DATAI_7_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n5909), .ZN(n5234) );
  NAND2_X1 U6396 ( .A1(n3004), .A2(DATAI_23_), .ZN(n5233) );
  OAI211_X1 U6397 ( .C1(n5235), .C2(n5666), .A(n5234), .B(n5233), .ZN(U2868)
         );
  AOI22_X1 U6398 ( .A1(n5915), .A2(DATAI_6_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n5909), .ZN(n5237) );
  NAND2_X1 U6399 ( .A1(n3004), .A2(DATAI_22_), .ZN(n5236) );
  OAI211_X1 U6400 ( .C1(n5623), .C2(n5666), .A(n5237), .B(n5236), .ZN(U2869)
         );
  AOI22_X1 U6401 ( .A1(n5915), .A2(DATAI_4_), .B1(EAX_REG_20__SCAN_IN), .B2(
        n5909), .ZN(n5239) );
  NAND2_X1 U6402 ( .A1(n3004), .A2(DATAI_20_), .ZN(n5238) );
  OAI211_X1 U6403 ( .C1(n5640), .C2(n5666), .A(n5239), .B(n5238), .ZN(U2871)
         );
  AOI22_X1 U6404 ( .A1(n5249), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n5909), .ZN(n5240) );
  OAI21_X1 U6405 ( .B1(n5813), .B2(n5666), .A(n5240), .ZN(U2876) );
  INV_X1 U6406 ( .A(DATAI_14_), .ZN(n6006) );
  INV_X1 U6407 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6626) );
  OAI222_X1 U6408 ( .A1(n5344), .A2(n5666), .B1(n5242), .B2(n6006), .C1(n5241), 
        .C2(n6626), .ZN(U2877) );
  AOI22_X1 U6409 ( .A1(n5249), .A2(DATAI_13_), .B1(EAX_REG_13__SCAN_IN), .B2(
        n5909), .ZN(n5243) );
  OAI21_X1 U6410 ( .B1(n5832), .B2(n5666), .A(n5243), .ZN(U2878) );
  AOI22_X1 U6411 ( .A1(n5249), .A2(DATAI_12_), .B1(EAX_REG_12__SCAN_IN), .B2(
        n5909), .ZN(n5244) );
  OAI21_X1 U6412 ( .B1(n5245), .B2(n5666), .A(n5244), .ZN(U2879) );
  AND2_X1 U6413 ( .A1(n5247), .A2(n5246), .ZN(n5248) );
  OR2_X1 U6414 ( .A1(n5248), .A2(n3015), .ZN(n6014) );
  AOI22_X1 U6415 ( .A1(n5249), .A2(DATAI_11_), .B1(EAX_REG_11__SCAN_IN), .B2(
        n5909), .ZN(n5250) );
  OAI21_X1 U6416 ( .B1(n6014), .B2(n5666), .A(n5250), .ZN(U2880) );
  INV_X1 U6417 ( .A(n5252), .ZN(n5254) );
  OAI21_X1 U6418 ( .B1(n5251), .B2(n5254), .A(n5253), .ZN(n5255) );
  XNOR2_X1 U6419 ( .A(n5255), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5406)
         );
  AND2_X1 U6420 ( .A1(n5705), .A2(REIP_REG_30__SCAN_IN), .ZN(n5398) );
  AOI21_X1 U6421 ( .B1(n6047), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5398), 
        .ZN(n5256) );
  OAI21_X1 U6422 ( .B1(n6040), .B2(n5257), .A(n5256), .ZN(n5258) );
  AOI21_X1 U6423 ( .B1(n5259), .B2(n6035), .A(n5258), .ZN(n5260) );
  OAI21_X1 U6424 ( .B1(n5406), .B2(n6041), .A(n5260), .ZN(U2956) );
  INV_X1 U6425 ( .A(n5261), .ZN(n5262) );
  OAI21_X1 U6426 ( .B1(n5251), .B2(n5263), .A(n5262), .ZN(n5264) );
  XNOR2_X1 U6427 ( .A(n5264), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5415)
         );
  AND2_X1 U6428 ( .A1(n5705), .A2(REIP_REG_29__SCAN_IN), .ZN(n5409) );
  AOI21_X1 U6429 ( .B1(n6047), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5409), 
        .ZN(n5265) );
  OAI21_X1 U6430 ( .B1(n6040), .B2(n5266), .A(n5265), .ZN(n5267) );
  AOI21_X1 U6431 ( .B1(n5268), .B2(n6035), .A(n5267), .ZN(n5269) );
  OAI21_X1 U6432 ( .B1(n5415), .B2(n6041), .A(n5269), .ZN(U2957) );
  NAND3_X1 U6433 ( .A1(n5251), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5686), .ZN(n5271) );
  AOI22_X1 U6434 ( .A1(n5271), .A2(n5277), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5437), .ZN(n5272) );
  XNOR2_X1 U6435 ( .A(n5272), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5425)
         );
  INV_X1 U6436 ( .A(n5588), .ZN(n5274) );
  AND2_X1 U6437 ( .A1(n5705), .A2(REIP_REG_28__SCAN_IN), .ZN(n5421) );
  AOI21_X1 U6438 ( .B1(n6047), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5421), 
        .ZN(n5273) );
  OAI21_X1 U6439 ( .B1(n6040), .B2(n5274), .A(n5273), .ZN(n5275) );
  AOI21_X1 U6440 ( .B1(n5591), .B2(n6035), .A(n5275), .ZN(n5276) );
  OAI21_X1 U6441 ( .B1(n5425), .B2(n6041), .A(n5276), .ZN(U2958) );
  NAND2_X1 U6442 ( .A1(n5278), .A2(n5277), .ZN(n5279) );
  XNOR2_X1 U6443 ( .A(n5279), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5434)
         );
  INV_X1 U6444 ( .A(n5280), .ZN(n5284) );
  AND2_X1 U6445 ( .A1(n5705), .A2(REIP_REG_27__SCAN_IN), .ZN(n5426) );
  AOI21_X1 U6446 ( .B1(n6047), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5426), 
        .ZN(n5281) );
  OAI21_X1 U6447 ( .B1(n6040), .B2(n5282), .A(n5281), .ZN(n5283) );
  AOI21_X1 U6448 ( .B1(n5284), .B2(n6035), .A(n5283), .ZN(n5285) );
  OAI21_X1 U6449 ( .B1(n5434), .B2(n6041), .A(n5285), .ZN(U2959) );
  INV_X1 U6450 ( .A(n5286), .ZN(n5287) );
  NOR2_X1 U6451 ( .A1(n5288), .A2(n5287), .ZN(n5289) );
  XOR2_X1 U6452 ( .A(n5289), .B(n5251), .Z(n5444) );
  INV_X1 U6453 ( .A(n5603), .ZN(n5293) );
  INV_X1 U6454 ( .A(n5597), .ZN(n5291) );
  AND2_X1 U6455 ( .A1(n5705), .A2(REIP_REG_26__SCAN_IN), .ZN(n5439) );
  AOI21_X1 U6456 ( .B1(n6047), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5439), 
        .ZN(n5290) );
  OAI21_X1 U6457 ( .B1(n6040), .B2(n5291), .A(n5290), .ZN(n5292) );
  AOI21_X1 U6458 ( .B1(n5293), .B2(n6035), .A(n5292), .ZN(n5294) );
  OAI21_X1 U6459 ( .B1(n5444), .B2(n6041), .A(n5294), .ZN(U2960) );
  NAND4_X1 U6460 ( .A1(n5296), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .A3(n5297), .A4(n5686), .ZN(n5298) );
  NAND2_X1 U6461 ( .A1(n5295), .A2(n5298), .ZN(n5299) );
  XNOR2_X1 U6462 ( .A(n5299), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5458)
         );
  NAND2_X1 U6463 ( .A1(n5705), .A2(REIP_REG_23__SCAN_IN), .ZN(n5453) );
  NAND2_X1 U6464 ( .A1(n6047), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5300)
         );
  OAI211_X1 U6465 ( .C1(n6040), .C2(n5610), .A(n5453), .B(n5300), .ZN(n5301)
         );
  AOI21_X1 U6466 ( .B1(n5614), .B2(n6035), .A(n5301), .ZN(n5302) );
  OAI21_X1 U6467 ( .B1(n5458), .B2(n6041), .A(n5302), .ZN(U2963) );
  AOI21_X1 U6468 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5686), .A(n5304), 
        .ZN(n5305) );
  XNOR2_X1 U6469 ( .A(n5303), .B(n5305), .ZN(n5467) );
  INV_X1 U6470 ( .A(n6047), .ZN(n5393) );
  NAND2_X1 U6471 ( .A1(n5705), .A2(REIP_REG_22__SCAN_IN), .ZN(n5462) );
  OAI21_X1 U6472 ( .B1(n5393), .B2(n6634), .A(n5462), .ZN(n5307) );
  NOR2_X1 U6473 ( .A1(n5623), .A2(n6043), .ZN(n5306) );
  AOI211_X1 U6474 ( .C1(n5395), .C2(n5621), .A(n5307), .B(n5306), .ZN(n5308)
         );
  OAI21_X1 U6475 ( .B1(n5467), .B2(n6041), .A(n5308), .ZN(U2964) );
  NAND2_X1 U6476 ( .A1(n5310), .A2(n5309), .ZN(n5311) );
  NAND2_X1 U6477 ( .A1(n5312), .A2(n5311), .ZN(n5665) );
  OAI21_X1 U6478 ( .B1(n5313), .B2(n2987), .A(n4086), .ZN(n5468) );
  NAND2_X1 U6479 ( .A1(n5468), .A2(n6036), .ZN(n5317) );
  NAND2_X1 U6480 ( .A1(n6112), .A2(REIP_REG_21__SCAN_IN), .ZN(n5474) );
  OAI21_X1 U6481 ( .B1(n5393), .B2(n6664), .A(n5474), .ZN(n5314) );
  AOI21_X1 U6482 ( .B1(n5315), .B2(n5395), .A(n5314), .ZN(n5316) );
  OAI211_X1 U6483 ( .C1(n6043), .C2(n5665), .A(n5317), .B(n5316), .ZN(U2965)
         );
  XNOR2_X1 U6484 ( .A(n5686), .B(n5318), .ZN(n5319) );
  XNOR2_X1 U6485 ( .A(n5296), .B(n5319), .ZN(n5699) );
  NAND2_X1 U6486 ( .A1(n5699), .A2(n6036), .ZN(n5322) );
  OAI22_X1 U6487 ( .A1(n5393), .A2(n5646), .B1(n6071), .B2(n6458), .ZN(n5320)
         );
  AOI21_X1 U6488 ( .B1(n5395), .B2(n5638), .A(n5320), .ZN(n5321) );
  OAI211_X1 U6489 ( .C1(n6043), .C2(n5640), .A(n5322), .B(n5321), .ZN(U2966)
         );
  NAND3_X1 U6490 ( .A1(n5686), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5325) );
  NAND4_X1 U6491 ( .A1(n5323), .A2(n5508), .A3(n5726), .A4(n6557), .ZN(n5324)
         );
  OAI21_X1 U6492 ( .B1(n5323), .B2(n5325), .A(n5324), .ZN(n5326) );
  XNOR2_X1 U6493 ( .A(n5326), .B(n3504), .ZN(n5716) );
  NAND2_X1 U6494 ( .A1(n5716), .A2(n6036), .ZN(n5330) );
  NAND2_X1 U6495 ( .A1(n6112), .A2(REIP_REG_18__SCAN_IN), .ZN(n5712) );
  OAI21_X1 U6496 ( .B1(n5393), .B2(n5327), .A(n5712), .ZN(n5328) );
  AOI21_X1 U6497 ( .B1(n5395), .B2(n5783), .A(n5328), .ZN(n5329) );
  OAI211_X1 U6498 ( .C1(n6043), .C2(n5907), .A(n5330), .B(n5329), .ZN(U2968)
         );
  XNOR2_X1 U6499 ( .A(n5686), .B(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5331)
         );
  XNOR2_X1 U6500 ( .A(n5323), .B(n5331), .ZN(n5735) );
  NAND2_X1 U6501 ( .A1(n5735), .A2(n6036), .ZN(n5335) );
  OAI22_X1 U6502 ( .A1(n5393), .A2(n5332), .B1(n6071), .B2(n6452), .ZN(n5333)
         );
  AOI21_X1 U6503 ( .B1(n5804), .B2(n5395), .A(n5333), .ZN(n5334) );
  OAI211_X1 U6504 ( .C1(n6043), .C2(n5336), .A(n5335), .B(n5334), .ZN(U2970)
         );
  XNOR2_X1 U6505 ( .A(n5686), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5337)
         );
  XNOR2_X1 U6506 ( .A(n3001), .B(n5337), .ZN(n5740) );
  AOI22_X1 U6507 ( .A1(n6047), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n5705), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U6508 ( .A1(n5395), .A2(n5815), .ZN(n5338) );
  OAI211_X1 U6509 ( .C1(n5813), .C2(n6043), .A(n5339), .B(n5338), .ZN(n5340)
         );
  AOI21_X1 U6510 ( .B1(n5740), .B2(n6036), .A(n5340), .ZN(n5341) );
  INV_X1 U6511 ( .A(n5341), .ZN(U2971) );
  XNOR2_X1 U6512 ( .A(n5686), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5342)
         );
  XNOR2_X1 U6513 ( .A(n5343), .B(n5342), .ZN(n5494) );
  INV_X1 U6514 ( .A(n5344), .ZN(n5349) );
  INV_X1 U6515 ( .A(n5345), .ZN(n5347) );
  NOR2_X1 U6516 ( .A1(n6071), .A2(n6449), .ZN(n5491) );
  AOI21_X1 U6517 ( .B1(n6047), .B2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n5491), 
        .ZN(n5346) );
  OAI21_X1 U6518 ( .B1(n6040), .B2(n5347), .A(n5346), .ZN(n5348) );
  AOI21_X1 U6519 ( .B1(n5349), .B2(n6035), .A(n5348), .ZN(n5350) );
  OAI21_X1 U6520 ( .B1(n5494), .B2(n6041), .A(n5350), .ZN(U2972) );
  XNOR2_X1 U6521 ( .A(n5352), .B(n5351), .ZN(n5747) );
  NAND2_X1 U6522 ( .A1(n5747), .A2(n6036), .ZN(n5356) );
  NOR2_X1 U6523 ( .A1(n6071), .A2(n6607), .ZN(n5744) );
  NOR2_X1 U6524 ( .A1(n6040), .A2(n5353), .ZN(n5354) );
  AOI211_X1 U6525 ( .C1(n6047), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5744), 
        .B(n5354), .ZN(n5355) );
  OAI211_X1 U6526 ( .C1(n6043), .C2(n5832), .A(n5356), .B(n5355), .ZN(U2973)
         );
  NOR2_X1 U6527 ( .A1(n5357), .A2(n3008), .ZN(n5358) );
  XNOR2_X1 U6528 ( .A(n5359), .B(n5358), .ZN(n5505) );
  AND2_X1 U6529 ( .A1(n5705), .A2(REIP_REG_12__SCAN_IN), .ZN(n5502) );
  AOI21_X1 U6530 ( .B1(n6047), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n5502), 
        .ZN(n5360) );
  OAI21_X1 U6531 ( .B1(n6040), .B2(n5361), .A(n5360), .ZN(n5362) );
  AOI21_X1 U6532 ( .B1(n5363), .B2(n6035), .A(n5362), .ZN(n5364) );
  OAI21_X1 U6533 ( .B1(n5505), .B2(n6041), .A(n5364), .ZN(U2974) );
  XNOR2_X1 U6534 ( .A(n5686), .B(n5365), .ZN(n5366) );
  XNOR2_X1 U6535 ( .A(n5507), .B(n5366), .ZN(n6060) );
  NAND2_X1 U6536 ( .A1(n6060), .A2(n6036), .ZN(n5371) );
  INV_X1 U6537 ( .A(REIP_REG_10__SCAN_IN), .ZN(n5367) );
  NOR2_X1 U6538 ( .A1(n6071), .A2(n5367), .ZN(n6051) );
  NOR2_X1 U6539 ( .A1(n6040), .A2(n5368), .ZN(n5369) );
  AOI211_X1 U6540 ( .C1(n6047), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6051), 
        .B(n5369), .ZN(n5370) );
  OAI211_X1 U6541 ( .C1(n6043), .C2(n5372), .A(n5371), .B(n5370), .ZN(U2976)
         );
  NOR2_X1 U6542 ( .A1(n5375), .A2(n3010), .ZN(n5376) );
  XNOR2_X1 U6543 ( .A(n5374), .B(n5376), .ZN(n6067) );
  NAND2_X1 U6544 ( .A1(n6067), .A2(n6036), .ZN(n5380) );
  NOR2_X1 U6545 ( .A1(n6071), .A2(n6442), .ZN(n6064) );
  NOR2_X1 U6546 ( .A1(n6040), .A2(n5377), .ZN(n5378) );
  AOI211_X1 U6547 ( .C1(n6047), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6064), 
        .B(n5378), .ZN(n5379) );
  OAI211_X1 U6548 ( .C1(n6043), .C2(n5849), .A(n5380), .B(n5379), .ZN(U2977)
         );
  AOI21_X1 U6549 ( .B1(n5382), .B2(n3009), .A(n5381), .ZN(n6074) );
  INV_X1 U6550 ( .A(n6074), .ZN(n5389) );
  INV_X1 U6551 ( .A(n5383), .ZN(n5387) );
  AOI22_X1 U6552 ( .A1(n6047), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n5705), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n5384) );
  OAI21_X1 U6553 ( .B1(n6040), .B2(n5385), .A(n5384), .ZN(n5386) );
  AOI21_X1 U6554 ( .B1(n5387), .B2(n6035), .A(n5386), .ZN(n5388) );
  OAI21_X1 U6555 ( .B1(n5389), .B2(n6041), .A(n5388), .ZN(U2978) );
  AOI21_X1 U6556 ( .B1(n5392), .B2(n5391), .A(n5390), .ZN(n6083) );
  NAND2_X1 U6557 ( .A1(n6083), .A2(n6036), .ZN(n5397) );
  INV_X1 U6558 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5860) );
  NAND2_X1 U6559 ( .A1(n6112), .A2(REIP_REG_7__SCAN_IN), .ZN(n6079) );
  OAI21_X1 U6560 ( .B1(n5393), .B2(n5860), .A(n6079), .ZN(n5394) );
  AOI21_X1 U6561 ( .B1(n5857), .B2(n5395), .A(n5394), .ZN(n5396) );
  OAI211_X1 U6562 ( .C1(n5862), .C2(n6043), .A(n5397), .B(n5396), .ZN(U2979)
         );
  AOI21_X1 U6563 ( .B1(n5400), .B2(n5399), .A(n5398), .ZN(n5401) );
  OAI21_X1 U6564 ( .B1(n5402), .B2(n6116), .A(n5401), .ZN(n5403) );
  AOI21_X1 U6565 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n5404), .A(n5403), 
        .ZN(n5405) );
  OAI21_X1 U6566 ( .B1(n5406), .B2(n5519), .A(n5405), .ZN(U2988) );
  INV_X1 U6567 ( .A(n5407), .ZN(n5410) );
  NOR3_X1 U6568 ( .A1(n5428), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5417), 
        .ZN(n5408) );
  AOI211_X1 U6569 ( .C1(n5410), .C2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5409), .B(n5408), .ZN(n5414) );
  INV_X1 U6570 ( .A(n5411), .ZN(n5412) );
  NAND2_X1 U6571 ( .A1(n5412), .A2(n6100), .ZN(n5413) );
  OAI211_X1 U6572 ( .C1(n5415), .C2(n5519), .A(n5414), .B(n5413), .ZN(U2989)
         );
  INV_X1 U6573 ( .A(n5416), .ZN(n5419) );
  INV_X1 U6574 ( .A(n5417), .ZN(n5418) );
  NOR3_X1 U6575 ( .A1(n5428), .A2(n5419), .A3(n5418), .ZN(n5420) );
  AOI211_X1 U6576 ( .C1(n5422), .C2(n6100), .A(n5421), .B(n5420), .ZN(n5424)
         );
  NAND2_X1 U6577 ( .A1(n5431), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5423) );
  OAI211_X1 U6578 ( .C1(n5425), .C2(n5519), .A(n5424), .B(n5423), .ZN(U2990)
         );
  INV_X1 U6579 ( .A(n5426), .ZN(n5427) );
  OAI21_X1 U6580 ( .B1(n5428), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5427), 
        .ZN(n5429) );
  AOI21_X1 U6581 ( .B1(n5430), .B2(n6100), .A(n5429), .ZN(n5433) );
  NAND2_X1 U6582 ( .A1(n5431), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5432) );
  OAI211_X1 U6583 ( .C1(n5434), .C2(n5519), .A(n5433), .B(n5432), .ZN(U2991)
         );
  INV_X1 U6584 ( .A(n5602), .ZN(n5440) );
  AOI211_X1 U6585 ( .C1(n5694), .C2(n5437), .A(n5436), .B(n5435), .ZN(n5438)
         );
  AOI211_X1 U6586 ( .C1(n5440), .C2(n6100), .A(n5439), .B(n5438), .ZN(n5443)
         );
  INV_X1 U6587 ( .A(n5695), .ZN(n5441) );
  NAND2_X1 U6588 ( .A1(n5441), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5442) );
  OAI211_X1 U6589 ( .C1(n5444), .C2(n5519), .A(n5443), .B(n5442), .ZN(U2992)
         );
  NAND2_X1 U6590 ( .A1(n5445), .A2(n6119), .ZN(n5452) );
  INV_X1 U6591 ( .A(n5455), .ZN(n5446) );
  AOI21_X1 U6592 ( .B1(n5446), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5447) );
  NOR2_X1 U6593 ( .A1(n5695), .A2(n5447), .ZN(n5448) );
  AOI211_X1 U6594 ( .C1(n6100), .C2(n5450), .A(n5449), .B(n5448), .ZN(n5451)
         );
  NAND2_X1 U6595 ( .A1(n5452), .A2(n5451), .ZN(U2994) );
  NAND2_X1 U6596 ( .A1(n5613), .A2(n6100), .ZN(n5454) );
  OAI211_X1 U6597 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n5455), .A(n5454), .B(n5453), .ZN(n5456) );
  AOI21_X1 U6598 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5465), .A(n5456), 
        .ZN(n5457) );
  OAI21_X1 U6599 ( .B1(n5458), .B2(n5519), .A(n5457), .ZN(U2995) );
  OAI21_X1 U6600 ( .B1(n5461), .B2(n5460), .A(n5459), .ZN(n5464) );
  OAI21_X1 U6601 ( .B1(n5622), .B2(n6116), .A(n5462), .ZN(n5463) );
  AOI21_X1 U6602 ( .B1(n5465), .B2(n5464), .A(n5463), .ZN(n5466) );
  OAI21_X1 U6603 ( .B1(n5467), .B2(n5519), .A(n5466), .ZN(U2996) );
  INV_X1 U6604 ( .A(n5468), .ZN(n5478) );
  OR2_X1 U6605 ( .A1(n5470), .A2(n5469), .ZN(n5471) );
  NAND2_X1 U6606 ( .A1(n5472), .A2(n5471), .ZN(n5660) );
  OAI211_X1 U6607 ( .C1(n5660), .C2(n6116), .A(n5474), .B(n5473), .ZN(n5475)
         );
  AOI21_X1 U6608 ( .B1(n5476), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5475), 
        .ZN(n5477) );
  OAI21_X1 U6609 ( .B1(n5478), .B2(n5519), .A(n5477), .ZN(U2997) );
  INV_X1 U6610 ( .A(n5511), .ZN(n5751) );
  NOR2_X1 U6611 ( .A1(n5751), .A2(n5483), .ZN(n5489) );
  NAND3_X1 U6612 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n3502), .ZN(n5750) );
  AOI21_X1 U6613 ( .B1(n5480), .B2(n5479), .A(n5750), .ZN(n5487) );
  NAND2_X1 U6614 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5481) );
  AOI22_X1 U6615 ( .A1(n5484), .A2(n5483), .B1(n5482), .B2(n5481), .ZN(n5485)
         );
  NAND2_X1 U6616 ( .A1(n5486), .A2(n5485), .ZN(n5746) );
  OR2_X1 U6617 ( .A1(n5487), .A2(n5746), .ZN(n5488) );
  MUX2_X1 U6618 ( .A(n5489), .B(n5488), .S(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .Z(n5490) );
  AOI211_X1 U6619 ( .C1(n6100), .C2(n5492), .A(n5491), .B(n5490), .ZN(n5493)
         );
  OAI21_X1 U6620 ( .B1(n5494), .B2(n5519), .A(n5493), .ZN(U3004) );
  INV_X1 U6621 ( .A(n5495), .ZN(n5503) );
  NOR2_X1 U6622 ( .A1(n5751), .A2(n3098), .ZN(n5500) );
  NAND2_X1 U6623 ( .A1(n6088), .A2(n5496), .ZN(n5697) );
  OAI22_X1 U6624 ( .A1(n3098), .A2(n5728), .B1(n5497), .B2(n5697), .ZN(n5498)
         );
  INV_X1 U6625 ( .A(n5498), .ZN(n5499) );
  MUX2_X1 U6626 ( .A(n5500), .B(n5499), .S(INSTADDRPOINTER_REG_12__SCAN_IN), 
        .Z(n5501) );
  AOI211_X1 U6627 ( .C1(n6100), .C2(n5503), .A(n5502), .B(n5501), .ZN(n5504)
         );
  OAI21_X1 U6628 ( .B1(n5505), .B2(n5519), .A(n5504), .ZN(U3006) );
  AOI22_X1 U6629 ( .A1(n5507), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .B1(n5508), .B2(n5506), .ZN(n5510) );
  XNOR2_X1 U6630 ( .A(n5508), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5509)
         );
  XNOR2_X1 U6631 ( .A(n5510), .B(n5509), .ZN(n6018) );
  AOI22_X1 U6632 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n5728), .B1(n5511), .B2(n3098), .ZN(n5518) );
  AOI21_X1 U6633 ( .B1(n5514), .B2(n5513), .A(n5512), .ZN(n5515) );
  OR2_X1 U6634 ( .A1(n5516), .A2(n5515), .ZN(n5900) );
  INV_X1 U6635 ( .A(n5900), .ZN(n5844) );
  AOI22_X1 U6636 ( .A1(n5844), .A2(n6100), .B1(n6112), .B2(
        REIP_REG_11__SCAN_IN), .ZN(n5517) );
  OAI211_X1 U6637 ( .C1(n6018), .C2(n5519), .A(n5518), .B(n5517), .ZN(U3007)
         );
  OAI211_X1 U6638 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n5521), .A(n5520), .B(
        n6245), .ZN(n5522) );
  OAI21_X1 U6639 ( .B1(n5525), .B2(n5523), .A(n5522), .ZN(n5524) );
  MUX2_X1 U6640 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5524), .S(n6124), 
        .Z(U3464) );
  XNOR2_X1 U6641 ( .A(n3566), .B(n6204), .ZN(n5527) );
  OAI22_X1 U6642 ( .A1(n5527), .A2(n6295), .B1(n5526), .B2(n5525), .ZN(n5528)
         );
  MUX2_X1 U6643 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5528), .S(n6124), 
        .Z(U3463) );
  OAI22_X1 U6644 ( .A1(n5530), .A2(n6494), .B1(n6395), .B2(n5529), .ZN(n5532)
         );
  MUX2_X1 U6645 ( .A(n5532), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n5531), 
        .Z(U3456) );
  NOR2_X1 U6646 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5533), .ZN(n5567)
         );
  INV_X1 U6647 ( .A(n5567), .ZN(n5577) );
  INV_X1 U6648 ( .A(n6137), .ZN(n5534) );
  OAI21_X1 U6649 ( .B1(n5573), .B2(n5534), .A(n6248), .ZN(n5535) );
  NAND2_X1 U6650 ( .A1(n5535), .A2(n5538), .ZN(n5537) );
  OAI221_X1 U6651 ( .B1(n5567), .B2(n6487), .C1(n5567), .C2(n5537), .A(n5536), 
        .ZN(n5570) );
  NAND2_X1 U6652 ( .A1(n5570), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5543) );
  OR2_X1 U6653 ( .A1(n5538), .A2(n6295), .ZN(n5540) );
  NAND3_X1 U6654 ( .A1(n6147), .A2(n6140), .A3(n6201), .ZN(n5539) );
  OAI22_X1 U6655 ( .A1(n6137), .A2(n6156), .B1(n5571), .B2(n6301), .ZN(n5541)
         );
  AOI21_X1 U6656 ( .B1(n6153), .B2(n5573), .A(n5541), .ZN(n5542) );
  OAI211_X1 U6657 ( .C1(n5544), .C2(n5577), .A(n5543), .B(n5542), .ZN(U3036)
         );
  NAND2_X1 U6658 ( .A1(n5570), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5547) );
  OAI22_X1 U6659 ( .A1(n6137), .A2(n6160), .B1(n5571), .B2(n6308), .ZN(n5545)
         );
  AOI21_X1 U6660 ( .B1(n6157), .B2(n5573), .A(n5545), .ZN(n5546) );
  OAI211_X1 U6661 ( .C1(n5577), .C2(n5548), .A(n5547), .B(n5546), .ZN(U3037)
         );
  NAND2_X1 U6662 ( .A1(n5570), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5551) );
  OAI22_X1 U6663 ( .A1(n6137), .A2(n6164), .B1(n5571), .B2(n6315), .ZN(n5549)
         );
  AOI21_X1 U6664 ( .B1(n6161), .B2(n5573), .A(n5549), .ZN(n5550) );
  OAI211_X1 U6665 ( .C1(n5577), .C2(n5552), .A(n5551), .B(n5550), .ZN(U3038)
         );
  NAND2_X1 U6666 ( .A1(n5570), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5555) );
  OAI22_X1 U6667 ( .A1(n6137), .A2(n6223), .B1(n5571), .B2(n6323), .ZN(n5553)
         );
  AOI21_X1 U6668 ( .B1(n6220), .B2(n5573), .A(n5553), .ZN(n5554) );
  OAI211_X1 U6669 ( .C1(n5577), .C2(n5556), .A(n5555), .B(n5554), .ZN(U3039)
         );
  NAND2_X1 U6670 ( .A1(n5570), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5559) );
  OAI22_X1 U6671 ( .A1(n6137), .A2(n6332), .B1(n5571), .B2(n6331), .ZN(n5557)
         );
  AOI21_X1 U6672 ( .B1(n6329), .B2(n5573), .A(n5557), .ZN(n5558) );
  OAI211_X1 U6673 ( .C1(n5577), .C2(n5560), .A(n5559), .B(n5558), .ZN(U3040)
         );
  NAND2_X1 U6674 ( .A1(n5570), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5563) );
  OAI22_X1 U6675 ( .A1(n6137), .A2(n6340), .B1(n5571), .B2(n6339), .ZN(n5561)
         );
  AOI21_X1 U6676 ( .B1(n6337), .B2(n5573), .A(n5561), .ZN(n5562) );
  OAI211_X1 U6677 ( .C1(n5577), .C2(n5564), .A(n5563), .B(n5562), .ZN(U3041)
         );
  NAND2_X1 U6678 ( .A1(n5570), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5569) );
  OAI22_X1 U6679 ( .A1(n5565), .A2(n6277), .B1(n6173), .B2(n6137), .ZN(n5566)
         );
  AOI21_X1 U6680 ( .B1(n6347), .B2(n5567), .A(n5566), .ZN(n5568) );
  OAI211_X1 U6681 ( .C1(n5571), .C2(n5585), .A(n5569), .B(n5568), .ZN(U3042)
         );
  NAND2_X1 U6682 ( .A1(n5570), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5575) );
  OAI22_X1 U6683 ( .A1(n6137), .A2(n6181), .B1(n5571), .B2(n6358), .ZN(n5572)
         );
  AOI21_X1 U6684 ( .B1(n6177), .B2(n5573), .A(n5572), .ZN(n5574) );
  OAI211_X1 U6685 ( .C1(n5577), .C2(n5576), .A(n5575), .B(n5574), .ZN(U3043)
         );
  INV_X1 U6686 ( .A(n5578), .ZN(n5579) );
  NAND2_X1 U6687 ( .A1(n5579), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5584) );
  OAI22_X1 U6688 ( .A1(n5580), .A2(n6173), .B1(n6277), .B2(n6126), .ZN(n5581)
         );
  AOI21_X1 U6689 ( .B1(n6347), .B2(n5582), .A(n5581), .ZN(n5583) );
  OAI211_X1 U6690 ( .C1(n5586), .C2(n5585), .A(n5584), .B(n5583), .ZN(U3058)
         );
  AND2_X1 U6691 ( .A1(n5934), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI22_X1 U6692 ( .A1(EBX_REG_28__SCAN_IN), .A2(n5865), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n5876), .ZN(n5596) );
  AOI22_X1 U6693 ( .A1(n5588), .A2(n5870), .B1(REIP_REG_28__SCAN_IN), .B2(
        n5587), .ZN(n5595) );
  NOR2_X1 U6694 ( .A1(n5589), .A2(n5873), .ZN(n5590) );
  AOI21_X1 U6695 ( .B1(n5591), .B2(n5880), .A(n5590), .ZN(n5594) );
  NAND3_X1 U6696 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5592), .A3(n6470), .ZN(
        n5593) );
  NAND4_X1 U6697 ( .A1(n5596), .A2(n5595), .A3(n5594), .A4(n5593), .ZN(U2799)
         );
  AOI22_X1 U6698 ( .A1(EBX_REG_26__SCAN_IN), .A2(n5865), .B1(n5597), .B2(n5870), .ZN(n5608) );
  INV_X1 U6699 ( .A(n5598), .ZN(n5606) );
  INV_X1 U6700 ( .A(REIP_REG_26__SCAN_IN), .ZN(n5599) );
  OAI21_X1 U6701 ( .B1(n5601), .B2(n5600), .A(n5599), .ZN(n5605) );
  OAI22_X1 U6702 ( .A1(n5603), .A2(n5861), .B1(n5602), .B2(n5873), .ZN(n5604)
         );
  AOI21_X1 U6703 ( .B1(n5606), .B2(n5605), .A(n5604), .ZN(n5607) );
  OAI211_X1 U6704 ( .C1(n6668), .C2(n5890), .A(n5608), .B(n5607), .ZN(U2801)
         );
  NOR2_X1 U6705 ( .A1(REIP_REG_23__SCAN_IN), .A2(n5609), .ZN(n5618) );
  INV_X1 U6706 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5611) );
  OAI22_X1 U6707 ( .A1(n5611), .A2(n5890), .B1(n5610), .B2(n5889), .ZN(n5612)
         );
  AOI21_X1 U6708 ( .B1(EBX_REG_23__SCAN_IN), .B2(n5865), .A(n5612), .ZN(n5616)
         );
  AOI22_X1 U6709 ( .A1(n5614), .A2(n5880), .B1(n5613), .B2(n5886), .ZN(n5615)
         );
  OAI211_X1 U6710 ( .C1(n5618), .C2(n5617), .A(n5616), .B(n5615), .ZN(U2804)
         );
  AOI22_X1 U6711 ( .A1(EBX_REG_22__SCAN_IN), .A2(n5865), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n5876), .ZN(n5630) );
  NOR2_X1 U6712 ( .A1(n5620), .A2(n5619), .ZN(n5643) );
  AOI22_X1 U6713 ( .A1(n5621), .A2(n5870), .B1(REIP_REG_22__SCAN_IN), .B2(
        n5643), .ZN(n5629) );
  OAI22_X1 U6714 ( .A1(n5623), .A2(n5861), .B1(n5622), .B2(n5873), .ZN(n5624)
         );
  INV_X1 U6715 ( .A(n5624), .ZN(n5628) );
  INV_X1 U6716 ( .A(n5637), .ZN(n5626) );
  OAI211_X1 U6717 ( .C1(REIP_REG_22__SCAN_IN), .C2(REIP_REG_21__SCAN_IN), .A(
        n5626), .B(n5625), .ZN(n5627) );
  NAND4_X1 U6718 ( .A1(n5630), .A2(n5629), .A3(n5628), .A4(n5627), .ZN(U2805)
         );
  AOI22_X1 U6719 ( .A1(EBX_REG_21__SCAN_IN), .A2(n5865), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n5876), .ZN(n5631) );
  OAI21_X1 U6720 ( .B1(n5632), .B2(n5889), .A(n5631), .ZN(n5633) );
  AOI21_X1 U6721 ( .B1(REIP_REG_21__SCAN_IN), .B2(n5643), .A(n5633), .ZN(n5636) );
  OAI22_X1 U6722 ( .A1(n5665), .A2(n5861), .B1(n5660), .B2(n5873), .ZN(n5634)
         );
  INV_X1 U6723 ( .A(n5634), .ZN(n5635) );
  OAI211_X1 U6724 ( .C1(REIP_REG_21__SCAN_IN), .C2(n5637), .A(n5636), .B(n5635), .ZN(U2806) );
  AOI22_X1 U6725 ( .A1(EBX_REG_20__SCAN_IN), .A2(n5865), .B1(n5638), .B2(n5870), .ZN(n5645) );
  OAI22_X1 U6726 ( .A1(n5640), .A2(n5861), .B1(n5639), .B2(n5873), .ZN(n5641)
         );
  AOI221_X1 U6727 ( .B1(REIP_REG_20__SCAN_IN), .B2(n5643), .C1(n5642), .C2(
        n5643), .A(n5641), .ZN(n5644) );
  OAI211_X1 U6728 ( .C1(n5646), .C2(n5890), .A(n5645), .B(n5644), .ZN(U2807)
         );
  OAI21_X1 U6729 ( .B1(REIP_REG_19__SCAN_IN), .B2(REIP_REG_18__SCAN_IN), .A(
        n5647), .ZN(n5659) );
  AND2_X1 U6730 ( .A1(n5887), .A2(n5648), .ZN(n5796) );
  INV_X1 U6731 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n6602) );
  OAI21_X1 U6732 ( .B1(n5890), .B2(n6602), .A(n5858), .ZN(n5650) );
  OAI22_X1 U6733 ( .A1(n5664), .A2(n5894), .B1(n5684), .B2(n5889), .ZN(n5649)
         );
  AOI211_X1 U6734 ( .C1(REIP_REG_19__SCAN_IN), .C2(n5796), .A(n5650), .B(n5649), .ZN(n5658) );
  OR2_X1 U6735 ( .A1(n5652), .A2(n5651), .ZN(n5653) );
  AND2_X1 U6736 ( .A1(n5175), .A2(n5653), .ZN(n5681) );
  NOR2_X1 U6737 ( .A1(n2990), .A2(n5654), .ZN(n5656) );
  XNOR2_X1 U6738 ( .A(n5656), .B(n5655), .ZN(n5706) );
  AOI22_X1 U6739 ( .A1(n5681), .A2(n5880), .B1(n5886), .B2(n5706), .ZN(n5657)
         );
  OAI211_X1 U6740 ( .C1(n5790), .C2(n5659), .A(n5658), .B(n5657), .ZN(U2808)
         );
  INV_X1 U6741 ( .A(EBX_REG_21__SCAN_IN), .ZN(n6553) );
  OAI22_X1 U6742 ( .A1(n5665), .A2(n5902), .B1(n5660), .B2(n5901), .ZN(n5661)
         );
  INV_X1 U6743 ( .A(n5661), .ZN(n5662) );
  OAI21_X1 U6744 ( .B1(n6553), .B2(n5905), .A(n5662), .ZN(U2838) );
  AOI22_X1 U6745 ( .A1(n5681), .A2(n6519), .B1(n6518), .B2(n5706), .ZN(n5663)
         );
  OAI21_X1 U6746 ( .B1(n5664), .B2(n5905), .A(n5663), .ZN(U2840) );
  INV_X1 U6747 ( .A(n5665), .ZN(n5667) );
  INV_X1 U6748 ( .A(n5666), .ZN(n5916) );
  AOI22_X1 U6749 ( .A1(n5667), .A2(n5916), .B1(n5915), .B2(DATAI_5_), .ZN(
        n5669) );
  AOI22_X1 U6750 ( .A1(EAX_REG_21__SCAN_IN), .A2(n5909), .B1(n3004), .B2(
        DATAI_21_), .ZN(n5668) );
  NAND2_X1 U6751 ( .A1(n5669), .A2(n5668), .ZN(U2870) );
  AOI22_X1 U6752 ( .A1(n5681), .A2(n5916), .B1(n5915), .B2(DATAI_3_), .ZN(
        n5671) );
  AOI22_X1 U6753 ( .A1(EAX_REG_19__SCAN_IN), .A2(n5909), .B1(n3004), .B2(
        DATAI_19_), .ZN(n5670) );
  NAND2_X1 U6754 ( .A1(n5671), .A2(n5670), .ZN(U2872) );
  AOI22_X1 U6755 ( .A1(n6112), .A2(REIP_REG_25__SCAN_IN), .B1(n6047), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5676) );
  OAI21_X1 U6756 ( .B1(n5673), .B2(n5672), .A(n3514), .ZN(n5691) );
  AOI22_X1 U6757 ( .A1(n5691), .A2(n6036), .B1(n6035), .B2(n6520), .ZN(n5675)
         );
  OAI211_X1 U6758 ( .C1(n6040), .C2(n5677), .A(n5676), .B(n5675), .ZN(U2961)
         );
  AOI22_X1 U6759 ( .A1(n6112), .A2(REIP_REG_19__SCAN_IN), .B1(n6047), .B2(
        PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5683) );
  XNOR2_X1 U6760 ( .A(n5686), .B(n5678), .ZN(n5679) );
  XNOR2_X1 U6761 ( .A(n5680), .B(n5679), .ZN(n5708) );
  AOI22_X1 U6762 ( .A1(n5708), .A2(n6036), .B1(n6035), .B2(n5681), .ZN(n5682)
         );
  OAI211_X1 U6763 ( .C1(n6040), .C2(n5684), .A(n5683), .B(n5682), .ZN(U2967)
         );
  AOI22_X1 U6764 ( .A1(n6112), .A2(REIP_REG_17__SCAN_IN), .B1(n6047), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5689) );
  MUX2_X1 U6765 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .B(n5508), .S(n5323), 
        .Z(n5685) );
  OAI21_X1 U6766 ( .B1(n6557), .B2(n5686), .A(n5685), .ZN(n5687) );
  XNOR2_X1 U6767 ( .A(n5687), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5723)
         );
  AOI22_X1 U6768 ( .A1(n5723), .A2(n6036), .B1(n6035), .B2(n5912), .ZN(n5688)
         );
  OAI211_X1 U6769 ( .C1(n6040), .C2(n5791), .A(n5689), .B(n5688), .ZN(U2969)
         );
  AOI22_X1 U6770 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6112), .B1(n5690), .B2(
        n5694), .ZN(n5693) );
  AOI22_X1 U6771 ( .A1(n5691), .A2(n6119), .B1(n6100), .B2(n3006), .ZN(n5692)
         );
  OAI211_X1 U6772 ( .C1(n5695), .C2(n5694), .A(n5693), .B(n5692), .ZN(U2993)
         );
  INV_X1 U6773 ( .A(n5727), .ZN(n5696) );
  AOI21_X1 U6774 ( .B1(n5726), .B2(n5697), .A(n5696), .ZN(n5719) );
  OAI21_X1 U6775 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n6059), .A(n5719), 
        .ZN(n5707) );
  AOI22_X1 U6776 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n5707), .B1(n6112), .B2(REIP_REG_20__SCAN_IN), .ZN(n5704) );
  AOI22_X1 U6777 ( .A1(n5699), .A2(n6119), .B1(n6100), .B2(n5698), .ZN(n5703)
         );
  INV_X1 U6778 ( .A(n5711), .ZN(n5701) );
  OAI211_X1 U6779 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .A(n5701), .B(n5700), .ZN(n5702) );
  NAND3_X1 U6780 ( .A1(n5704), .A2(n5703), .A3(n5702), .ZN(U2998) );
  AOI22_X1 U6781 ( .A1(n5706), .A2(n6100), .B1(n5705), .B2(
        REIP_REG_19__SCAN_IN), .ZN(n5710) );
  AOI22_X1 U6782 ( .A1(n5708), .A2(n6119), .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n5707), .ZN(n5709) );
  OAI211_X1 U6783 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n5711), .A(n5710), .B(n5709), .ZN(U2999) );
  INV_X1 U6784 ( .A(n5786), .ZN(n5714) );
  INV_X1 U6785 ( .A(n5712), .ZN(n5713) );
  AOI21_X1 U6786 ( .B1(n5714), .B2(n6100), .A(n5713), .ZN(n5718) );
  NOR2_X1 U6787 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n5726), .ZN(n5715)
         );
  AOI22_X1 U6788 ( .A1(n5716), .A2(n6119), .B1(n5722), .B2(n5715), .ZN(n5717)
         );
  OAI211_X1 U6789 ( .C1(n5719), .C2(n3504), .A(n5718), .B(n5717), .ZN(U3000)
         );
  INV_X1 U6790 ( .A(REIP_REG_17__SCAN_IN), .ZN(n5720) );
  OAI22_X1 U6791 ( .A1(n5794), .A2(n6116), .B1(n6071), .B2(n5720), .ZN(n5721)
         );
  INV_X1 U6792 ( .A(n5721), .ZN(n5725) );
  AOI22_X1 U6793 ( .A1(n5723), .A2(n6119), .B1(n5722), .B2(n5726), .ZN(n5724)
         );
  OAI211_X1 U6794 ( .C1(n5727), .C2(n5726), .A(n5725), .B(n5724), .ZN(U3001)
         );
  AOI21_X1 U6795 ( .B1(n5730), .B2(n5729), .A(n5728), .ZN(n5743) );
  INV_X1 U6796 ( .A(n5731), .ZN(n5732) );
  AOI211_X1 U6797 ( .C1(n6557), .C2(n5742), .A(n5732), .B(n5737), .ZN(n5734)
         );
  OAI22_X1 U6798 ( .A1(n5810), .A2(n6116), .B1(n6452), .B2(n6071), .ZN(n5733)
         );
  AOI211_X1 U6799 ( .C1(n5735), .C2(n6119), .A(n5734), .B(n5733), .ZN(n5736)
         );
  OAI21_X1 U6800 ( .B1(n5743), .B2(n6557), .A(n5736), .ZN(U3002) );
  NOR2_X1 U6801 ( .A1(n5737), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5739)
         );
  INV_X1 U6802 ( .A(REIP_REG_15__SCAN_IN), .ZN(n5824) );
  OAI22_X1 U6803 ( .A1(n5818), .A2(n6116), .B1(n5824), .B2(n6071), .ZN(n5738)
         );
  AOI211_X1 U6804 ( .C1(n5740), .C2(n6119), .A(n5739), .B(n5738), .ZN(n5741)
         );
  OAI21_X1 U6805 ( .B1(n5743), .B2(n5742), .A(n5741), .ZN(U3003) );
  INV_X1 U6806 ( .A(n5829), .ZN(n5745) );
  AOI21_X1 U6807 ( .B1(n5745), .B2(n6100), .A(n5744), .ZN(n5749) );
  AOI22_X1 U6808 ( .A1(n5747), .A2(n6119), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5746), .ZN(n5748) );
  OAI211_X1 U6809 ( .C1(n5751), .C2(n5750), .A(n5749), .B(n5748), .ZN(U3005)
         );
  INV_X1 U6810 ( .A(n5752), .ZN(n5756) );
  NAND4_X1 U6811 ( .A1(n5756), .A2(n5755), .A3(n5754), .A4(n5753), .ZN(n5757)
         );
  OAI21_X1 U6812 ( .B1(n6490), .B2(n5758), .A(n5757), .ZN(U3455) );
  INV_X1 U6813 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6428) );
  AOI21_X1 U6814 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6428), .A(n6420), .ZN(n5764) );
  INV_X1 U6815 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5759) );
  INV_X1 U6816 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6598) );
  AOI21_X1 U6817 ( .B1(n5764), .B2(n5759), .A(n6516), .ZN(U2789) );
  INV_X1 U6818 ( .A(n5760), .ZN(n5761) );
  OAI21_X1 U6819 ( .B1(n5761), .B2(n6400), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5762) );
  OAI21_X1 U6820 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6401), .A(n5762), .ZN(
        U2790) );
  INV_X2 U6821 ( .A(n6516), .ZN(n6505) );
  NOR2_X1 U6822 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n5765) );
  OAI21_X1 U6823 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5765), .A(n6505), .ZN(n5763)
         );
  OAI21_X1 U6824 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6505), .A(n5763), .ZN(
        U2791) );
  NOR2_X1 U6825 ( .A1(n6516), .A2(n5764), .ZN(n6484) );
  OAI21_X1 U6826 ( .B1(BS16_N), .B2(n5765), .A(n6484), .ZN(n6482) );
  OAI21_X1 U6827 ( .B1(n6484), .B2(n6638), .A(n6482), .ZN(U2792) );
  OAI21_X1 U6828 ( .B1(n5767), .B2(n5766), .A(n6041), .ZN(U2793) );
  NOR4_X1 U6829 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n5771) );
  NOR4_X1 U6830 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(
        DATAWIDTH_REG_16__SCAN_IN), .A3(DATAWIDTH_REG_17__SCAN_IN), .A4(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n5770) );
  NOR4_X1 U6831 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5769) );
  NOR4_X1 U6832 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n5768) );
  NAND4_X1 U6833 ( .A1(n5771), .A2(n5770), .A3(n5769), .A4(n5768), .ZN(n5777)
         );
  NOR4_X1 U6834 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_18__SCAN_IN), .A4(DATAWIDTH_REG_3__SCAN_IN), .ZN(
        n5775) );
  AOI211_X1 U6835 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_12__SCAN_IN), .B(
        DATAWIDTH_REG_5__SCAN_IN), .ZN(n5774) );
  NOR4_X1 U6836 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(
        DATAWIDTH_REG_11__SCAN_IN), .A3(DATAWIDTH_REG_13__SCAN_IN), .A4(
        DATAWIDTH_REG_14__SCAN_IN), .ZN(n5773) );
  NOR4_X1 U6837 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(DATAWIDTH_REG_7__SCAN_IN), 
        .A3(DATAWIDTH_REG_8__SCAN_IN), .A4(DATAWIDTH_REG_9__SCAN_IN), .ZN(
        n5772) );
  NAND4_X1 U6838 ( .A1(n5775), .A2(n5774), .A3(n5773), .A4(n5772), .ZN(n5776)
         );
  NOR2_X1 U6839 ( .A1(n5777), .A2(n5776), .ZN(n6503) );
  INV_X1 U6840 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5779) );
  NOR3_X1 U6841 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5780) );
  OAI21_X1 U6842 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5780), .A(n6503), .ZN(n5778)
         );
  OAI21_X1 U6843 ( .B1(n6503), .B2(n5779), .A(n5778), .ZN(U2794) );
  INV_X1 U6844 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6483) );
  AOI21_X1 U6845 ( .B1(n6496), .B2(n6483), .A(n5780), .ZN(n5782) );
  INV_X1 U6846 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n5781) );
  INV_X1 U6847 ( .A(n6503), .ZN(n6498) );
  AOI22_X1 U6848 ( .A1(n6503), .A2(n5782), .B1(n5781), .B2(n6498), .ZN(U2795)
         );
  AOI22_X1 U6849 ( .A1(n5783), .A2(n5870), .B1(REIP_REG_18__SCAN_IN), .B2(
        n5796), .ZN(n5784) );
  OAI21_X1 U6850 ( .B1(n5183), .B2(n5894), .A(n5784), .ZN(n5785) );
  AOI211_X1 U6851 ( .C1(n5876), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n5875), 
        .B(n5785), .ZN(n5789) );
  OAI22_X1 U6852 ( .A1(n5907), .A2(n5861), .B1(n5786), .B2(n5873), .ZN(n5787)
         );
  INV_X1 U6853 ( .A(n5787), .ZN(n5788) );
  OAI211_X1 U6854 ( .C1(REIP_REG_18__SCAN_IN), .C2(n5790), .A(n5789), .B(n5788), .ZN(U2809) );
  INV_X1 U6855 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5792) );
  OAI22_X1 U6856 ( .A1(n5792), .A2(n5890), .B1(n5791), .B2(n5889), .ZN(n5793)
         );
  AOI211_X1 U6857 ( .C1(n5865), .C2(EBX_REG_17__SCAN_IN), .A(n5875), .B(n5793), 
        .ZN(n5800) );
  NOR2_X1 U6858 ( .A1(n5794), .A2(n5873), .ZN(n5795) );
  AOI21_X1 U6859 ( .B1(n5912), .B2(n5880), .A(n5795), .ZN(n5799) );
  OAI21_X1 U6860 ( .B1(REIP_REG_17__SCAN_IN), .B2(n5797), .A(n5796), .ZN(n5798) );
  NAND3_X1 U6861 ( .A1(n5800), .A2(n5799), .A3(n5798), .ZN(U2810) );
  NAND3_X1 U6862 ( .A1(n5802), .A2(n5824), .A3(n5801), .ZN(n5816) );
  INV_X1 U6863 ( .A(n5803), .ZN(n5808) );
  AOI22_X1 U6864 ( .A1(PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n5876), .B1(n5804), 
        .B2(n5870), .ZN(n5805) );
  OAI211_X1 U6865 ( .C1(n5894), .C2(n5806), .A(n5805), .B(n5858), .ZN(n5807)
         );
  AOI21_X1 U6866 ( .B1(n5808), .B2(n6452), .A(n5807), .ZN(n5809) );
  OAI21_X1 U6867 ( .B1(n5810), .B2(n5873), .A(n5809), .ZN(n5811) );
  AOI21_X1 U6868 ( .B1(n5917), .B2(n5880), .A(n5811), .ZN(n5812) );
  OAI221_X1 U6869 ( .B1(n6452), .B2(n5823), .C1(n6452), .C2(n5816), .A(n5812), 
        .ZN(U2811) );
  INV_X1 U6870 ( .A(n5813), .ZN(n5821) );
  OAI22_X1 U6871 ( .A1(n6639), .A2(n5894), .B1(n5814), .B2(n5890), .ZN(n5820)
         );
  AOI21_X1 U6872 ( .B1(n5815), .B2(n5870), .A(n5875), .ZN(n5817) );
  OAI211_X1 U6873 ( .C1(n5818), .C2(n5873), .A(n5817), .B(n5816), .ZN(n5819)
         );
  AOI211_X1 U6874 ( .C1(n5821), .C2(n5880), .A(n5820), .B(n5819), .ZN(n5822)
         );
  OAI21_X1 U6875 ( .B1(n5824), .B2(n5823), .A(n5822), .ZN(U2812) );
  NOR3_X1 U6876 ( .A1(n5826), .A2(REIP_REG_13__SCAN_IN), .A3(n5825), .ZN(n5827) );
  AOI21_X1 U6877 ( .B1(n5870), .B2(n5828), .A(n5827), .ZN(n5836) );
  NOR2_X1 U6878 ( .A1(n5829), .A2(n5873), .ZN(n5830) );
  AOI211_X1 U6879 ( .C1(n5876), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5875), 
        .B(n5830), .ZN(n5831) );
  OAI21_X1 U6880 ( .B1(n5832), .B2(n5861), .A(n5831), .ZN(n5833) );
  AOI221_X1 U6881 ( .B1(n5837), .B2(REIP_REG_13__SCAN_IN), .C1(n5834), .C2(
        REIP_REG_13__SCAN_IN), .A(n5833), .ZN(n5835) );
  OAI211_X1 U6882 ( .C1(n6621), .C2(n5894), .A(n5836), .B(n5835), .ZN(U2814)
         );
  AOI22_X1 U6883 ( .A1(n5838), .A2(n5870), .B1(REIP_REG_11__SCAN_IN), .B2(
        n5837), .ZN(n5846) );
  OR3_X1 U6884 ( .A1(n5883), .A2(REIP_REG_11__SCAN_IN), .A3(n5839), .ZN(n5841)
         );
  AOI21_X1 U6885 ( .B1(n5876), .B2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n5875), 
        .ZN(n5840) );
  OAI211_X1 U6886 ( .C1(n5906), .C2(n5894), .A(n5841), .B(n5840), .ZN(n5843)
         );
  NOR2_X1 U6887 ( .A1(n6014), .A2(n5861), .ZN(n5842) );
  AOI211_X1 U6888 ( .C1(n5844), .C2(n5886), .A(n5843), .B(n5842), .ZN(n5845)
         );
  NAND2_X1 U6889 ( .A1(n5846), .A2(n5845), .ZN(U2816) );
  AOI22_X1 U6890 ( .A1(n5848), .A2(n5870), .B1(REIP_REG_9__SCAN_IN), .B2(n5847), .ZN(n5855) );
  AOI22_X1 U6891 ( .A1(n6065), .A2(n5886), .B1(PHYADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n5876), .ZN(n5854) );
  AOI21_X1 U6892 ( .B1(n5865), .B2(EBX_REG_9__SCAN_IN), .A(n5875), .ZN(n5853)
         );
  INV_X1 U6893 ( .A(n5849), .ZN(n5851) );
  AOI22_X1 U6894 ( .A1(n5851), .A2(n5880), .B1(n5850), .B2(n6442), .ZN(n5852)
         );
  NAND4_X1 U6895 ( .A1(n5855), .A2(n5854), .A3(n5853), .A4(n5852), .ZN(U2818)
         );
  OAI21_X1 U6896 ( .B1(REIP_REG_7__SCAN_IN), .B2(REIP_REG_6__SCAN_IN), .A(
        n5856), .ZN(n5868) );
  AOI22_X1 U6897 ( .A1(n5857), .A2(n5870), .B1(REIP_REG_7__SCAN_IN), .B2(n5869), .ZN(n5867) );
  NAND2_X1 U6898 ( .A1(n5886), .A2(n6081), .ZN(n5859) );
  OAI211_X1 U6899 ( .C1(n5890), .C2(n5860), .A(n5859), .B(n5858), .ZN(n5864)
         );
  NOR2_X1 U6900 ( .A1(n5862), .A2(n5861), .ZN(n5863) );
  AOI211_X1 U6901 ( .C1(n5865), .C2(EBX_REG_7__SCAN_IN), .A(n5864), .B(n5863), 
        .ZN(n5866) );
  OAI211_X1 U6902 ( .C1(n5883), .C2(n5868), .A(n5867), .B(n5866), .ZN(U2820)
         );
  INV_X1 U6903 ( .A(n6023), .ZN(n5871) );
  AOI22_X1 U6904 ( .A1(n5871), .A2(n5870), .B1(REIP_REG_6__SCAN_IN), .B2(n5869), .ZN(n5882) );
  NOR2_X1 U6905 ( .A1(n5873), .A2(n5872), .ZN(n5874) );
  AOI211_X1 U6906 ( .C1(n5876), .C2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n5875), 
        .B(n5874), .ZN(n5877) );
  OAI21_X1 U6907 ( .B1(n5894), .B2(n5878), .A(n5877), .ZN(n5879) );
  AOI21_X1 U6908 ( .B1(n6019), .B2(n5880), .A(n5879), .ZN(n5881) );
  OAI211_X1 U6909 ( .C1(REIP_REG_6__SCAN_IN), .C2(n5883), .A(n5882), .B(n5881), 
        .ZN(U2821) );
  INV_X1 U6910 ( .A(n5884), .ZN(n5885) );
  AOI22_X1 U6911 ( .A1(REIP_REG_0__SCAN_IN), .A2(n5887), .B1(n5886), .B2(n5885), .ZN(n5898) );
  NAND2_X1 U6912 ( .A1(n5888), .A2(n6369), .ZN(n5893) );
  NAND2_X1 U6913 ( .A1(n5890), .A2(n5889), .ZN(n5891) );
  NAND2_X1 U6914 ( .A1(n5891), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n5892)
         );
  OAI211_X1 U6915 ( .C1(n5895), .C2(n5894), .A(n5893), .B(n5892), .ZN(n5896)
         );
  INV_X1 U6916 ( .A(n5896), .ZN(n5897) );
  OAI211_X1 U6917 ( .C1(n5899), .C2(n6044), .A(n5898), .B(n5897), .ZN(U2827)
         );
  OAI22_X1 U6918 ( .A1(n6014), .A2(n5902), .B1(n5901), .B2(n5900), .ZN(n5903)
         );
  INV_X1 U6919 ( .A(n5903), .ZN(n5904) );
  OAI21_X1 U6920 ( .B1(n5906), .B2(n5905), .A(n5904), .ZN(U2848) );
  INV_X1 U6921 ( .A(n5907), .ZN(n5908) );
  AOI22_X1 U6922 ( .A1(n5908), .A2(n5916), .B1(n5915), .B2(DATAI_2_), .ZN(
        n5911) );
  AOI22_X1 U6923 ( .A1(EAX_REG_18__SCAN_IN), .A2(n5909), .B1(n3004), .B2(
        DATAI_18_), .ZN(n5910) );
  NAND2_X1 U6924 ( .A1(n5911), .A2(n5910), .ZN(U2873) );
  AOI22_X1 U6925 ( .A1(n5912), .A2(n5916), .B1(n5915), .B2(DATAI_1_), .ZN(
        n5914) );
  AOI22_X1 U6926 ( .A1(EAX_REG_17__SCAN_IN), .A2(n5909), .B1(n3004), .B2(
        DATAI_17_), .ZN(n5913) );
  NAND2_X1 U6927 ( .A1(n5914), .A2(n5913), .ZN(U2874) );
  AOI22_X1 U6928 ( .A1(n5917), .A2(n5916), .B1(n5915), .B2(DATAI_0_), .ZN(
        n5919) );
  AOI22_X1 U6929 ( .A1(EAX_REG_16__SCAN_IN), .A2(n5909), .B1(n3004), .B2(
        DATAI_16_), .ZN(n5918) );
  NAND2_X1 U6930 ( .A1(n5919), .A2(n5918), .ZN(U2875) );
  INV_X1 U6931 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6012) );
  AOI22_X1 U6932 ( .A1(n5943), .A2(LWORD_REG_15__SCAN_IN), .B1(n5934), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n5921) );
  OAI21_X1 U6933 ( .B1(n6012), .B2(n5945), .A(n5921), .ZN(U2908) );
  AOI22_X1 U6934 ( .A1(n5943), .A2(LWORD_REG_14__SCAN_IN), .B1(n5934), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n5922) );
  OAI21_X1 U6935 ( .B1(n6626), .B2(n5945), .A(n5922), .ZN(U2909) );
  INV_X1 U6936 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6003) );
  AOI22_X1 U6937 ( .A1(n5943), .A2(LWORD_REG_13__SCAN_IN), .B1(n5934), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n5923) );
  OAI21_X1 U6938 ( .B1(n6003), .B2(n5945), .A(n5923), .ZN(U2910) );
  INV_X1 U6939 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5999) );
  AOI22_X1 U6940 ( .A1(n5943), .A2(LWORD_REG_12__SCAN_IN), .B1(n5934), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n5924) );
  OAI21_X1 U6941 ( .B1(n5999), .B2(n5945), .A(n5924), .ZN(U2911) );
  INV_X1 U6942 ( .A(EAX_REG_11__SCAN_IN), .ZN(n5996) );
  AOI22_X1 U6943 ( .A1(n5943), .A2(LWORD_REG_11__SCAN_IN), .B1(n5934), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n5925) );
  OAI21_X1 U6944 ( .B1(n5996), .B2(n5945), .A(n5925), .ZN(U2912) );
  AOI22_X1 U6945 ( .A1(n5943), .A2(LWORD_REG_10__SCAN_IN), .B1(n5934), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n5926) );
  OAI21_X1 U6946 ( .B1(n6601), .B2(n5945), .A(n5926), .ZN(U2913) );
  INV_X1 U6947 ( .A(EAX_REG_9__SCAN_IN), .ZN(n5991) );
  AOI22_X1 U6948 ( .A1(n5943), .A2(LWORD_REG_9__SCAN_IN), .B1(n5934), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n5927) );
  OAI21_X1 U6949 ( .B1(n5991), .B2(n5945), .A(n5927), .ZN(U2914) );
  AOI22_X1 U6950 ( .A1(DATAO_REG_8__SCAN_IN), .A2(n5934), .B1(n5943), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n5928) );
  OAI21_X1 U6951 ( .B1(n6550), .B2(n5945), .A(n5928), .ZN(U2915) );
  AOI22_X1 U6952 ( .A1(n5943), .A2(LWORD_REG_7__SCAN_IN), .B1(n5934), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n5929) );
  OAI21_X1 U6953 ( .B1(n5930), .B2(n5945), .A(n5929), .ZN(U2916) );
  AOI22_X1 U6954 ( .A1(n5943), .A2(LWORD_REG_6__SCAN_IN), .B1(n5934), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n5931) );
  OAI21_X1 U6955 ( .B1(n5000), .B2(n5945), .A(n5931), .ZN(U2917) );
  AOI22_X1 U6956 ( .A1(n5943), .A2(LWORD_REG_5__SCAN_IN), .B1(n5934), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n5932) );
  OAI21_X1 U6957 ( .B1(n5933), .B2(n5945), .A(n5932), .ZN(U2918) );
  AOI22_X1 U6958 ( .A1(n5943), .A2(LWORD_REG_4__SCAN_IN), .B1(n5934), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n5935) );
  OAI21_X1 U6959 ( .B1(n5936), .B2(n5945), .A(n5935), .ZN(U2919) );
  AOI22_X1 U6960 ( .A1(n5943), .A2(LWORD_REG_3__SCAN_IN), .B1(n5934), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n5937) );
  OAI21_X1 U6961 ( .B1(n5938), .B2(n5945), .A(n5937), .ZN(U2920) );
  AOI22_X1 U6962 ( .A1(n5943), .A2(LWORD_REG_2__SCAN_IN), .B1(n5934), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n5939) );
  OAI21_X1 U6963 ( .B1(n5940), .B2(n5945), .A(n5939), .ZN(U2921) );
  AOI22_X1 U6964 ( .A1(LWORD_REG_1__SCAN_IN), .A2(n5943), .B1(n5934), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n5941) );
  OAI21_X1 U6965 ( .B1(n5942), .B2(n5945), .A(n5941), .ZN(U2922) );
  AOI22_X1 U6966 ( .A1(n5943), .A2(LWORD_REG_0__SCAN_IN), .B1(n5934), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n5944) );
  OAI21_X1 U6967 ( .B1(n5946), .B2(n5945), .A(n5944), .ZN(U2923) );
  AOI22_X1 U6968 ( .A1(n6009), .A2(UWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_16__SCAN_IN), .B2(n6004), .ZN(n5948) );
  OAI21_X1 U6969 ( .B1(n6007), .B2(n5972), .A(n5948), .ZN(U2924) );
  AOI22_X1 U6970 ( .A1(n6009), .A2(UWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_17__SCAN_IN), .B2(n6004), .ZN(n5949) );
  OAI21_X1 U6971 ( .B1(n6007), .B2(n5974), .A(n5949), .ZN(U2925) );
  AOI22_X1 U6972 ( .A1(n6009), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n6004), .ZN(n5950) );
  OAI21_X1 U6973 ( .B1(n6007), .B2(n5976), .A(n5950), .ZN(U2926) );
  AOI22_X1 U6974 ( .A1(n6009), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n6004), .ZN(n5951) );
  OAI21_X1 U6975 ( .B1(n6007), .B2(n5978), .A(n5951), .ZN(U2927) );
  AOI22_X1 U6976 ( .A1(n6009), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n6004), .ZN(n5952) );
  OAI21_X1 U6977 ( .B1(n6007), .B2(n5980), .A(n5952), .ZN(U2928) );
  AOI22_X1 U6978 ( .A1(n6009), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n6004), .ZN(n5953) );
  OAI21_X1 U6979 ( .B1(n6007), .B2(n5982), .A(n5953), .ZN(U2929) );
  AOI22_X1 U6980 ( .A1(n6009), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n6004), .ZN(n5954) );
  OAI21_X1 U6981 ( .B1(n6007), .B2(n5984), .A(n5954), .ZN(U2930) );
  AOI22_X1 U6982 ( .A1(n6009), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n6004), .ZN(n5955) );
  OAI21_X1 U6983 ( .B1(n6007), .B2(n5986), .A(n5955), .ZN(U2931) );
  AOI22_X1 U6984 ( .A1(n6009), .A2(UWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_24__SCAN_IN), .B2(n6004), .ZN(n5956) );
  OAI21_X1 U6985 ( .B1(n6007), .B2(n5988), .A(n5956), .ZN(U2932) );
  INV_X1 U6986 ( .A(DATAI_9_), .ZN(n5957) );
  NOR2_X1 U6987 ( .A1(n6007), .A2(n5957), .ZN(n5989) );
  AOI21_X1 U6988 ( .B1(UWORD_REG_9__SCAN_IN), .B2(n6001), .A(n5989), .ZN(n5958) );
  OAI21_X1 U6989 ( .B1(n5959), .B2(n6011), .A(n5958), .ZN(U2933) );
  AOI22_X1 U6990 ( .A1(n6009), .A2(UWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_26__SCAN_IN), .B2(n6004), .ZN(n5960) );
  OAI21_X1 U6991 ( .B1(n6007), .B2(n5993), .A(n5960), .ZN(U2934) );
  INV_X1 U6992 ( .A(DATAI_11_), .ZN(n5961) );
  NOR2_X1 U6993 ( .A1(n6007), .A2(n5961), .ZN(n5994) );
  AOI21_X1 U6994 ( .B1(UWORD_REG_11__SCAN_IN), .B2(n6009), .A(n5994), .ZN(
        n5962) );
  OAI21_X1 U6995 ( .B1(n5963), .B2(n6011), .A(n5962), .ZN(U2935) );
  INV_X1 U6996 ( .A(DATAI_12_), .ZN(n5964) );
  NOR2_X1 U6997 ( .A1(n6007), .A2(n5964), .ZN(n5997) );
  AOI21_X1 U6998 ( .B1(UWORD_REG_12__SCAN_IN), .B2(n6009), .A(n5997), .ZN(
        n5965) );
  OAI21_X1 U6999 ( .B1(n5966), .B2(n6011), .A(n5965), .ZN(U2936) );
  INV_X1 U7000 ( .A(DATAI_13_), .ZN(n5967) );
  NOR2_X1 U7001 ( .A1(n6007), .A2(n5967), .ZN(n6000) );
  AOI21_X1 U7002 ( .B1(UWORD_REG_13__SCAN_IN), .B2(n6001), .A(n6000), .ZN(
        n5968) );
  OAI21_X1 U7003 ( .B1(n5969), .B2(n6011), .A(n5968), .ZN(U2937) );
  AOI22_X1 U7004 ( .A1(n6009), .A2(UWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_30__SCAN_IN), .B2(n6004), .ZN(n5970) );
  OAI21_X1 U7005 ( .B1(n6007), .B2(n6006), .A(n5970), .ZN(U2938) );
  AOI22_X1 U7006 ( .A1(n6009), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n6004), .ZN(n5971) );
  OAI21_X1 U7007 ( .B1(n6007), .B2(n5972), .A(n5971), .ZN(U2939) );
  AOI22_X1 U7008 ( .A1(n6009), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n6004), .ZN(n5973) );
  OAI21_X1 U7009 ( .B1(n6007), .B2(n5974), .A(n5973), .ZN(U2940) );
  AOI22_X1 U7010 ( .A1(n6009), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n6004), .ZN(n5975) );
  OAI21_X1 U7011 ( .B1(n6007), .B2(n5976), .A(n5975), .ZN(U2941) );
  AOI22_X1 U7012 ( .A1(n6009), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n6004), .ZN(n5977) );
  OAI21_X1 U7013 ( .B1(n6007), .B2(n5978), .A(n5977), .ZN(U2942) );
  AOI22_X1 U7014 ( .A1(n6009), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n6004), .ZN(n5979) );
  OAI21_X1 U7015 ( .B1(n6007), .B2(n5980), .A(n5979), .ZN(U2943) );
  AOI22_X1 U7016 ( .A1(n6009), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n6004), .ZN(n5981) );
  OAI21_X1 U7017 ( .B1(n6007), .B2(n5982), .A(n5981), .ZN(U2944) );
  AOI22_X1 U7018 ( .A1(n6009), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n6004), .ZN(n5983) );
  OAI21_X1 U7019 ( .B1(n6007), .B2(n5984), .A(n5983), .ZN(U2945) );
  AOI22_X1 U7020 ( .A1(n6009), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n6004), .ZN(n5985) );
  OAI21_X1 U7021 ( .B1(n6007), .B2(n5986), .A(n5985), .ZN(U2946) );
  AOI22_X1 U7022 ( .A1(n6009), .A2(LWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_8__SCAN_IN), .B2(n6004), .ZN(n5987) );
  OAI21_X1 U7023 ( .B1(n6007), .B2(n5988), .A(n5987), .ZN(U2947) );
  AOI21_X1 U7024 ( .B1(LWORD_REG_9__SCAN_IN), .B2(n6009), .A(n5989), .ZN(n5990) );
  OAI21_X1 U7025 ( .B1(n5991), .B2(n6011), .A(n5990), .ZN(U2948) );
  AOI22_X1 U7026 ( .A1(n6009), .A2(LWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_10__SCAN_IN), .B2(n6004), .ZN(n5992) );
  OAI21_X1 U7027 ( .B1(n6007), .B2(n5993), .A(n5992), .ZN(U2949) );
  AOI21_X1 U7028 ( .B1(LWORD_REG_11__SCAN_IN), .B2(n6001), .A(n5994), .ZN(
        n5995) );
  OAI21_X1 U7029 ( .B1(n5996), .B2(n6011), .A(n5995), .ZN(U2950) );
  AOI21_X1 U7030 ( .B1(LWORD_REG_12__SCAN_IN), .B2(n6001), .A(n5997), .ZN(
        n5998) );
  OAI21_X1 U7031 ( .B1(n5999), .B2(n6011), .A(n5998), .ZN(U2951) );
  AOI21_X1 U7032 ( .B1(LWORD_REG_13__SCAN_IN), .B2(n6001), .A(n6000), .ZN(
        n6002) );
  OAI21_X1 U7033 ( .B1(n6003), .B2(n6011), .A(n6002), .ZN(U2952) );
  AOI22_X1 U7034 ( .A1(n6009), .A2(LWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_14__SCAN_IN), .B2(n6004), .ZN(n6005) );
  OAI21_X1 U7035 ( .B1(n6007), .B2(n6006), .A(n6005), .ZN(U2953) );
  INV_X1 U7036 ( .A(n6007), .ZN(n6008) );
  AOI22_X1 U7037 ( .A1(n6009), .A2(LWORD_REG_15__SCAN_IN), .B1(n6008), .B2(
        DATAI_15_), .ZN(n6010) );
  OAI21_X1 U7038 ( .B1(n6012), .B2(n6011), .A(n6010), .ZN(U2954) );
  AOI22_X1 U7039 ( .A1(n6112), .A2(REIP_REG_11__SCAN_IN), .B1(n6047), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6017) );
  OAI22_X1 U7040 ( .A1(n6014), .A2(n6043), .B1(n6013), .B2(n6040), .ZN(n6015)
         );
  INV_X1 U7041 ( .A(n6015), .ZN(n6016) );
  OAI211_X1 U7042 ( .C1(n6018), .C2(n6041), .A(n6017), .B(n6016), .ZN(U2975)
         );
  AOI22_X1 U7043 ( .A1(n6112), .A2(REIP_REG_6__SCAN_IN), .B1(n6047), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6022) );
  AOI22_X1 U7044 ( .A1(n6020), .A2(n6036), .B1(n6035), .B2(n6019), .ZN(n6021)
         );
  OAI211_X1 U7045 ( .C1(n6040), .C2(n6023), .A(n6022), .B(n6021), .ZN(U2980)
         );
  AOI22_X1 U7046 ( .A1(n6112), .A2(REIP_REG_4__SCAN_IN), .B1(n6047), .B2(
        PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6029) );
  AOI21_X1 U7047 ( .B1(n6026), .B2(n6025), .A(n6024), .ZN(n6089) );
  AOI22_X1 U7048 ( .A1(n6089), .A2(n6036), .B1(n6035), .B2(n6027), .ZN(n6028)
         );
  OAI211_X1 U7049 ( .C1(n6040), .C2(n6030), .A(n6029), .B(n6028), .ZN(U2982)
         );
  AOI22_X1 U7050 ( .A1(n6112), .A2(REIP_REG_2__SCAN_IN), .B1(n6047), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6038) );
  XNOR2_X1 U7051 ( .A(n6032), .B(n3422), .ZN(n6033) );
  XNOR2_X1 U7052 ( .A(n6031), .B(n6033), .ZN(n6120) );
  AOI22_X1 U7053 ( .A1(n6120), .A2(n6036), .B1(n6035), .B2(n6034), .ZN(n6037)
         );
  OAI211_X1 U7054 ( .C1(n6040), .C2(n6039), .A(n6038), .B(n6037), .ZN(U2984)
         );
  OAI22_X1 U7055 ( .A1(n6044), .A2(n6043), .B1(n6042), .B2(n6041), .ZN(n6045)
         );
  AOI221_X1 U7056 ( .B1(n6047), .B2(PHYADDRPOINTER_REG_0__SCAN_IN), .C1(n6046), 
        .C2(PHYADDRPOINTER_REG_0__SCAN_IN), .A(n6045), .ZN(n6049) );
  NAND2_X1 U7057 ( .A1(n6049), .A2(n6048), .ZN(U2986) );
  NOR2_X1 U7058 ( .A1(n6058), .A2(n6092), .ZN(n6082) );
  NAND2_X1 U7059 ( .A1(n6075), .A2(n6082), .ZN(n6070) );
  INV_X1 U7060 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6050) );
  AOI22_X1 U7061 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n6050), .B1(
        INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n5365), .ZN(n6063) );
  AOI21_X1 U7062 ( .B1(n6052), .B2(n6100), .A(n6051), .ZN(n6062) );
  INV_X1 U7063 ( .A(n6053), .ZN(n6055) );
  OAI21_X1 U7064 ( .B1(n6056), .B2(n6055), .A(n6054), .ZN(n6057) );
  AOI21_X1 U7065 ( .B1(n6111), .B2(n6058), .A(n6057), .ZN(n6087) );
  OAI21_X1 U7066 ( .B1(n6059), .B2(n6075), .A(n6087), .ZN(n6066) );
  AOI22_X1 U7067 ( .A1(n6060), .A2(n6119), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6066), .ZN(n6061) );
  OAI211_X1 U7068 ( .C1(n6070), .C2(n6063), .A(n6062), .B(n6061), .ZN(U3008)
         );
  AOI21_X1 U7069 ( .B1(n6065), .B2(n6100), .A(n6064), .ZN(n6069) );
  AOI22_X1 U7070 ( .A1(n6067), .A2(n6119), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6066), .ZN(n6068) );
  OAI211_X1 U7071 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6070), .A(n6069), 
        .B(n6068), .ZN(U3009) );
  OAI22_X1 U7072 ( .A1(n6072), .A2(n6116), .B1(n6439), .B2(n6071), .ZN(n6073)
         );
  AOI21_X1 U7073 ( .B1(n6074), .B2(n6119), .A(n6073), .ZN(n6078) );
  INV_X1 U7074 ( .A(n6075), .ZN(n6076) );
  OAI211_X1 U7075 ( .C1(INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .A(n6082), .B(n6076), .ZN(n6077) );
  OAI211_X1 U7076 ( .C1(n6087), .C2(n3496), .A(n6078), .B(n6077), .ZN(U3010)
         );
  INV_X1 U7077 ( .A(n6079), .ZN(n6080) );
  AOI21_X1 U7078 ( .B1(n6081), .B2(n6100), .A(n6080), .ZN(n6085) );
  AOI22_X1 U7079 ( .A1(n6083), .A2(n6119), .B1(n6082), .B2(n6086), .ZN(n6084)
         );
  OAI211_X1 U7080 ( .C1(n6087), .C2(n6086), .A(n6085), .B(n6084), .ZN(U3011)
         );
  NOR2_X1 U7081 ( .A1(n6088), .A2(n6091), .ZN(n6117) );
  NOR2_X1 U7082 ( .A1(n6117), .A2(n6109), .ZN(n6107) );
  AOI222_X1 U7083 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6112), .B1(n6100), .B2(
        n6090), .C1(n6119), .C2(n6089), .ZN(n6096) );
  INV_X1 U7084 ( .A(n6091), .ZN(n6093) );
  NOR2_X1 U7085 ( .A1(n6093), .A2(n6092), .ZN(n6103) );
  OAI211_X1 U7086 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A(n6103), .B(n6094), .ZN(n6095) );
  OAI211_X1 U7087 ( .C1(n6107), .C2(n6097), .A(n6096), .B(n6095), .ZN(U3014)
         );
  AOI21_X1 U7088 ( .B1(n6100), .B2(n6099), .A(n6098), .ZN(n6105) );
  INV_X1 U7089 ( .A(n6101), .ZN(n6102) );
  AOI22_X1 U7090 ( .A1(n6103), .A2(n6106), .B1(n6102), .B2(n6119), .ZN(n6104)
         );
  OAI211_X1 U7091 ( .C1(n6107), .C2(n6106), .A(n6105), .B(n6104), .ZN(U3015)
         );
  NAND2_X1 U7092 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6108), .ZN(n6123)
         );
  INV_X1 U7093 ( .A(n6109), .ZN(n6122) );
  NAND3_X1 U7094 ( .A1(n6111), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .A3(n6110), 
        .ZN(n6114) );
  NAND2_X1 U7095 ( .A1(n6112), .A2(REIP_REG_2__SCAN_IN), .ZN(n6113) );
  OAI211_X1 U7096 ( .C1(n6116), .C2(n6115), .A(n6114), .B(n6113), .ZN(n6118)
         );
  AOI211_X1 U7097 ( .C1(n6120), .C2(n6119), .A(n6118), .B(n6117), .ZN(n6121)
         );
  OAI221_X1 U7098 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6123), .C1(n3422), .C2(n6122), .A(n6121), .ZN(U3016) );
  NOR2_X1 U7099 ( .A1(n6125), .A2(n6124), .ZN(U3019) );
  INV_X1 U7100 ( .A(n6126), .ZN(n6131) );
  AOI22_X1 U7101 ( .A1(n6314), .A2(n6132), .B1(n6313), .B2(n6131), .ZN(n6128)
         );
  AOI22_X1 U7102 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6134), .B1(n6259), 
        .B2(n6133), .ZN(n6127) );
  OAI211_X1 U7103 ( .C1(n6137), .C2(n6316), .A(n6128), .B(n6127), .ZN(U3046)
         );
  AOI22_X1 U7104 ( .A1(n6347), .A2(n6132), .B1(n6348), .B2(n6131), .ZN(n6130)
         );
  AOI22_X1 U7105 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6134), .B1(n6350), 
        .B2(n6133), .ZN(n6129) );
  OAI211_X1 U7106 ( .C1(n6137), .C2(n6277), .A(n6130), .B(n6129), .ZN(U3050)
         );
  AOI22_X1 U7107 ( .A1(n6357), .A2(n6132), .B1(n6355), .B2(n6131), .ZN(n6136)
         );
  AOI22_X1 U7108 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6134), .B1(n6279), 
        .B2(n6133), .ZN(n6135) );
  OAI211_X1 U7109 ( .C1(n6137), .C2(n6360), .A(n6136), .B(n6135), .ZN(U3051)
         );
  NOR2_X1 U7110 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6138), .ZN(n6175)
         );
  INV_X1 U7111 ( .A(n6139), .ZN(n6144) );
  NAND3_X1 U7112 ( .A1(n6141), .A2(n6140), .A3(n6201), .ZN(n6142) );
  OAI21_X1 U7113 ( .B1(n6144), .B2(n6143), .A(n6142), .ZN(n6174) );
  AOI22_X1 U7114 ( .A1(n6294), .A2(n6175), .B1(n6243), .B2(n6174), .ZN(n6155)
         );
  AOI21_X1 U7115 ( .B1(n6152), .B2(n6200), .A(n6638), .ZN(n6151) );
  NAND2_X1 U7116 ( .A1(n6245), .A2(n6145), .ZN(n6150) );
  INV_X1 U7117 ( .A(n6175), .ZN(n6148) );
  AOI211_X1 U7118 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6148), .A(n6147), .B(
        n6146), .ZN(n6149) );
  OAI211_X1 U7119 ( .C1(n6151), .C2(n6150), .A(n6149), .B(n6201), .ZN(n6178)
         );
  AOI22_X1 U7120 ( .A1(n6178), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6153), 
        .B2(n6176), .ZN(n6154) );
  OAI211_X1 U7121 ( .C1(n6156), .C2(n6200), .A(n6155), .B(n6154), .ZN(U3068)
         );
  AOI22_X1 U7122 ( .A1(n6307), .A2(n6175), .B1(n6256), .B2(n6174), .ZN(n6159)
         );
  AOI22_X1 U7123 ( .A1(n6178), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6157), 
        .B2(n6176), .ZN(n6158) );
  OAI211_X1 U7124 ( .C1(n6160), .C2(n6200), .A(n6159), .B(n6158), .ZN(U3069)
         );
  AOI22_X1 U7125 ( .A1(n6314), .A2(n6175), .B1(n6259), .B2(n6174), .ZN(n6163)
         );
  AOI22_X1 U7126 ( .A1(n6178), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6161), 
        .B2(n6176), .ZN(n6162) );
  OAI211_X1 U7127 ( .C1(n6164), .C2(n6200), .A(n6163), .B(n6162), .ZN(U3070)
         );
  AOI22_X1 U7128 ( .A1(n6322), .A2(n6175), .B1(n6262), .B2(n6174), .ZN(n6166)
         );
  AOI22_X1 U7129 ( .A1(n6178), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6220), 
        .B2(n6176), .ZN(n6165) );
  OAI211_X1 U7130 ( .C1(n6223), .C2(n6200), .A(n6166), .B(n6165), .ZN(U3071)
         );
  AOI22_X1 U7131 ( .A1(n6330), .A2(n6175), .B1(n6265), .B2(n6174), .ZN(n6168)
         );
  AOI22_X1 U7132 ( .A1(n6178), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6329), 
        .B2(n6176), .ZN(n6167) );
  OAI211_X1 U7133 ( .C1(n6332), .C2(n6200), .A(n6168), .B(n6167), .ZN(U3072)
         );
  AOI22_X1 U7134 ( .A1(n6338), .A2(n6175), .B1(n6270), .B2(n6174), .ZN(n6170)
         );
  AOI22_X1 U7135 ( .A1(n6178), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6337), 
        .B2(n6176), .ZN(n6169) );
  OAI211_X1 U7136 ( .C1(n6340), .C2(n6200), .A(n6170), .B(n6169), .ZN(U3073)
         );
  AOI22_X1 U7137 ( .A1(n6350), .A2(n6174), .B1(n6347), .B2(n6175), .ZN(n6172)
         );
  AOI22_X1 U7138 ( .A1(n6178), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6346), 
        .B2(n6176), .ZN(n6171) );
  OAI211_X1 U7139 ( .C1(n6173), .C2(n6200), .A(n6172), .B(n6171), .ZN(U3074)
         );
  AOI22_X1 U7140 ( .A1(n6357), .A2(n6175), .B1(n6279), .B2(n6174), .ZN(n6180)
         );
  AOI22_X1 U7141 ( .A1(n6178), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6177), 
        .B2(n6176), .ZN(n6179) );
  OAI211_X1 U7142 ( .C1(n6181), .C2(n6200), .A(n6180), .B(n6179), .ZN(U3075)
         );
  AOI22_X1 U7143 ( .A1(n6307), .A2(n6195), .B1(n6306), .B2(n6194), .ZN(n6183)
         );
  AOI22_X1 U7144 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6197), .B1(n6256), 
        .B2(n6196), .ZN(n6182) );
  OAI211_X1 U7145 ( .C1(n6309), .C2(n6200), .A(n6183), .B(n6182), .ZN(U3077)
         );
  AOI22_X1 U7146 ( .A1(n6314), .A2(n6195), .B1(n6313), .B2(n6194), .ZN(n6185)
         );
  AOI22_X1 U7147 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6197), .B1(n6259), 
        .B2(n6196), .ZN(n6184) );
  OAI211_X1 U7148 ( .C1(n6316), .C2(n6200), .A(n6185), .B(n6184), .ZN(U3078)
         );
  AOI22_X1 U7149 ( .A1(n6322), .A2(n6195), .B1(n6321), .B2(n6194), .ZN(n6187)
         );
  AOI22_X1 U7150 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6197), .B1(n6262), 
        .B2(n6196), .ZN(n6186) );
  OAI211_X1 U7151 ( .C1(n6324), .C2(n6200), .A(n6187), .B(n6186), .ZN(U3079)
         );
  AOI22_X1 U7152 ( .A1(n6330), .A2(n6195), .B1(n6266), .B2(n6194), .ZN(n6189)
         );
  AOI22_X1 U7153 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6197), .B1(n6265), 
        .B2(n6196), .ZN(n6188) );
  OAI211_X1 U7154 ( .C1(n6269), .C2(n6200), .A(n6189), .B(n6188), .ZN(U3080)
         );
  AOI22_X1 U7155 ( .A1(n6338), .A2(n6195), .B1(n6271), .B2(n6194), .ZN(n6191)
         );
  AOI22_X1 U7156 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6197), .B1(n6270), 
        .B2(n6196), .ZN(n6190) );
  OAI211_X1 U7157 ( .C1(n6274), .C2(n6200), .A(n6191), .B(n6190), .ZN(U3081)
         );
  AOI22_X1 U7158 ( .A1(n6347), .A2(n6195), .B1(n6348), .B2(n6194), .ZN(n6193)
         );
  AOI22_X1 U7159 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6197), .B1(n6350), 
        .B2(n6196), .ZN(n6192) );
  OAI211_X1 U7160 ( .C1(n6277), .C2(n6200), .A(n6193), .B(n6192), .ZN(U3082)
         );
  AOI22_X1 U7161 ( .A1(n6357), .A2(n6195), .B1(n6355), .B2(n6194), .ZN(n6199)
         );
  AOI22_X1 U7162 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6197), .B1(n6279), 
        .B2(n6196), .ZN(n6198) );
  OAI211_X1 U7163 ( .C1(n6360), .C2(n6200), .A(n6199), .B(n6198), .ZN(U3083)
         );
  NOR2_X1 U7164 ( .A1(n6202), .A2(n6201), .ZN(n6232) );
  INV_X1 U7165 ( .A(n6284), .ZN(n6231) );
  AOI22_X1 U7166 ( .A1(n6294), .A2(n6232), .B1(n6293), .B2(n6231), .ZN(n6215)
         );
  AOI21_X1 U7167 ( .B1(n6205), .B2(n6204), .A(n6295), .ZN(n6209) );
  AOI21_X1 U7168 ( .B1(n6206), .B2(n6369), .A(n6232), .ZN(n6212) );
  AOI22_X1 U7169 ( .A1(n6209), .A2(n6212), .B1(n6211), .B2(n6295), .ZN(n6207)
         );
  NAND2_X1 U7170 ( .A1(n6208), .A2(n6207), .ZN(n6234) );
  INV_X1 U7171 ( .A(n6209), .ZN(n6213) );
  OAI22_X1 U7172 ( .A1(n6213), .A2(n6212), .B1(n6211), .B2(n6210), .ZN(n6233)
         );
  AOI22_X1 U7173 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6234), .B1(n6243), 
        .B2(n6233), .ZN(n6214) );
  OAI211_X1 U7174 ( .C1(n6302), .C2(n6237), .A(n6215), .B(n6214), .ZN(U3108)
         );
  AOI22_X1 U7175 ( .A1(n6307), .A2(n6232), .B1(n6306), .B2(n6231), .ZN(n6217)
         );
  AOI22_X1 U7176 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6234), .B1(n6256), 
        .B2(n6233), .ZN(n6216) );
  OAI211_X1 U7177 ( .C1(n6309), .C2(n6237), .A(n6217), .B(n6216), .ZN(U3109)
         );
  AOI22_X1 U7178 ( .A1(n6314), .A2(n6232), .B1(n6313), .B2(n6231), .ZN(n6219)
         );
  AOI22_X1 U7179 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6234), .B1(n6259), 
        .B2(n6233), .ZN(n6218) );
  OAI211_X1 U7180 ( .C1(n6316), .C2(n6237), .A(n6219), .B(n6218), .ZN(U3110)
         );
  INV_X1 U7181 ( .A(n6237), .ZN(n6226) );
  AOI22_X1 U7182 ( .A1(n6322), .A2(n6232), .B1(n6226), .B2(n6220), .ZN(n6222)
         );
  AOI22_X1 U7183 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6234), .B1(n6262), 
        .B2(n6233), .ZN(n6221) );
  OAI211_X1 U7184 ( .C1(n6223), .C2(n6284), .A(n6222), .B(n6221), .ZN(U3111)
         );
  AOI22_X1 U7185 ( .A1(n6330), .A2(n6232), .B1(n6226), .B2(n6329), .ZN(n6225)
         );
  AOI22_X1 U7186 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6234), .B1(n6265), 
        .B2(n6233), .ZN(n6224) );
  OAI211_X1 U7187 ( .C1(n6332), .C2(n6284), .A(n6225), .B(n6224), .ZN(U3112)
         );
  AOI22_X1 U7188 ( .A1(n6338), .A2(n6232), .B1(n6226), .B2(n6337), .ZN(n6228)
         );
  AOI22_X1 U7189 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6234), .B1(n6270), 
        .B2(n6233), .ZN(n6227) );
  OAI211_X1 U7190 ( .C1(n6340), .C2(n6284), .A(n6228), .B(n6227), .ZN(U3113)
         );
  AOI22_X1 U7191 ( .A1(n6347), .A2(n6232), .B1(n6348), .B2(n6231), .ZN(n6230)
         );
  AOI22_X1 U7192 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6234), .B1(n6350), 
        .B2(n6233), .ZN(n6229) );
  OAI211_X1 U7193 ( .C1(n6277), .C2(n6237), .A(n6230), .B(n6229), .ZN(U3114)
         );
  AOI22_X1 U7194 ( .A1(n6357), .A2(n6232), .B1(n6355), .B2(n6231), .ZN(n6236)
         );
  AOI22_X1 U7195 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6234), .B1(n6279), 
        .B2(n6233), .ZN(n6235) );
  OAI211_X1 U7196 ( .C1(n6360), .C2(n6237), .A(n6236), .B(n6235), .ZN(U3115)
         );
  NAND3_X1 U7197 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6373), .ZN(n6297) );
  NOR2_X1 U7198 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6297), .ZN(n6280)
         );
  INV_X1 U7199 ( .A(n6238), .ZN(n6242) );
  OAI22_X1 U7200 ( .A1(n6242), .A2(n6241), .B1(n6240), .B2(n6239), .ZN(n6278)
         );
  AOI22_X1 U7201 ( .A1(n6294), .A2(n6280), .B1(n6243), .B2(n6278), .ZN(n6255)
         );
  OR2_X1 U7202 ( .A1(n6244), .A2(n3574), .ZN(n6361) );
  NAND3_X1 U7203 ( .A1(n6284), .A2(n6245), .A3(n6361), .ZN(n6249) );
  INV_X1 U7204 ( .A(n6246), .ZN(n6285) );
  AOI22_X1 U7205 ( .A1(n6249), .A2(n6248), .B1(n6285), .B2(n6247), .ZN(n6253)
         );
  OAI211_X1 U7206 ( .C1(n6280), .C2(n6487), .A(n6251), .B(n6250), .ZN(n6252)
         );
  AOI22_X1 U7207 ( .A1(n6281), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n6293), 
        .B2(n6345), .ZN(n6254) );
  OAI211_X1 U7208 ( .C1(n6302), .C2(n6284), .A(n6255), .B(n6254), .ZN(U3116)
         );
  AOI22_X1 U7209 ( .A1(n6307), .A2(n6280), .B1(n6256), .B2(n6278), .ZN(n6258)
         );
  AOI22_X1 U7210 ( .A1(n6281), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n6306), 
        .B2(n6345), .ZN(n6257) );
  OAI211_X1 U7211 ( .C1(n6309), .C2(n6284), .A(n6258), .B(n6257), .ZN(U3117)
         );
  AOI22_X1 U7212 ( .A1(n6314), .A2(n6280), .B1(n6259), .B2(n6278), .ZN(n6261)
         );
  AOI22_X1 U7213 ( .A1(n6281), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n6313), 
        .B2(n6345), .ZN(n6260) );
  OAI211_X1 U7214 ( .C1(n6316), .C2(n6284), .A(n6261), .B(n6260), .ZN(U3118)
         );
  AOI22_X1 U7215 ( .A1(n6322), .A2(n6280), .B1(n6262), .B2(n6278), .ZN(n6264)
         );
  AOI22_X1 U7216 ( .A1(n6281), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n6321), 
        .B2(n6345), .ZN(n6263) );
  OAI211_X1 U7217 ( .C1(n6324), .C2(n6284), .A(n6264), .B(n6263), .ZN(U3119)
         );
  AOI22_X1 U7218 ( .A1(n6330), .A2(n6280), .B1(n6265), .B2(n6278), .ZN(n6268)
         );
  AOI22_X1 U7219 ( .A1(n6281), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n6266), 
        .B2(n6345), .ZN(n6267) );
  OAI211_X1 U7220 ( .C1(n6269), .C2(n6284), .A(n6268), .B(n6267), .ZN(U3120)
         );
  AOI22_X1 U7221 ( .A1(n6338), .A2(n6280), .B1(n6270), .B2(n6278), .ZN(n6273)
         );
  AOI22_X1 U7222 ( .A1(n6281), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n6271), 
        .B2(n6345), .ZN(n6272) );
  OAI211_X1 U7223 ( .C1(n6274), .C2(n6284), .A(n6273), .B(n6272), .ZN(U3121)
         );
  AOI22_X1 U7224 ( .A1(n6350), .A2(n6278), .B1(n6347), .B2(n6280), .ZN(n6276)
         );
  AOI22_X1 U7225 ( .A1(n6281), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n6348), 
        .B2(n6345), .ZN(n6275) );
  OAI211_X1 U7226 ( .C1(n6277), .C2(n6284), .A(n6276), .B(n6275), .ZN(U3122)
         );
  AOI22_X1 U7227 ( .A1(n6357), .A2(n6280), .B1(n6279), .B2(n6278), .ZN(n6283)
         );
  AOI22_X1 U7228 ( .A1(n6281), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n6355), 
        .B2(n6345), .ZN(n6282) );
  OAI211_X1 U7229 ( .C1(n6360), .C2(n6284), .A(n6283), .B(n6282), .ZN(U3123)
         );
  NAND2_X1 U7230 ( .A1(n6286), .A2(n6285), .ZN(n6289) );
  NOR2_X1 U7231 ( .A1(n6287), .A2(n6297), .ZN(n6356) );
  INV_X1 U7232 ( .A(n6356), .ZN(n6288) );
  NAND2_X1 U7233 ( .A1(n6289), .A2(n6288), .ZN(n6296) );
  NOR3_X1 U7234 ( .A1(n6290), .A2(n6295), .A3(n6296), .ZN(n6292) );
  INV_X1 U7235 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n6605) );
  AOI22_X1 U7236 ( .A1(n6294), .A2(n6356), .B1(n6293), .B2(n6354), .ZN(n6305)
         );
  NAND2_X1 U7237 ( .A1(n6296), .A2(n6245), .ZN(n6300) );
  INV_X1 U7238 ( .A(n6297), .ZN(n6298) );
  NAND2_X1 U7239 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6298), .ZN(n6299) );
  NAND2_X1 U7240 ( .A1(n6300), .A2(n6299), .ZN(n6349) );
  INV_X1 U7241 ( .A(n6349), .ZN(n6359) );
  OAI22_X1 U7242 ( .A1(n6361), .A2(n6302), .B1(n6359), .B2(n6301), .ZN(n6303)
         );
  INV_X1 U7243 ( .A(n6303), .ZN(n6304) );
  OAI211_X1 U7244 ( .C1(n6366), .C2(n6605), .A(n6305), .B(n6304), .ZN(U3124)
         );
  INV_X1 U7245 ( .A(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n6658) );
  AOI22_X1 U7246 ( .A1(n6307), .A2(n6356), .B1(n6306), .B2(n6354), .ZN(n6312)
         );
  OAI22_X1 U7247 ( .A1(n6361), .A2(n6309), .B1(n6359), .B2(n6308), .ZN(n6310)
         );
  INV_X1 U7248 ( .A(n6310), .ZN(n6311) );
  OAI211_X1 U7249 ( .C1(n6366), .C2(n6658), .A(n6312), .B(n6311), .ZN(U3125)
         );
  INV_X1 U7250 ( .A(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n6320) );
  AOI22_X1 U7251 ( .A1(n6314), .A2(n6356), .B1(n6313), .B2(n6354), .ZN(n6319)
         );
  OAI22_X1 U7252 ( .A1(n6361), .A2(n6316), .B1(n6359), .B2(n6315), .ZN(n6317)
         );
  INV_X1 U7253 ( .A(n6317), .ZN(n6318) );
  OAI211_X1 U7254 ( .C1(n6366), .C2(n6320), .A(n6319), .B(n6318), .ZN(U3126)
         );
  INV_X1 U7255 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n6328) );
  AOI22_X1 U7256 ( .A1(n6322), .A2(n6356), .B1(n6321), .B2(n6354), .ZN(n6327)
         );
  OAI22_X1 U7257 ( .A1(n6361), .A2(n6324), .B1(n6359), .B2(n6323), .ZN(n6325)
         );
  INV_X1 U7258 ( .A(n6325), .ZN(n6326) );
  OAI211_X1 U7259 ( .C1(n6366), .C2(n6328), .A(n6327), .B(n6326), .ZN(U3127)
         );
  INV_X1 U7260 ( .A(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n6336) );
  AOI22_X1 U7261 ( .A1(n6330), .A2(n6356), .B1(n6329), .B2(n6345), .ZN(n6335)
         );
  OAI22_X1 U7262 ( .A1(n6341), .A2(n6332), .B1(n6359), .B2(n6331), .ZN(n6333)
         );
  INV_X1 U7263 ( .A(n6333), .ZN(n6334) );
  OAI211_X1 U7264 ( .C1(n6366), .C2(n6336), .A(n6335), .B(n6334), .ZN(U3128)
         );
  AOI22_X1 U7265 ( .A1(n6338), .A2(n6356), .B1(n6337), .B2(n6345), .ZN(n6344)
         );
  OAI22_X1 U7266 ( .A1(n6341), .A2(n6340), .B1(n6359), .B2(n6339), .ZN(n6342)
         );
  INV_X1 U7267 ( .A(n6342), .ZN(n6343) );
  OAI211_X1 U7268 ( .C1(n6366), .C2(n6665), .A(n6344), .B(n6343), .ZN(U3129)
         );
  INV_X1 U7269 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n6353) );
  AOI22_X1 U7270 ( .A1(n6347), .A2(n6356), .B1(n6346), .B2(n6345), .ZN(n6352)
         );
  AOI22_X1 U7271 ( .A1(n6350), .A2(n6349), .B1(n6348), .B2(n6354), .ZN(n6351)
         );
  OAI211_X1 U7272 ( .C1(n6366), .C2(n6353), .A(n6352), .B(n6351), .ZN(U3130)
         );
  INV_X1 U7273 ( .A(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n6365) );
  AOI22_X1 U7274 ( .A1(n6357), .A2(n6356), .B1(n6355), .B2(n6354), .ZN(n6364)
         );
  OAI22_X1 U7275 ( .A1(n6361), .A2(n6360), .B1(n6359), .B2(n6358), .ZN(n6362)
         );
  INV_X1 U7276 ( .A(n6362), .ZN(n6363) );
  OAI211_X1 U7277 ( .C1(n6366), .C2(n6365), .A(n6364), .B(n6363), .ZN(U3131)
         );
  AOI22_X1 U7278 ( .A1(n6369), .A2(n6368), .B1(n6367), .B2(n3114), .ZN(n6489)
         );
  NAND2_X1 U7279 ( .A1(n6370), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6495) );
  NAND3_X1 U7280 ( .A1(n6489), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6495), .ZN(n6374) );
  OAI211_X1 U7281 ( .C1(n6374), .C2(n6373), .A(n6372), .B(n6371), .ZN(n6376)
         );
  NAND2_X1 U7282 ( .A1(n6374), .A2(n6373), .ZN(n6375) );
  NAND2_X1 U7283 ( .A1(n6376), .A2(n6375), .ZN(n6377) );
  AOI222_X1 U7284 ( .A1(n6589), .A2(n6378), .B1(n6589), .B2(n6377), .C1(n6378), 
        .C2(n6377), .ZN(n6380) );
  OAI21_X1 U7285 ( .B1(n6380), .B2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n6379), 
        .ZN(n6388) );
  AOI21_X1 U7286 ( .B1(n6380), .B2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6387) );
  NOR2_X1 U7287 ( .A1(FLUSH_REG_SCAN_IN), .A2(MORE_REG_SCAN_IN), .ZN(n6383) );
  OAI211_X1 U7288 ( .C1(n6384), .C2(n6383), .A(n6382), .B(n6381), .ZN(n6385)
         );
  AOI211_X1 U7289 ( .C1(n6388), .C2(n6387), .A(n6386), .B(n6385), .ZN(n6398)
         );
  INV_X1 U7290 ( .A(n6398), .ZN(n6389) );
  OAI22_X1 U7291 ( .A1(n6389), .A2(n6400), .B1(n6599), .B2(n6513), .ZN(n6390)
         );
  OAI21_X1 U7292 ( .B1(n6392), .B2(n6391), .A(n6390), .ZN(n6486) );
  OAI21_X1 U7293 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6599), .A(n6486), .ZN(
        n6399) );
  AOI221_X1 U7294 ( .B1(n6394), .B2(STATE2_REG_0__SCAN_IN), .C1(n6399), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6393), .ZN(n6397) );
  OAI211_X1 U7295 ( .C1(n6508), .C2(n6395), .A(n6509), .B(n6486), .ZN(n6396)
         );
  OAI211_X1 U7296 ( .C1(n6398), .C2(n6400), .A(n6397), .B(n6396), .ZN(U3148)
         );
  OAI211_X1 U7297 ( .C1(STATE2_REG_0__SCAN_IN), .C2(STATE2_REG_2__SCAN_IN), 
        .A(STATE2_REG_1__SCAN_IN), .B(n6399), .ZN(n6405) );
  OAI21_X1 U7298 ( .B1(READY_N), .B2(n6401), .A(n6400), .ZN(n6403) );
  AOI21_X1 U7299 ( .B1(n6403), .B2(n6486), .A(n6402), .ZN(n6404) );
  NAND2_X1 U7300 ( .A1(n6405), .A2(n6404), .ZN(U3149) );
  OAI221_X1 U7301 ( .B1(STATE2_REG_2__SCAN_IN), .B2(STATE2_REG_0__SCAN_IN), 
        .C1(STATE2_REG_2__SCAN_IN), .C2(n6599), .A(n6485), .ZN(n6407) );
  OAI21_X1 U7302 ( .B1(n6408), .B2(n6407), .A(n6406), .ZN(U3150) );
  AND2_X1 U7303 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6480), .ZN(U3151) );
  AND2_X1 U7304 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6480), .ZN(U3152) );
  AND2_X1 U7305 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6480), .ZN(U3153) );
  AND2_X1 U7306 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6480), .ZN(U3154) );
  AND2_X1 U7307 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6480), .ZN(U3155) );
  AND2_X1 U7308 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6480), .ZN(U3156) );
  AND2_X1 U7309 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6480), .ZN(U3157) );
  AND2_X1 U7310 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6480), .ZN(U3158) );
  AND2_X1 U7311 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6480), .ZN(U3159) );
  AND2_X1 U7312 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6480), .ZN(U3160) );
  AND2_X1 U7313 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6480), .ZN(U3161) );
  AND2_X1 U7314 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6480), .ZN(U3162) );
  AND2_X1 U7315 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6480), .ZN(U3163) );
  AND2_X1 U7316 ( .A1(n6480), .A2(DATAWIDTH_REG_18__SCAN_IN), .ZN(U3164) );
  AND2_X1 U7317 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6480), .ZN(U3165) );
  AND2_X1 U7318 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6480), .ZN(U3166) );
  AND2_X1 U7319 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6480), .ZN(U3167) );
  AND2_X1 U7320 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6480), .ZN(U3168) );
  AND2_X1 U7321 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6480), .ZN(U3169) );
  AND2_X1 U7322 ( .A1(n6480), .A2(DATAWIDTH_REG_12__SCAN_IN), .ZN(U3170) );
  AND2_X1 U7323 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6480), .ZN(U3171) );
  AND2_X1 U7324 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6480), .ZN(U3172) );
  AND2_X1 U7325 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6480), .ZN(U3173) );
  AND2_X1 U7326 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6480), .ZN(U3174) );
  AND2_X1 U7327 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6480), .ZN(U3175) );
  AND2_X1 U7328 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6480), .ZN(U3176) );
  AND2_X1 U7329 ( .A1(n6480), .A2(DATAWIDTH_REG_5__SCAN_IN), .ZN(U3177) );
  AND2_X1 U7330 ( .A1(n6480), .A2(DATAWIDTH_REG_4__SCAN_IN), .ZN(U3178) );
  AND2_X1 U7331 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6480), .ZN(U3179) );
  AND2_X1 U7332 ( .A1(n6480), .A2(DATAWIDTH_REG_2__SCAN_IN), .ZN(U3180) );
  NOR2_X1 U7333 ( .A1(n6598), .A2(n6428), .ZN(n6423) );
  NOR2_X1 U7334 ( .A1(n6599), .A2(n6598), .ZN(n6416) );
  AOI21_X1 U7335 ( .B1(HOLD), .B2(STATE_REG_2__SCAN_IN), .A(n6416), .ZN(n6427)
         );
  OAI21_X1 U7336 ( .B1(NA_N), .B2(n6428), .A(n6420), .ZN(n6422) );
  INV_X1 U7337 ( .A(HOLD), .ZN(n6419) );
  NOR2_X1 U7338 ( .A1(n6598), .A2(n6419), .ZN(n6411) );
  INV_X1 U7339 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6409) );
  OAI21_X1 U7340 ( .B1(n6411), .B2(n6409), .A(n6505), .ZN(n6410) );
  OAI221_X1 U7341 ( .B1(n6423), .B2(n6427), .C1(n6423), .C2(n6422), .A(n6410), 
        .ZN(U3181) );
  NOR2_X1 U7342 ( .A1(n6428), .A2(n6419), .ZN(n6415) );
  AOI21_X1 U7343 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(STATE_REG_0__SCAN_IN), 
        .A(n6411), .ZN(n6414) );
  INV_X1 U7344 ( .A(n6416), .ZN(n6412) );
  OAI211_X1 U7345 ( .C1(n6415), .C2(n6414), .A(n6413), .B(n6412), .ZN(U3182)
         );
  INV_X1 U7346 ( .A(n6423), .ZN(n6426) );
  INV_X1 U7347 ( .A(NA_N), .ZN(n6417) );
  NAND4_X1 U7348 ( .A1(REQUESTPENDING_REG_SCAN_IN), .A2(STATE_REG_0__SCAN_IN), 
        .A3(n6416), .A4(n6417), .ZN(n6425) );
  AOI21_X1 U7349 ( .B1(READY_N), .B2(n6417), .A(n6598), .ZN(n6418) );
  AOI211_X1 U7350 ( .C1(n6428), .C2(REQUESTPENDING_REG_SCAN_IN), .A(n6419), 
        .B(n6418), .ZN(n6421) );
  OAI22_X1 U7351 ( .A1(n6423), .A2(n6422), .B1(n6421), .B2(n6420), .ZN(n6424)
         );
  OAI211_X1 U7352 ( .C1(n6427), .C2(n6426), .A(n6425), .B(n6424), .ZN(U3183)
         );
  NAND2_X1 U7353 ( .A1(n6516), .A2(n6428), .ZN(n6477) );
  NOR2_X2 U7354 ( .A1(n6428), .A2(n6505), .ZN(n6475) );
  AOI22_X1 U7355 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6475), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6505), .ZN(n6429) );
  OAI21_X1 U7356 ( .B1(n6633), .B2(n6477), .A(n6429), .ZN(U3184) );
  AOI22_X1 U7357 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6475), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6505), .ZN(n6430) );
  OAI21_X1 U7358 ( .B1(n6431), .B2(n6477), .A(n6430), .ZN(U3185) );
  AOI22_X1 U7359 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6475), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6505), .ZN(n6432) );
  OAI21_X1 U7360 ( .B1(n6433), .B2(n6477), .A(n6432), .ZN(U3186) );
  AOI22_X1 U7361 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6475), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6505), .ZN(n6434) );
  OAI21_X1 U7362 ( .B1(n6436), .B2(n6477), .A(n6434), .ZN(U3187) );
  AOI22_X1 U7363 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6471), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6505), .ZN(n6435) );
  OAI21_X1 U7364 ( .B1(n6436), .B2(n6473), .A(n6435), .ZN(U3188) );
  AOI22_X1 U7365 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6471), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6505), .ZN(n6437) );
  OAI21_X1 U7366 ( .B1(n4950), .B2(n6473), .A(n6437), .ZN(U3189) );
  AOI22_X1 U7367 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6475), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6505), .ZN(n6438) );
  OAI21_X1 U7368 ( .B1(n6439), .B2(n6477), .A(n6438), .ZN(U3190) );
  AOI22_X1 U7369 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6475), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6505), .ZN(n6440) );
  OAI21_X1 U7370 ( .B1(n6442), .B2(n6477), .A(n6440), .ZN(U3191) );
  AOI22_X1 U7371 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6471), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6505), .ZN(n6441) );
  OAI21_X1 U7372 ( .B1(n6442), .B2(n6473), .A(n6441), .ZN(U3192) );
  AOI22_X1 U7373 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6475), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6505), .ZN(n6443) );
  OAI21_X1 U7374 ( .B1(n6445), .B2(n6477), .A(n6443), .ZN(U3193) );
  AOI22_X1 U7375 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6471), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6505), .ZN(n6444) );
  OAI21_X1 U7376 ( .B1(n6445), .B2(n6473), .A(n6444), .ZN(U3194) );
  AOI22_X1 U7377 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6475), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6505), .ZN(n6446) );
  OAI21_X1 U7378 ( .B1(n6607), .B2(n6477), .A(n6446), .ZN(U3195) );
  AOI22_X1 U7379 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6471), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6505), .ZN(n6447) );
  OAI21_X1 U7380 ( .B1(n6607), .B2(n6473), .A(n6447), .ZN(U3196) );
  AOI22_X1 U7381 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6471), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6505), .ZN(n6448) );
  OAI21_X1 U7382 ( .B1(n6449), .B2(n6473), .A(n6448), .ZN(U3197) );
  AOI22_X1 U7383 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6475), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6505), .ZN(n6450) );
  OAI21_X1 U7384 ( .B1(n6452), .B2(n6477), .A(n6450), .ZN(U3198) );
  AOI22_X1 U7385 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6471), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6505), .ZN(n6451) );
  OAI21_X1 U7386 ( .B1(n6452), .B2(n6473), .A(n6451), .ZN(U3199) );
  INV_X1 U7387 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6455) );
  AOI22_X1 U7388 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6475), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6505), .ZN(n6453) );
  OAI21_X1 U7389 ( .B1(n6455), .B2(n6477), .A(n6453), .ZN(U3200) );
  AOI22_X1 U7390 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6471), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6505), .ZN(n6454) );
  OAI21_X1 U7391 ( .B1(n6455), .B2(n6473), .A(n6454), .ZN(U3201) );
  AOI22_X1 U7392 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6475), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6505), .ZN(n6456) );
  OAI21_X1 U7393 ( .B1(n6458), .B2(n6477), .A(n6456), .ZN(U3202) );
  AOI22_X1 U7394 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6471), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6505), .ZN(n6457) );
  OAI21_X1 U7395 ( .B1(n6458), .B2(n6473), .A(n6457), .ZN(U3203) );
  INV_X1 U7396 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6460) );
  AOI22_X1 U7397 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6471), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6505), .ZN(n6459) );
  OAI21_X1 U7398 ( .B1(n6460), .B2(n6473), .A(n6459), .ZN(U3204) );
  INV_X1 U7399 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6673) );
  AOI22_X1 U7400 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6475), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6505), .ZN(n6461) );
  OAI21_X1 U7401 ( .B1(n6673), .B2(n6477), .A(n6461), .ZN(U3205) );
  AOI22_X1 U7402 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6475), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6505), .ZN(n6462) );
  OAI21_X1 U7403 ( .B1(n4092), .B2(n6477), .A(n6462), .ZN(U3206) );
  AOI22_X1 U7404 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6471), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6505), .ZN(n6463) );
  OAI21_X1 U7405 ( .B1(n4092), .B2(n6473), .A(n6463), .ZN(U3207) );
  AOI22_X1 U7406 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6471), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6505), .ZN(n6464) );
  OAI21_X1 U7407 ( .B1(n6465), .B2(n6473), .A(n6464), .ZN(U3208) );
  AOI22_X1 U7408 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6475), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6505), .ZN(n6466) );
  OAI21_X1 U7409 ( .B1(n6468), .B2(n6477), .A(n6466), .ZN(U3209) );
  AOI22_X1 U7410 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6471), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6505), .ZN(n6467) );
  OAI21_X1 U7411 ( .B1(n6468), .B2(n6473), .A(n6467), .ZN(U3210) );
  AOI22_X1 U7412 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6471), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6505), .ZN(n6469) );
  OAI21_X1 U7413 ( .B1(n6470), .B2(n6473), .A(n6469), .ZN(U3211) );
  AOI22_X1 U7414 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6471), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6505), .ZN(n6472) );
  OAI21_X1 U7415 ( .B1(n6474), .B2(n6473), .A(n6472), .ZN(U3212) );
  INV_X1 U7416 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6478) );
  AOI22_X1 U7417 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6475), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6505), .ZN(n6476) );
  OAI21_X1 U7418 ( .B1(n6478), .B2(n6477), .A(n6476), .ZN(U3213) );
  MUX2_X1 U7419 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6516), .Z(U3445) );
  MUX2_X1 U7420 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6516), .Z(U3446) );
  MUX2_X1 U7421 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6516), .Z(U3447) );
  MUX2_X1 U7422 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6516), .Z(U3448) );
  INV_X1 U7423 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6481) );
  INV_X1 U7424 ( .A(n6482), .ZN(n6479) );
  AOI21_X1 U7425 ( .B1(n6481), .B2(n6480), .A(n6479), .ZN(U3451) );
  OAI21_X1 U7426 ( .B1(n6484), .B2(n6483), .A(n6482), .ZN(U3452) );
  OAI221_X1 U7427 ( .B1(n6487), .B2(STATE2_REG_0__SCAN_IN), .C1(n6487), .C2(
        n6486), .A(n6485), .ZN(U3453) );
  OAI22_X1 U7428 ( .A1(n6489), .A2(n6494), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n6488), .ZN(n6492) );
  OAI22_X1 U7429 ( .A1(n6492), .A2(n6491), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6490), .ZN(n6493) );
  OAI21_X1 U7430 ( .B1(n6495), .B2(n6494), .A(n6493), .ZN(U3461) );
  AOI21_X1 U7431 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6497) );
  AOI22_X1 U7432 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6497), .B2(n6496), .ZN(n6500) );
  INV_X1 U7433 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6499) );
  AOI22_X1 U7434 ( .A1(n6503), .A2(n6500), .B1(n6499), .B2(n6498), .ZN(U3468)
         );
  INV_X1 U7435 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6502) );
  OAI21_X1 U7436 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6503), .ZN(n6501) );
  OAI21_X1 U7437 ( .B1(n6503), .B2(n6502), .A(n6501), .ZN(U3469) );
  NAND2_X1 U7438 ( .A1(n6505), .A2(W_R_N_REG_SCAN_IN), .ZN(n6504) );
  OAI21_X1 U7439 ( .B1(n6505), .B2(READREQUEST_REG_SCAN_IN), .A(n6504), .ZN(
        U3470) );
  AOI211_X1 U7440 ( .C1(n6507), .C2(n6638), .A(n6210), .B(n6506), .ZN(n6510)
         );
  OAI21_X1 U7441 ( .B1(n6510), .B2(n6509), .A(n6508), .ZN(n6515) );
  OAI211_X1 U7442 ( .C1(READY_N), .C2(n6513), .A(n6512), .B(n6511), .ZN(n6514)
         );
  MUX2_X1 U7443 ( .A(REQUESTPENDING_REG_SCAN_IN), .B(n6515), .S(n6514), .Z(
        U3472) );
  MUX2_X1 U7444 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6516), .Z(U3473) );
  AOI222_X1 U7445 ( .A1(n6520), .A2(n6519), .B1(n3006), .B2(n6518), .C1(n6517), 
        .C2(EBX_REG_25__SCAN_IN), .ZN(n6687) );
  NOR2_X1 U7446 ( .A1(keyinput16), .A2(keyinput36), .ZN(n6521) );
  NAND3_X1 U7447 ( .A1(keyinput27), .A2(keyinput58), .A3(n6521), .ZN(n6526) );
  NAND3_X1 U7448 ( .A1(keyinput20), .A2(keyinput24), .A3(keyinput39), .ZN(
        n6525) );
  NOR2_X1 U7449 ( .A1(keyinput22), .A2(keyinput46), .ZN(n6523) );
  NOR4_X1 U7450 ( .A1(keyinput8), .A2(keyinput26), .A3(keyinput32), .A4(
        keyinput49), .ZN(n6522) );
  NAND4_X1 U7451 ( .A1(keyinput10), .A2(keyinput59), .A3(n6523), .A4(n6522), 
        .ZN(n6524) );
  NOR4_X1 U7452 ( .A1(keyinput21), .A2(n6526), .A3(n6525), .A4(n6524), .ZN(
        n6685) );
  NAND3_X1 U7453 ( .A1(keyinput47), .A2(keyinput54), .A3(keyinput55), .ZN(
        n6548) );
  NOR3_X1 U7454 ( .A1(keyinput0), .A2(keyinput40), .A3(keyinput33), .ZN(n6531)
         );
  NAND2_X1 U7455 ( .A1(keyinput13), .A2(keyinput45), .ZN(n6527) );
  NOR3_X1 U7456 ( .A1(keyinput29), .A2(keyinput42), .A3(n6527), .ZN(n6530) );
  NAND2_X1 U7457 ( .A1(keyinput12), .A2(keyinput15), .ZN(n6528) );
  NOR3_X1 U7458 ( .A1(keyinput30), .A2(keyinput44), .A3(n6528), .ZN(n6529) );
  NAND4_X1 U7459 ( .A1(keyinput31), .A2(n6531), .A3(n6530), .A4(n6529), .ZN(
        n6547) );
  INV_X1 U7460 ( .A(keyinput1), .ZN(n6532) );
  NOR3_X1 U7461 ( .A1(keyinput7), .A2(keyinput56), .A3(n6532), .ZN(n6545) );
  NAND2_X1 U7462 ( .A1(keyinput34), .A2(keyinput37), .ZN(n6536) );
  NOR3_X1 U7463 ( .A1(keyinput3), .A2(keyinput19), .A3(keyinput28), .ZN(n6534)
         );
  NOR3_X1 U7464 ( .A1(keyinput35), .A2(keyinput53), .A3(keyinput18), .ZN(n6533) );
  NAND4_X1 U7465 ( .A1(keyinput9), .A2(n6534), .A3(keyinput5), .A4(n6533), 
        .ZN(n6535) );
  NOR4_X1 U7466 ( .A1(keyinput63), .A2(keyinput11), .A3(n6536), .A4(n6535), 
        .ZN(n6544) );
  NAND2_X1 U7467 ( .A1(keyinput50), .A2(keyinput23), .ZN(n6542) );
  NOR2_X1 U7468 ( .A1(keyinput4), .A2(keyinput51), .ZN(n6540) );
  NAND3_X1 U7469 ( .A1(keyinput25), .A2(keyinput41), .A3(keyinput57), .ZN(
        n6538) );
  INV_X1 U7470 ( .A(keyinput61), .ZN(n6657) );
  NAND3_X1 U7471 ( .A1(keyinput14), .A2(keyinput2), .A3(n6657), .ZN(n6537) );
  NOR4_X1 U7472 ( .A1(keyinput17), .A2(keyinput6), .A3(n6538), .A4(n6537), 
        .ZN(n6539) );
  NAND4_X1 U7473 ( .A1(keyinput62), .A2(keyinput60), .A3(n6540), .A4(n6539), 
        .ZN(n6541) );
  NOR4_X1 U7474 ( .A1(keyinput52), .A2(keyinput43), .A3(n6542), .A4(n6541), 
        .ZN(n6543) );
  NAND4_X1 U7475 ( .A1(keyinput48), .A2(n6545), .A3(n6544), .A4(n6543), .ZN(
        n6546) );
  NOR4_X1 U7476 ( .A1(keyinput38), .A2(n6548), .A3(n6547), .A4(n6546), .ZN(
        n6684) );
  INV_X1 U7477 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n6551) );
  AOI22_X1 U7478 ( .A1(n6551), .A2(keyinput27), .B1(keyinput36), .B2(n6550), 
        .ZN(n6549) );
  OAI221_X1 U7479 ( .B1(n6551), .B2(keyinput27), .C1(n6550), .C2(keyinput36), 
        .A(n6549), .ZN(n6564) );
  INV_X1 U7480 ( .A(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n6554) );
  AOI22_X1 U7481 ( .A1(n6554), .A2(keyinput16), .B1(keyinput58), .B2(n6553), 
        .ZN(n6552) );
  OAI221_X1 U7482 ( .B1(n6554), .B2(keyinput16), .C1(n6553), .C2(keyinput58), 
        .A(n6552), .ZN(n6563) );
  INV_X1 U7483 ( .A(keyinput24), .ZN(n6556) );
  AOI22_X1 U7484 ( .A1(n6557), .A2(keyinput20), .B1(DATAWIDTH_REG_12__SCAN_IN), 
        .B2(n6556), .ZN(n6555) );
  OAI221_X1 U7485 ( .B1(n6557), .B2(keyinput20), .C1(n6556), .C2(
        DATAWIDTH_REG_12__SCAN_IN), .A(n6555), .ZN(n6562) );
  INV_X1 U7486 ( .A(keyinput39), .ZN(n6559) );
  AOI22_X1 U7487 ( .A1(n6560), .A2(keyinput21), .B1(UWORD_REG_12__SCAN_IN), 
        .B2(n6559), .ZN(n6558) );
  OAI221_X1 U7488 ( .B1(n6560), .B2(keyinput21), .C1(n6559), .C2(
        UWORD_REG_12__SCAN_IN), .A(n6558), .ZN(n6561) );
  NOR4_X1 U7489 ( .A1(n6564), .A2(n6563), .A3(n6562), .A4(n6561), .ZN(n6616)
         );
  INV_X1 U7490 ( .A(keyinput22), .ZN(n6567) );
  INV_X1 U7491 ( .A(keyinput46), .ZN(n6566) );
  AOI22_X1 U7492 ( .A1(n6567), .A2(DATAO_REG_16__SCAN_IN), .B1(
        DATAWIDTH_REG_5__SCAN_IN), .B2(n6566), .ZN(n6565) );
  OAI221_X1 U7493 ( .B1(n6567), .B2(DATAO_REG_16__SCAN_IN), .C1(n6566), .C2(
        DATAWIDTH_REG_5__SCAN_IN), .A(n6565), .ZN(n6580) );
  INV_X1 U7494 ( .A(keyinput10), .ZN(n6569) );
  AOI22_X1 U7495 ( .A1(n6570), .A2(keyinput59), .B1(DATAO_REG_18__SCAN_IN), 
        .B2(n6569), .ZN(n6568) );
  OAI221_X1 U7496 ( .B1(n6570), .B2(keyinput59), .C1(n6569), .C2(
        DATAO_REG_18__SCAN_IN), .A(n6568), .ZN(n6579) );
  INV_X1 U7497 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6573) );
  INV_X1 U7498 ( .A(keyinput8), .ZN(n6572) );
  AOI22_X1 U7499 ( .A1(n6573), .A2(keyinput26), .B1(DATAWIDTH_REG_4__SCAN_IN), 
        .B2(n6572), .ZN(n6571) );
  OAI221_X1 U7500 ( .B1(n6573), .B2(keyinput26), .C1(n6572), .C2(
        DATAWIDTH_REG_4__SCAN_IN), .A(n6571), .ZN(n6578) );
  INV_X1 U7501 ( .A(keyinput32), .ZN(n6575) );
  AOI22_X1 U7502 ( .A1(n6576), .A2(keyinput49), .B1(REQUESTPENDING_REG_SCAN_IN), .B2(n6575), .ZN(n6574) );
  OAI221_X1 U7503 ( .B1(n6576), .B2(keyinput49), .C1(n6575), .C2(
        REQUESTPENDING_REG_SCAN_IN), .A(n6574), .ZN(n6577) );
  NOR4_X1 U7504 ( .A1(n6580), .A2(n6579), .A3(n6578), .A4(n6577), .ZN(n6615)
         );
  INV_X1 U7505 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n6583) );
  INV_X1 U7506 ( .A(keyinput31), .ZN(n6582) );
  AOI22_X1 U7507 ( .A1(n6583), .A2(keyinput0), .B1(DATAWIDTH_REG_18__SCAN_IN), 
        .B2(n6582), .ZN(n6581) );
  OAI221_X1 U7508 ( .B1(n6583), .B2(keyinput0), .C1(n6582), .C2(
        DATAWIDTH_REG_18__SCAN_IN), .A(n6581), .ZN(n6596) );
  INV_X1 U7509 ( .A(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n6586) );
  INV_X1 U7510 ( .A(keyinput33), .ZN(n6585) );
  AOI22_X1 U7511 ( .A1(n6586), .A2(keyinput40), .B1(BYTEENABLE_REG_0__SCAN_IN), 
        .B2(n6585), .ZN(n6584) );
  OAI221_X1 U7512 ( .B1(n6586), .B2(keyinput40), .C1(n6585), .C2(
        BYTEENABLE_REG_0__SCAN_IN), .A(n6584), .ZN(n6595) );
  INV_X1 U7513 ( .A(keyinput38), .ZN(n6588) );
  AOI22_X1 U7514 ( .A1(n6589), .A2(keyinput47), .B1(DATAI_26_), .B2(n6588), 
        .ZN(n6587) );
  OAI221_X1 U7515 ( .B1(n6589), .B2(keyinput47), .C1(n6588), .C2(DATAI_26_), 
        .A(n6587), .ZN(n6594) );
  INV_X1 U7516 ( .A(keyinput54), .ZN(n6592) );
  INV_X1 U7517 ( .A(keyinput55), .ZN(n6591) );
  AOI22_X1 U7518 ( .A1(n6592), .A2(ADDRESS_REG_9__SCAN_IN), .B1(
        LWORD_REG_1__SCAN_IN), .B2(n6591), .ZN(n6590) );
  OAI221_X1 U7519 ( .B1(n6592), .B2(ADDRESS_REG_9__SCAN_IN), .C1(n6591), .C2(
        LWORD_REG_1__SCAN_IN), .A(n6590), .ZN(n6593) );
  NOR4_X1 U7520 ( .A1(n6596), .A2(n6595), .A3(n6594), .A4(n6593), .ZN(n6614)
         );
  AOI22_X1 U7521 ( .A1(n6599), .A2(keyinput29), .B1(keyinput45), .B2(n6598), 
        .ZN(n6597) );
  OAI221_X1 U7522 ( .B1(n6599), .B2(keyinput29), .C1(n6598), .C2(keyinput45), 
        .A(n6597), .ZN(n6612) );
  AOI22_X1 U7523 ( .A1(n6602), .A2(keyinput13), .B1(keyinput42), .B2(n6601), 
        .ZN(n6600) );
  OAI221_X1 U7524 ( .B1(n6602), .B2(keyinput13), .C1(n6601), .C2(keyinput42), 
        .A(n6600), .ZN(n6611) );
  INV_X1 U7525 ( .A(keyinput15), .ZN(n6604) );
  AOI22_X1 U7526 ( .A1(n6605), .A2(keyinput44), .B1(DATAI_3_), .B2(n6604), 
        .ZN(n6603) );
  OAI221_X1 U7527 ( .B1(n6605), .B2(keyinput44), .C1(n6604), .C2(DATAI_3_), 
        .A(n6603), .ZN(n6610) );
  INV_X1 U7528 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n6608) );
  AOI22_X1 U7529 ( .A1(n6608), .A2(keyinput30), .B1(keyinput12), .B2(n6607), 
        .ZN(n6606) );
  OAI221_X1 U7530 ( .B1(n6608), .B2(keyinput30), .C1(n6607), .C2(keyinput12), 
        .A(n6606), .ZN(n6609) );
  NOR4_X1 U7531 ( .A1(n6612), .A2(n6611), .A3(n6610), .A4(n6609), .ZN(n6613)
         );
  NAND4_X1 U7532 ( .A1(n6616), .A2(n6615), .A3(n6614), .A4(n6613), .ZN(n6683)
         );
  INV_X1 U7533 ( .A(keyinput19), .ZN(n6618) );
  AOI22_X1 U7534 ( .A1(n5078), .A2(keyinput28), .B1(REIP_REG_0__SCAN_IN), .B2(
        n6618), .ZN(n6617) );
  OAI221_X1 U7535 ( .B1(n5078), .B2(keyinput28), .C1(n6618), .C2(
        REIP_REG_0__SCAN_IN), .A(n6617), .ZN(n6631) );
  INV_X1 U7536 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n6620) );
  AOI22_X1 U7537 ( .A1(n6621), .A2(keyinput9), .B1(n6620), .B2(keyinput3), 
        .ZN(n6619) );
  OAI221_X1 U7538 ( .B1(n6621), .B2(keyinput9), .C1(n6620), .C2(keyinput3), 
        .A(n6619), .ZN(n6630) );
  INV_X1 U7539 ( .A(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n6624) );
  INV_X1 U7540 ( .A(keyinput53), .ZN(n6623) );
  AOI22_X1 U7541 ( .A1(n6624), .A2(keyinput18), .B1(DATAO_REG_8__SCAN_IN), 
        .B2(n6623), .ZN(n6622) );
  OAI221_X1 U7542 ( .B1(n6624), .B2(keyinput18), .C1(n6623), .C2(
        DATAO_REG_8__SCAN_IN), .A(n6622), .ZN(n6629) );
  INV_X1 U7543 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n6627) );
  AOI22_X1 U7544 ( .A1(n6627), .A2(keyinput35), .B1(keyinput5), .B2(n6626), 
        .ZN(n6625) );
  OAI221_X1 U7545 ( .B1(n6627), .B2(keyinput35), .C1(n6626), .C2(keyinput5), 
        .A(n6625), .ZN(n6628) );
  NOR4_X1 U7546 ( .A1(n6631), .A2(n6630), .A3(n6629), .A4(n6628), .ZN(n6681)
         );
  AOI22_X1 U7547 ( .A1(n6634), .A2(keyinput56), .B1(keyinput1), .B2(n6633), 
        .ZN(n6632) );
  OAI221_X1 U7548 ( .B1(n6634), .B2(keyinput56), .C1(n6633), .C2(keyinput1), 
        .A(n6632), .ZN(n6646) );
  AOI22_X1 U7549 ( .A1(n3761), .A2(keyinput7), .B1(n6636), .B2(keyinput48), 
        .ZN(n6635) );
  OAI221_X1 U7550 ( .B1(n3761), .B2(keyinput7), .C1(n6636), .C2(keyinput48), 
        .A(n6635), .ZN(n6645) );
  AOI22_X1 U7551 ( .A1(n6639), .A2(keyinput37), .B1(keyinput11), .B2(n6638), 
        .ZN(n6637) );
  OAI221_X1 U7552 ( .B1(n6639), .B2(keyinput37), .C1(n6638), .C2(keyinput11), 
        .A(n6637), .ZN(n6644) );
  INV_X1 U7553 ( .A(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n6642) );
  INV_X1 U7554 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n6641) );
  AOI22_X1 U7555 ( .A1(n6642), .A2(keyinput34), .B1(n6641), .B2(keyinput63), 
        .ZN(n6640) );
  OAI221_X1 U7556 ( .B1(n6642), .B2(keyinput34), .C1(n6641), .C2(keyinput63), 
        .A(n6640), .ZN(n6643) );
  NOR4_X1 U7557 ( .A1(n6646), .A2(n6645), .A3(n6644), .A4(n6643), .ZN(n6680)
         );
  INV_X1 U7558 ( .A(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n6649) );
  INV_X1 U7559 ( .A(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n6648) );
  AOI22_X1 U7560 ( .A1(n6649), .A2(keyinput51), .B1(keyinput60), .B2(n6648), 
        .ZN(n6647) );
  OAI221_X1 U7561 ( .B1(n6649), .B2(keyinput51), .C1(n6648), .C2(keyinput60), 
        .A(n6647), .ZN(n6662) );
  INV_X1 U7562 ( .A(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n6652) );
  INV_X1 U7563 ( .A(keyinput4), .ZN(n6651) );
  AOI22_X1 U7564 ( .A1(n6652), .A2(keyinput62), .B1(DATAWIDTH_REG_2__SCAN_IN), 
        .B2(n6651), .ZN(n6650) );
  OAI221_X1 U7565 ( .B1(n6652), .B2(keyinput62), .C1(n6651), .C2(
        DATAWIDTH_REG_2__SCAN_IN), .A(n6650), .ZN(n6661) );
  INV_X1 U7566 ( .A(keyinput2), .ZN(n6654) );
  AOI22_X1 U7567 ( .A1(n6655), .A2(keyinput14), .B1(UWORD_REG_10__SCAN_IN), 
        .B2(n6654), .ZN(n6653) );
  OAI221_X1 U7568 ( .B1(n6655), .B2(keyinput14), .C1(n6654), .C2(
        UWORD_REG_10__SCAN_IN), .A(n6653), .ZN(n6660) );
  AOI22_X1 U7569 ( .A1(n6658), .A2(keyinput6), .B1(UWORD_REG_3__SCAN_IN), .B2(
        n6657), .ZN(n6656) );
  OAI221_X1 U7570 ( .B1(n6658), .B2(keyinput6), .C1(n6657), .C2(
        UWORD_REG_3__SCAN_IN), .A(n6656), .ZN(n6659) );
  NOR4_X1 U7571 ( .A1(n6662), .A2(n6661), .A3(n6660), .A4(n6659), .ZN(n6679)
         );
  AOI22_X1 U7572 ( .A1(n6665), .A2(keyinput57), .B1(keyinput17), .B2(n6664), 
        .ZN(n6663) );
  OAI221_X1 U7573 ( .B1(n6665), .B2(keyinput57), .C1(n6664), .C2(keyinput17), 
        .A(n6663), .ZN(n6677) );
  AOI22_X1 U7574 ( .A1(n6668), .A2(keyinput25), .B1(n6667), .B2(keyinput41), 
        .ZN(n6666) );
  OAI221_X1 U7575 ( .B1(n6668), .B2(keyinput25), .C1(n6667), .C2(keyinput41), 
        .A(n6666), .ZN(n6676) );
  INV_X1 U7576 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n6671) );
  INV_X1 U7577 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n6670) );
  AOI22_X1 U7578 ( .A1(n6671), .A2(keyinput43), .B1(keyinput23), .B2(n6670), 
        .ZN(n6669) );
  OAI221_X1 U7579 ( .B1(n6671), .B2(keyinput43), .C1(n6670), .C2(keyinput23), 
        .A(n6669), .ZN(n6675) );
  AOI22_X1 U7580 ( .A1(n4092), .A2(keyinput52), .B1(keyinput50), .B2(n6673), 
        .ZN(n6672) );
  OAI221_X1 U7581 ( .B1(n4092), .B2(keyinput52), .C1(n6673), .C2(keyinput50), 
        .A(n6672), .ZN(n6674) );
  NOR4_X1 U7582 ( .A1(n6677), .A2(n6676), .A3(n6675), .A4(n6674), .ZN(n6678)
         );
  NAND4_X1 U7583 ( .A1(n6681), .A2(n6680), .A3(n6679), .A4(n6678), .ZN(n6682)
         );
  AOI211_X1 U7584 ( .C1(n6685), .C2(n6684), .A(n6683), .B(n6682), .ZN(n6686)
         );
  XNOR2_X1 U7585 ( .A(n6687), .B(n6686), .ZN(U2834) );
  CLKBUF_X1 U3438 ( .A(n3302), .Z(n4020) );
  CLKBUF_X1 U34530 ( .A(n5167), .Z(n5310) );
  OR2_X1 U3704 ( .A1(n5476), .A2(n4256), .ZN(n5465) );
  AOI211_X2 U5246 ( .C1(n6295), .C2(n6297), .A(n6292), .B(n6291), .ZN(n6366)
         );
endmodule

