

module b15_C_gen_AntiSAT_k_256_2 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, 
        keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, 
        keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, 
        keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, 
        keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, 
        keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, 
        keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, 
        keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101, 
        keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105, 
        keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109, 
        keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113, 
        keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117, 
        keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121, 
        keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125, 
        keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67, 
        keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72, 
        keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77, 
        keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82, 
        keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87, 
        keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92, 
        keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97, 
        keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, U3445, U3446, U3447, U3448, U3213, U3212, 
        U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, 
        U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, 
        U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, 
        U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, 
        U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, 
        U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, 
        U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, 
        U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, 
        U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, 
        U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, 
        U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, 
        U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, 
        U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, 
        U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, 
        U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, 
        U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, 
        U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, 
        U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, 
        U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, 
        U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, 
        U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, 
        U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, 
        U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, 
        U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, 
        U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, 
        U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, 
        U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, 
        U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, 
        U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, 
        U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, 
        U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, 
        U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, 
        U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, 
        U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, 
        U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, 
        U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, 
        U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, 
        U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, 
        U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, 
        U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, 
        U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, 
        U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, 
        U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, 
        U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, 
        U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1,
         keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6,
         keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11,
         keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16,
         keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21,
         keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26,
         keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31,
         keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36,
         keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41,
         keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46,
         keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51,
         keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56,
         keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61,
         keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66,
         keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71,
         keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76,
         keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81,
         keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86,
         keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91,
         keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96,
         keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100,
         keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104,
         keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108,
         keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112,
         keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116,
         keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120,
         keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124,
         keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1,
         keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6,
         keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11,
         keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16,
         keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21,
         keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26,
         keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31,
         keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36,
         keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41,
         keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46,
         keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51,
         keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56,
         keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61,
         keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66,
         keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71,
         keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76,
         keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81,
         keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86,
         keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91,
         keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96,
         keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100,
         keyinput_g101, keyinput_g102, keyinput_g103, keyinput_g104,
         keyinput_g105, keyinput_g106, keyinput_g107, keyinput_g108,
         keyinput_g109, keyinput_g110, keyinput_g111, keyinput_g112,
         keyinput_g113, keyinput_g114, keyinput_g115, keyinput_g116,
         keyinput_g117, keyinput_g118, keyinput_g119, keyinput_g120,
         keyinput_g121, keyinput_g122, keyinput_g123, keyinput_g124,
         keyinput_g125, keyinput_g126, keyinput_g127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096;

  AND2_X1 U3606 ( .A1(n4056), .A2(n4608), .ZN(n3404) );
  INV_X2 U3608 ( .A(n3398), .ZN(n4620) );
  AND2_X1 U3609 ( .A1(n5395), .A2(n4545), .ZN(n3421) );
  OR2_X1 U3610 ( .A1(n3539), .A2(n3538), .ZN(n3537) );
  CLKBUF_X2 U3611 ( .A(n3374), .Z(n4028) );
  CLKBUF_X2 U3612 ( .A(n3421), .Z(n3413) );
  NAND2_X1 U3613 ( .A1(n3479), .A2(n3478), .ZN(n3539) );
  AND2_X2 U3614 ( .A1(n4553), .A2(n4545), .ZN(n3351) );
  OR2_X1 U3615 ( .A1(n3405), .A2(n3404), .ZN(n4128) );
  XNOR2_X1 U3616 ( .A(n3539), .B(n3538), .ZN(n3483) );
  AND4_X1 U3617 ( .A1(n3360), .A2(n3359), .A3(n3358), .A4(n3357), .ZN(n3361)
         );
  INV_X1 U3618 ( .A(n4150), .ZN(n5557) );
  AND2_X1 U3619 ( .A1(n4313), .A2(n4312), .ZN(n4314) );
  INV_X1 U3621 ( .A(n3386), .ZN(n4608) );
  INV_X1 U3622 ( .A(n4490), .ZN(n4159) );
  INV_X1 U3623 ( .A(n6162), .ZN(n6150) );
  INV_X1 U3625 ( .A(n6211), .ZN(n6205) );
  INV_X2 U3627 ( .A(n4117), .ZN(n3445) );
  AND4_X2 U3628 ( .A1(n3338), .A2(n3337), .A3(n3336), .A4(n3335), .ZN(n3255)
         );
  NAND2_X2 U3629 ( .A1(n3180), .A2(n3298), .ZN(n3365) );
  AND4_X2 U3630 ( .A1(n3309), .A2(n3310), .A3(n3308), .A4(n3307), .ZN(n3311)
         );
  NOR2_X2 U3631 ( .A1(n4442), .A2(n3158), .ZN(n4410) );
  AND2_X1 U3632 ( .A1(n4553), .A2(n4545), .ZN(n3157) );
  XNOR2_X2 U3633 ( .A(n5766), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4464)
         );
  NAND2_X2 U3634 ( .A1(n5767), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5766)
         );
  OR2_X1 U3635 ( .A1(n3543), .A2(n3542), .ZN(n3544) );
  AND2_X1 U3637 ( .A1(n5608), .A2(n3185), .ZN(n5597) );
  OR2_X1 U3638 ( .A1(n5349), .A2(n3179), .ZN(n5568) );
  OR2_X1 U3639 ( .A1(n5465), .A2(n4232), .ZN(n4235) );
  NAND2_X1 U3640 ( .A1(n4540), .A2(n4585), .ZN(n4584) );
  NOR2_X2 U3641 ( .A1(n4521), .A2(n4539), .ZN(n4540) );
  NAND2_X1 U3642 ( .A1(n5617), .A2(n3191), .ZN(n5834) );
  CLKBUF_X2 U3643 ( .A(n6283), .Z(n6344) );
  NAND2_X1 U3644 ( .A1(n3387), .A2(n4608), .ZN(n4117) );
  NAND2_X2 U3645 ( .A1(n4244), .A2(n3398), .ZN(n4150) );
  INV_X1 U3646 ( .A(n4244), .ZN(n4612) );
  INV_X2 U3647 ( .A(n3436), .ZN(n3158) );
  CLKBUF_X2 U3648 ( .A(n3427), .Z(n4026) );
  BUF_X2 U3649 ( .A(n3407), .Z(n4006) );
  BUF_X2 U3650 ( .A(n3465), .Z(n4034) );
  BUF_X2 U3651 ( .A(n3408), .Z(n4037) );
  BUF_X2 U3652 ( .A(n3471), .Z(n4033) );
  AND2_X1 U3653 ( .A1(n3215), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3273)
         );
  OR2_X1 U3654 ( .A1(n5701), .A2(n4367), .ZN(n4370) );
  OAI211_X1 U3655 ( .C1(n5476), .C2(n6162), .A(n3200), .B(n5474), .ZN(n3199)
         );
  AND2_X1 U3656 ( .A1(n4382), .A2(n4381), .ZN(n5634) );
  AND2_X1 U3657 ( .A1(n4376), .A2(n4375), .ZN(n4377) );
  OAI21_X1 U3658 ( .B1(n5501), .B2(n5487), .A(n4378), .ZN(n5667) );
  CLKBUF_X1 U3659 ( .A(n5486), .Z(n5501) );
  CLKBUF_X1 U3660 ( .A(n5499), .Z(n5500) );
  AND2_X1 U3661 ( .A1(n3163), .A2(n3164), .ZN(n4328) );
  NOR2_X1 U3662 ( .A1(n3249), .A2(n5309), .ZN(n3248) );
  NOR2_X1 U3663 ( .A1(n5256), .A2(n3210), .ZN(n3209) );
  NAND2_X1 U3664 ( .A1(n4288), .A2(n4287), .ZN(n4888) );
  NOR2_X1 U3665 ( .A1(n3253), .A2(n5309), .ZN(n3246) );
  NAND2_X1 U3666 ( .A1(n3243), .A2(n3240), .ZN(n3250) );
  NOR2_X1 U3667 ( .A1(n3251), .A2(n3242), .ZN(n3241) );
  XNOR2_X1 U3668 ( .A(n5468), .B(n3201), .ZN(n5772) );
  INV_X2 U3670 ( .A(n4314), .ZN(n5729) );
  AOI21_X1 U3671 ( .B1(n5467), .B2(n5466), .A(n5465), .ZN(n5468) );
  OR2_X1 U3672 ( .A1(n5467), .A2(n4389), .ZN(n5480) );
  AOI21_X1 U3673 ( .B1(n4289), .B2(n3766), .A(n3646), .ZN(n5013) );
  AND2_X1 U3674 ( .A1(n3620), .A2(n5210), .ZN(n3229) );
  XNOR2_X1 U3675 ( .A(n4313), .B(n3649), .ZN(n4301) );
  AND2_X1 U3676 ( .A1(n4313), .A2(n3640), .ZN(n4289) );
  NAND2_X1 U3677 ( .A1(n3637), .A2(n3636), .ZN(n4313) );
  NOR2_X1 U3678 ( .A1(n6095), .A2(n6109), .ZN(n6079) );
  NOR2_X1 U3679 ( .A1(n6659), .A2(n5411), .ZN(n6113) );
  NOR2_X1 U3680 ( .A1(n6190), .A2(n5275), .ZN(n6123) );
  NAND2_X1 U3681 ( .A1(n3569), .A2(n3568), .ZN(n3577) );
  NAND2_X1 U3682 ( .A1(n5231), .A2(n5230), .ZN(n6190) );
  AND2_X1 U3683 ( .A1(n5471), .A2(n5239), .ZN(n5229) );
  CLKBUF_X1 U3684 ( .A(n4589), .Z(n5902) );
  XNOR2_X1 U3685 ( .A(n4565), .B(n4852), .ZN(n4550) );
  NAND2_X1 U3686 ( .A1(n3532), .A2(n3531), .ZN(n3535) );
  INV_X1 U3687 ( .A(n5240), .ZN(n5471) );
  BUF_X1 U3688 ( .A(n6261), .Z(n6266) );
  NAND2_X1 U3689 ( .A1(n3551), .A2(n3550), .ZN(n4565) );
  NAND2_X1 U3690 ( .A1(n6215), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5240) );
  NOR2_X1 U3691 ( .A1(n6111), .A2(n6112), .ZN(n6110) );
  OR2_X2 U3692 ( .A1(n6690), .A2(n5225), .ZN(n6215) );
  NOR2_X1 U3693 ( .A1(n5213), .A2(n5215), .ZN(n5147) );
  AND2_X2 U3694 ( .A1(n4471), .A2(n4505), .ZN(n4515) );
  AND2_X2 U3695 ( .A1(n4115), .A2(n4114), .ZN(n4471) );
  NAND2_X1 U3696 ( .A1(n4112), .A2(n4111), .ZN(n4115) );
  OR2_X1 U3697 ( .A1(n4103), .A2(n4102), .ZN(n4112) );
  AND2_X1 U3698 ( .A1(n4129), .A2(n4064), .ZN(n4504) );
  INV_X1 U3699 ( .A(n3448), .ZN(n3369) );
  NAND2_X1 U3700 ( .A1(n4490), .A2(n5557), .ZN(n4224) );
  NOR2_X1 U3701 ( .A1(n3420), .A2(n3557), .ZN(n4309) );
  CLKBUF_X1 U3702 ( .A(n4118), .Z(n6271) );
  AND2_X1 U3703 ( .A1(n3444), .A2(n3452), .ZN(n3446) );
  AND2_X1 U3704 ( .A1(n3366), .A2(n4244), .ZN(n3444) );
  NAND2_X1 U3705 ( .A1(n3366), .A2(n3365), .ZN(n4473) );
  OR2_X1 U3706 ( .A1(n3419), .A2(n3418), .ZN(n4315) );
  NAND2_X1 U3707 ( .A1(n3333), .A2(n3332), .ZN(n4465) );
  NAND2_X2 U3708 ( .A1(n3279), .A2(n3278), .ZN(n3366) );
  NAND3_X1 U3709 ( .A1(n3255), .A2(n3263), .A3(n3342), .ZN(n4244) );
  AND2_X1 U3710 ( .A1(n3324), .A2(n3323), .ZN(n3333) );
  AND4_X1 U3711 ( .A1(n3346), .A2(n3345), .A3(n3344), .A4(n3343), .ZN(n3364)
         );
  AND4_X1 U3712 ( .A1(n3316), .A2(n3315), .A3(n3314), .A4(n3313), .ZN(n3254)
         );
  AND4_X1 U3713 ( .A1(n3297), .A2(n3296), .A3(n3295), .A4(n3294), .ZN(n3298)
         );
  AND2_X1 U3714 ( .A1(n3322), .A2(n3321), .ZN(n3323) );
  AND4_X1 U3715 ( .A1(n3271), .A2(n3270), .A3(n3269), .A4(n3268), .ZN(n3279)
         );
  AND4_X1 U3716 ( .A1(n3277), .A2(n3276), .A3(n3275), .A4(n3274), .ZN(n3278)
         );
  INV_X2 U3717 ( .A(n6359), .ZN(n6379) );
  NAND2_X2 U3718 ( .A1(STATE_REG_2__SCAN_IN), .A2(n7094), .ZN(n6671) );
  BUF_X2 U3719 ( .A(n3659), .Z(n3911) );
  BUF_X2 U3720 ( .A(n3380), .Z(n4012) );
  BUF_X2 U3721 ( .A(n3373), .Z(n5396) );
  BUF_X2 U3722 ( .A(n3379), .Z(n4025) );
  BUF_X2 U3723 ( .A(n3356), .Z(n4035) );
  BUF_X2 U3724 ( .A(n4027), .Z(n4011) );
  BUF_X2 U3725 ( .A(n3422), .Z(n3285) );
  AND2_X2 U3726 ( .A1(n5395), .A2(n3273), .ZN(n3407) );
  AND2_X2 U3727 ( .A1(n5395), .A2(n4563), .ZN(n3427) );
  AND2_X2 U3728 ( .A1(n3273), .A2(n4542), .ZN(n3465) );
  AND2_X2 U3729 ( .A1(n3273), .A2(n4553), .ZN(n3471) );
  NAND2_X2 U3730 ( .A1(n6683), .A2(n4969), .ZN(n6519) );
  AND2_X2 U3731 ( .A1(n4563), .A2(n4542), .ZN(n3422) );
  AND2_X2 U3732 ( .A1(n5458), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5395)
         );
  CLKBUF_X1 U3734 ( .A(n4053), .Z(n4002) );
  AND2_X2 U3735 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4542) );
  CLKBUF_X1 U3736 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n4559) );
  NOR2_X1 U3737 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n6027) );
  OAI21_X2 U3738 ( .B1(n4850), .B2(n4310), .A(n4247), .ZN(n5767) );
  NOR2_X1 U3739 ( .A1(n4122), .A2(n3391), .ZN(n3399) );
  AOI211_X2 U3740 ( .C1(n5424), .C2(REIP_REG_30__SCAN_IN), .A(n5423), .B(n5422), .ZN(n5425) );
  NOR2_X2 U3741 ( .A1(n5834), .A2(n4209), .ZN(n5593) );
  CLKBUF_X1 U3742 ( .A(n6375), .Z(n3159) );
  CLKBUF_X1 U3743 ( .A(n4575), .Z(n3160) );
  CLKBUF_X1 U3744 ( .A(n5141), .Z(n3161) );
  CLKBUF_X1 U3745 ( .A(n4998), .Z(n3162) );
  NAND2_X1 U3746 ( .A1(n5331), .A2(n3166), .ZN(n3163) );
  OR2_X1 U3747 ( .A1(n3165), .A2(n4325), .ZN(n3164) );
  INV_X1 U3748 ( .A(n4326), .ZN(n3165) );
  AND2_X1 U3749 ( .A1(n5330), .A2(n4326), .ZN(n3166) );
  CLKBUF_X1 U3750 ( .A(n5754), .Z(n3167) );
  INV_X1 U3751 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3168) );
  XNOR2_X1 U3753 ( .A(n3464), .B(n3507), .ZN(n4591) );
  NAND2_X1 U3754 ( .A1(n3394), .A2(n3365), .ZN(n3387) );
  NAND2_X1 U3755 ( .A1(n3510), .A2(n3463), .ZN(n3507) );
  NAND2_X2 U3756 ( .A1(n5660), .A2(n5687), .ZN(n4394) );
  NAND2_X2 U3757 ( .A1(n4323), .A2(n4322), .ZN(n5280) );
  AND2_X2 U3758 ( .A1(n4260), .A2(n6376), .ZN(n4526) );
  AND2_X2 U3759 ( .A1(n3776), .A2(n3398), .ZN(n4056) );
  INV_X1 U3760 ( .A(n3365), .ZN(n3334) );
  AND2_X4 U3761 ( .A1(n3272), .A2(n4553), .ZN(n4027) );
  NAND2_X1 U3762 ( .A1(n3334), .A2(n3776), .ZN(n3389) );
  NAND2_X2 U3763 ( .A1(n4361), .A2(n4335), .ZN(n4360) );
  NAND2_X2 U3764 ( .A1(n4333), .A2(n3190), .ZN(n4361) );
  AND2_X1 U3765 ( .A1(n3272), .A2(n3267), .ZN(n3172) );
  AND2_X4 U3766 ( .A1(n3272), .A2(n4542), .ZN(n3379) );
  NAND2_X4 U3767 ( .A1(n3181), .A2(n3262), .ZN(n3436) );
  AND2_X1 U3768 ( .A1(n4563), .A2(n4553), .ZN(n3175) );
  AND2_X1 U3769 ( .A1(n4563), .A2(n4553), .ZN(n4036) );
  AND2_X2 U3770 ( .A1(n4563), .A2(n4553), .ZN(n3174) );
  AND2_X2 U3771 ( .A1(n3544), .A2(n3578), .ZN(n4586) );
  AND2_X4 U3772 ( .A1(n5395), .A2(n3272), .ZN(n3408) );
  AND2_X1 U3773 ( .A1(n5395), .A2(n4545), .ZN(n3173) );
  AOI21_X2 U3774 ( .B1(n4360), .B2(n4339), .A(n4338), .ZN(n5660) );
  XNOR2_X2 U3775 ( .A(n3406), .B(n3442), .ZN(n3491) );
  NAND2_X2 U3776 ( .A1(n3446), .A2(n3445), .ZN(n4442) );
  AND2_X4 U3777 ( .A1(n3272), .A2(n3267), .ZN(n3659) );
  AND2_X1 U3778 ( .A1(n3635), .A2(n3634), .ZN(n3639) );
  INV_X1 U3779 ( .A(n5598), .ZN(n3206) );
  AND2_X1 U3780 ( .A1(n5745), .A2(n4334), .ZN(n4335) );
  NAND2_X1 U3781 ( .A1(n5732), .A2(n3235), .ZN(n5730) );
  AND2_X1 U3782 ( .A1(n4331), .A2(n4330), .ZN(n3235) );
  INV_X1 U3783 ( .A(n5747), .ZN(n4331) );
  INV_X1 U3784 ( .A(n3250), .ZN(n3249) );
  NAND2_X1 U3785 ( .A1(n4157), .A2(n4150), .ZN(n5464) );
  AND2_X1 U3786 ( .A1(n4199), .A2(n5615), .ZN(n3203) );
  INV_X1 U3787 ( .A(n5716), .ZN(n4363) );
  INV_X1 U3788 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4057) );
  AND2_X1 U3789 ( .A1(n3457), .A2(n3456), .ZN(n3459) );
  INV_X1 U3790 ( .A(n3638), .ZN(n3637) );
  NAND2_X1 U3791 ( .A1(n3221), .A2(n3436), .ZN(n3220) );
  OAI211_X1 U3792 ( .C1(n3512), .C2(n4057), .A(n3458), .B(n3459), .ZN(n3510)
         );
  NAND2_X1 U3793 ( .A1(n3385), .A2(n3158), .ZN(n3405) );
  AOI22_X1 U3794 ( .A1(n3421), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3422), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3328) );
  AOI22_X1 U3795 ( .A1(n3408), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3659), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3329) );
  NAND2_X1 U3796 ( .A1(n4143), .A2(n3204), .ZN(n4147) );
  NOR2_X1 U3797 ( .A1(n4465), .A2(n3776), .ZN(n3452) );
  OR2_X1 U3798 ( .A1(n3225), .A2(n5527), .ZN(n3224) );
  AND2_X1 U3799 ( .A1(n3852), .A2(n5609), .ZN(n3207) );
  NOR2_X1 U3800 ( .A1(n5711), .A2(n3238), .ZN(n3237) );
  INV_X1 U3801 ( .A(n4365), .ZN(n3238) );
  NOR2_X1 U3802 ( .A1(n5260), .A2(n3197), .ZN(n3196) );
  INV_X1 U3803 ( .A(n5148), .ZN(n3197) );
  NAND2_X1 U3804 ( .A1(n4550), .A2(n6613), .ZN(n3569) );
  AND2_X1 U3805 ( .A1(n4446), .A2(n4064), .ZN(n4543) );
  NOR2_X1 U3806 ( .A1(n4052), .A2(n5445), .ZN(n4401) );
  NAND2_X1 U3807 ( .A1(n4515), .A2(n4509), .ZN(n6272) );
  AND2_X1 U3808 ( .A1(n4508), .A2(n7066), .ZN(n4509) );
  NAND2_X1 U3809 ( .A1(n5486), .A2(n3231), .ZN(n4400) );
  AND2_X1 U3810 ( .A1(n4055), .A2(n3232), .ZN(n3231) );
  NAND2_X1 U3811 ( .A1(n4373), .A2(n3226), .ZN(n3225) );
  INV_X1 U3812 ( .A(n5590), .ZN(n3226) );
  AOI21_X1 U3813 ( .B1(n4586), .B2(n3766), .A(n3545), .ZN(n4523) );
  NAND2_X1 U3814 ( .A1(n3486), .A2(n3674), .ZN(n3213) );
  INV_X1 U3815 ( .A(n3486), .ZN(n3214) );
  INV_X1 U3816 ( .A(n5600), .ZN(n3202) );
  AND2_X1 U3817 ( .A1(n4195), .A2(n5612), .ZN(n5611) );
  NAND2_X1 U3818 ( .A1(n4361), .A2(n3189), .ZN(n5723) );
  NAND2_X1 U3819 ( .A1(n5629), .A2(n5630), .ZN(n5628) );
  AND2_X1 U3820 ( .A1(n5729), .A2(n5734), .ZN(n5747) );
  NAND2_X1 U3821 ( .A1(n4328), .A2(n4327), .ZN(n5754) );
  NAND2_X1 U3822 ( .A1(n4314), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4326) );
  NAND2_X1 U3823 ( .A1(n3247), .A2(n3245), .ZN(n5331) );
  AOI21_X1 U3824 ( .B1(n3246), .B2(n3250), .A(n3192), .ZN(n3245) );
  NAND2_X1 U3825 ( .A1(n4478), .A2(n4477), .ZN(n4495) );
  INV_X1 U3826 ( .A(n6620), .ZN(n4505) );
  NAND2_X1 U3827 ( .A1(n5475), .A2(REIP_REG_31__SCAN_IN), .ZN(n3200) );
  AND2_X1 U3828 ( .A1(n5244), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5245) );
  AND2_X1 U3829 ( .A1(n6215), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6212) );
  OAI21_X1 U3830 ( .B1(n4380), .B2(n4055), .A(n4400), .ZN(n4356) );
  AOI21_X1 U3831 ( .B1(n5792), .B2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n5777), 
        .ZN(n5778) );
  NAND2_X1 U3832 ( .A1(n3592), .A2(n3591), .ZN(n3622) );
  OR2_X1 U3833 ( .A1(n3633), .A2(n3632), .ZN(n4293) );
  INV_X1 U3834 ( .A(n4315), .ZN(n3420) );
  OR2_X1 U3835 ( .A1(n3477), .A2(n3476), .ZN(n4239) );
  OR2_X1 U3836 ( .A1(n3529), .A2(n3528), .ZN(n4249) );
  OR2_X1 U3837 ( .A1(n3386), .A2(n6613), .ZN(n3557) );
  OR2_X1 U3838 ( .A1(n3436), .A2(n6613), .ZN(n3556) );
  AND2_X1 U3839 ( .A1(n4097), .A2(n4096), .ZN(n4413) );
  AOI22_X1 U3840 ( .A1(n3407), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3465), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3303) );
  AOI22_X1 U3841 ( .A1(n3427), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3292) );
  AOI22_X1 U3842 ( .A1(n3471), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3422), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3290) );
  AOI22_X1 U3843 ( .A1(n3407), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3422), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3275) );
  NOR2_X1 U3844 ( .A1(n4379), .A2(n3233), .ZN(n3232) );
  INV_X1 U3845 ( .A(n5487), .ZN(n3233) );
  NAND2_X1 U3846 ( .A1(n3223), .A2(n5512), .ZN(n3222) );
  INV_X1 U3847 ( .A(n3224), .ZN(n3223) );
  NAND2_X1 U3848 ( .A1(n3211), .A2(n5306), .ZN(n3210) );
  INV_X1 U3849 ( .A(n3729), .ZN(n3211) );
  NAND2_X1 U3850 ( .A1(n3728), .A2(n3727), .ZN(n3743) );
  NOR2_X1 U3851 ( .A1(n5256), .A2(n3258), .ZN(n3728) );
  NAND2_X1 U3852 ( .A1(n3670), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3675)
         );
  INV_X1 U3853 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3676) );
  INV_X1 U3854 ( .A(n3642), .ZN(n3264) );
  INV_X1 U3855 ( .A(n5013), .ZN(n3230) );
  INV_X1 U3856 ( .A(n3504), .ZN(n3506) );
  NOR2_X1 U3857 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4053) );
  NOR2_X1 U3858 ( .A1(n5503), .A2(n3195), .ZN(n3194) );
  INV_X1 U3859 ( .A(n5515), .ZN(n3195) );
  AND3_X1 U3860 ( .A1(n3386), .A2(n3436), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n4098) );
  OAI21_X1 U3861 ( .B1(n3512), .B2(n4061), .A(n3397), .ZN(n3443) );
  NAND2_X1 U3862 ( .A1(n4128), .A2(n3216), .ZN(n3442) );
  INV_X1 U3863 ( .A(n3217), .ZN(n3216) );
  OAI211_X1 U3864 ( .C1(n3399), .C2(n4620), .A(n3218), .B(n3401), .ZN(n3217)
         );
  NAND2_X1 U3865 ( .A1(n3462), .A2(n3461), .ZN(n3463) );
  OR2_X1 U3866 ( .A1(n3460), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3461)
         );
  AND3_X1 U3867 ( .A1(n4445), .A2(n4126), .A3(n4125), .ZN(n4127) );
  AOI21_X1 U3868 ( .B1(n4109), .B2(n4108), .A(n4107), .ZN(n4418) );
  NAND2_X1 U3869 ( .A1(n3519), .A2(n3518), .ZN(n3550) );
  OR2_X1 U3870 ( .A1(n3512), .A2(n3168), .ZN(n3519) );
  NOR2_X1 U3871 ( .A1(n3331), .A2(n3330), .ZN(n3332) );
  AOI21_X1 U3872 ( .B1(n6615), .B2(n4570), .A(n5927), .ZN(n4601) );
  AND2_X1 U3873 ( .A1(n4346), .A2(n4345), .ZN(n4446) );
  INV_X1 U3874 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6590) );
  INV_X1 U3875 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6586) );
  NOR2_X1 U3876 ( .A1(n4483), .A2(n4470), .ZN(n4544) );
  INV_X1 U3877 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5297) );
  INV_X1 U3878 ( .A(n4064), .ZN(n5227) );
  OR2_X1 U3879 ( .A1(n4192), .A2(n4191), .ZN(n5630) );
  NOR2_X1 U3880 ( .A1(n5337), .A2(n5338), .ZN(n5351) );
  OR2_X1 U3881 ( .A1(n4189), .A2(n4188), .ZN(n5352) );
  NOR2_X1 U3882 ( .A1(n4149), .A2(n6209), .ZN(n4645) );
  AND2_X1 U3883 ( .A1(n4517), .A2(n5234), .ZN(n6249) );
  AND2_X1 U3884 ( .A1(n3997), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3998)
         );
  AND2_X1 U3885 ( .A1(n3960), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3961)
         );
  NAND2_X1 U3886 ( .A1(n3961), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3996)
         );
  AND2_X1 U3887 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n3882), .ZN(n3883)
         );
  NAND2_X1 U3888 ( .A1(n3883), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3922)
         );
  NOR2_X1 U3889 ( .A1(n3848), .A2(n5971), .ZN(n3849) );
  NAND2_X1 U3890 ( .A1(n3849), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3881)
         );
  NOR2_X1 U3891 ( .A1(n3804), .A2(n5573), .ZN(n3805) );
  NAND2_X1 U3892 ( .A1(n3805), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3848)
         );
  NAND2_X1 U3893 ( .A1(n3790), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3804)
         );
  INV_X1 U3894 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5573) );
  NOR2_X1 U3895 ( .A1(n3774), .A2(n5755), .ZN(n3790) );
  OR2_X1 U3896 ( .A1(n3757), .A2(n6081), .ZN(n3774) );
  AND2_X1 U3897 ( .A1(n3722), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3723)
         );
  NOR2_X1 U3898 ( .A1(n3691), .A2(n6115), .ZN(n3722) );
  NOR2_X1 U3899 ( .A1(n5256), .A2(n3729), .ZN(n5307) );
  INV_X1 U3900 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6115) );
  NOR2_X1 U3901 ( .A1(n3675), .A2(n3676), .ZN(n3707) );
  CLKBUF_X1 U3902 ( .A(n5208), .Z(n5209) );
  AND2_X1 U3903 ( .A1(n3641), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3670)
         );
  INV_X1 U3904 ( .A(n3656), .ZN(n3657) );
  NAND2_X1 U3905 ( .A1(n4301), .A2(n3766), .ZN(n3658) );
  OAI21_X1 U3906 ( .B1(n4020), .B2(n3655), .A(n3654), .ZN(n3656) );
  INV_X1 U3907 ( .A(n3598), .ZN(n3616) );
  NAND2_X1 U3908 ( .A1(n3616), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3642)
         );
  NAND2_X1 U3909 ( .A1(n3599), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3598)
         );
  NAND2_X1 U3910 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3571) );
  OR2_X1 U3911 ( .A1(n5491), .A2(n4387), .ZN(n4385) );
  AND2_X1 U3912 ( .A1(n4385), .A2(n4150), .ZN(n5465) );
  NAND2_X1 U3913 ( .A1(n5514), .A2(n3193), .ZN(n5491) );
  AND2_X1 U3914 ( .A1(n3194), .A2(n5489), .ZN(n3193) );
  NAND2_X1 U3915 ( .A1(n5514), .A2(n5515), .ZN(n5517) );
  NAND2_X1 U3916 ( .A1(n5692), .A2(n3188), .ZN(n5693) );
  NAND2_X1 U3917 ( .A1(n5351), .A2(n5352), .ZN(n5357) );
  NOR2_X1 U3918 ( .A1(n5357), .A2(n5358), .ZN(n5629) );
  OR2_X1 U3919 ( .A1(n4183), .A2(n4182), .ZN(n5314) );
  NAND2_X1 U3920 ( .A1(n6110), .A2(n5314), .ZN(n5337) );
  NAND2_X1 U3921 ( .A1(n5281), .A2(n5282), .ZN(n3239) );
  NAND2_X1 U3922 ( .A1(n3244), .A2(n6349), .ZN(n3243) );
  NAND2_X1 U3923 ( .A1(n5281), .A2(n3241), .ZN(n3240) );
  NAND2_X1 U3924 ( .A1(n6348), .A2(n3242), .ZN(n3244) );
  NAND2_X1 U3925 ( .A1(n5147), .A2(n3187), .ZN(n6111) );
  AND2_X1 U3926 ( .A1(n5147), .A2(n3196), .ZN(n5271) );
  NAND2_X1 U3927 ( .A1(n5141), .A2(n5142), .ZN(n3234) );
  NAND2_X1 U3928 ( .A1(n5147), .A2(n5148), .ZN(n5259) );
  XNOR2_X1 U3929 ( .A(n4306), .B(n4305), .ZN(n5212) );
  AND2_X1 U3930 ( .A1(n4528), .A2(n6451), .ZN(n5381) );
  OR2_X1 U3931 ( .A1(n4167), .A2(n4166), .ZN(n4892) );
  OR2_X1 U3932 ( .A1(n4162), .A2(n4161), .ZN(n4579) );
  NAND2_X1 U3933 ( .A1(n4578), .A2(n4579), .ZN(n4768) );
  NAND2_X1 U3934 ( .A1(n4645), .A2(n4644), .ZN(n4646) );
  NOR2_X1 U3935 ( .A1(n4646), .A2(n4530), .ZN(n4578) );
  NAND2_X1 U3936 ( .A1(n3491), .A2(n6613), .ZN(n3487) );
  CLKBUF_X1 U3937 ( .A(n4546), .Z(n4547) );
  CLKBUF_X1 U3938 ( .A(n4411), .Z(n4412) );
  INV_X1 U3939 ( .A(n4899), .ZN(n4901) );
  NOR2_X1 U3940 ( .A1(n4735), .A2(n5902), .ZN(n4697) );
  AND2_X1 U3941 ( .A1(n5902), .A2(n4962), .ZN(n4773) );
  OR2_X1 U3942 ( .A1(n6514), .A2(n5902), .ZN(n4961) );
  AND2_X1 U3943 ( .A1(n4965), .A2(n5154), .ZN(n4967) );
  NAND2_X1 U3944 ( .A1(n4651), .A2(n4587), .ZN(n6514) );
  OR2_X1 U3945 ( .A1(n3512), .A2(n5398), .ZN(n3555) );
  NOR2_X1 U3946 ( .A1(n4849), .A2(n5902), .ZN(n4931) );
  INV_X1 U3947 ( .A(n4850), .ZN(n4962) );
  INV_X1 U3948 ( .A(n5023), .ZN(n4813) );
  INV_X1 U3949 ( .A(n4773), .ZN(n4848) );
  OR2_X1 U3950 ( .A1(n6681), .A2(n4601), .ZN(n4630) );
  OR2_X1 U3951 ( .A1(n4587), .A2(n4588), .ZN(n4849) );
  AOI21_X1 U3952 ( .B1(n6580), .B2(STATE2_REG_3__SCAN_IN), .A(n4813), .ZN(
        n6521) );
  AND2_X1 U3953 ( .A1(n5454), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4131) );
  NOR2_X1 U3954 ( .A1(n5412), .A2(n6078), .ZN(n6056) );
  NAND2_X1 U3955 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6079), .ZN(n6078) );
  AND2_X1 U3956 ( .A1(n5238), .A2(n5471), .ZN(n6156) );
  INV_X1 U3957 ( .A(n6212), .ZN(n6198) );
  INV_X1 U3958 ( .A(n6202), .ZN(n6178) );
  INV_X1 U3959 ( .A(n6156), .ZN(n6224) );
  AND2_X1 U3960 ( .A1(n4491), .A2(n4490), .ZN(n6209) );
  INV_X1 U3961 ( .A(n5449), .ZN(n6245) );
  AND2_X1 U3962 ( .A1(n5449), .A2(n4513), .ZN(n6246) );
  NAND2_X1 U3963 ( .A1(n4510), .A2(n6272), .ZN(n5449) );
  OAI21_X1 U3964 ( .B1(n4507), .B2(n4506), .A(n4505), .ZN(n4510) );
  OAI21_X1 U3965 ( .B1(n6271), .B2(n7066), .A(n6270), .ZN(n6283) );
  INV_X1 U3966 ( .A(n6609), .ZN(n4514) );
  XNOR2_X1 U3967 ( .A(n4405), .B(n4404), .ZN(n5244) );
  OR2_X1 U3968 ( .A1(n5589), .A2(n3225), .ZN(n5526) );
  AND2_X1 U3969 ( .A1(n5550), .A2(n5553), .ZN(n5990) );
  INV_X1 U3970 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5971) );
  INV_X1 U3971 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5755) );
  INV_X1 U3972 ( .A(n6391), .ZN(n6366) );
  NAND2_X1 U3973 ( .A1(n6372), .A2(n5768), .ZN(n6391) );
  NAND2_X1 U3974 ( .A1(n3212), .A2(n3486), .ZN(n4536) );
  NAND2_X1 U3975 ( .A1(n4589), .A2(n3766), .ZN(n3212) );
  INV_X1 U3976 ( .A(n6372), .ZN(n6383) );
  NAND2_X1 U3977 ( .A1(n5617), .A2(n3203), .ZN(n5601) );
  NAND2_X1 U3978 ( .A1(n5692), .A2(n4365), .ZN(n5710) );
  AND2_X1 U3979 ( .A1(n5617), .A2(n5615), .ZN(n5556) );
  INV_X1 U3980 ( .A(n4360), .ZN(n5724) );
  NAND2_X1 U3981 ( .A1(n5732), .A2(n4330), .ZN(n5746) );
  INV_X1 U3982 ( .A(n6427), .ZN(n6392) );
  INV_X1 U3983 ( .A(n5385), .ZN(n6424) );
  OR2_X1 U3984 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n4496), .ZN(n4529)
         );
  OR2_X1 U3985 ( .A1(n5858), .A2(n6425), .ZN(n6403) );
  INV_X1 U3986 ( .A(n6394), .ZN(n6439) );
  INV_X1 U3988 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6454) );
  NOR2_X1 U3989 ( .A1(n4412), .A2(n4620), .ZN(n6581) );
  INV_X1 U3990 ( .A(n4559), .ZN(n5398) );
  INV_X1 U3991 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6031) );
  INV_X1 U3992 ( .A(n4659), .ZN(n4687) );
  AND2_X1 U3993 ( .A1(n4663), .A2(n4662), .ZN(n4686) );
  INV_X1 U3994 ( .A(n6497), .ZN(n4723) );
  INV_X1 U3995 ( .A(n6460), .ZN(n6495) );
  INV_X1 U3996 ( .A(n6506), .ZN(n4758) );
  NAND2_X1 U3997 ( .A1(n5910), .A2(n4773), .ZN(n6503) );
  OAI211_X1 U3998 ( .C1(n5163), .C2(n6518), .A(n5162), .B(n5161), .ZN(n5199)
         );
  AOI22_X1 U3999 ( .A1(n5159), .A2(n6518), .B1(n5158), .B2(n5157), .ZN(n5207)
         );
  INV_X1 U4000 ( .A(n6512), .ZN(n5195) );
  INV_X1 U4001 ( .A(n6536), .ZN(n5165) );
  INV_X1 U4002 ( .A(n6544), .ZN(n5201) );
  AND2_X1 U4003 ( .A1(n4931), .A2(n4962), .ZN(n5936) );
  INV_X1 U4004 ( .A(n6532), .ZN(n5189) );
  INV_X1 U4005 ( .A(n6539), .ZN(n5169) );
  INV_X1 U4006 ( .A(n6546), .ZN(n5206) );
  INV_X1 U4007 ( .A(n6552), .ZN(n5174) );
  INV_X1 U4008 ( .A(n6564), .ZN(n5194) );
  INV_X1 U4009 ( .A(n6573), .ZN(n5184) );
  NOR2_X1 U4010 ( .A1(n4630), .A2(n3158), .ZN(n6512) );
  NOR2_X1 U4011 ( .A1(n6897), .A2(n4813), .ZN(n6526) );
  NOR2_X1 U4012 ( .A1(n4619), .A2(n4813), .ZN(n6532) );
  NOR2_X1 U4013 ( .A1(n4624), .A2(n4813), .ZN(n6539) );
  NOR2_X1 U4014 ( .A1(n4630), .A2(n4612), .ZN(n6544) );
  NOR2_X1 U4015 ( .A1(n7034), .A2(n4813), .ZN(n6546) );
  NOR2_X1 U4016 ( .A1(n6899), .A2(n4813), .ZN(n6552) );
  NOR2_X1 U4017 ( .A1(n5016), .A2(n4813), .ZN(n6564) );
  NOR2_X1 U4018 ( .A1(n4849), .A2(n4848), .ZN(n4659) );
  NOR2_X1 U4019 ( .A1(n4849), .A2(n5153), .ZN(n5935) );
  NOR2_X1 U4020 ( .A1(n4630), .A2(n5450), .ZN(n6569) );
  INV_X1 U4021 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6613) );
  INV_X1 U4022 ( .A(n6694), .ZN(n6615) );
  NAND2_X1 U4023 ( .A1(n4131), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6620) );
  INV_X1 U4024 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6683) );
  OAI21_X1 U4025 ( .B1(n5772), .B2(n6202), .A(n3198), .ZN(U2796) );
  INV_X1 U4026 ( .A(n3199), .ZN(n3198) );
  OR2_X1 U4027 ( .A1(n5790), .A2(n6233), .ZN(n4237) );
  AOI21_X1 U4028 ( .B1(n4391), .B2(n5980), .A(n4390), .ZN(n4392) );
  NOR2_X1 U4029 ( .A1(n6230), .A2(n5479), .ZN(n4390) );
  AOI21_X1 U4030 ( .B1(n5781), .B2(n6445), .A(n5780), .ZN(n5782) );
  NAND2_X1 U4031 ( .A1(n5779), .A2(n5778), .ZN(n5780) );
  INV_X1 U4032 ( .A(n3227), .ZN(n5567) );
  NOR2_X1 U4033 ( .A1(n5589), .A2(n5590), .ZN(n4372) );
  INV_X1 U4034 ( .A(n3776), .ZN(n3394) );
  AND2_X1 U4035 ( .A1(n3158), .A2(n4620), .ZN(n4064) );
  AND3_X1 U4036 ( .A1(n3449), .A2(n3448), .A3(n3158), .ZN(n3176) );
  OR2_X1 U4037 ( .A1(n5733), .A2(n6422), .ZN(n3177) );
  OR2_X1 U4038 ( .A1(n5355), .A2(n5631), .ZN(n3178) );
  OR2_X1 U4039 ( .A1(n3178), .A2(n3228), .ZN(n3179) );
  NAND2_X1 U4040 ( .A1(n3396), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3512) );
  NOR2_X1 U4041 ( .A1(n5589), .A2(n3224), .ZN(n5511) );
  NAND2_X1 U4042 ( .A1(n5608), .A2(n5609), .ZN(n5551) );
  INV_X1 U4043 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5458) );
  AND4_X1 U4044 ( .A1(n3293), .A2(n3292), .A3(n3291), .A4(n3290), .ZN(n3180)
         );
  AND4_X1 U4045 ( .A1(n3378), .A2(n3377), .A3(n3376), .A4(n3375), .ZN(n3181)
         );
  INV_X1 U4046 ( .A(n5282), .ZN(n3242) );
  NOR2_X1 U4047 ( .A1(n5568), .A2(n3819), .ZN(n5608) );
  OR3_X1 U4048 ( .A1(n5429), .A2(n5428), .A3(n5438), .ZN(n3182) );
  INV_X1 U4049 ( .A(n6349), .ZN(n3251) );
  NAND2_X1 U4050 ( .A1(n3334), .A2(n3366), .ZN(n3448) );
  INV_X1 U4051 ( .A(n3253), .ZN(n3252) );
  AND2_X1 U4052 ( .A1(n3239), .A2(n6348), .ZN(n3253) );
  OAI211_X1 U4053 ( .C1(n4589), .C2(n3214), .A(n3213), .B(n4535), .ZN(n3504)
         );
  INV_X1 U4054 ( .A(n3236), .ZN(n5709) );
  NAND2_X1 U4055 ( .A1(n5692), .A2(n3237), .ZN(n3236) );
  NAND2_X1 U4056 ( .A1(n4364), .A2(n4363), .ZN(n5692) );
  NAND2_X1 U4057 ( .A1(n3615), .A2(n3614), .ZN(n3623) );
  AND2_X1 U4058 ( .A1(n4321), .A2(n3177), .ZN(n3183) );
  AND2_X1 U4059 ( .A1(n3623), .A2(n3591), .ZN(n3184) );
  NAND2_X2 U4060 ( .A1(n4612), .A2(n3436), .ZN(n4157) );
  OR2_X1 U4061 ( .A1(n5208), .A2(n5257), .ZN(n5256) );
  NAND2_X1 U4062 ( .A1(n3261), .A2(n3388), .ZN(n4122) );
  OR2_X1 U4063 ( .A1(n5349), .A2(n5355), .ZN(n5354) );
  AND2_X1 U4064 ( .A1(n3207), .A2(n3206), .ZN(n3185) );
  AND3_X1 U4065 ( .A1(n3621), .A2(n3230), .A3(n3620), .ZN(n5014) );
  AND2_X1 U4066 ( .A1(n5014), .A2(n5093), .ZN(n5092) );
  OAI21_X1 U4067 ( .B1(n5280), .B2(n3252), .A(n3250), .ZN(n5308) );
  NAND2_X1 U4068 ( .A1(n3234), .A2(n4321), .ZN(n5263) );
  AND2_X1 U4069 ( .A1(n5593), .A2(n4216), .ZN(n5514) );
  NAND2_X1 U4070 ( .A1(n3621), .A2(n3620), .ZN(n4765) );
  AND2_X1 U4071 ( .A1(n5514), .A2(n3194), .ZN(n3186) );
  NAND2_X1 U4072 ( .A1(n3731), .A2(n3208), .ZN(n5326) );
  AND2_X1 U4073 ( .A1(n5272), .A2(n3196), .ZN(n3187) );
  OR2_X1 U4074 ( .A1(n5349), .A2(n3178), .ZN(n3227) );
  AND2_X1 U4075 ( .A1(n3237), .A2(n5702), .ZN(n3188) );
  AND2_X1 U4076 ( .A1(n4335), .A2(n5874), .ZN(n3189) );
  NAND2_X1 U4077 ( .A1(n5729), .A2(n4332), .ZN(n3190) );
  AND2_X1 U4078 ( .A1(n3203), .A2(n3202), .ZN(n3191) );
  NOR2_X1 U4079 ( .A1(n4768), .A2(n4770), .ZN(n4890) );
  AND2_X1 U4080 ( .A1(n5729), .A2(n4324), .ZN(n3192) );
  INV_X1 U4081 ( .A(n5566), .ZN(n3228) );
  INV_X1 U4082 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6081) );
  INV_X1 U4083 ( .A(n5469), .ZN(n3201) );
  NAND2_X1 U4084 ( .A1(n3389), .A2(n4244), .ZN(n3449) );
  XNOR2_X1 U4085 ( .A(n4148), .B(n4147), .ZN(n4491) );
  NAND3_X1 U4086 ( .A1(n5557), .A2(n4490), .A3(n3205), .ZN(n3204) );
  INV_X1 U4087 ( .A(EBX_REG_1__SCAN_IN), .ZN(n3205) );
  NAND2_X1 U4088 ( .A1(n5608), .A2(n3207), .ZN(n5550) );
  NAND2_X1 U4089 ( .A1(n3743), .A2(n3209), .ZN(n3208) );
  NAND2_X1 U4090 ( .A1(n5326), .A2(n5328), .ZN(n5327) );
  INV_X1 U4091 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3215) );
  INV_X1 U4092 ( .A(n3219), .ZN(n3218) );
  OAI211_X1 U4093 ( .C1(n3403), .C2(n3221), .A(n3220), .B(n3400), .ZN(n3219)
         );
  INV_X1 U4094 ( .A(n4625), .ZN(n3221) );
  OR2_X2 U4095 ( .A1(n5589), .A2(n3222), .ZN(n5499) );
  NAND4_X1 U4096 ( .A1(n3230), .A2(n5093), .A3(n3621), .A4(n3229), .ZN(n5208)
         );
  NAND2_X1 U4097 ( .A1(n5486), .A2(n5487), .ZN(n4378) );
  AND2_X1 U4098 ( .A1(n5486), .A2(n3232), .ZN(n4380) );
  XNOR2_X2 U4099 ( .A(n4400), .B(n4399), .ZN(n5462) );
  NAND2_X1 U4100 ( .A1(n3234), .A2(n3183), .ZN(n4323) );
  NAND2_X1 U4101 ( .A1(n3592), .A2(n3184), .ZN(n3638) );
  NAND2_X2 U4102 ( .A1(n5754), .A2(n5753), .ZN(n5732) );
  NAND2_X1 U4103 ( .A1(n5280), .A2(n3248), .ZN(n3247) );
  OAI21_X1 U4104 ( .B1(n5280), .B2(n5281), .A(n5282), .ZN(n6350) );
  NAND2_X1 U4105 ( .A1(n3743), .A2(n3727), .ZN(n3731) );
  NAND2_X1 U4106 ( .A1(n4368), .A2(n5825), .ZN(n4369) );
  NAND2_X1 U4107 ( .A1(n3369), .A2(n3386), .ZN(n3402) );
  AND2_X1 U4108 ( .A1(n4620), .A2(n3436), .ZN(n4118) );
  NAND2_X1 U4109 ( .A1(n4586), .A2(n4056), .ZN(n4256) );
  INV_X1 U4110 ( .A(n4465), .ZN(n4625) );
  NAND2_X1 U4111 ( .A1(n3511), .A2(n3169), .ZN(n3549) );
  INV_X1 U4112 ( .A(n6445), .ZN(n6431) );
  AND2_X1 U4113 ( .A1(n4495), .A2(n4489), .ZN(n6445) );
  INV_X1 U4114 ( .A(n4586), .ZN(n4587) );
  NOR2_X1 U4115 ( .A1(n4547), .A2(n3170), .ZN(n3256) );
  NOR2_X2 U4116 ( .A1(n4651), .A2(n5020), .ZN(n3257) );
  OR2_X1 U4117 ( .A1(n3259), .A2(n5270), .ZN(n3258) );
  OR2_X1 U4118 ( .A1(n5302), .A2(n3706), .ZN(n3259) );
  AND4_X1 U4119 ( .A1(n3320), .A2(n3319), .A3(n3318), .A4(n3317), .ZN(n3260)
         );
  AND2_X2 U4120 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4545) );
  NAND2_X1 U4121 ( .A1(n3334), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3674) );
  INV_X1 U4122 ( .A(n6230), .ZN(n5605) );
  INV_X1 U4123 ( .A(n5605), .ZN(n6238) );
  AND2_X1 U4124 ( .A1(n6238), .A2(n5450), .ZN(n5980) );
  NAND2_X1 U4125 ( .A1(n6238), .A2(n3366), .ZN(n6226) );
  INV_X1 U4126 ( .A(n6226), .ZN(n4383) );
  OR2_X1 U4127 ( .A1(n3389), .A2(n3386), .ZN(n3261) );
  AND4_X1 U4128 ( .A1(n3384), .A2(n3383), .A3(n3382), .A4(n3381), .ZN(n3262)
         );
  AND3_X1 U4129 ( .A1(n3341), .A2(n3340), .A3(n3339), .ZN(n3263) );
  NOR2_X1 U4130 ( .A1(n3366), .A2(n4969), .ZN(n3492) );
  OR2_X1 U4131 ( .A1(n4073), .A2(n4072), .ZN(n4075) );
  AND2_X1 U4132 ( .A1(n4089), .A2(n4076), .ZN(n4079) );
  NAND2_X1 U4133 ( .A1(n3387), .A2(n3366), .ZN(n3392) );
  AND2_X1 U4134 ( .A1(n3449), .A2(n4620), .ZN(n3371) );
  AND2_X2 U4135 ( .A1(n4061), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3272)
         );
  OR2_X1 U4136 ( .A1(n3613), .A2(n3612), .ZN(n4290) );
  AOI22_X1 U4137 ( .A1(n3421), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3422), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3307) );
  NAND2_X1 U4138 ( .A1(n4098), .A2(n4056), .ZN(n4104) );
  OR2_X1 U4139 ( .A1(n3567), .A2(n3566), .ZN(n4269) );
  AOI22_X1 U4140 ( .A1(n3465), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3374), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3274) );
  INV_X1 U4141 ( .A(n5552), .ZN(n3852) );
  INV_X1 U4142 ( .A(n3639), .ZN(n3636) );
  NAND2_X1 U4143 ( .A1(n3590), .A2(n3589), .ZN(n3591) );
  NAND2_X1 U4144 ( .A1(n3326), .A2(n3325), .ZN(n3331) );
  INV_X1 U4145 ( .A(n5621), .ZN(n3819) );
  INV_X1 U4146 ( .A(n3492), .ZN(n4020) );
  INV_X1 U4147 ( .A(n3881), .ZN(n3882) );
  INV_X1 U4148 ( .A(n4766), .ZN(n3620) );
  INV_X1 U4149 ( .A(n3923), .ZN(n3545) );
  NOR2_X1 U4150 ( .A1(n4311), .A2(n4310), .ZN(n4312) );
  OR2_X1 U4151 ( .A1(n3588), .A2(n3587), .ZN(n4273) );
  NAND2_X1 U4152 ( .A1(n4490), .A2(n4150), .ZN(n4219) );
  NAND2_X1 U4153 ( .A1(n3557), .A2(n3556), .ZN(n4113) );
  OR2_X1 U4154 ( .A1(n3433), .A2(n3432), .ZN(n4245) );
  OR2_X1 U4155 ( .A1(n6384), .A2(n6622), .ZN(n5224) );
  AND2_X1 U4156 ( .A1(n3436), .A2(n5229), .ZN(n5230) );
  INV_X1 U4157 ( .A(n4053), .ZN(n3924) );
  INV_X1 U4158 ( .A(n4020), .ZN(n4048) );
  OR2_X1 U4159 ( .A1(n4403), .A2(n4402), .ZN(n4405) );
  OR2_X1 U4160 ( .A1(n5919), .A2(n6613), .ZN(n4050) );
  NAND2_X1 U4161 ( .A1(n3707), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3691)
         );
  OR4_X1 U4162 ( .A1(n5729), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_26__SCAN_IN), .A4(INSTADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n4395) );
  NAND2_X1 U4163 ( .A1(n5733), .A2(n5844), .ZN(n4366) );
  NAND2_X1 U4164 ( .A1(n4213), .A2(n4159), .ZN(n4193) );
  NAND2_X1 U4165 ( .A1(n4504), .A2(n4512), .ZN(n4488) );
  NAND2_X1 U4166 ( .A1(n3555), .A2(n3554), .ZN(n4852) );
  NAND2_X1 U4167 ( .A1(n3998), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4052)
         );
  NOR2_X1 U4168 ( .A1(n3922), .A2(n5697), .ZN(n3943) );
  OR2_X1 U4169 ( .A1(n6611), .A2(n5224), .ZN(n5225) );
  AND2_X1 U4170 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n3264), .ZN(n3641)
         );
  INV_X1 U4171 ( .A(n4133), .ZN(n4490) );
  INV_X1 U4172 ( .A(n3674), .ZN(n3766) );
  NAND2_X1 U4173 ( .A1(n5723), .A2(n4362), .ZN(n5717) );
  NAND2_X1 U4174 ( .A1(n4589), .A2(n4056), .ZN(n4243) );
  NOR2_X1 U4175 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4601), .ZN(n5023) );
  OR2_X1 U4176 ( .A1(n4651), .A2(n4653), .ZN(n4899) );
  AND2_X1 U4177 ( .A1(n3455), .A2(n3514), .ZN(n5065) );
  INV_X1 U4178 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6594) );
  AND2_X1 U4179 ( .A1(n5067), .A2(n5066), .ZN(n5933) );
  INV_X1 U4180 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n5454) );
  NAND2_X1 U4181 ( .A1(n4435), .A2(n4436), .ZN(n6690) );
  OR2_X1 U4182 ( .A1(n5960), .A2(n5406), .ZN(n5529) );
  AND2_X1 U4183 ( .A1(n5405), .A2(n6062), .ZN(n5960) );
  NAND2_X1 U4184 ( .A1(n3723), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3757)
         );
  NOR2_X1 U4185 ( .A1(n5244), .A2(n5454), .ZN(n5226) );
  INV_X1 U4186 ( .A(n6181), .ZN(n6169) );
  NOR2_X1 U4187 ( .A1(n3571), .A2(n5297), .ZN(n3599) );
  AND2_X1 U4188 ( .A1(n6215), .A2(n5245), .ZN(n6211) );
  NOR2_X1 U4189 ( .A1(n6267), .A2(n6249), .ZN(n6261) );
  INV_X1 U4190 ( .A(n6272), .ZN(n6343) );
  INV_X1 U4191 ( .A(n5705), .ZN(n5984) );
  INV_X1 U4192 ( .A(n5993), .ZN(n6239) );
  AND2_X1 U4193 ( .A1(n4446), .A2(n4348), .ZN(n6597) );
  INV_X1 U4194 ( .A(n6357), .ZN(n6387) );
  OAI211_X1 U4195 ( .C1(n5431), .C2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5430), .B(n3182), .ZN(n5432) );
  AND2_X1 U4196 ( .A1(n5836), .A2(n5843), .ZN(n5826) );
  AND2_X1 U4197 ( .A1(n6027), .A2(n4351), .ZN(n6427) );
  INV_X1 U4198 ( .A(n5853), .ZN(n6425) );
  INV_X1 U4199 ( .A(n6392), .ZN(n6384) );
  AND2_X1 U4200 ( .A1(n4471), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5927) );
  NOR2_X1 U4201 ( .A1(n4899), .A2(n4962), .ZN(n4924) );
  OAI21_X1 U4202 ( .B1(n5024), .B2(n5025), .A(n5162), .ZN(n5049) );
  OAI21_X1 U4203 ( .B1(n5107), .B2(n5106), .A(n5105), .ZN(n5131) );
  OAI21_X1 U4204 ( .B1(n4701), .B2(n4700), .A(n4699), .ZN(n4725) );
  AND2_X1 U4205 ( .A1(n4697), .A2(n4962), .ZN(n6497) );
  INV_X1 U4206 ( .A(n4735), .ZN(n5910) );
  OR2_X1 U4207 ( .A1(n4816), .A2(n4815), .ZN(n4842) );
  INV_X1 U4208 ( .A(n4972), .ZN(n4990) );
  INV_X1 U4209 ( .A(n5152), .ZN(n5203) );
  INV_X1 U4210 ( .A(n6542), .ZN(n6571) );
  OR2_X1 U4211 ( .A1(n4856), .A2(n4855), .ZN(n4882) );
  INV_X1 U4212 ( .A(n4857), .ZN(n4951) );
  NOR2_X1 U4213 ( .A1(n4630), .A2(n4625), .ZN(n6536) );
  NOR2_X1 U4214 ( .A1(n6941), .A2(n4813), .ZN(n6558) );
  NOR2_X1 U4215 ( .A1(n6950), .A2(n4813), .ZN(n6573) );
  INV_X1 U4216 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6961) );
  AND2_X1 U4217 ( .A1(n5523), .A2(n5410), .ZN(n5488) );
  OR2_X1 U4218 ( .A1(n4159), .A2(n6206), .ZN(n6202) );
  NAND2_X1 U4219 ( .A1(n6215), .A2(n5226), .ZN(n6162) );
  AND2_X1 U4220 ( .A1(n4237), .A2(n4236), .ZN(n4238) );
  AND2_X1 U4221 ( .A1(n4132), .A2(n4505), .ZN(n6230) );
  INV_X1 U4222 ( .A(n6249), .ZN(n6269) );
  NAND2_X2 U4223 ( .A1(n4515), .A2(n4514), .ZN(n6346) );
  OR2_X1 U4224 ( .A1(n6627), .A2(n6519), .ZN(n6359) );
  NAND2_X1 U4225 ( .A1(n6357), .A2(n4350), .ZN(n6372) );
  NAND2_X1 U4226 ( .A1(n4515), .A2(n6597), .ZN(n6357) );
  AND2_X1 U4227 ( .A1(n5824), .A2(n5388), .ZN(n6002) );
  NAND2_X1 U4228 ( .A1(n4495), .A2(n4482), .ZN(n6394) );
  INV_X1 U4229 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6580) );
  INV_X1 U4230 ( .A(n4924), .ZN(n4692) );
  NAND2_X1 U4231 ( .A1(n4901), .A2(n4962), .ZN(n5056) );
  OR2_X1 U4232 ( .A1(n4651), .A2(n4774), .ZN(n5128) );
  NAND2_X1 U4233 ( .A1(n5910), .A2(n5019), .ZN(n6510) );
  OR2_X1 U4234 ( .A1(n4961), .A2(n4962), .ZN(n4972) );
  NAND2_X1 U4235 ( .A1(n4963), .A2(n4962), .ZN(n5152) );
  INV_X1 U4236 ( .A(n6526), .ZN(n5932) );
  INV_X1 U4237 ( .A(n6558), .ZN(n5179) );
  OR2_X1 U4238 ( .A1(n6514), .A2(n5153), .ZN(n6577) );
  OR2_X1 U4239 ( .A1(n6514), .A2(n4848), .ZN(n6542) );
  INV_X1 U4240 ( .A(n6569), .ZN(n5180) );
  INV_X1 U4241 ( .A(n5936), .ZN(n5091) );
  AOI21_X1 U4242 ( .B1(n4595), .B2(n4596), .A(n4594), .ZN(n4635) );
  OAI21_X1 U4243 ( .B1(n4356), .B2(n6226), .A(n4238), .ZN(U2829) );
  INV_X1 U4244 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3265) );
  XNOR2_X1 U4245 ( .A(n3722), .B(n3265), .ZN(n6105) );
  NOR2_X4 U4246 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4563) );
  INV_X1 U4247 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3266) );
  NOR2_X2 U4248 ( .A1(n3266), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3267)
         );
  AND2_X2 U4249 ( .A1(n3267), .A2(n3273), .ZN(n3380) );
  AOI22_X1 U4250 ( .A1(n3427), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3271) );
  NOR2_X4 U4251 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4553) );
  AND2_X2 U4252 ( .A1(n3267), .A2(n4545), .ZN(n3373) );
  AOI22_X1 U4253 ( .A1(n3471), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3373), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3270) );
  AND2_X2 U4254 ( .A1(n3267), .A2(n4563), .ZN(n3356) );
  AOI22_X1 U4255 ( .A1(n3659), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3356), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3269) );
  AOI22_X1 U4256 ( .A1(n3408), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3175), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3268) );
  AOI22_X1 U4257 ( .A1(n4027), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3173), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3277) );
  AOI22_X1 U4258 ( .A1(n3379), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3276) );
  AOI22_X1 U4259 ( .A1(n4048), .A2(EAX_REG_12__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n4969), .ZN(n3280) );
  MUX2_X1 U4260 ( .A(n6105), .B(n3280), .S(n3924), .Z(n3302) );
  AOI22_X1 U4261 ( .A1(n4026), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3284) );
  AOI22_X1 U4262 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n4006), .B1(n4033), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3283) );
  AOI22_X1 U4263 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n3911), .B1(n5396), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3282) );
  AOI22_X1 U4264 ( .A1(n4037), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4028), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3281) );
  NAND4_X1 U4265 ( .A1(n3284), .A2(n3283), .A3(n3282), .A4(n3281), .ZN(n3300)
         );
  AOI22_X1 U4266 ( .A1(n4011), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3413), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3289) );
  AOI22_X1 U4267 ( .A1(n4025), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3288) );
  AOI22_X1 U4268 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n4035), .B1(n3174), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3287) );
  AOI22_X1 U4269 ( .A1(n4034), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3286) );
  NAND4_X1 U4270 ( .A1(n3289), .A2(n3288), .A3(n3287), .A4(n3286), .ZN(n3299)
         );
  AOI22_X1 U4271 ( .A1(n3465), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3373), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3293) );
  AOI22_X1 U4272 ( .A1(n3408), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3175), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3291) );
  AOI22_X1 U4273 ( .A1(n4027), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3173), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3297) );
  AOI22_X1 U4274 ( .A1(n3659), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3374), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3296) );
  AOI22_X1 U4275 ( .A1(n3407), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3356), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3295) );
  AOI22_X1 U4276 ( .A1(n3380), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3379), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3294) );
  OAI21_X1 U4277 ( .B1(n3300), .B2(n3299), .A(n3766), .ZN(n3301) );
  NAND2_X1 U4278 ( .A1(n3302), .A2(n3301), .ZN(n5306) );
  AOI22_X1 U4279 ( .A1(n3408), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3172), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3306) );
  AOI22_X1 U4280 ( .A1(n4036), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3374), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3305) );
  AOI22_X1 U4281 ( .A1(n3373), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3356), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3304) );
  AND4_X2 U4282 ( .A1(n3306), .A2(n3305), .A3(n3304), .A4(n3303), .ZN(n3312)
         );
  AOI22_X1 U4283 ( .A1(n4027), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3471), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3310) );
  AOI22_X1 U4284 ( .A1(n3427), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3379), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3309) );
  AOI22_X1 U4285 ( .A1(n3380), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3308) );
  NAND2_X4 U4286 ( .A1(n3312), .A2(n3311), .ZN(n3776) );
  AOI22_X1 U4287 ( .A1(n3427), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3316) );
  AOI22_X1 U4288 ( .A1(n4027), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3379), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3315) );
  AOI22_X1 U4289 ( .A1(n3408), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3465), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3314) );
  AOI22_X1 U4290 ( .A1(n3173), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3422), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3313) );
  AOI22_X1 U4291 ( .A1(n3407), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3373), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3320) );
  AOI22_X1 U4292 ( .A1(n3659), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3356), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3319) );
  AOI22_X1 U4293 ( .A1(n3471), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3318) );
  AOI22_X1 U4294 ( .A1(n3175), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3374), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3317) );
  NAND2_X2 U4295 ( .A1(n3254), .A2(n3260), .ZN(n3386) );
  AOI22_X1 U4296 ( .A1(n4036), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3374), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3324) );
  AOI22_X1 U4297 ( .A1(n3373), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3356), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3322) );
  AOI22_X1 U4298 ( .A1(n3407), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3465), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3321) );
  AOI22_X1 U4299 ( .A1(n3427), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3379), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3326) );
  AOI22_X1 U4300 ( .A1(n4027), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3471), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3325) );
  AOI22_X1 U4301 ( .A1(n3380), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3327) );
  NAND3_X1 U4302 ( .A1(n3329), .A2(n3328), .A3(n3327), .ZN(n3330) );
  OAI21_X1 U4303 ( .B1(n4117), .B2(n3369), .A(n4465), .ZN(n3372) );
  AOI22_X1 U4304 ( .A1(n3427), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3379), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3338) );
  AOI22_X1 U4305 ( .A1(n3408), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3659), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3337) );
  AOI22_X1 U4306 ( .A1(n3465), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3373), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3336) );
  AOI22_X1 U4307 ( .A1(n4027), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3422), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3335) );
  AOI22_X1 U4308 ( .A1(n3175), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3374), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3342) );
  AOI22_X1 U4309 ( .A1(n3407), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3356), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3341) );
  AOI22_X1 U4310 ( .A1(n3380), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3340) );
  AOI22_X1 U4311 ( .A1(n3421), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3471), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3339) );
  NAND2_X1 U4312 ( .A1(n3427), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3346) );
  NAND2_X1 U4313 ( .A1(n3380), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3345) );
  NAND2_X1 U4314 ( .A1(n4027), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3344) );
  NAND2_X1 U4315 ( .A1(n3471), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3343) );
  NAND2_X1 U4316 ( .A1(n3173), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3350)
         );
  NAND2_X1 U4317 ( .A1(n3407), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3349) );
  NAND2_X1 U4318 ( .A1(n3659), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3348) );
  NAND2_X1 U4319 ( .A1(n3422), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3347)
         );
  AND4_X2 U4320 ( .A1(n3350), .A2(n3349), .A3(n3348), .A4(n3347), .ZN(n3363)
         );
  NAND2_X1 U4321 ( .A1(n3379), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3355)
         );
  NAND2_X1 U4322 ( .A1(n3465), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3354)
         );
  NAND2_X1 U4323 ( .A1(n3373), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3353) );
  NAND2_X1 U4324 ( .A1(n3351), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3352) );
  AND4_X2 U4325 ( .A1(n3355), .A2(n3354), .A3(n3353), .A4(n3352), .ZN(n3362)
         );
  NAND2_X1 U4326 ( .A1(n3408), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3360)
         );
  NAND2_X1 U4327 ( .A1(n3356), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3359) );
  NAND2_X1 U4328 ( .A1(n4036), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3358) );
  NAND2_X1 U4329 ( .A1(n3374), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3357)
         );
  NAND4_X4 U4330 ( .A1(n3364), .A2(n3363), .A3(n3362), .A4(n3361), .ZN(n3398)
         );
  NAND2_X1 U4331 ( .A1(n4465), .A2(n3366), .ZN(n3367) );
  OAI21_X1 U4332 ( .B1(n4473), .B2(n3776), .A(n3367), .ZN(n3368) );
  INV_X1 U4333 ( .A(n3368), .ZN(n3370) );
  NAND2_X1 U4334 ( .A1(n3370), .A2(n3402), .ZN(n3450) );
  NAND3_X1 U4335 ( .A1(n3372), .A2(n3371), .A3(n3450), .ZN(n3385) );
  AOI22_X1 U4336 ( .A1(n3407), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3465), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3378) );
  AOI22_X1 U4337 ( .A1(n3408), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3659), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3377) );
  AOI22_X1 U4338 ( .A1(n3373), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3356), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3376) );
  AOI22_X1 U4339 ( .A1(n4036), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3374), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3375) );
  AOI22_X1 U4340 ( .A1(n3427), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3379), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3384) );
  AOI22_X1 U4341 ( .A1(n4027), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3471), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3383) );
  AOI22_X1 U4342 ( .A1(n3380), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3382) );
  AOI22_X1 U4343 ( .A1(n3421), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3422), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3381) );
  INV_X1 U4344 ( .A(n3392), .ZN(n3388) );
  NAND2_X1 U4345 ( .A1(n3389), .A2(n3386), .ZN(n3390) );
  NAND2_X1 U4346 ( .A1(n3390), .A2(n4244), .ZN(n3391) );
  OAI21_X1 U4347 ( .B1(n3392), .B2(n3386), .A(n4118), .ZN(n3393) );
  NAND2_X1 U4348 ( .A1(n3404), .A2(n4244), .ZN(n4485) );
  AND2_X2 U4349 ( .A1(n3393), .A2(n4485), .ZN(n3401) );
  NAND2_X1 U4350 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_1__SCAN_IN), .ZN(
        n6632) );
  OAI21_X1 U4351 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .A(
        n6632), .ZN(n4420) );
  NAND2_X1 U4352 ( .A1(n4620), .A2(n4420), .ZN(n3447) );
  AOI21_X1 U4353 ( .B1(n3447), .B2(n3394), .A(n4465), .ZN(n3395) );
  NAND4_X1 U4354 ( .A1(n3405), .A2(n3399), .A3(n3401), .A4(n3395), .ZN(n3396)
         );
  INV_X1 U4355 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4061) );
  NAND2_X1 U4356 ( .A1(n6027), .A2(n6613), .ZN(n4349) );
  MUX2_X1 U4357 ( .A(n4131), .B(n4349), .S(n6580), .Z(n3397) );
  INV_X1 U4358 ( .A(n3443), .ZN(n3406) );
  NAND2_X1 U4359 ( .A1(n6027), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6621) );
  AOI21_X1 U4360 ( .B1(n3449), .B2(n4118), .A(n6621), .ZN(n3400) );
  INV_X1 U4361 ( .A(n3402), .ZN(n3775) );
  NAND2_X1 U4362 ( .A1(n3775), .A2(n4612), .ZN(n3403) );
  AOI22_X1 U4363 ( .A1(n4006), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4034), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3412) );
  AOI22_X1 U4364 ( .A1(n4037), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3172), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3411) );
  AOI22_X1 U4365 ( .A1(n3373), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3356), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3410) );
  AOI22_X1 U4366 ( .A1(n3174), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4028), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3409) );
  NAND4_X1 U4367 ( .A1(n3412), .A2(n3411), .A3(n3410), .A4(n3409), .ZN(n3419)
         );
  AOI22_X1 U4368 ( .A1(n3427), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3417) );
  AOI22_X1 U4369 ( .A1(n4011), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3416) );
  AOI22_X1 U4370 ( .A1(n4012), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3415) );
  AOI22_X1 U4371 ( .A1(n3413), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3422), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3414) );
  NAND4_X1 U4372 ( .A1(n3417), .A2(n3416), .A3(n3415), .A4(n3414), .ZN(n3418)
         );
  INV_X1 U4373 ( .A(n3557), .ZN(n3530) );
  NAND2_X1 U4374 ( .A1(n3530), .A2(n3420), .ZN(n3481) );
  INV_X1 U4375 ( .A(n3481), .ZN(n3434) );
  AOI22_X1 U4376 ( .A1(n4012), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3426) );
  AOI22_X1 U4377 ( .A1(n4011), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3413), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3425) );
  AOI22_X1 U4378 ( .A1(n4034), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3422), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3424) );
  AOI22_X1 U4379 ( .A1(n4037), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3374), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3423) );
  NAND4_X1 U4380 ( .A1(n3426), .A2(n3425), .A3(n3424), .A4(n3423), .ZN(n3433)
         );
  AOI22_X1 U4381 ( .A1(n4006), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3431) );
  AOI22_X1 U4382 ( .A1(n3373), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3356), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3430) );
  AOI22_X1 U4383 ( .A1(n3659), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3429) );
  AOI22_X1 U4384 ( .A1(n3427), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3428) );
  NAND4_X1 U4385 ( .A1(n3431), .A2(n3430), .A3(n3429), .A4(n3428), .ZN(n3432)
         );
  MUX2_X1 U4386 ( .A(n4309), .B(n3434), .S(n4245), .Z(n3488) );
  INV_X1 U4387 ( .A(n3488), .ZN(n3435) );
  NAND2_X1 U4388 ( .A1(n3487), .A2(n3435), .ZN(n3440) );
  INV_X1 U4389 ( .A(n4245), .ZN(n3439) );
  AOI21_X1 U4390 ( .B1(n4608), .B2(n4315), .A(n6613), .ZN(n3438) );
  NAND2_X1 U4391 ( .A1(n4098), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3437) );
  OAI211_X1 U4392 ( .C1(n3439), .C2(n3436), .A(n3438), .B(n3437), .ZN(n3489)
         );
  AOI21_X1 U4393 ( .B1(n3440), .B2(n3489), .A(n4309), .ZN(n3441) );
  INV_X1 U4394 ( .A(n3441), .ZN(n3536) );
  NAND2_X1 U4395 ( .A1(n3443), .A2(n3442), .ZN(n3508) );
  INV_X1 U4396 ( .A(n3508), .ZN(n3464) );
  NAND2_X1 U4397 ( .A1(n4410), .A2(n3447), .ZN(n3453) );
  NAND3_X1 U4398 ( .A1(n3176), .A2(n3450), .A3(n3445), .ZN(n4411) );
  INV_X1 U4399 ( .A(n4411), .ZN(n3451) );
  NAND2_X1 U4400 ( .A1(n3451), .A2(n4620), .ZN(n4438) );
  AND2_X1 U4401 ( .A1(n3452), .A2(n4612), .ZN(n4129) );
  INV_X1 U4402 ( .A(n4473), .ZN(n4512) );
  NAND3_X1 U4403 ( .A1(n3453), .A2(n4438), .A3(n4488), .ZN(n3454) );
  NAND2_X1 U4404 ( .A1(n3454), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3458) );
  INV_X1 U4405 ( .A(n4349), .ZN(n3517) );
  NAND2_X1 U4406 ( .A1(n6580), .A2(n6586), .ZN(n3455) );
  NAND2_X1 U4407 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3514) );
  NAND2_X1 U4408 ( .A1(n3517), .A2(n5065), .ZN(n3457) );
  INV_X1 U4409 ( .A(n4131), .ZN(n3516) );
  NAND2_X1 U4410 ( .A1(n3516), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3456) );
  INV_X1 U4411 ( .A(n3458), .ZN(n3462) );
  INV_X1 U4412 ( .A(n3459), .ZN(n3460) );
  NAND2_X1 U4413 ( .A1(n4591), .A2(n6613), .ZN(n3479) );
  AOI22_X1 U4414 ( .A1(n4011), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3413), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3469) );
  AOI22_X1 U4415 ( .A1(n4006), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4034), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3468) );
  AOI22_X1 U4416 ( .A1(n4037), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4035), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3467) );
  AOI22_X1 U4417 ( .A1(n3174), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3374), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3466) );
  NAND4_X1 U4418 ( .A1(n3469), .A2(n3468), .A3(n3467), .A4(n3466), .ZN(n3477)
         );
  AOI22_X1 U4419 ( .A1(n3427), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3475) );
  AOI22_X1 U4420 ( .A1(n3659), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3474) );
  AOI22_X1 U4421 ( .A1(n4012), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3473) );
  AOI22_X1 U4422 ( .A1(n4033), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3422), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3472) );
  NAND4_X1 U4423 ( .A1(n3475), .A2(n3474), .A3(n3473), .A4(n3472), .ZN(n3476)
         );
  NAND2_X1 U4424 ( .A1(n3530), .A2(n4239), .ZN(n3478) );
  INV_X1 U4425 ( .A(n4239), .ZN(n3482) );
  NAND2_X1 U4426 ( .A1(n4098), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3480) );
  OAI211_X1 U4427 ( .C1(n3482), .C2(n3556), .A(n3481), .B(n3480), .ZN(n3538)
         );
  XNOR2_X2 U4428 ( .A(n3536), .B(n3483), .ZN(n4589) );
  AOI22_X1 U4429 ( .A1(n3492), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n4969), .ZN(n3485) );
  AND2_X1 U4430 ( .A1(n4512), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3570) );
  NAND2_X1 U4431 ( .A1(n3570), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3484) );
  AND2_X1 U4432 ( .A1(n3485), .A2(n3484), .ZN(n3486) );
  NAND2_X1 U4433 ( .A1(n3487), .A2(n3489), .ZN(n3490) );
  MUX2_X2 U4434 ( .A(n3490), .B(n3489), .S(n3488), .Z(n4850) );
  NAND2_X1 U4435 ( .A1(n4850), .A2(n3369), .ZN(n4499) );
  NAND2_X1 U4436 ( .A1(n3491), .A2(n3766), .ZN(n3496) );
  AOI22_X1 U4437 ( .A1(n3492), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n4969), .ZN(n3494) );
  NAND2_X1 U4438 ( .A1(n3570), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3493) );
  AND2_X1 U4439 ( .A1(n3494), .A2(n3493), .ZN(n3495) );
  NAND2_X1 U4440 ( .A1(n3496), .A2(n3495), .ZN(n4501) );
  AND2_X1 U4441 ( .A1(n4501), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3497) );
  NAND2_X1 U4442 ( .A1(n4499), .A2(n3497), .ZN(n4500) );
  INV_X1 U4443 ( .A(n4501), .ZN(n3498) );
  NAND2_X1 U4444 ( .A1(n3498), .A2(n4053), .ZN(n3499) );
  NAND2_X1 U4445 ( .A1(n4500), .A2(n3499), .ZN(n4535) );
  NAND2_X1 U4446 ( .A1(n3570), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3503) );
  INV_X1 U4447 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6197) );
  NAND2_X1 U4448 ( .A1(n4969), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3923) );
  OAI21_X1 U4449 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3571), .ZN(n6382) );
  NAND2_X1 U4450 ( .A1(n4053), .A2(n6382), .ZN(n3500) );
  OAI21_X1 U4451 ( .B1(n6197), .B2(n3923), .A(n3500), .ZN(n3501) );
  AOI21_X1 U4452 ( .B1(n3492), .B2(EAX_REG_2__SCAN_IN), .A(n3501), .ZN(n3502)
         );
  AND2_X1 U4453 ( .A1(n3503), .A2(n3502), .ZN(n4522) );
  NAND2_X1 U4454 ( .A1(n3504), .A2(n4522), .ZN(n3548) );
  INV_X1 U4455 ( .A(n4522), .ZN(n3505) );
  NAND2_X1 U4456 ( .A1(n3506), .A2(n3505), .ZN(n3546) );
  INV_X1 U4457 ( .A(n3507), .ZN(n3509) );
  NAND2_X1 U4458 ( .A1(n3509), .A2(n3508), .ZN(n3511) );
  INV_X1 U4459 ( .A(n3514), .ZN(n3513) );
  NAND2_X1 U4460 ( .A1(n3513), .A2(n6590), .ZN(n6511) );
  NAND2_X1 U4461 ( .A1(n3514), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3515) );
  NAND2_X1 U4462 ( .A1(n6511), .A2(n3515), .ZN(n4661) );
  AOI22_X1 U4463 ( .A1(n3517), .A2(n4661), .B1(n3516), .B2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3518) );
  XNOR2_X1 U4464 ( .A(n3549), .B(n3550), .ZN(n4546) );
  NAND2_X1 U4465 ( .A1(n4546), .A2(n6613), .ZN(n3532) );
  AOI22_X1 U4466 ( .A1(n4006), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4034), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3523) );
  AOI22_X1 U4467 ( .A1(n4037), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3659), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3522) );
  AOI22_X1 U4468 ( .A1(n5396), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4035), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3521) );
  AOI22_X1 U4469 ( .A1(n3174), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4028), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3520) );
  NAND4_X1 U4470 ( .A1(n3523), .A2(n3522), .A3(n3521), .A4(n3520), .ZN(n3529)
         );
  AOI22_X1 U4471 ( .A1(n4026), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3527) );
  AOI22_X1 U4472 ( .A1(n4011), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3526) );
  AOI22_X1 U4473 ( .A1(n4012), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3525) );
  AOI22_X1 U4474 ( .A1(n3413), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3524) );
  NAND4_X1 U4475 ( .A1(n3527), .A2(n3526), .A3(n3525), .A4(n3524), .ZN(n3528)
         );
  NAND2_X1 U4476 ( .A1(n3530), .A2(n4249), .ZN(n3531) );
  INV_X1 U4477 ( .A(n3556), .ZN(n3533) );
  AOI22_X1 U4478 ( .A1(n4098), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3533), 
        .B2(n4249), .ZN(n3534) );
  XNOR2_X2 U4479 ( .A(n3535), .B(n3534), .ZN(n3543) );
  NAND2_X1 U4480 ( .A1(n3537), .A2(n3536), .ZN(n3541) );
  NAND2_X1 U4481 ( .A1(n3539), .A2(n3538), .ZN(n3540) );
  NAND2_X1 U4482 ( .A1(n3541), .A2(n3540), .ZN(n3542) );
  NAND2_X2 U4483 ( .A1(n3543), .A2(n3542), .ZN(n3578) );
  NAND2_X1 U4484 ( .A1(n3546), .A2(n4523), .ZN(n3547) );
  NAND2_X1 U4485 ( .A1(n3548), .A2(n3547), .ZN(n4521) );
  INV_X1 U4486 ( .A(n3549), .ZN(n3551) );
  NOR3_X1 U4487 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6590), .A3(n6586), 
        .ZN(n6455) );
  NAND2_X1 U4488 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6455), .ZN(n4754) );
  NAND2_X1 U4489 ( .A1(n6594), .A2(n4754), .ZN(n3552) );
  NOR3_X1 U4490 ( .A1(n6594), .A2(n6590), .A3(n6586), .ZN(n5059) );
  NAND2_X1 U4491 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5059), .ZN(n4592) );
  NAND2_X1 U4492 ( .A1(n3552), .A2(n4592), .ZN(n4812) );
  OAI22_X1 U4493 ( .A1(n4349), .A2(n4812), .B1(n4131), .B2(n6594), .ZN(n3553)
         );
  INV_X1 U4494 ( .A(n3553), .ZN(n3554) );
  AOI22_X1 U4495 ( .A1(n4026), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3561) );
  AOI22_X1 U4496 ( .A1(n4011), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3413), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3560) );
  AOI22_X1 U4497 ( .A1(n4006), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3559) );
  AOI22_X1 U4498 ( .A1(n4037), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4028), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3558) );
  NAND4_X1 U4499 ( .A1(n3561), .A2(n3560), .A3(n3559), .A4(n3558), .ZN(n3567)
         );
  AOI22_X1 U4500 ( .A1(n4034), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3565) );
  AOI22_X1 U4501 ( .A1(n5396), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4035), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3564) );
  AOI22_X1 U4502 ( .A1(n3172), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3563) );
  AOI22_X1 U4503 ( .A1(n4025), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3562) );
  NAND4_X1 U4504 ( .A1(n3565), .A2(n3564), .A3(n3563), .A4(n3562), .ZN(n3566)
         );
  AOI22_X1 U4505 ( .A1(n4113), .A2(n4269), .B1(n4098), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3568) );
  XNOR2_X2 U4506 ( .A(n3578), .B(n3577), .ZN(n4650) );
  INV_X1 U4507 ( .A(n3570), .ZN(n3597) );
  INV_X1 U4508 ( .A(n3571), .ZN(n3573) );
  INV_X1 U4509 ( .A(n3599), .ZN(n3572) );
  OAI21_X1 U4510 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3573), .A(n3572), 
        .ZN(n5296) );
  AOI22_X1 U4511 ( .A1(n4002), .A2(n5296), .B1(n3545), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3575) );
  NAND2_X1 U4512 ( .A1(n4048), .A2(EAX_REG_3__SCAN_IN), .ZN(n3574) );
  OAI211_X1 U4513 ( .C1(n3597), .C2(n5398), .A(n3575), .B(n3574), .ZN(n3576)
         );
  AOI21_X1 U4514 ( .B1(n4650), .B2(n3766), .A(n3576), .ZN(n4539) );
  INV_X1 U4515 ( .A(n3577), .ZN(n4588) );
  NOR2_X2 U4516 ( .A1(n3578), .A2(n4588), .ZN(n3592) );
  AOI22_X1 U4517 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n4006), .B1(n4034), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3582) );
  AOI22_X1 U4518 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n4037), .B1(n3911), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3581) );
  AOI22_X1 U4519 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n5396), .B1(n4035), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3580) );
  AOI22_X1 U4520 ( .A1(n3174), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4028), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3579) );
  NAND4_X1 U4521 ( .A1(n3582), .A2(n3581), .A3(n3580), .A4(n3579), .ZN(n3588)
         );
  AOI22_X1 U4522 ( .A1(n4026), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3586) );
  AOI22_X1 U4523 ( .A1(n4011), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3585) );
  AOI22_X1 U4524 ( .A1(n4012), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3584) );
  AOI22_X1 U4525 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n3413), .B1(n3285), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3583) );
  NAND4_X1 U4526 ( .A1(n3586), .A2(n3585), .A3(n3584), .A4(n3583), .ZN(n3587)
         );
  NAND2_X1 U4527 ( .A1(n4113), .A2(n4273), .ZN(n3590) );
  NAND2_X1 U4528 ( .A1(n4098), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3589) );
  OR2_X1 U4529 ( .A1(n3592), .A2(n3591), .ZN(n3593) );
  NAND2_X1 U4530 ( .A1(n3593), .A2(n3622), .ZN(n4276) );
  INV_X1 U4531 ( .A(n4276), .ZN(n3594) );
  NAND2_X1 U4532 ( .A1(n3594), .A2(n3766), .ZN(n3603) );
  NAND2_X1 U4533 ( .A1(n4969), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3596)
         );
  NAND2_X1 U4534 ( .A1(n4048), .A2(EAX_REG_4__SCAN_IN), .ZN(n3595) );
  OAI211_X1 U4535 ( .C1(n3597), .C2(n6031), .A(n3596), .B(n3595), .ZN(n3600)
         );
  OAI21_X1 U4536 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n3599), .A(n3598), 
        .ZN(n6189) );
  MUX2_X1 U4537 ( .A(n3600), .B(n6189), .S(n4053), .Z(n3601) );
  INV_X1 U4538 ( .A(n3601), .ZN(n3602) );
  NAND2_X1 U4539 ( .A1(n3603), .A2(n3602), .ZN(n4585) );
  INV_X1 U4540 ( .A(n4584), .ZN(n3621) );
  AOI22_X1 U4541 ( .A1(n4012), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3607) );
  AOI22_X1 U4542 ( .A1(n4006), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4034), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3606) );
  AOI22_X1 U4543 ( .A1(n4011), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3605) );
  AOI22_X1 U4544 ( .A1(n5396), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3604) );
  NAND4_X1 U4545 ( .A1(n3607), .A2(n3606), .A3(n3605), .A4(n3604), .ZN(n3613)
         );
  AOI22_X1 U4546 ( .A1(n4025), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3413), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3611) );
  AOI22_X1 U4547 ( .A1(n3911), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4035), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3610) );
  AOI22_X1 U4548 ( .A1(n4026), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3609) );
  AOI22_X1 U4549 ( .A1(n4037), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4028), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3608) );
  NAND4_X1 U4550 ( .A1(n3611), .A2(n3610), .A3(n3609), .A4(n3608), .ZN(n3612)
         );
  NAND2_X1 U4551 ( .A1(n4113), .A2(n4290), .ZN(n3615) );
  NAND2_X1 U4552 ( .A1(n4098), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3614) );
  XNOR2_X1 U4553 ( .A(n3622), .B(n3623), .ZN(n4281) );
  INV_X1 U4554 ( .A(EAX_REG_5__SCAN_IN), .ZN(n3618) );
  OAI21_X1 U4555 ( .B1(PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n3616), .A(n3642), 
        .ZN(n6365) );
  AOI22_X1 U4556 ( .A1(n4002), .A2(n6365), .B1(n3545), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3617) );
  OAI21_X1 U4557 ( .B1(n4020), .B2(n3618), .A(n3617), .ZN(n3619) );
  AOI21_X1 U4558 ( .B1(n4281), .B2(n3766), .A(n3619), .ZN(n4766) );
  AOI22_X1 U4559 ( .A1(n4006), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4034), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3627) );
  AOI22_X1 U4560 ( .A1(n4037), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3626) );
  AOI22_X1 U4561 ( .A1(n5396), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4035), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3625) );
  AOI22_X1 U4562 ( .A1(n3174), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4028), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3624) );
  NAND4_X1 U4563 ( .A1(n3627), .A2(n3626), .A3(n3625), .A4(n3624), .ZN(n3633)
         );
  AOI22_X1 U4564 ( .A1(n4026), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3631) );
  AOI22_X1 U4565 ( .A1(n4011), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3630) );
  AOI22_X1 U4566 ( .A1(n4012), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3629) );
  AOI22_X1 U4567 ( .A1(n3413), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3628) );
  NAND4_X1 U4568 ( .A1(n3631), .A2(n3630), .A3(n3629), .A4(n3628), .ZN(n3632)
         );
  NAND2_X1 U4569 ( .A1(n4113), .A2(n4293), .ZN(n3635) );
  NAND2_X1 U4570 ( .A1(n4098), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3634) );
  NAND2_X1 U4571 ( .A1(n3638), .A2(n3639), .ZN(n3640) );
  INV_X1 U4572 ( .A(n3641), .ZN(n3651) );
  INV_X1 U4573 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3644) );
  NAND2_X1 U4574 ( .A1(n3644), .A2(n3642), .ZN(n3643) );
  NAND2_X1 U4575 ( .A1(n3651), .A2(n3643), .ZN(n6165) );
  INV_X1 U4576 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6319) );
  OAI22_X1 U4577 ( .A1(n4020), .A2(n6319), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3644), .ZN(n3645) );
  MUX2_X1 U4578 ( .A(n6165), .B(n3645), .S(n3924), .Z(n3646) );
  NAND2_X1 U4579 ( .A1(n4113), .A2(n4315), .ZN(n3648) );
  NAND2_X1 U4580 ( .A1(n4098), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3647) );
  NAND2_X1 U4581 ( .A1(n3648), .A2(n3647), .ZN(n3649) );
  INV_X1 U4582 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3655) );
  INV_X1 U4583 ( .A(n3670), .ZN(n3653) );
  INV_X1 U4584 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3650) );
  NAND2_X1 U4585 ( .A1(n3651), .A2(n3650), .ZN(n3652) );
  NAND2_X1 U4586 ( .A1(n3653), .A2(n3652), .ZN(n6358) );
  AOI22_X1 U4587 ( .A1(n6358), .A2(n4002), .B1(n3545), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3654) );
  NAND2_X1 U4588 ( .A1(n3658), .A2(n3657), .ZN(n5093) );
  AOI22_X1 U4589 ( .A1(n4025), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3663) );
  AOI22_X1 U4590 ( .A1(n4011), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3413), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3662) );
  AOI22_X1 U4591 ( .A1(n4006), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3661) );
  AOI22_X1 U4592 ( .A1(n4037), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3660) );
  NAND4_X1 U4593 ( .A1(n3663), .A2(n3662), .A3(n3661), .A4(n3660), .ZN(n3669)
         );
  AOI22_X1 U4594 ( .A1(n4034), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3667) );
  AOI22_X1 U4595 ( .A1(n4012), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3666) );
  AOI22_X1 U4596 ( .A1(n4026), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3665) );
  AOI22_X1 U4597 ( .A1(n4035), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4028), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3664) );
  NAND4_X1 U4598 ( .A1(n3667), .A2(n3666), .A3(n3665), .A4(n3664), .ZN(n3668)
         );
  NOR2_X1 U4599 ( .A1(n3669), .A2(n3668), .ZN(n3673) );
  XNOR2_X1 U4600 ( .A(n3670), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n6137) );
  AOI22_X1 U4601 ( .A1(n6137), .A2(n4002), .B1(n3545), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3672) );
  NAND2_X1 U4602 ( .A1(n4048), .A2(EAX_REG_8__SCAN_IN), .ZN(n3671) );
  OAI211_X1 U4603 ( .C1(n3674), .C2(n3673), .A(n3672), .B(n3671), .ZN(n5210)
         );
  XOR2_X1 U4604 ( .A(n3676), .B(n3675), .Z(n6124) );
  INV_X1 U4605 ( .A(n6124), .ZN(n5266) );
  AOI22_X1 U4606 ( .A1(n4026), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3680) );
  AOI22_X1 U4607 ( .A1(n4011), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3413), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3679) );
  AOI22_X1 U4608 ( .A1(n4037), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3678) );
  AOI22_X1 U4609 ( .A1(n4034), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3677) );
  NAND4_X1 U4610 ( .A1(n3680), .A2(n3679), .A3(n3678), .A4(n3677), .ZN(n3686)
         );
  AOI22_X1 U4611 ( .A1(n4006), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3684) );
  AOI22_X1 U4612 ( .A1(n3911), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4035), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3683) );
  AOI22_X1 U4613 ( .A1(n4025), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3682) );
  AOI22_X1 U4614 ( .A1(n3174), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4028), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3681) );
  NAND4_X1 U4615 ( .A1(n3684), .A2(n3683), .A3(n3682), .A4(n3681), .ZN(n3685)
         );
  OAI21_X1 U4616 ( .B1(n3686), .B2(n3685), .A(n3766), .ZN(n3689) );
  NAND2_X1 U4617 ( .A1(n4048), .A2(EAX_REG_9__SCAN_IN), .ZN(n3688) );
  NAND2_X1 U4618 ( .A1(n3545), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3687)
         );
  NAND3_X1 U4619 ( .A1(n3689), .A2(n3688), .A3(n3687), .ZN(n3690) );
  AOI21_X1 U4620 ( .B1(n5266), .B2(n4002), .A(n3690), .ZN(n5257) );
  XNOR2_X1 U4621 ( .A(n6115), .B(n3691), .ZN(n6352) );
  AOI22_X1 U4622 ( .A1(n4026), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3695) );
  AOI22_X1 U4623 ( .A1(n3413), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3694) );
  AOI22_X1 U4624 ( .A1(n4034), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3693) );
  AOI22_X1 U4625 ( .A1(n4035), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3692) );
  NAND4_X1 U4626 ( .A1(n3695), .A2(n3694), .A3(n3693), .A4(n3692), .ZN(n3701)
         );
  AOI22_X1 U4627 ( .A1(n4006), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4011), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3699) );
  AOI22_X1 U4628 ( .A1(n3911), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3698) );
  AOI22_X1 U4629 ( .A1(n4012), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3697) );
  AOI22_X1 U4630 ( .A1(n4037), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4028), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3696) );
  NAND4_X1 U4631 ( .A1(n3699), .A2(n3698), .A3(n3697), .A4(n3696), .ZN(n3700)
         );
  OAI21_X1 U4632 ( .B1(n3701), .B2(n3700), .A(n3766), .ZN(n3704) );
  NAND2_X1 U4633 ( .A1(n4048), .A2(EAX_REG_11__SCAN_IN), .ZN(n3703) );
  NAND2_X1 U4634 ( .A1(n3545), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3702)
         );
  NAND3_X1 U4635 ( .A1(n3704), .A2(n3703), .A3(n3702), .ZN(n3705) );
  AOI21_X1 U4636 ( .B1(n6352), .B2(n4002), .A(n3705), .ZN(n5302) );
  INV_X1 U4637 ( .A(n5306), .ZN(n3706) );
  XNOR2_X1 U4638 ( .A(n3707), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5286)
         );
  AOI22_X1 U4639 ( .A1(n4026), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3413), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3711) );
  AOI22_X1 U4640 ( .A1(n4006), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4034), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3710) );
  AOI22_X1 U4641 ( .A1(n3911), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3709) );
  AOI22_X1 U4642 ( .A1(n4037), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4028), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3708) );
  NAND4_X1 U4643 ( .A1(n3711), .A2(n3710), .A3(n3709), .A4(n3708), .ZN(n3717)
         );
  AOI22_X1 U4644 ( .A1(n4025), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3715) );
  AOI22_X1 U4645 ( .A1(n4012), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3714) );
  AOI22_X1 U4646 ( .A1(n4035), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3713) );
  AOI22_X1 U4647 ( .A1(n4011), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3712) );
  NAND4_X1 U4648 ( .A1(n3715), .A2(n3714), .A3(n3713), .A4(n3712), .ZN(n3716)
         );
  OAI21_X1 U4649 ( .B1(n3717), .B2(n3716), .A(n3766), .ZN(n3720) );
  NAND2_X1 U4650 ( .A1(n4048), .A2(EAX_REG_10__SCAN_IN), .ZN(n3719) );
  NAND2_X1 U4651 ( .A1(n3545), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3718)
         );
  NAND3_X1 U4652 ( .A1(n3720), .A2(n3719), .A3(n3718), .ZN(n3721) );
  AOI21_X1 U4653 ( .B1(n5286), .B2(n4002), .A(n3721), .ZN(n5270) );
  INV_X1 U4654 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3725) );
  OAI21_X1 U4655 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n3723), .A(n3757), 
        .ZN(n6100) );
  NAND2_X1 U4656 ( .A1(n6100), .A2(n4002), .ZN(n3724) );
  OAI21_X1 U4657 ( .B1(n3725), .B2(n3923), .A(n3724), .ZN(n3726) );
  AOI21_X1 U4658 ( .B1(n4048), .B2(EAX_REG_13__SCAN_IN), .A(n3726), .ZN(n3730)
         );
  INV_X1 U4659 ( .A(n3730), .ZN(n3727) );
  OR2_X1 U4660 ( .A1(n5270), .A2(n5302), .ZN(n3729) );
  AOI22_X1 U4661 ( .A1(n4026), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3735) );
  AOI22_X1 U4662 ( .A1(n3413), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3734) );
  AOI22_X1 U4663 ( .A1(n4006), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3733) );
  AOI22_X1 U4664 ( .A1(n4037), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4035), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3732) );
  NAND4_X1 U4665 ( .A1(n3735), .A2(n3734), .A3(n3733), .A4(n3732), .ZN(n3741)
         );
  AOI22_X1 U4666 ( .A1(n4034), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3739) );
  AOI22_X1 U4667 ( .A1(n4025), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3738) );
  AOI22_X1 U4668 ( .A1(n4011), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3737) );
  AOI22_X1 U4669 ( .A1(n3174), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4028), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3736) );
  NAND4_X1 U4670 ( .A1(n3739), .A2(n3738), .A3(n3737), .A4(n3736), .ZN(n3740)
         );
  OR2_X1 U4671 ( .A1(n3741), .A2(n3740), .ZN(n3742) );
  AND2_X1 U4672 ( .A1(n3766), .A2(n3742), .ZN(n5328) );
  NAND2_X1 U4673 ( .A1(n5327), .A2(n3743), .ZN(n5348) );
  XOR2_X1 U4674 ( .A(n6081), .B(n3757), .Z(n6084) );
  AOI22_X1 U4675 ( .A1(n4025), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3413), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3747) );
  AOI22_X1 U4676 ( .A1(n4037), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3746) );
  AOI22_X1 U4677 ( .A1(n4034), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4035), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3745) );
  AOI22_X1 U4678 ( .A1(n4026), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3744) );
  NAND4_X1 U4679 ( .A1(n3747), .A2(n3746), .A3(n3745), .A4(n3744), .ZN(n3753)
         );
  AOI22_X1 U4680 ( .A1(n4012), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3751) );
  AOI22_X1 U4681 ( .A1(n4006), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3750) );
  AOI22_X1 U4682 ( .A1(n4011), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3749) );
  AOI22_X1 U4683 ( .A1(n3174), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4028), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3748) );
  NAND4_X1 U4684 ( .A1(n3751), .A2(n3750), .A3(n3749), .A4(n3748), .ZN(n3752)
         );
  OR2_X1 U4685 ( .A1(n3753), .A2(n3752), .ZN(n3754) );
  AOI22_X1 U4686 ( .A1(n3766), .A2(n3754), .B1(n3545), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3756) );
  NAND2_X1 U4687 ( .A1(n4048), .A2(EAX_REG_14__SCAN_IN), .ZN(n3755) );
  OAI211_X1 U4688 ( .C1(n6084), .C2(n3924), .A(n3756), .B(n3755), .ZN(n5347)
         );
  NAND2_X1 U4689 ( .A1(n5348), .A2(n5347), .ZN(n5349) );
  XNOR2_X1 U4690 ( .A(n3774), .B(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6071)
         );
  INV_X1 U4691 ( .A(n6071), .ZN(n3773) );
  AOI22_X1 U4692 ( .A1(n4011), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3761) );
  AOI22_X1 U4693 ( .A1(n4006), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3760) );
  AOI22_X1 U4694 ( .A1(n4037), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4035), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3759) );
  AOI22_X1 U4695 ( .A1(n3413), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3758) );
  NAND4_X1 U4696 ( .A1(n3761), .A2(n3760), .A3(n3759), .A4(n3758), .ZN(n3768)
         );
  AOI22_X1 U4697 ( .A1(n4026), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3765) );
  AOI22_X1 U4698 ( .A1(n4034), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3764) );
  AOI22_X1 U4699 ( .A1(n4012), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3763) );
  AOI22_X1 U4700 ( .A1(n3174), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4028), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3762) );
  NAND4_X1 U4701 ( .A1(n3765), .A2(n3764), .A3(n3763), .A4(n3762), .ZN(n3767)
         );
  OAI21_X1 U4702 ( .B1(n3768), .B2(n3767), .A(n3766), .ZN(n3771) );
  NAND2_X1 U4703 ( .A1(n4048), .A2(EAX_REG_15__SCAN_IN), .ZN(n3770) );
  NAND2_X1 U4704 ( .A1(n3545), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3769)
         );
  NAND3_X1 U4705 ( .A1(n3771), .A2(n3770), .A3(n3769), .ZN(n3772) );
  AOI21_X1 U4706 ( .B1(n3773), .B2(n4053), .A(n3772), .ZN(n5355) );
  XNOR2_X1 U4707 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3790), .ZN(n6065)
         );
  NAND2_X1 U4708 ( .A1(n3775), .A2(n3776), .ZN(n5919) );
  AOI22_X1 U4709 ( .A1(n4011), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3780) );
  AOI22_X1 U4710 ( .A1(n4006), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3413), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3779) );
  AOI22_X1 U4711 ( .A1(n4025), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4712 ( .A1(n4034), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3777) );
  NAND4_X1 U4713 ( .A1(n3780), .A2(n3779), .A3(n3778), .A4(n3777), .ZN(n3786)
         );
  AOI22_X1 U4714 ( .A1(n4026), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3784) );
  AOI22_X1 U4715 ( .A1(n3911), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4035), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3783) );
  AOI22_X1 U4716 ( .A1(n5396), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3782) );
  AOI22_X1 U4717 ( .A1(n4037), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4028), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3781) );
  NAND4_X1 U4718 ( .A1(n3784), .A2(n3783), .A3(n3782), .A4(n3781), .ZN(n3785)
         );
  NOR2_X1 U4719 ( .A1(n3786), .A2(n3785), .ZN(n3788) );
  AOI22_X1 U4720 ( .A1(n4048), .A2(EAX_REG_16__SCAN_IN), .B1(n3545), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3787) );
  OAI21_X1 U4721 ( .B1(n4050), .B2(n3788), .A(n3787), .ZN(n3789) );
  AOI21_X1 U4722 ( .B1(n6065), .B2(n4002), .A(n3789), .ZN(n5631) );
  XNOR2_X1 U4723 ( .A(n3804), .B(n5573), .ZN(n5741) );
  AOI22_X1 U4724 ( .A1(n4026), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4725 ( .A1(n4011), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4726 ( .A1(n4035), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4727 ( .A1(n3911), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4028), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3791) );
  NAND4_X1 U4728 ( .A1(n3794), .A2(n3793), .A3(n3792), .A4(n3791), .ZN(n3800)
         );
  AOI22_X1 U4729 ( .A1(n4006), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3413), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3798) );
  AOI22_X1 U4730 ( .A1(n4034), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3797) );
  AOI22_X1 U4731 ( .A1(n4037), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3796) );
  AOI22_X1 U4732 ( .A1(n4025), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3795) );
  NAND4_X1 U4733 ( .A1(n3798), .A2(n3797), .A3(n3796), .A4(n3795), .ZN(n3799)
         );
  NOR2_X1 U4734 ( .A1(n3800), .A2(n3799), .ZN(n3802) );
  AOI22_X1 U4735 ( .A1(n4048), .A2(EAX_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n4969), .ZN(n3801) );
  OAI21_X1 U4736 ( .B1(n4050), .B2(n3802), .A(n3801), .ZN(n3803) );
  MUX2_X1 U4737 ( .A(n5741), .B(n3803), .S(n3924), .Z(n5566) );
  OAI21_X1 U4738 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n3805), .A(n3848), 
        .ZN(n6054) );
  AOI22_X1 U4739 ( .A1(n4026), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4740 ( .A1(n4006), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4011), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3808) );
  AOI22_X1 U4741 ( .A1(n4034), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4742 ( .A1(n4037), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4028), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3806) );
  NAND4_X1 U4743 ( .A1(n3809), .A2(n3808), .A3(n3807), .A4(n3806), .ZN(n3815)
         );
  AOI22_X1 U4744 ( .A1(n3413), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3813) );
  AOI22_X1 U4745 ( .A1(n4025), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3812) );
  AOI22_X1 U4746 ( .A1(n4035), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3811) );
  AOI22_X1 U4747 ( .A1(n5396), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3810) );
  NAND4_X1 U4748 ( .A1(n3813), .A2(n3812), .A3(n3811), .A4(n3810), .ZN(n3814)
         );
  NOR2_X1 U4749 ( .A1(n3815), .A2(n3814), .ZN(n3817) );
  AOI22_X1 U4750 ( .A1(n4048), .A2(EAX_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n4969), .ZN(n3816) );
  OAI21_X1 U4751 ( .B1(n4050), .B2(n3817), .A(n3816), .ZN(n3818) );
  MUX2_X1 U4752 ( .A(n6054), .B(n3818), .S(n3924), .Z(n5621) );
  XNOR2_X1 U4753 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .B(n3848), .ZN(n5969)
         );
  INV_X1 U4754 ( .A(n5969), .ZN(n3833) );
  AOI22_X1 U4755 ( .A1(n4025), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3823) );
  AOI22_X1 U4756 ( .A1(n4006), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3413), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4757 ( .A1(n4034), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4035), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4758 ( .A1(n4037), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4028), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3820) );
  NAND4_X1 U4759 ( .A1(n3823), .A2(n3822), .A3(n3821), .A4(n3820), .ZN(n3829)
         );
  AOI22_X1 U4760 ( .A1(n4026), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4011), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4761 ( .A1(n4012), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4762 ( .A1(n3911), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4763 ( .A1(n5396), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3824) );
  NAND4_X1 U4764 ( .A1(n3827), .A2(n3826), .A3(n3825), .A4(n3824), .ZN(n3828)
         );
  NOR2_X1 U4765 ( .A1(n3829), .A2(n3828), .ZN(n3831) );
  AOI22_X1 U4766 ( .A1(n4048), .A2(EAX_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n4969), .ZN(n3830) );
  OAI21_X1 U4767 ( .B1(n4050), .B2(n3831), .A(n3830), .ZN(n3832) );
  MUX2_X1 U4768 ( .A(n3833), .B(n3832), .S(n3924), .Z(n5609) );
  AOI22_X1 U4769 ( .A1(n4026), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3837) );
  AOI22_X1 U4770 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n4011), .B1(n4033), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3836) );
  AOI22_X1 U4771 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n4006), .B1(n5396), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3835) );
  AOI22_X1 U4772 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n4035), .B1(n3174), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3834) );
  NAND4_X1 U4773 ( .A1(n3837), .A2(n3836), .A3(n3835), .A4(n3834), .ZN(n3843)
         );
  AOI22_X1 U4774 ( .A1(n4034), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3841) );
  AOI22_X1 U4775 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n4012), .B1(n3470), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4776 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n3413), .B1(n3285), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3839) );
  AOI22_X1 U4777 ( .A1(n4037), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4028), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3838) );
  NAND4_X1 U4778 ( .A1(n3841), .A2(n3840), .A3(n3839), .A4(n3838), .ZN(n3842)
         );
  NOR2_X1 U4779 ( .A1(n3843), .A2(n3842), .ZN(n3847) );
  INV_X1 U4780 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6786) );
  OAI21_X1 U4781 ( .B1(PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6786), .A(n4969), 
        .ZN(n3844) );
  INV_X1 U4782 ( .A(n3844), .ZN(n3845) );
  AOI21_X1 U4783 ( .B1(n4048), .B2(EAX_REG_20__SCAN_IN), .A(n3845), .ZN(n3846)
         );
  OAI21_X1 U4784 ( .B1(n4050), .B2(n3847), .A(n3846), .ZN(n3851) );
  OAI21_X1 U4785 ( .B1(PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n3849), .A(n3881), 
        .ZN(n5720) );
  OR2_X1 U4786 ( .A1(n3924), .A2(n5720), .ZN(n3850) );
  NAND2_X1 U4787 ( .A1(n3851), .A2(n3850), .ZN(n5552) );
  AOI22_X1 U4788 ( .A1(n4026), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3856) );
  AOI22_X1 U4789 ( .A1(n4011), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4790 ( .A1(n4012), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4791 ( .A1(n3413), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3853) );
  NAND4_X1 U4792 ( .A1(n3856), .A2(n3855), .A3(n3854), .A4(n3853), .ZN(n3862)
         );
  AOI22_X1 U4793 ( .A1(n4006), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4034), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4794 ( .A1(n4037), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4795 ( .A1(n5396), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4035), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4796 ( .A1(n3174), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4028), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3857) );
  NAND4_X1 U4797 ( .A1(n3860), .A2(n3859), .A3(n3858), .A4(n3857), .ZN(n3861)
         );
  NOR2_X1 U4798 ( .A1(n3862), .A2(n3861), .ZN(n3866) );
  INV_X1 U4799 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3863) );
  AOI21_X1 U4800 ( .B1(n3863), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3864) );
  AOI21_X1 U4801 ( .B1(n4048), .B2(EAX_REG_21__SCAN_IN), .A(n3864), .ZN(n3865)
         );
  OAI21_X1 U4802 ( .B1(n4050), .B2(n3866), .A(n3865), .ZN(n3868) );
  XNOR2_X1 U4803 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .B(n3881), .ZN(n5961)
         );
  NAND2_X1 U4804 ( .A1(n5961), .A2(n4002), .ZN(n3867) );
  NAND2_X1 U4805 ( .A1(n3868), .A2(n3867), .ZN(n5598) );
  AOI22_X1 U4806 ( .A1(n4011), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3872) );
  AOI22_X1 U4807 ( .A1(n4034), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3871) );
  AOI22_X1 U4808 ( .A1(n4012), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3870) );
  AOI22_X1 U4809 ( .A1(n4037), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4028), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3869) );
  NAND4_X1 U4810 ( .A1(n3872), .A2(n3871), .A3(n3870), .A4(n3869), .ZN(n3878)
         );
  AOI22_X1 U4811 ( .A1(n4026), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3876) );
  AOI22_X1 U4812 ( .A1(n4006), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4035), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3875) );
  AOI22_X1 U4813 ( .A1(n3911), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3874) );
  AOI22_X1 U4814 ( .A1(n3413), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3873) );
  NAND4_X1 U4815 ( .A1(n3876), .A2(n3875), .A3(n3874), .A4(n3873), .ZN(n3877)
         );
  NOR2_X1 U4816 ( .A1(n3878), .A2(n3877), .ZN(n3880) );
  AOI22_X1 U4817 ( .A1(n4048), .A2(EAX_REG_22__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n4969), .ZN(n3879) );
  OAI21_X1 U4818 ( .B1(n4050), .B2(n3880), .A(n3879), .ZN(n3884) );
  OAI21_X1 U4819 ( .B1(n3883), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n3922), 
        .ZN(n5952) );
  MUX2_X1 U4820 ( .A(n3884), .B(n5952), .S(n4002), .Z(n5704) );
  NAND2_X1 U4821 ( .A1(n5597), .A2(n5704), .ZN(n5589) );
  AOI22_X1 U4822 ( .A1(n4026), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3888) );
  AOI22_X1 U4823 ( .A1(n4034), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4035), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3887) );
  AOI22_X1 U4824 ( .A1(n3911), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3886) );
  AOI22_X1 U4825 ( .A1(n4011), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3885) );
  NAND4_X1 U4826 ( .A1(n3888), .A2(n3887), .A3(n3886), .A4(n3885), .ZN(n3894)
         );
  AOI22_X1 U4827 ( .A1(n3413), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4828 ( .A1(n4006), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4829 ( .A1(n4025), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4830 ( .A1(n4037), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4028), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3889) );
  NAND4_X1 U4831 ( .A1(n3892), .A2(n3891), .A3(n3890), .A4(n3889), .ZN(n3893)
         );
  NOR2_X1 U4832 ( .A1(n3894), .A2(n3893), .ZN(n3909) );
  AOI22_X1 U4833 ( .A1(n4026), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3898) );
  AOI22_X1 U4834 ( .A1(n4011), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3897) );
  AOI22_X1 U4835 ( .A1(n4012), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3896) );
  AOI22_X1 U4836 ( .A1(n3413), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3895) );
  NAND4_X1 U4837 ( .A1(n3898), .A2(n3897), .A3(n3896), .A4(n3895), .ZN(n3904)
         );
  AOI22_X1 U4838 ( .A1(n4006), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4034), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3902) );
  AOI22_X1 U4839 ( .A1(n4037), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3901) );
  AOI22_X1 U4840 ( .A1(n5396), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4035), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3900) );
  AOI22_X1 U4841 ( .A1(n3174), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4028), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3899) );
  NAND4_X1 U4842 ( .A1(n3902), .A2(n3901), .A3(n3900), .A4(n3899), .ZN(n3903)
         );
  NOR2_X1 U4843 ( .A1(n3904), .A2(n3903), .ZN(n3910) );
  XOR2_X1 U4844 ( .A(n3909), .B(n3910), .Z(n3907) );
  INV_X1 U4845 ( .A(n4050), .ZN(n4022) );
  INV_X1 U4846 ( .A(EAX_REG_23__SCAN_IN), .ZN(n3905) );
  INV_X1 U4847 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5697) );
  OAI22_X1 U4848 ( .A1(n4020), .A2(n3905), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5697), .ZN(n3906) );
  AOI21_X1 U4849 ( .B1(n3907), .B2(n4022), .A(n3906), .ZN(n3908) );
  XNOR2_X1 U4850 ( .A(n3922), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5942)
         );
  MUX2_X1 U4851 ( .A(n3908), .B(n5942), .S(n4002), .Z(n5590) );
  OR2_X1 U4852 ( .A1(n3910), .A2(n3909), .ZN(n3929) );
  AOI22_X1 U4853 ( .A1(n4034), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4035), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4854 ( .A1(n4037), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3914) );
  AOI22_X1 U4855 ( .A1(n4026), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3913) );
  AOI22_X1 U4856 ( .A1(n3174), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4028), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3912) );
  NAND4_X1 U4857 ( .A1(n3915), .A2(n3914), .A3(n3913), .A4(n3912), .ZN(n3921)
         );
  AOI22_X1 U4858 ( .A1(n4012), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3919) );
  AOI22_X1 U4859 ( .A1(n4006), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3413), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3918) );
  AOI22_X1 U4860 ( .A1(n4025), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3917) );
  AOI22_X1 U4861 ( .A1(n4011), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3916) );
  NAND4_X1 U4862 ( .A1(n3919), .A2(n3918), .A3(n3917), .A4(n3916), .ZN(n3920)
         );
  NOR2_X1 U4863 ( .A1(n3921), .A2(n3920), .ZN(n3928) );
  XNOR2_X1 U4864 ( .A(n3929), .B(n3928), .ZN(n3927) );
  INV_X1 U4865 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5544) );
  XNOR2_X1 U4866 ( .A(n3943), .B(n5544), .ZN(n5547) );
  OAI22_X1 U4867 ( .A1(n5547), .A2(n3924), .B1(n5544), .B2(n3923), .ZN(n3925)
         );
  AOI21_X1 U4868 ( .B1(n4048), .B2(EAX_REG_24__SCAN_IN), .A(n3925), .ZN(n3926)
         );
  OAI21_X1 U4869 ( .B1(n4050), .B2(n3927), .A(n3926), .ZN(n4373) );
  OR2_X1 U4870 ( .A1(n3929), .A2(n3928), .ZN(n3945) );
  AOI22_X1 U4871 ( .A1(n4025), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4872 ( .A1(n4011), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3413), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3932) );
  AOI22_X1 U4873 ( .A1(n5396), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4035), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3931) );
  AOI22_X1 U4874 ( .A1(n3911), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4028), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3930) );
  NAND4_X1 U4875 ( .A1(n3933), .A2(n3932), .A3(n3931), .A4(n3930), .ZN(n3939)
         );
  AOI22_X1 U4876 ( .A1(n4006), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4034), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3937) );
  AOI22_X1 U4877 ( .A1(n4012), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3936) );
  AOI22_X1 U4878 ( .A1(n4037), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3935) );
  AOI22_X1 U4879 ( .A1(n4026), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3934) );
  NAND4_X1 U4880 ( .A1(n3937), .A2(n3936), .A3(n3935), .A4(n3934), .ZN(n3938)
         );
  NOR2_X1 U4881 ( .A1(n3939), .A2(n3938), .ZN(n3946) );
  XOR2_X1 U4882 ( .A(n3945), .B(n3946), .Z(n3942) );
  INV_X1 U4883 ( .A(EAX_REG_25__SCAN_IN), .ZN(n3940) );
  INV_X1 U4884 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5684) );
  OAI22_X1 U4885 ( .A1(n4020), .A2(n3940), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5684), .ZN(n3941) );
  AOI21_X1 U4886 ( .B1(n3942), .B2(n4022), .A(n3941), .ZN(n3944) );
  NAND2_X1 U4887 ( .A1(n3943), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3959)
         );
  XNOR2_X1 U4888 ( .A(n3959), .B(n5684), .ZN(n5534) );
  INV_X1 U4889 ( .A(n5534), .ZN(n5686) );
  MUX2_X1 U4890 ( .A(n3944), .B(n5686), .S(n4002), .Z(n5527) );
  NOR2_X1 U4891 ( .A1(n3946), .A2(n3945), .ZN(n3967) );
  AOI22_X1 U4892 ( .A1(n4006), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4034), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3950) );
  AOI22_X1 U4893 ( .A1(n4037), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3949) );
  AOI22_X1 U4894 ( .A1(n5396), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4035), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3948) );
  AOI22_X1 U4895 ( .A1(n3174), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4028), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3947) );
  NAND4_X1 U4896 ( .A1(n3950), .A2(n3949), .A3(n3948), .A4(n3947), .ZN(n3956)
         );
  AOI22_X1 U4897 ( .A1(n4026), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3954) );
  AOI22_X1 U4898 ( .A1(n4011), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3953) );
  AOI22_X1 U4899 ( .A1(n4012), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3952) );
  AOI22_X1 U4900 ( .A1(n3413), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3951) );
  NAND4_X1 U4901 ( .A1(n3954), .A2(n3953), .A3(n3952), .A4(n3951), .ZN(n3955)
         );
  OR2_X1 U4902 ( .A1(n3956), .A2(n3955), .ZN(n3966) );
  XNOR2_X1 U4903 ( .A(n3967), .B(n3966), .ZN(n3958) );
  AOI22_X1 U4904 ( .A1(n4048), .A2(EAX_REG_26__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n4969), .ZN(n3957) );
  OAI21_X1 U4905 ( .B1(n3958), .B2(n4050), .A(n3957), .ZN(n3965) );
  INV_X1 U4906 ( .A(n3959), .ZN(n3960) );
  INV_X1 U4907 ( .A(n3961), .ZN(n3963) );
  INV_X1 U4908 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3962) );
  NAND2_X1 U4909 ( .A1(n3963), .A2(n3962), .ZN(n3964) );
  NAND2_X1 U4910 ( .A1(n3996), .A2(n3964), .ZN(n5677) );
  MUX2_X1 U4911 ( .A(n3965), .B(n5677), .S(n4002), .Z(n5512) );
  NAND2_X1 U4912 ( .A1(n3967), .A2(n3966), .ZN(n3982) );
  AOI22_X1 U4913 ( .A1(n4026), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3971) );
  AOI22_X1 U4914 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4006), .B1(n4033), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3970) );
  AOI22_X1 U4915 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n3911), .B1(n4034), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3969) );
  AOI22_X1 U4916 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n4037), .B1(n3174), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3968) );
  NAND4_X1 U4917 ( .A1(n3971), .A2(n3970), .A3(n3969), .A4(n3968), .ZN(n3977)
         );
  AOI22_X1 U4918 ( .A1(n4011), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3413), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3975) );
  AOI22_X1 U4919 ( .A1(n4025), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3974) );
  AOI22_X1 U4920 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n5396), .B1(n3285), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3973) );
  AOI22_X1 U4921 ( .A1(n4035), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4028), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3972) );
  NAND4_X1 U4922 ( .A1(n3975), .A2(n3974), .A3(n3973), .A4(n3972), .ZN(n3976)
         );
  NOR2_X1 U4923 ( .A1(n3977), .A2(n3976), .ZN(n3983) );
  XOR2_X1 U4924 ( .A(n3982), .B(n3983), .Z(n3980) );
  INV_X1 U4925 ( .A(EAX_REG_27__SCAN_IN), .ZN(n3978) );
  INV_X1 U4926 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5673) );
  OAI22_X1 U4927 ( .A1(n4020), .A2(n3978), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5673), .ZN(n3979) );
  AOI21_X1 U4928 ( .B1(n3980), .B2(n4022), .A(n3979), .ZN(n3981) );
  XNOR2_X1 U4929 ( .A(n3996), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5671)
         );
  MUX2_X1 U4930 ( .A(n3981), .B(n5671), .S(n4002), .Z(n5502) );
  NOR2_X2 U4931 ( .A1(n5499), .A2(n5502), .ZN(n5486) );
  NOR2_X1 U4932 ( .A1(n3983), .A2(n3982), .ZN(n4005) );
  AOI22_X1 U4933 ( .A1(n4006), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4034), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3987) );
  AOI22_X1 U4934 ( .A1(n4037), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3986) );
  AOI22_X1 U4935 ( .A1(n5396), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4035), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3985) );
  AOI22_X1 U4936 ( .A1(n3174), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4028), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3984) );
  NAND4_X1 U4937 ( .A1(n3987), .A2(n3986), .A3(n3985), .A4(n3984), .ZN(n3993)
         );
  AOI22_X1 U4938 ( .A1(n4026), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3991) );
  AOI22_X1 U4939 ( .A1(n4011), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3990) );
  AOI22_X1 U4940 ( .A1(n4012), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3989) );
  AOI22_X1 U4941 ( .A1(n3413), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3988) );
  NAND4_X1 U4942 ( .A1(n3991), .A2(n3990), .A3(n3989), .A4(n3988), .ZN(n3992)
         );
  OR2_X1 U4943 ( .A1(n3993), .A2(n3992), .ZN(n4004) );
  XNOR2_X1 U4944 ( .A(n4005), .B(n4004), .ZN(n3995) );
  AOI22_X1 U4945 ( .A1(n4048), .A2(EAX_REG_28__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n4969), .ZN(n3994) );
  OAI21_X1 U4946 ( .B1(n3995), .B2(n4050), .A(n3994), .ZN(n4003) );
  INV_X1 U4947 ( .A(n3996), .ZN(n3997) );
  INV_X1 U4948 ( .A(n3998), .ZN(n4000) );
  INV_X1 U4949 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n3999) );
  NAND2_X1 U4950 ( .A1(n4000), .A2(n3999), .ZN(n4001) );
  NAND2_X1 U4951 ( .A1(n4052), .A2(n4001), .ZN(n5657) );
  MUX2_X1 U4952 ( .A(n4003), .B(n5657), .S(n4002), .Z(n5487) );
  NAND2_X1 U4953 ( .A1(n4005), .A2(n4004), .ZN(n4044) );
  AOI22_X1 U4954 ( .A1(n4026), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4010) );
  AOI22_X1 U4955 ( .A1(n4034), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4009) );
  AOI22_X1 U4956 ( .A1(n3911), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4035), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U4957 ( .A1(n4006), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4007) );
  NAND4_X1 U4958 ( .A1(n4010), .A2(n4009), .A3(n4008), .A4(n4007), .ZN(n4018)
         );
  AOI22_X1 U4959 ( .A1(n4011), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4016) );
  AOI22_X1 U4960 ( .A1(n4037), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3413), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4015) );
  AOI22_X1 U4961 ( .A1(n4012), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4014) );
  AOI22_X1 U4962 ( .A1(n3174), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4028), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4013) );
  NAND4_X1 U4963 ( .A1(n4016), .A2(n4015), .A3(n4014), .A4(n4013), .ZN(n4017)
         );
  NOR2_X1 U4964 ( .A1(n4018), .A2(n4017), .ZN(n4045) );
  XOR2_X1 U4965 ( .A(n4044), .B(n4045), .Z(n4023) );
  INV_X1 U4966 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4019) );
  INV_X1 U4967 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5445) );
  OAI22_X1 U4968 ( .A1(n4020), .A2(n4019), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5445), .ZN(n4021) );
  AOI21_X1 U4969 ( .B1(n4023), .B2(n4022), .A(n4021), .ZN(n4024) );
  XNOR2_X1 U4970 ( .A(n4052), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5483)
         );
  MUX2_X1 U4971 ( .A(n4024), .B(n5483), .S(n4053), .Z(n4379) );
  AOI22_X1 U4972 ( .A1(n4026), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4032) );
  AOI22_X1 U4973 ( .A1(n4012), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4031) );
  AOI22_X1 U4974 ( .A1(n4027), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4030) );
  AOI22_X1 U4975 ( .A1(n4006), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4028), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4029) );
  NAND4_X1 U4976 ( .A1(n4032), .A2(n4031), .A3(n4030), .A4(n4029), .ZN(n4043)
         );
  AOI22_X1 U4977 ( .A1(n3413), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4041) );
  AOI22_X1 U4978 ( .A1(n4034), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4040) );
  AOI22_X1 U4979 ( .A1(n3911), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4035), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4039) );
  AOI22_X1 U4980 ( .A1(n4037), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4038) );
  NAND4_X1 U4981 ( .A1(n4041), .A2(n4040), .A3(n4039), .A4(n4038), .ZN(n4042)
         );
  NOR2_X1 U4982 ( .A1(n4043), .A2(n4042), .ZN(n4047) );
  NOR2_X1 U4983 ( .A1(n4045), .A2(n4044), .ZN(n4046) );
  XOR2_X1 U4984 ( .A(n4047), .B(n4046), .Z(n4051) );
  AOI22_X1 U4985 ( .A1(n4048), .A2(EAX_REG_30__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n4969), .ZN(n4049) );
  OAI21_X1 U4986 ( .B1(n4051), .B2(n4050), .A(n4049), .ZN(n4054) );
  XNOR2_X1 U4987 ( .A(n4401), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5421)
         );
  MUX2_X1 U4988 ( .A(n4054), .B(n5421), .S(n4053), .Z(n4055) );
  NAND2_X1 U4989 ( .A1(n6586), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4074) );
  NAND2_X1 U4990 ( .A1(n4057), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4058) );
  NAND2_X1 U4991 ( .A1(n4074), .A2(n4058), .ZN(n4073) );
  NAND2_X1 U4992 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6580), .ZN(n4072) );
  INV_X1 U4993 ( .A(n4072), .ZN(n4060) );
  XNOR2_X1 U4994 ( .A(n4073), .B(n4060), .ZN(n4414) );
  NAND2_X1 U4995 ( .A1(n4113), .A2(n3398), .ZN(n4059) );
  NAND2_X1 U4996 ( .A1(n4059), .A2(n3776), .ZN(n4069) );
  AOI21_X1 U4997 ( .B1(n4061), .B2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n4060), 
        .ZN(n4063) );
  NAND2_X1 U4998 ( .A1(n4113), .A2(n4063), .ZN(n4062) );
  NAND2_X1 U4999 ( .A1(n4104), .A2(n4062), .ZN(n4068) );
  NAND2_X1 U5000 ( .A1(n4608), .A2(n3776), .ZN(n4347) );
  AOI21_X1 U5001 ( .B1(n4347), .B2(n4063), .A(n3158), .ZN(n4066) );
  NAND2_X1 U5002 ( .A1(n4620), .A2(n3776), .ZN(n4065) );
  NAND2_X1 U5003 ( .A1(n5227), .A2(n4065), .ZN(n4087) );
  OR2_X1 U5004 ( .A1(n4066), .A2(n4087), .ZN(n4067) );
  OAI211_X1 U5005 ( .C1(n4069), .C2(n4414), .A(n4068), .B(n4067), .ZN(n4071)
         );
  NAND3_X1 U5006 ( .A1(n4069), .A2(STATE2_REG_0__SCAN_IN), .A3(n4414), .ZN(
        n4070) );
  OAI211_X1 U5007 ( .C1(n4104), .C2(n4414), .A(n4071), .B(n4070), .ZN(n4085)
         );
  NAND2_X1 U5008 ( .A1(n4075), .A2(n4074), .ZN(n4080) );
  INV_X1 U5009 ( .A(n4080), .ZN(n4078) );
  NAND2_X1 U5010 ( .A1(n6590), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4089) );
  NAND2_X1 U5011 ( .A1(n3168), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4076) );
  INV_X1 U5012 ( .A(n4079), .ZN(n4077) );
  NAND2_X1 U5013 ( .A1(n4078), .A2(n4077), .ZN(n4081) );
  NAND2_X1 U5014 ( .A1(n4080), .A2(n4079), .ZN(n4090) );
  AND2_X1 U5015 ( .A1(n4081), .A2(n4090), .ZN(n4416) );
  INV_X1 U5016 ( .A(n4098), .ZN(n4083) );
  INV_X1 U5017 ( .A(n4087), .ZN(n4082) );
  NAND2_X1 U5018 ( .A1(n4113), .A2(n4416), .ZN(n4086) );
  OAI211_X1 U5019 ( .C1(n4416), .C2(n4083), .A(n4082), .B(n4086), .ZN(n4084)
         );
  NAND2_X1 U5020 ( .A1(n4085), .A2(n4084), .ZN(n4101) );
  INV_X1 U5021 ( .A(n4086), .ZN(n4088) );
  NAND2_X1 U5022 ( .A1(n4088), .A2(n4087), .ZN(n4100) );
  NAND2_X1 U5023 ( .A1(n4090), .A2(n4089), .ZN(n4095) );
  XNOR2_X1 U5024 ( .A(n4559), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4093)
         );
  NAND2_X1 U5025 ( .A1(n4095), .A2(n4093), .ZN(n4092) );
  NAND2_X1 U5026 ( .A1(n6594), .A2(n4559), .ZN(n4091) );
  NAND2_X1 U5027 ( .A1(n4092), .A2(n4091), .ZN(n4105) );
  NAND2_X1 U5028 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n6031), .ZN(n4106) );
  OR2_X1 U5029 ( .A1(n4105), .A2(n4106), .ZN(n4097) );
  INV_X1 U5030 ( .A(n4093), .ZN(n4094) );
  XNOR2_X1 U5031 ( .A(n4095), .B(n4094), .ZN(n4096) );
  NOR2_X1 U5032 ( .A1(n4413), .A2(n4098), .ZN(n4099) );
  AOI21_X1 U5033 ( .B1(n4101), .B2(n4100), .A(n4099), .ZN(n4103) );
  OAI22_X1 U5034 ( .A1(n4104), .A2(n4413), .B1(STATE2_REG_0__SCAN_IN), .B2(
        n6031), .ZN(n4102) );
  INV_X1 U5035 ( .A(n4104), .ZN(n4110) );
  INV_X1 U5036 ( .A(n4105), .ZN(n4109) );
  NAND2_X1 U5037 ( .A1(n6454), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4108) );
  INV_X1 U5038 ( .A(n4106), .ZN(n4107) );
  NAND2_X1 U5039 ( .A1(n4110), .A2(n4418), .ZN(n4111) );
  NAND2_X1 U5040 ( .A1(n4418), .A2(n4113), .ZN(n4114) );
  INV_X1 U5041 ( .A(n4471), .ZN(n4423) );
  AND2_X1 U5042 ( .A1(n3394), .A2(n3366), .ZN(n4513) );
  INV_X1 U5043 ( .A(n4513), .ZN(n4116) );
  AND2_X1 U5044 ( .A1(n4473), .A2(n4116), .ZN(n4511) );
  OR2_X1 U5045 ( .A1(n4511), .A2(n4117), .ZN(n4121) );
  INV_X1 U5046 ( .A(n6271), .ZN(n6693) );
  NAND2_X1 U5047 ( .A1(n3389), .A2(n3436), .ZN(n4119) );
  NAND2_X1 U5048 ( .A1(n6693), .A2(n4119), .ZN(n4120) );
  NAND2_X1 U5049 ( .A1(n4121), .A2(n4120), .ZN(n4445) );
  NAND2_X1 U5050 ( .A1(n4122), .A2(n5557), .ZN(n4126) );
  NAND2_X1 U5051 ( .A1(n3158), .A2(n3398), .ZN(n5232) );
  OR2_X1 U5052 ( .A1(n5232), .A2(n4465), .ZN(n4448) );
  NOR2_X1 U5053 ( .A1(n4473), .A2(n3436), .ZN(n4123) );
  NAND2_X1 U5054 ( .A1(n4448), .A2(n4123), .ZN(n4124) );
  NAND2_X1 U5055 ( .A1(n4625), .A2(n4244), .ZN(n4344) );
  NAND2_X1 U5056 ( .A1(n4124), .A2(n4344), .ZN(n4125) );
  NAND2_X1 U5057 ( .A1(n4128), .A2(n4127), .ZN(n4483) );
  OR2_X1 U5058 ( .A1(n5919), .A2(n4620), .ZN(n4470) );
  NAND2_X1 U5059 ( .A1(n4423), .A2(n4544), .ZN(n4451) );
  NAND2_X1 U5060 ( .A1(n3436), .A2(n3398), .ZN(n4133) );
  INV_X1 U5061 ( .A(n3366), .ZN(n5450) );
  AND3_X1 U5062 ( .A1(n3365), .A2(n5450), .A3(n4608), .ZN(n4503) );
  NAND3_X1 U5063 ( .A1(n4129), .A2(n4490), .A3(n4503), .ZN(n4130) );
  NAND2_X1 U5064 ( .A1(n4451), .A2(n4130), .ZN(n4132) );
  OR2_X1 U5065 ( .A1(n4219), .A2(EBX_REG_17__SCAN_IN), .ZN(n4136) );
  NAND2_X1 U5066 ( .A1(n4150), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4134) );
  OAI211_X1 U5067 ( .C1(n4159), .C2(EBX_REG_17__SCAN_IN), .A(n4157), .B(n4134), 
        .ZN(n4135) );
  NAND2_X1 U5068 ( .A1(n4136), .A2(n4135), .ZN(n5571) );
  OR2_X1 U5069 ( .A1(n4219), .A2(EBX_REG_15__SCAN_IN), .ZN(n4139) );
  NAND2_X1 U5070 ( .A1(n4150), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4137) );
  OAI211_X1 U5071 ( .C1(n4159), .C2(EBX_REG_15__SCAN_IN), .A(n4157), .B(n4137), 
        .ZN(n4138) );
  NAND2_X1 U5072 ( .A1(n4139), .A2(n4138), .ZN(n5358) );
  NAND2_X1 U5073 ( .A1(n5557), .A2(EBX_REG_9__SCAN_IN), .ZN(n4141) );
  OR2_X1 U5074 ( .A1(n4219), .A2(EBX_REG_9__SCAN_IN), .ZN(n4140) );
  OAI211_X1 U5075 ( .C1(n5464), .C2(INSTADDRPOINTER_REG_9__SCAN_IN), .A(n4141), 
        .B(n4140), .ZN(n5260) );
  INV_X1 U5076 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5453) );
  NAND2_X1 U5077 ( .A1(n4157), .A2(n5453), .ZN(n4142) );
  OAI211_X1 U5078 ( .C1(n4133), .C2(EBX_REG_1__SCAN_IN), .A(n4142), .B(n4150), 
        .ZN(n4143) );
  INV_X1 U5079 ( .A(n4147), .ZN(n4149) );
  NAND2_X1 U5080 ( .A1(n4157), .A2(EBX_REG_0__SCAN_IN), .ZN(n4146) );
  INV_X1 U5081 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4144) );
  NAND2_X1 U5082 ( .A1(n4150), .A2(n4144), .ZN(n4145) );
  AND2_X1 U5083 ( .A1(n4146), .A2(n4145), .ZN(n4534) );
  INV_X1 U5084 ( .A(n4534), .ZN(n4148) );
  OR2_X1 U5085 ( .A1(n4224), .A2(EBX_REG_2__SCAN_IN), .ZN(n4153) );
  INV_X1 U5086 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4258) );
  NAND2_X1 U5087 ( .A1(n4157), .A2(n4258), .ZN(n4151) );
  OAI211_X1 U5088 ( .C1(n4159), .C2(EBX_REG_2__SCAN_IN), .A(n4151), .B(n4150), 
        .ZN(n4152) );
  NAND2_X1 U5089 ( .A1(n4153), .A2(n4152), .ZN(n4644) );
  OR2_X1 U5090 ( .A1(n4219), .A2(EBX_REG_3__SCAN_IN), .ZN(n4156) );
  NAND2_X1 U5091 ( .A1(n4150), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4154)
         );
  OAI211_X1 U5092 ( .C1(n4159), .C2(EBX_REG_3__SCAN_IN), .A(n4157), .B(n4154), 
        .ZN(n4155) );
  NAND2_X1 U5093 ( .A1(n4156), .A2(n4155), .ZN(n4530) );
  INV_X1 U5094 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4158) );
  INV_X1 U5095 ( .A(n4157), .ZN(n4213) );
  OAI21_X1 U5096 ( .B1(n4157), .B2(n4158), .A(n4193), .ZN(n4162) );
  NAND2_X1 U5097 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n4159), .ZN(n4160)
         );
  OAI21_X1 U5098 ( .B1(n4224), .B2(EBX_REG_4__SCAN_IN), .A(n4160), .ZN(n4161)
         );
  NAND2_X1 U5099 ( .A1(n5557), .A2(EBX_REG_5__SCAN_IN), .ZN(n4164) );
  OR2_X1 U5100 ( .A1(n4219), .A2(EBX_REG_5__SCAN_IN), .ZN(n4163) );
  OAI211_X1 U5101 ( .C1(n5464), .C2(INSTADDRPOINTER_REG_5__SCAN_IN), .A(n4164), 
        .B(n4163), .ZN(n4770) );
  INV_X1 U5102 ( .A(EBX_REG_6__SCAN_IN), .ZN(n5018) );
  OAI21_X1 U5103 ( .B1(n4157), .B2(n5018), .A(n4193), .ZN(n4167) );
  NAND2_X1 U5104 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4159), .ZN(n4165)
         );
  OAI21_X1 U5105 ( .B1(n4224), .B2(EBX_REG_6__SCAN_IN), .A(n4165), .ZN(n4166)
         );
  NAND2_X1 U5106 ( .A1(n4890), .A2(n4892), .ZN(n5213) );
  OR2_X1 U5107 ( .A1(n4219), .A2(EBX_REG_7__SCAN_IN), .ZN(n4170) );
  NAND2_X1 U5108 ( .A1(n4150), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4168)
         );
  OAI211_X1 U5109 ( .C1(n4159), .C2(EBX_REG_7__SCAN_IN), .A(n4157), .B(n4168), 
        .ZN(n4169) );
  NAND2_X1 U5110 ( .A1(n4170), .A2(n4169), .ZN(n5215) );
  OR2_X1 U5111 ( .A1(n4224), .A2(EBX_REG_8__SCAN_IN), .ZN(n4173) );
  INV_X1 U5112 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4319) );
  NAND2_X1 U5113 ( .A1(n4157), .A2(n4319), .ZN(n4171) );
  OAI211_X1 U5114 ( .C1(n4159), .C2(EBX_REG_8__SCAN_IN), .A(n4171), .B(n4150), 
        .ZN(n4172) );
  NAND2_X1 U5115 ( .A1(n4173), .A2(n4172), .ZN(n5148) );
  INV_X1 U5116 ( .A(n4193), .ZN(n4174) );
  AOI21_X1 U5117 ( .B1(n4213), .B2(EBX_REG_10__SCAN_IN), .A(n4174), .ZN(n4176)
         );
  NAND2_X1 U5118 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n4159), .ZN(n4175) );
  OAI211_X1 U5119 ( .C1(EBX_REG_10__SCAN_IN), .C2(n4224), .A(n4176), .B(n4175), 
        .ZN(n5272) );
  OR2_X1 U5120 ( .A1(n4219), .A2(EBX_REG_11__SCAN_IN), .ZN(n4179) );
  NAND2_X1 U5121 ( .A1(n4150), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4177) );
  OAI211_X1 U5122 ( .C1(n4159), .C2(EBX_REG_11__SCAN_IN), .A(n4157), .B(n4177), 
        .ZN(n4178) );
  NAND2_X1 U5123 ( .A1(n4179), .A2(n4178), .ZN(n6112) );
  INV_X1 U5124 ( .A(EBX_REG_12__SCAN_IN), .ZN(n4180) );
  OAI21_X1 U5125 ( .B1(n4157), .B2(n4180), .A(n4193), .ZN(n4183) );
  NAND2_X1 U5126 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n4159), .ZN(n4181) );
  OAI21_X1 U5127 ( .B1(n4224), .B2(EBX_REG_12__SCAN_IN), .A(n4181), .ZN(n4182)
         );
  OR2_X1 U5128 ( .A1(n4219), .A2(EBX_REG_13__SCAN_IN), .ZN(n4186) );
  NAND2_X1 U5129 ( .A1(n4150), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4184) );
  OAI211_X1 U5130 ( .C1(n4159), .C2(EBX_REG_13__SCAN_IN), .A(n4157), .B(n4184), 
        .ZN(n4185) );
  NAND2_X1 U5131 ( .A1(n4186), .A2(n4185), .ZN(n5338) );
  INV_X1 U5132 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5353) );
  OAI21_X1 U5133 ( .B1(n4157), .B2(n5353), .A(n4193), .ZN(n4189) );
  NAND2_X1 U5134 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n4159), .ZN(n4187) );
  OAI21_X1 U5135 ( .B1(n4224), .B2(EBX_REG_14__SCAN_IN), .A(n4187), .ZN(n4188)
         );
  INV_X1 U5136 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5633) );
  OAI21_X1 U5137 ( .B1(n4157), .B2(n5633), .A(n4193), .ZN(n4192) );
  NAND2_X1 U5138 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n4159), .ZN(n4190) );
  OAI21_X1 U5139 ( .B1(n4224), .B2(EBX_REG_16__SCAN_IN), .A(n4190), .ZN(n4191)
         );
  NOR2_X4 U5140 ( .A1(n5571), .A2(n5628), .ZN(n5617) );
  AOI22_X1 U5141 ( .A1(n4213), .A2(EBX_REG_19__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n4159), .ZN(n4194) );
  OAI211_X1 U5142 ( .C1(EBX_REG_19__SCAN_IN), .C2(n4224), .A(n4194), .B(n4193), 
        .ZN(n5615) );
  OR2_X1 U5143 ( .A1(n5464), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4195)
         );
  INV_X1 U5144 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5623) );
  NAND2_X1 U5145 ( .A1(n4490), .A2(n5623), .ZN(n5612) );
  OAI22_X1 U5146 ( .A1(n5464), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        EBX_REG_20__SCAN_IN), .B2(n4159), .ZN(n5558) );
  NAND2_X1 U5147 ( .A1(n5611), .A2(n5558), .ZN(n4197) );
  NAND2_X1 U5148 ( .A1(n5557), .A2(EBX_REG_20__SCAN_IN), .ZN(n4196) );
  OAI211_X1 U5149 ( .C1(n5611), .C2(n5557), .A(n4197), .B(n4196), .ZN(n4198)
         );
  INV_X1 U5150 ( .A(n4198), .ZN(n4199) );
  INV_X1 U5151 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5603) );
  OR2_X1 U5152 ( .A1(n4219), .A2(EBX_REG_21__SCAN_IN), .ZN(n4201) );
  OR2_X1 U5153 ( .A1(n5464), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4200)
         );
  OAI211_X1 U5154 ( .C1(n5603), .C2(n4150), .A(n4201), .B(n4200), .ZN(n5600)
         );
  OR2_X1 U5155 ( .A1(n4219), .A2(EBX_REG_23__SCAN_IN), .ZN(n4204) );
  NAND2_X1 U5156 ( .A1(n4150), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4202) );
  OAI211_X1 U5157 ( .C1(n4159), .C2(EBX_REG_23__SCAN_IN), .A(n4157), .B(n4202), 
        .ZN(n4203) );
  AND2_X1 U5158 ( .A1(n4204), .A2(n4203), .ZN(n5591) );
  INV_X1 U5159 ( .A(n4224), .ZN(n4384) );
  INV_X1 U5160 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5982) );
  NAND2_X1 U5161 ( .A1(n4384), .A2(n5982), .ZN(n4208) );
  INV_X1 U5162 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4205) );
  NAND2_X1 U5163 ( .A1(n4157), .A2(n4205), .ZN(n4206) );
  OAI211_X1 U5164 ( .C1(n4133), .C2(EBX_REG_22__SCAN_IN), .A(n4206), .B(n4150), 
        .ZN(n4207) );
  NAND2_X1 U5165 ( .A1(n4208), .A2(n4207), .ZN(n5833) );
  NAND2_X1 U5166 ( .A1(n5591), .A2(n5833), .ZN(n4209) );
  OR2_X1 U5167 ( .A1(n4219), .A2(EBX_REG_25__SCAN_IN), .ZN(n4212) );
  NAND2_X1 U5168 ( .A1(n4150), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4210) );
  OAI211_X1 U5169 ( .C1(n4159), .C2(EBX_REG_25__SCAN_IN), .A(n4157), .B(n4210), 
        .ZN(n4211) );
  AND2_X1 U5170 ( .A1(n4212), .A2(n4211), .ZN(n5531) );
  AOI22_X1 U5171 ( .A1(n4213), .A2(EBX_REG_24__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n4159), .ZN(n4215) );
  INV_X1 U5172 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5587) );
  NAND2_X1 U5173 ( .A1(n4384), .A2(n5587), .ZN(n4214) );
  NAND2_X1 U5174 ( .A1(n4215), .A2(n4214), .ZN(n5532) );
  AND2_X1 U5175 ( .A1(n5531), .A2(n5532), .ZN(n4216) );
  INV_X1 U5176 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5823) );
  NAND2_X1 U5177 ( .A1(n4157), .A2(n5823), .ZN(n4217) );
  OAI211_X1 U5178 ( .C1(EBX_REG_26__SCAN_IN), .C2(n4159), .A(n4217), .B(n4150), 
        .ZN(n4218) );
  OAI21_X1 U5179 ( .B1(n4224), .B2(EBX_REG_26__SCAN_IN), .A(n4218), .ZN(n5515)
         );
  INV_X1 U5180 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5581) );
  OR2_X1 U5181 ( .A1(n4219), .A2(EBX_REG_27__SCAN_IN), .ZN(n4221) );
  OR2_X1 U5182 ( .A1(n5464), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4220)
         );
  OAI211_X1 U5183 ( .C1(n5581), .C2(n4150), .A(n4221), .B(n4220), .ZN(n5503)
         );
  INV_X1 U5184 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5796) );
  NAND2_X1 U5185 ( .A1(n4157), .A2(n5796), .ZN(n4222) );
  OAI211_X1 U5186 ( .C1(EBX_REG_28__SCAN_IN), .C2(n4133), .A(n4222), .B(n4150), 
        .ZN(n4223) );
  OAI21_X1 U5187 ( .B1(n4224), .B2(EBX_REG_28__SCAN_IN), .A(n4223), .ZN(n5489)
         );
  OR2_X1 U5188 ( .A1(n5464), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4226)
         );
  INV_X1 U5189 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5479) );
  NAND2_X1 U5190 ( .A1(n4490), .A2(n5479), .ZN(n4225) );
  NAND2_X1 U5191 ( .A1(n4226), .A2(n4225), .ZN(n4387) );
  INV_X1 U5192 ( .A(n5491), .ZN(n4227) );
  NAND2_X1 U5193 ( .A1(n4385), .A2(n4227), .ZN(n4231) );
  NAND2_X1 U5194 ( .A1(n5464), .A2(EBX_REG_30__SCAN_IN), .ZN(n4229) );
  NAND2_X1 U5195 ( .A1(n4159), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4228) );
  AND2_X1 U5196 ( .A1(n4229), .A2(n4228), .ZN(n5466) );
  INV_X1 U5197 ( .A(n5466), .ZN(n4230) );
  NAND2_X1 U5198 ( .A1(n4231), .A2(n4230), .ZN(n4232) );
  NAND2_X1 U5199 ( .A1(n5491), .A2(n5557), .ZN(n4233) );
  NAND3_X1 U5200 ( .A1(n4385), .A2(n5466), .A3(n4233), .ZN(n4234) );
  NAND2_X1 U5201 ( .A1(n4235), .A2(n4234), .ZN(n5790) );
  INV_X2 U5202 ( .A(n5980), .ZN(n6233) );
  INV_X1 U5203 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5417) );
  OR2_X1 U5204 ( .A1(n6238), .A2(n5417), .ZN(n4236) );
  NOR2_X1 U5205 ( .A1(n4344), .A2(n3394), .ZN(n4241) );
  NAND2_X1 U5206 ( .A1(n4239), .A2(n4245), .ZN(n4250) );
  OAI211_X1 U5207 ( .C1(n4239), .C2(n4245), .A(n6271), .B(n4250), .ZN(n4240)
         );
  AND2_X1 U5208 ( .A1(n4241), .A2(n4240), .ZN(n4242) );
  NAND2_X1 U5209 ( .A1(n4243), .A2(n4242), .ZN(n4463) );
  INV_X1 U5210 ( .A(n4056), .ZN(n4310) );
  NAND2_X1 U5211 ( .A1(n3158), .A2(n4244), .ZN(n4252) );
  OAI21_X1 U5212 ( .B1(n6693), .B2(n4245), .A(n4252), .ZN(n4246) );
  INV_X1 U5213 ( .A(n4246), .ZN(n4247) );
  NAND2_X1 U5214 ( .A1(n4463), .A2(n4464), .ZN(n4462) );
  OR2_X1 U5215 ( .A1(n5766), .A2(n5453), .ZN(n4248) );
  INV_X1 U5216 ( .A(n4249), .ZN(n4251) );
  NAND2_X1 U5217 ( .A1(n4250), .A2(n4251), .ZN(n4270) );
  OAI21_X1 U5218 ( .B1(n4251), .B2(n4250), .A(n4270), .ZN(n4254) );
  INV_X1 U5219 ( .A(n4252), .ZN(n4253) );
  AOI21_X1 U5220 ( .B1(n4254), .B2(n6271), .A(n4253), .ZN(n4255) );
  NAND2_X1 U5221 ( .A1(n4256), .A2(n4255), .ZN(n4257) );
  NAND2_X1 U5222 ( .A1(n4257), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6375)
         );
  NAND2_X1 U5223 ( .A1(n6374), .A2(n6375), .ZN(n4260) );
  INV_X1 U5224 ( .A(n4257), .ZN(n4259) );
  NAND2_X1 U5225 ( .A1(n4259), .A2(n4258), .ZN(n6376) );
  NAND2_X1 U5226 ( .A1(n4650), .A2(n4056), .ZN(n4264) );
  INV_X1 U5227 ( .A(n4269), .ZN(n4261) );
  XNOR2_X1 U5228 ( .A(n4270), .B(n4261), .ZN(n4262) );
  NAND2_X1 U5229 ( .A1(n4262), .A2(n6271), .ZN(n4263) );
  INV_X1 U5230 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4265) );
  XNOR2_X1 U5231 ( .A(n4266), .B(n4265), .ZN(n4527) );
  NAND2_X1 U5232 ( .A1(n4526), .A2(n4527), .ZN(n4268) );
  NAND2_X1 U5233 ( .A1(n4266), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4267)
         );
  NAND2_X1 U5234 ( .A1(n4268), .A2(n4267), .ZN(n4575) );
  NAND2_X1 U5235 ( .A1(n4270), .A2(n4269), .ZN(n4272) );
  INV_X1 U5236 ( .A(n4272), .ZN(n4274) );
  INV_X1 U5237 ( .A(n4273), .ZN(n4271) );
  OR2_X1 U5238 ( .A1(n4272), .A2(n4271), .ZN(n4292) );
  OAI211_X1 U5239 ( .C1(n4274), .C2(n4273), .A(n6271), .B(n4292), .ZN(n4275)
         );
  OAI21_X2 U5240 ( .B1(n4276), .B2(n4310), .A(n4275), .ZN(n4278) );
  INV_X1 U5241 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4277) );
  XNOR2_X1 U5242 ( .A(n4278), .B(n4277), .ZN(n4576) );
  NAND2_X1 U5243 ( .A1(n4575), .A2(n4576), .ZN(n4280) );
  NAND2_X1 U5244 ( .A1(n4278), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4279)
         );
  NAND2_X1 U5245 ( .A1(n4280), .A2(n4279), .ZN(n4998) );
  NAND2_X1 U5246 ( .A1(n4281), .A2(n4056), .ZN(n4284) );
  XNOR2_X1 U5247 ( .A(n4292), .B(n4290), .ZN(n4282) );
  NAND2_X1 U5248 ( .A1(n4282), .A2(n6271), .ZN(n4283) );
  NAND2_X1 U5249 ( .A1(n4284), .A2(n4283), .ZN(n4286) );
  INV_X1 U5250 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4285) );
  XNOR2_X1 U5251 ( .A(n4286), .B(n4285), .ZN(n4999) );
  NAND2_X1 U5252 ( .A1(n4998), .A2(n4999), .ZN(n4288) );
  NAND2_X1 U5253 ( .A1(n4286), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4287)
         );
  NAND2_X1 U5254 ( .A1(n4289), .A2(n4056), .ZN(n4296) );
  INV_X1 U5255 ( .A(n4290), .ZN(n4291) );
  NOR2_X1 U5256 ( .A1(n4292), .A2(n4291), .ZN(n4294) );
  NAND2_X1 U5257 ( .A1(n4294), .A2(n4293), .ZN(n4317) );
  OAI211_X1 U5258 ( .C1(n4294), .C2(n4293), .A(n4317), .B(n6271), .ZN(n4295)
         );
  NAND2_X1 U5259 ( .A1(n4296), .A2(n4295), .ZN(n4298) );
  INV_X1 U5260 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4297) );
  XNOR2_X1 U5261 ( .A(n4298), .B(n4297), .ZN(n4889) );
  NAND2_X1 U5262 ( .A1(n4888), .A2(n4889), .ZN(n4300) );
  NAND2_X1 U5263 ( .A1(n4298), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4299)
         );
  NAND2_X1 U5264 ( .A1(n4300), .A2(n4299), .ZN(n5211) );
  NAND2_X1 U5265 ( .A1(n4301), .A2(n4056), .ZN(n4304) );
  XNOR2_X1 U5266 ( .A(n4317), .B(n4315), .ZN(n4302) );
  NAND2_X1 U5267 ( .A1(n4302), .A2(n6271), .ZN(n4303) );
  NAND2_X1 U5268 ( .A1(n4304), .A2(n4303), .ZN(n4306) );
  INV_X1 U5269 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4305) );
  NAND2_X1 U5270 ( .A1(n5211), .A2(n5212), .ZN(n4308) );
  NAND2_X1 U5271 ( .A1(n4306), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4307)
         );
  NAND2_X1 U5272 ( .A1(n4308), .A2(n4307), .ZN(n5141) );
  INV_X1 U5273 ( .A(n4309), .ZN(n4311) );
  NAND2_X1 U5274 ( .A1(n6271), .A2(n4315), .ZN(n4316) );
  OR2_X1 U5275 ( .A1(n4317), .A2(n4316), .ZN(n4318) );
  NAND2_X1 U5276 ( .A1(n5729), .A2(n4318), .ZN(n4320) );
  XNOR2_X1 U5277 ( .A(n4320), .B(n4319), .ZN(n5142) );
  NAND2_X1 U5278 ( .A1(n4320), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4321)
         );
  INV_X1 U5279 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6422) );
  NAND2_X1 U5280 ( .A1(n5729), .A2(n6422), .ZN(n4322) );
  INV_X1 U5281 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6414) );
  AND2_X1 U5282 ( .A1(n5729), .A2(n6414), .ZN(n5281) );
  NAND2_X1 U5283 ( .A1(n4314), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5282) );
  INV_X1 U5284 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6400) );
  NAND2_X1 U5285 ( .A1(n5729), .A2(n6400), .ZN(n6348) );
  NAND2_X1 U5286 ( .A1(n4314), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6349) );
  INV_X1 U5287 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4324) );
  NOR2_X1 U5288 ( .A1(n5733), .A2(n4324), .ZN(n5309) );
  XNOR2_X1 U5289 ( .A(n5733), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5330)
         );
  NAND2_X1 U5290 ( .A1(n5331), .A2(n5330), .ZN(n5329) );
  INV_X1 U5291 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5335) );
  NAND2_X1 U5292 ( .A1(n5729), .A2(n5335), .ZN(n4325) );
  NAND2_X1 U5293 ( .A1(n5329), .A2(n4325), .ZN(n5361) );
  INV_X1 U5294 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5367) );
  NAND2_X1 U5295 ( .A1(n5729), .A2(n5367), .ZN(n4327) );
  XNOR2_X1 U5296 ( .A(n5733), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5753)
         );
  INV_X1 U5297 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4329) );
  NAND2_X1 U5298 ( .A1(n5729), .A2(n4329), .ZN(n4330) );
  INV_X1 U5299 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5734) );
  INV_X1 U5300 ( .A(n5730), .ZN(n4333) );
  AND2_X1 U5301 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5863) );
  INV_X1 U5302 ( .A(n5863), .ZN(n4332) );
  NAND2_X1 U5303 ( .A1(n4314), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5745) );
  OAI21_X1 U5304 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .A(n4314), .ZN(n4334) );
  AND2_X1 U5305 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5435) );
  AND2_X1 U5306 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5836) );
  AND2_X1 U5307 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5864) );
  NAND3_X1 U5308 ( .A1(n5435), .A2(n5836), .A3(n5864), .ZN(n4336) );
  NAND2_X1 U5309 ( .A1(n5729), .A2(n4336), .ZN(n4339) );
  NOR2_X1 U5310 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5865) );
  NOR2_X1 U5311 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5837) );
  INV_X1 U5312 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5390) );
  INV_X1 U5313 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5825) );
  AND4_X1 U5314 ( .A1(n5865), .A2(n5837), .A3(n5390), .A4(n5825), .ZN(n4337)
         );
  NOR2_X1 U5315 ( .A1(n5729), .A2(n4337), .ZN(n4338) );
  XNOR2_X1 U5316 ( .A(n5733), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5687)
         );
  INV_X1 U5317 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U5318 ( .A1(n5729), .A2(n5661), .ZN(n4340) );
  NAND2_X1 U5319 ( .A1(n4394), .A2(n4340), .ZN(n4341) );
  OR3_X2 U5320 ( .A1(n4341), .A2(n4314), .A3(n5823), .ZN(n5669) );
  NAND2_X1 U5321 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5437) );
  NOR2_X4 U5322 ( .A1(n5669), .A2(n5437), .ZN(n5429) );
  BUF_X2 U5323 ( .A(n4341), .Z(n5680) );
  INV_X1 U5324 ( .A(n4395), .ZN(n4342) );
  NAND2_X2 U5325 ( .A1(n5680), .A2(n4342), .ZN(n5427) );
  NOR2_X1 U5326 ( .A1(n5427), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5426)
         );
  AOI21_X1 U5327 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5429), .A(n5426), 
        .ZN(n4343) );
  XNOR2_X2 U5328 ( .A(n4343), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5784)
         );
  NAND2_X1 U5329 ( .A1(n5919), .A2(n3158), .ZN(n4346) );
  NOR2_X1 U5330 ( .A1(n4122), .A2(n4344), .ZN(n4345) );
  INV_X1 U5331 ( .A(n4347), .ZN(n4348) );
  NAND2_X1 U5332 ( .A1(n5784), .A2(n6387), .ZN(n4359) );
  NAND3_X1 U5333 ( .A1(n6613), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6627) );
  NAND2_X1 U5334 ( .A1(n4349), .A2(n6519), .ZN(n6691) );
  NAND2_X1 U5335 ( .A1(n6691), .A2(n6613), .ZN(n4350) );
  NAND2_X1 U5336 ( .A1(n6613), .A2(n4969), .ZN(n6626) );
  INV_X1 U5337 ( .A(n6626), .ZN(n4351) );
  INV_X1 U5338 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6900) );
  NOR2_X1 U5339 ( .A1(n6392), .A2(n6900), .ZN(n5785) );
  NAND2_X1 U5340 ( .A1(n6613), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4353) );
  NAND2_X1 U5341 ( .A1(n6786), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4352) );
  NAND2_X1 U5342 ( .A1(n4353), .A2(n4352), .ZN(n5768) );
  NOR2_X1 U5343 ( .A1(n6391), .A2(n5421), .ZN(n4354) );
  AOI211_X1 U5344 ( .C1(n6383), .C2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5785), 
        .B(n4354), .ZN(n4355) );
  OAI21_X1 U5345 ( .B1(n4356), .B2(n6359), .A(n4355), .ZN(n4357) );
  INV_X1 U5346 ( .A(n4357), .ZN(n4358) );
  NAND2_X1 U5347 ( .A1(n4359), .A2(n4358), .ZN(U2956) );
  INV_X1 U5348 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5874) );
  OAI21_X1 U5349 ( .B1(n4361), .B2(n5874), .A(n5733), .ZN(n4362) );
  INV_X1 U5350 ( .A(n5717), .ZN(n4364) );
  INV_X1 U5351 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5861) );
  XNOR2_X1 U5352 ( .A(n5733), .B(n5861), .ZN(n5716) );
  NAND2_X1 U5353 ( .A1(n4314), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4365) );
  INV_X1 U5354 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5844) );
  XNOR2_X1 U5355 ( .A(n5733), .B(n5844), .ZN(n5711) );
  NAND2_X1 U5356 ( .A1(n3236), .A2(n4366), .ZN(n5701) );
  NAND3_X1 U5357 ( .A1(n5729), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4367) );
  NOR2_X1 U5358 ( .A1(n5733), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5702)
         );
  INV_X1 U5359 ( .A(n5693), .ZN(n4368) );
  NAND2_X1 U5360 ( .A1(n4370), .A2(n4369), .ZN(n4371) );
  XNOR2_X1 U5361 ( .A(n4371), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5394)
         );
  XOR2_X1 U5362 ( .A(n4373), .B(n4372), .Z(n5586) );
  NAND2_X1 U5363 ( .A1(n5586), .A2(n6379), .ZN(n4376) );
  INV_X1 U5364 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6922) );
  NOR2_X1 U5365 ( .A1(n6392), .A2(n6922), .ZN(n5392) );
  NOR2_X1 U5366 ( .A1(n6372), .A2(n5544), .ZN(n4374) );
  AOI211_X1 U5367 ( .C1(n5547), .C2(n6366), .A(n5392), .B(n4374), .ZN(n4375)
         );
  OAI21_X1 U5368 ( .B1(n5394), .B2(n6357), .A(n4377), .ZN(U2962) );
  NAND2_X1 U5369 ( .A1(n4378), .A2(n4379), .ZN(n4382) );
  INV_X1 U5370 ( .A(n4380), .ZN(n4381) );
  NAND2_X1 U5371 ( .A1(n5634), .A2(n4383), .ZN(n4393) );
  NAND2_X1 U5372 ( .A1(n4384), .A2(n5479), .ZN(n4386) );
  OAI22_X1 U5373 ( .A1(n4385), .A2(n5557), .B1(n4386), .B2(n5491), .ZN(n5467)
         );
  OAI211_X1 U5374 ( .C1(n5557), .C2(n4387), .A(n5491), .B(n4386), .ZN(n4388)
         );
  INV_X1 U5375 ( .A(n4388), .ZN(n4389) );
  INV_X1 U5376 ( .A(n5480), .ZN(n4391) );
  NAND2_X1 U5377 ( .A1(n4393), .A2(n4392), .ZN(U2830) );
  AND2_X1 U5378 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5775) );
  NOR4_X1 U5379 ( .A1(n4394), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_29__SCAN_IN), .A4(n4395), .ZN(n4396) );
  AOI21_X1 U5380 ( .B1(n5429), .B2(n5775), .A(n4396), .ZN(n4397) );
  INV_X1 U5381 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5773) );
  XNOR2_X1 U5382 ( .A(n4397), .B(n5773), .ZN(n5783) );
  AOI22_X1 U5383 ( .A1(n3492), .A2(EAX_REG_31__SCAN_IN), .B1(n3545), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4398) );
  INV_X1 U5384 ( .A(n4398), .ZN(n4399) );
  NAND2_X1 U5385 ( .A1(n5462), .A2(n6379), .ZN(n4409) );
  INV_X1 U5386 ( .A(n4401), .ZN(n4403) );
  INV_X1 U5387 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4402) );
  INV_X1 U5388 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4404) );
  NAND2_X1 U5389 ( .A1(n6427), .A2(REIP_REG_31__SCAN_IN), .ZN(n5776) );
  NAND2_X1 U5390 ( .A1(n6383), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4406)
         );
  OAI211_X1 U5391 ( .C1(n6391), .C2(n5244), .A(n5776), .B(n4406), .ZN(n4407)
         );
  INV_X1 U5392 ( .A(n4407), .ZN(n4408) );
  OAI211_X1 U5393 ( .C1(n5783), .C2(n6357), .A(n4409), .B(n4408), .ZN(U2955)
         );
  AND2_X1 U5394 ( .A1(n4414), .A2(n4413), .ZN(n4415) );
  AND2_X1 U5395 ( .A1(n4416), .A2(n4415), .ZN(n4417) );
  OR2_X1 U5396 ( .A1(n4418), .A2(n4417), .ZN(n4439) );
  NOR2_X1 U5397 ( .A1(n4412), .A2(n4439), .ZN(n4431) );
  OAI22_X1 U5398 ( .A1(n4471), .A2(n4064), .B1(n4410), .B2(n4431), .ZN(n6033)
         );
  INV_X1 U5399 ( .A(n5232), .ZN(n4419) );
  OR2_X1 U5400 ( .A1(n6271), .A2(n4419), .ZN(n4433) );
  OR2_X1 U5401 ( .A1(n4420), .A2(STATE_REG_0__SCAN_IN), .ZN(n6639) );
  AOI21_X1 U5402 ( .B1(n4433), .B2(n6639), .A(READY_N), .ZN(n6692) );
  NOR2_X1 U5403 ( .A1(n6033), .A2(n6692), .ZN(n6598) );
  NOR2_X1 U5404 ( .A1(n6598), .A2(n6620), .ZN(n6037) );
  INV_X1 U5405 ( .A(MORE_REG_SCAN_IN), .ZN(n4430) );
  NOR2_X1 U5406 ( .A1(n6597), .A2(n4543), .ZN(n4481) );
  INV_X1 U5407 ( .A(n4410), .ZN(n4421) );
  NAND2_X1 U5408 ( .A1(n4481), .A2(n4421), .ZN(n4422) );
  NAND2_X1 U5409 ( .A1(n4423), .A2(n4422), .ZN(n4427) );
  NAND2_X1 U5410 ( .A1(n4471), .A2(n4544), .ZN(n4426) );
  INV_X1 U5411 ( .A(n4439), .ZN(n4424) );
  OR2_X1 U5412 ( .A1(n4412), .A2(n4424), .ZN(n4425) );
  AND3_X1 U5413 ( .A1(n4427), .A2(n4426), .A3(n4425), .ZN(n6601) );
  INV_X1 U5414 ( .A(n6601), .ZN(n4428) );
  NAND2_X1 U5415 ( .A1(n6037), .A2(n4428), .ZN(n4429) );
  OAI21_X1 U5416 ( .B1(n6037), .B2(n4430), .A(n4429), .ZN(U3471) );
  NAND2_X1 U5417 ( .A1(n4515), .A2(n4410), .ZN(n4435) );
  NAND2_X1 U5418 ( .A1(n4431), .A2(n4505), .ZN(n4436) );
  INV_X1 U5419 ( .A(n6690), .ZN(n4434) );
  NOR2_X1 U5420 ( .A1(n6519), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5273) );
  OAI21_X1 U5421 ( .B1(n5273), .B2(READREQUEST_REG_SCAN_IN), .A(n4434), .ZN(
        n4432) );
  OAI21_X1 U5422 ( .B1(n4434), .B2(n4433), .A(n4432), .ZN(U3474) );
  INV_X1 U5423 ( .A(n4435), .ZN(n6270) );
  AOI211_X1 U5424 ( .C1(MEMORYFETCH_REG_SCAN_IN), .C2(n4436), .A(n5273), .B(
        n6270), .ZN(n4437) );
  INV_X1 U5425 ( .A(n4437), .ZN(U2788) );
  NAND2_X1 U5426 ( .A1(n4471), .A2(n4543), .ZN(n4441) );
  INV_X1 U5427 ( .A(n4438), .ZN(n6028) );
  NOR2_X1 U5428 ( .A1(READY_N), .A2(n4439), .ZN(n4466) );
  NAND2_X1 U5429 ( .A1(n6028), .A2(n4466), .ZN(n4440) );
  NAND2_X1 U5430 ( .A1(n4441), .A2(n4440), .ZN(n4507) );
  INV_X1 U5431 ( .A(n4507), .ZN(n4453) );
  INV_X1 U5432 ( .A(n4442), .ZN(n4487) );
  AOI21_X1 U5433 ( .B1(n4159), .B2(n6639), .A(READY_N), .ZN(n4443) );
  OAI21_X1 U5434 ( .B1(n6581), .B2(n4487), .A(n4443), .ZN(n4444) );
  INV_X1 U5435 ( .A(n4444), .ZN(n4450) );
  NAND2_X1 U5436 ( .A1(n4446), .A2(n4445), .ZN(n4447) );
  NAND2_X1 U5437 ( .A1(n4447), .A2(n4412), .ZN(n4468) );
  NAND2_X1 U5438 ( .A1(n4468), .A2(n4448), .ZN(n4449) );
  AOI21_X1 U5439 ( .B1(n4471), .B2(n4450), .A(n4449), .ZN(n4452) );
  NAND3_X1 U5440 ( .A1(n4453), .A2(n4452), .A3(n4451), .ZN(n6583) );
  NAND2_X1 U5441 ( .A1(n6583), .A2(n4505), .ZN(n4456) );
  NAND2_X1 U5442 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .ZN(n4570) );
  OR2_X1 U5443 ( .A1(n6613), .A2(n4570), .ZN(n6680) );
  INV_X1 U5444 ( .A(n6680), .ZN(n4454) );
  NAND2_X1 U5445 ( .A1(n4454), .A2(FLUSH_REG_SCAN_IN), .ZN(n4455) );
  NAND2_X1 U5446 ( .A1(n4456), .A2(n4455), .ZN(n6026) );
  NOR2_X1 U5447 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6683), .ZN(n4600) );
  OR2_X1 U5448 ( .A1(n6026), .A2(n4600), .ZN(n6032) );
  INV_X1 U5449 ( .A(n6032), .ZN(n5460) );
  AOI21_X1 U5450 ( .B1(n6581), .B2(n6027), .A(n5460), .ZN(n4461) );
  INV_X1 U5451 ( .A(n3491), .ZN(n5233) );
  INV_X1 U5452 ( .A(n4504), .ZN(n4457) );
  NAND4_X1 U5453 ( .A1(n4438), .A2(n4485), .A3(n4442), .A4(n4457), .ZN(n4458)
         );
  NOR2_X1 U5454 ( .A1(n4483), .A2(n4458), .ZN(n5916) );
  OAI22_X1 U5455 ( .A1(n5233), .A2(n5916), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n5919), .ZN(n6579) );
  INV_X1 U5456 ( .A(n5927), .ZN(n6614) );
  OAI22_X1 U5457 ( .A1(n6614), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n5454), .ZN(n4459) );
  AOI21_X1 U5458 ( .B1(n6027), .B2(n6579), .A(n4459), .ZN(n4460) );
  OAI22_X1 U5459 ( .A1(n4461), .A2(n4061), .B1(n5460), .B2(n4460), .ZN(U3461)
         );
  OAI21_X1 U5460 ( .B1(n4464), .B2(n4463), .A(n4462), .ZN(n6385) );
  NAND2_X1 U5461 ( .A1(n3398), .A2(n6639), .ZN(n4467) );
  NAND3_X1 U5462 ( .A1(n4467), .A2(n4466), .A3(n4465), .ZN(n4469) );
  OAI211_X1 U5463 ( .C1(n4471), .C2(n4470), .A(n4469), .B(n4468), .ZN(n4472)
         );
  NAND2_X1 U5464 ( .A1(n4472), .A2(n4505), .ZN(n4478) );
  NAND2_X1 U5465 ( .A1(n4620), .A2(n6639), .ZN(n5231) );
  INV_X1 U5466 ( .A(READY_N), .ZN(n7066) );
  NAND2_X1 U5467 ( .A1(n5231), .A2(n7066), .ZN(n4474) );
  OAI211_X1 U5468 ( .C1(n4442), .C2(n4474), .A(n3436), .B(n4473), .ZN(n4475)
         );
  AND2_X1 U5469 ( .A1(n4475), .A2(n4625), .ZN(n4476) );
  NAND2_X1 U5470 ( .A1(n4515), .A2(n4476), .ZN(n4477) );
  INV_X1 U5471 ( .A(n4488), .ZN(n4479) );
  NOR2_X1 U5472 ( .A1(n4442), .A2(n4133), .ZN(n4508) );
  AOI21_X1 U5473 ( .B1(n4479), .B2(n3386), .A(n4508), .ZN(n4480) );
  NAND3_X1 U5474 ( .A1(n4481), .A2(n4480), .A3(n4438), .ZN(n4482) );
  OR2_X1 U5475 ( .A1(n4495), .A2(n6384), .ZN(n6451) );
  NAND2_X1 U5476 ( .A1(n4495), .A2(n4544), .ZN(n5853) );
  INV_X1 U5477 ( .A(n4483), .ZN(n4484) );
  OAI21_X1 U5478 ( .B1(n3436), .B2(n4485), .A(n4484), .ZN(n4486) );
  NAND2_X1 U5479 ( .A1(n4495), .A2(n4486), .ZN(n5364) );
  NAND2_X1 U5480 ( .A1(n5853), .A2(n5364), .ZN(n5332) );
  INV_X1 U5481 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6452) );
  NAND2_X1 U5482 ( .A1(n5332), .A2(n6452), .ZN(n6446) );
  AOI21_X1 U5483 ( .B1(n6451), .B2(n6446), .A(n5453), .ZN(n4494) );
  NAND2_X1 U5484 ( .A1(n4487), .A2(n6271), .ZN(n6609) );
  OAI21_X1 U5485 ( .B1(n4488), .B2(n3386), .A(n6609), .ZN(n4489) );
  NOR2_X1 U5486 ( .A1(n4491), .A2(n4490), .ZN(n4492) );
  NOR2_X1 U5487 ( .A1(n6209), .A2(n4492), .ZN(n4641) );
  NOR2_X1 U5488 ( .A1(n6431), .A2(n4641), .ZN(n4493) );
  AOI211_X1 U5489 ( .C1(REIP_REG_1__SCAN_IN), .C2(n6384), .A(n4494), .B(n4493), 
        .ZN(n4498) );
  NAND2_X1 U5490 ( .A1(n4495), .A2(n6581), .ZN(n6450) );
  NAND2_X1 U5491 ( .A1(n6450), .A2(n5364), .ZN(n5858) );
  INV_X1 U5492 ( .A(n6450), .ZN(n4496) );
  NAND3_X1 U5493 ( .A1(n6403), .A2(n5453), .A3(n4529), .ZN(n4497) );
  OAI211_X1 U5494 ( .C1(n6385), .C2(n6394), .A(n4498), .B(n4497), .ZN(U3017)
         );
  AND2_X1 U5495 ( .A1(n4499), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4502) );
  OAI21_X1 U5496 ( .B1(n4502), .B2(n4501), .A(n4500), .ZN(n5764) );
  AND2_X1 U5497 ( .A1(n4504), .A2(n4503), .ZN(n4506) );
  NAND2_X2 U5498 ( .A1(n5449), .A2(n4511), .ZN(n5983) );
  AND2_X1 U5499 ( .A1(n5449), .A2(n4512), .ZN(n6242) );
  NOR2_X2 U5500 ( .A1(n6242), .A2(n6246), .ZN(n5360) );
  INV_X1 U5501 ( .A(DATAI_0_), .ZN(n6897) );
  INV_X1 U5502 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6302) );
  OAI222_X1 U5503 ( .A1(n5764), .A2(n5983), .B1(n5360), .B2(n6897), .C1(n5449), 
        .C2(n6302), .ZN(U2891) );
  NAND2_X1 U5504 ( .A1(n4515), .A2(n6581), .ZN(n4516) );
  NAND2_X1 U5505 ( .A1(n6346), .A2(n4516), .ZN(n4517) );
  INV_X1 U5506 ( .A(n6639), .ZN(n5234) );
  NAND2_X1 U5507 ( .A1(n6249), .A2(n3436), .ZN(n5012) );
  OR2_X1 U5508 ( .A1(n4570), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6606) );
  AOI22_X1 U5509 ( .A1(n6267), .A2(UWORD_REG_11__SCAN_IN), .B1(n6261), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4518) );
  OAI21_X1 U5510 ( .B1(n3978), .B2(n5012), .A(n4518), .ZN(U2896) );
  AOI22_X1 U5511 ( .A1(n6267), .A2(UWORD_REG_9__SCAN_IN), .B1(n6261), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4519) );
  OAI21_X1 U5512 ( .B1(n3940), .B2(n5012), .A(n4519), .ZN(U2898) );
  AOI22_X1 U5513 ( .A1(n6267), .A2(UWORD_REG_13__SCAN_IN), .B1(n6261), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4520) );
  OAI21_X1 U5514 ( .B1(n4019), .B2(n5012), .A(n4520), .ZN(U2894) );
  NAND3_X1 U5515 ( .A1(n4523), .A2(n4522), .A3(n3504), .ZN(n4524) );
  AND2_X1 U5516 ( .A1(n4521), .A2(n4524), .ZN(n6378) );
  INV_X1 U5517 ( .A(n6378), .ZN(n4525) );
  INV_X1 U5518 ( .A(DATAI_2_), .ZN(n4624) );
  INV_X1 U5519 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6308) );
  OAI222_X1 U5520 ( .A1(n4525), .A2(n5983), .B1(n5360), .B2(n4624), .C1(n5449), 
        .C2(n6308), .ZN(U2889) );
  XNOR2_X1 U5521 ( .A(n4527), .B(n4526), .ZN(n4640) );
  NOR2_X1 U5522 ( .A1(n4258), .A2(n5453), .ZN(n6426) );
  INV_X1 U5523 ( .A(n6426), .ZN(n4994) );
  OR2_X1 U5524 ( .A1(n5364), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4528)
         );
  INV_X1 U5525 ( .A(n5381), .ZN(n5855) );
  AOI21_X1 U5526 ( .B1(n5858), .B2(n4994), .A(n5855), .ZN(n6437) );
  AOI21_X1 U5527 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n4893) );
  NAND2_X1 U5528 ( .A1(n6425), .A2(n4893), .ZN(n6432) );
  NAND2_X1 U5529 ( .A1(n6437), .A2(n6432), .ZN(n4581) );
  NAND2_X1 U5530 ( .A1(n5858), .A2(n4529), .ZN(n5385) );
  AOI21_X1 U5531 ( .B1(n6426), .B2(n6424), .A(n6425), .ZN(n5144) );
  NOR2_X1 U5532 ( .A1(n4893), .A2(n5144), .ZN(n4577) );
  AOI22_X1 U5533 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n4581), .B1(n4577), 
        .B2(n4265), .ZN(n4532) );
  AOI21_X1 U5534 ( .B1(n4530), .B2(n4646), .A(n4578), .ZN(n6231) );
  AND2_X1 U5535 ( .A1(n6384), .A2(REIP_REG_3__SCAN_IN), .ZN(n4636) );
  AOI21_X1 U5536 ( .B1(n6445), .B2(n6231), .A(n4636), .ZN(n4531) );
  OAI211_X1 U5537 ( .C1(n4640), .C2(n6394), .A(n4532), .B(n4531), .ZN(U3015)
         );
  NOR2_X1 U5538 ( .A1(n5464), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4533)
         );
  OR2_X1 U5539 ( .A1(n4534), .A2(n4533), .ZN(n6441) );
  OAI222_X1 U5540 ( .A1(n6441), .A2(n6233), .B1(n6230), .B2(n4144), .C1(n5764), 
        .C2(n6226), .ZN(U2859) );
  OR2_X1 U5541 ( .A1(n4536), .A2(n4535), .ZN(n4537) );
  AND2_X1 U5542 ( .A1(n3504), .A2(n4537), .ZN(n6386) );
  INV_X1 U5543 ( .A(n6386), .ZN(n4538) );
  INV_X1 U5544 ( .A(DATAI_1_), .ZN(n4619) );
  INV_X1 U5545 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6305) );
  OAI222_X1 U5546 ( .A1(n4538), .A2(n5983), .B1(n5360), .B2(n4619), .C1(n5449), 
        .C2(n6305), .ZN(U2890) );
  AND2_X1 U5547 ( .A1(n4521), .A2(n4539), .ZN(n4541) );
  OR2_X1 U5548 ( .A1(n4541), .A2(n4540), .ZN(n6234) );
  INV_X1 U5549 ( .A(DATAI_3_), .ZN(n7034) );
  INV_X1 U5550 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6311) );
  OAI222_X1 U5551 ( .A1(n6234), .A2(n5983), .B1(n5360), .B2(n7034), .C1(n5449), 
        .C2(n6311), .ZN(U2888) );
  INV_X1 U5552 ( .A(FLUSH_REG_SCAN_IN), .ZN(n7063) );
  NAND2_X1 U5553 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n7063), .ZN(n4562) );
  INV_X1 U5554 ( .A(n4542), .ZN(n4561) );
  INV_X1 U5555 ( .A(n6581), .ZN(n5920) );
  XNOR2_X1 U5556 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4549) );
  NOR2_X1 U5557 ( .A1(n4544), .A2(n4543), .ZN(n4555) );
  XNOR2_X1 U5558 ( .A(n4545), .B(n3168), .ZN(n4548) );
  INV_X1 U5559 ( .A(n4547), .ZN(n6196) );
  OAI222_X1 U5560 ( .A1(n5920), .A2(n4549), .B1(n4555), .B2(n4548), .C1(n6196), 
        .C2(n5916), .ZN(n5455) );
  MUX2_X1 U5561 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n5455), .S(n6583), 
        .Z(n6591) );
  INV_X1 U5562 ( .A(n3171), .ZN(n6458) );
  NAND2_X1 U5563 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4551) );
  INV_X1 U5564 ( .A(n4551), .ZN(n4552) );
  MUX2_X1 U5565 ( .A(n4552), .B(n4551), .S(n4559), .Z(n4557) );
  MUX2_X1 U5566 ( .A(n4553), .B(n4559), .S(n4545), .Z(n4554) );
  NOR3_X1 U5567 ( .A1(n4555), .A2(n4542), .A3(n4554), .ZN(n4556) );
  AOI21_X1 U5568 ( .B1(n6581), .B2(n4557), .A(n4556), .ZN(n4558) );
  OAI21_X1 U5569 ( .B1(n6458), .B2(n5916), .A(n4558), .ZN(n5397) );
  MUX2_X1 U5570 ( .A(n4559), .B(n5397), .S(n6583), .Z(n6592) );
  NAND3_X1 U5571 ( .A1(n6591), .A2(n6592), .A3(n5454), .ZN(n4560) );
  OAI21_X1 U5572 ( .B1(n4562), .B2(n4561), .A(n4560), .ZN(n6604) );
  INV_X1 U5573 ( .A(n4563), .ZN(n5918) );
  NAND2_X1 U5574 ( .A1(n6604), .A2(n5918), .ZN(n4572) );
  INV_X1 U5575 ( .A(n6583), .ZN(n4564) );
  MUX2_X1 U5576 ( .A(n7063), .B(n4564), .S(n5454), .Z(n4568) );
  INV_X1 U5577 ( .A(n4852), .ZN(n4693) );
  OR2_X1 U5578 ( .A1(n4565), .A2(n4693), .ZN(n4566) );
  XNOR2_X1 U5579 ( .A(n4566), .B(n6031), .ZN(n6184) );
  NOR3_X1 U5580 ( .A1(n6184), .A2(STATE2_REG_1__SCAN_IN), .A3(n4438), .ZN(
        n4567) );
  AOI21_X1 U5581 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n4568), .A(n4567), 
        .ZN(n6602) );
  AND3_X1 U5582 ( .A1(n4572), .A2(n7063), .A3(n6602), .ZN(n4569) );
  NOR2_X1 U5583 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6694) );
  OAI21_X1 U5584 ( .B1(n4569), .B2(n6680), .A(n4813), .ZN(n6453) );
  INV_X1 U5585 ( .A(n4570), .ZN(n4571) );
  AND3_X1 U5586 ( .A1(n4572), .A2(n6602), .A3(n4571), .ZN(n6612) );
  AND2_X1 U5587 ( .A1(n6683), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5911) );
  OAI22_X1 U5588 ( .A1(n4850), .A2(n6519), .B1(n5233), .B2(n5911), .ZN(n4573)
         );
  OAI21_X1 U5589 ( .B1(n6612), .B2(n4573), .A(n6453), .ZN(n4574) );
  OAI21_X1 U5590 ( .B1(n6453), .B2(n6580), .A(n4574), .ZN(U3465) );
  XNOR2_X1 U5591 ( .A(n3160), .B(n4576), .ZN(n4764) );
  NAND2_X1 U5592 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4993) );
  OAI211_X1 U5593 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4577), .B(n4993), .ZN(n4583) );
  INV_X1 U5594 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6649) );
  NOR2_X1 U5595 ( .A1(n6392), .A2(n6649), .ZN(n4760) );
  OAI21_X1 U5596 ( .B1(n4579), .B2(n4578), .A(n4768), .ZN(n6175) );
  NOR2_X1 U5597 ( .A1(n6431), .A2(n6175), .ZN(n4580) );
  AOI211_X1 U5598 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n4581), .A(n4760), 
        .B(n4580), .ZN(n4582) );
  OAI211_X1 U5599 ( .C1(n6394), .C2(n4764), .A(n4583), .B(n4582), .ZN(U3014)
         );
  OAI21_X1 U5600 ( .B1(n4540), .B2(n4585), .A(n4584), .ZN(n4759) );
  INV_X1 U5601 ( .A(DATAI_4_), .ZN(n6899) );
  INV_X1 U5602 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6314) );
  OAI222_X1 U5603 ( .A1(n4759), .A2(n5983), .B1(n5360), .B2(n6899), .C1(n6314), 
        .C2(n5449), .ZN(U2887) );
  INV_X1 U5604 ( .A(n5902), .ZN(n4652) );
  OAI21_X1 U5605 ( .B1(n4849), .B2(n4652), .A(n6379), .ZN(n4590) );
  OR2_X1 U5606 ( .A1(n6519), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5914) );
  NAND2_X1 U5607 ( .A1(n4590), .A2(n5914), .ZN(n4595) );
  AND2_X1 U5608 ( .A1(n3171), .A2(n3491), .ZN(n4964) );
  NAND2_X1 U5609 ( .A1(n4547), .A2(n3170), .ZN(n5064) );
  INV_X1 U5610 ( .A(n5064), .ZN(n4593) );
  INV_X1 U5611 ( .A(n4592), .ZN(n4631) );
  AOI21_X1 U5612 ( .B1(n4964), .B2(n4593), .A(n4631), .ZN(n4596) );
  INV_X1 U5613 ( .A(n6519), .ZN(n5154) );
  OAI21_X1 U5614 ( .B1(n5154), .B2(n5059), .A(n6521), .ZN(n4594) );
  INV_X1 U5615 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4604) );
  NAND2_X1 U5616 ( .A1(n6379), .A2(DATAI_22_), .ZN(n6494) );
  INV_X1 U5617 ( .A(n6494), .ZN(n6563) );
  INV_X1 U5618 ( .A(DATAI_6_), .ZN(n5016) );
  INV_X1 U5619 ( .A(n4596), .ZN(n4597) );
  NAND2_X1 U5620 ( .A1(n4597), .A2(n5154), .ZN(n4599) );
  NAND2_X1 U5621 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5059), .ZN(n4598) );
  NAND2_X1 U5622 ( .A1(n4599), .A2(n4598), .ZN(n4629) );
  AOI22_X1 U5623 ( .A1(n4659), .A2(n6563), .B1(n6564), .B2(n4629), .ZN(n4603)
         );
  INV_X1 U5624 ( .A(n4600), .ZN(n6681) );
  NOR2_X1 U5625 ( .A1(n4630), .A2(n3334), .ZN(n6562) );
  NAND2_X1 U5626 ( .A1(n5902), .A2(n4850), .ZN(n5153) );
  NAND2_X1 U5627 ( .A1(n6379), .A2(DATAI_30_), .ZN(n6567) );
  INV_X1 U5628 ( .A(n6567), .ZN(n6491) );
  AOI22_X1 U5629 ( .A1(n6562), .A2(n4631), .B1(n5935), .B2(n6491), .ZN(n4602)
         );
  OAI211_X1 U5630 ( .C1(n4635), .C2(n4604), .A(n4603), .B(n4602), .ZN(U3146)
         );
  INV_X1 U5631 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4607) );
  NAND2_X1 U5632 ( .A1(n6379), .A2(DATAI_23_), .ZN(n6502) );
  INV_X1 U5633 ( .A(n6502), .ZN(n6570) );
  INV_X1 U5634 ( .A(DATAI_7_), .ZN(n6950) );
  AOI22_X1 U5635 ( .A1(n4659), .A2(n6570), .B1(n6573), .B2(n4629), .ZN(n4606)
         );
  NAND2_X1 U5636 ( .A1(n6379), .A2(DATAI_31_), .ZN(n6578) );
  INV_X1 U5637 ( .A(n6578), .ZN(n6498) );
  AOI22_X1 U5638 ( .A1(n6569), .A2(n4631), .B1(n5935), .B2(n6498), .ZN(n4605)
         );
  OAI211_X1 U5639 ( .C1(n4635), .C2(n4607), .A(n4606), .B(n4605), .ZN(U3147)
         );
  INV_X1 U5640 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4611) );
  NAND2_X1 U5641 ( .A1(n6379), .A2(DATAI_20_), .ZN(n6486) );
  INV_X1 U5642 ( .A(n6486), .ZN(n6551) );
  AOI22_X1 U5643 ( .A1(n4659), .A2(n6551), .B1(n6552), .B2(n4629), .ZN(n4610)
         );
  NOR2_X1 U5644 ( .A1(n4630), .A2(n4608), .ZN(n6550) );
  NAND2_X1 U5645 ( .A1(n6379), .A2(DATAI_28_), .ZN(n6555) );
  INV_X1 U5646 ( .A(n6555), .ZN(n6483) );
  AOI22_X1 U5647 ( .A1(n6550), .A2(n4631), .B1(n5935), .B2(n6483), .ZN(n4609)
         );
  OAI211_X1 U5648 ( .C1(n4635), .C2(n4611), .A(n4610), .B(n4609), .ZN(U3144)
         );
  INV_X1 U5649 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4615) );
  NAND2_X1 U5650 ( .A1(n6379), .A2(DATAI_19_), .ZN(n6482) );
  INV_X1 U5651 ( .A(n6482), .ZN(n6545) );
  AOI22_X1 U5652 ( .A1(n4659), .A2(n6545), .B1(n6546), .B2(n4629), .ZN(n4614)
         );
  NAND2_X1 U5653 ( .A1(n6379), .A2(DATAI_27_), .ZN(n6549) );
  INV_X1 U5654 ( .A(n6549), .ZN(n6479) );
  AOI22_X1 U5655 ( .A1(n6544), .A2(n4631), .B1(n5935), .B2(n6479), .ZN(n4613)
         );
  OAI211_X1 U5656 ( .C1(n4635), .C2(n4615), .A(n4614), .B(n4613), .ZN(U3143)
         );
  INV_X1 U5657 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4618) );
  NAND2_X1 U5658 ( .A1(n6379), .A2(DATAI_21_), .ZN(n6490) );
  INV_X1 U5659 ( .A(n6490), .ZN(n6557) );
  INV_X1 U5660 ( .A(DATAI_5_), .ZN(n6941) );
  AOI22_X1 U5661 ( .A1(n4659), .A2(n6557), .B1(n6558), .B2(n4629), .ZN(n4617)
         );
  NOR2_X1 U5662 ( .A1(n4630), .A2(n3394), .ZN(n6556) );
  NAND2_X1 U5663 ( .A1(n6379), .A2(DATAI_29_), .ZN(n6561) );
  INV_X1 U5664 ( .A(n6561), .ZN(n6487) );
  AOI22_X1 U5665 ( .A1(n6556), .A2(n4631), .B1(n5935), .B2(n6487), .ZN(n4616)
         );
  OAI211_X1 U5666 ( .C1(n4635), .C2(n4618), .A(n4617), .B(n4616), .ZN(U3145)
         );
  INV_X1 U5667 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4623) );
  NAND2_X1 U5668 ( .A1(n6379), .A2(DATAI_17_), .ZN(n6476) );
  INV_X1 U5669 ( .A(n6476), .ZN(n6531) );
  AOI22_X1 U5670 ( .A1(n4659), .A2(n6531), .B1(n6532), .B2(n4629), .ZN(n4622)
         );
  NOR2_X1 U5671 ( .A1(n4630), .A2(n4620), .ZN(n6530) );
  NAND2_X1 U5672 ( .A1(n6379), .A2(DATAI_25_), .ZN(n6535) );
  INV_X1 U5673 ( .A(n6535), .ZN(n6473) );
  AOI22_X1 U5674 ( .A1(n6530), .A2(n4631), .B1(n5935), .B2(n6473), .ZN(n4621)
         );
  OAI211_X1 U5675 ( .C1(n4635), .C2(n4623), .A(n4622), .B(n4621), .ZN(U3141)
         );
  INV_X1 U5676 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4628) );
  NAND2_X1 U5677 ( .A1(n6379), .A2(DATAI_18_), .ZN(n6543) );
  INV_X1 U5678 ( .A(n6543), .ZN(n5053) );
  AOI22_X1 U5679 ( .A1(n4659), .A2(n5053), .B1(n6539), .B2(n4629), .ZN(n4627)
         );
  INV_X1 U5680 ( .A(DATAI_26_), .ZN(n6965) );
  NOR2_X1 U5681 ( .A1(n6359), .A2(n6965), .ZN(n6537) );
  AOI22_X1 U5682 ( .A1(n6536), .A2(n4631), .B1(n5935), .B2(n6537), .ZN(n4626)
         );
  OAI211_X1 U5683 ( .C1(n4635), .C2(n4628), .A(n4627), .B(n4626), .ZN(U3142)
         );
  INV_X1 U5684 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4634) );
  NAND2_X1 U5685 ( .A1(n6379), .A2(DATAI_16_), .ZN(n6472) );
  INV_X1 U5686 ( .A(n6472), .ZN(n6513) );
  AOI22_X1 U5687 ( .A1(n4659), .A2(n6513), .B1(n6526), .B2(n4629), .ZN(n4633)
         );
  NAND2_X1 U5688 ( .A1(n6379), .A2(DATAI_24_), .ZN(n6529) );
  INV_X1 U5689 ( .A(n6529), .ZN(n6469) );
  AOI22_X1 U5690 ( .A1(n6512), .A2(n4631), .B1(n5935), .B2(n6469), .ZN(n4632)
         );
  OAI211_X1 U5691 ( .C1(n4635), .C2(n4634), .A(n4633), .B(n4632), .ZN(U3140)
         );
  INV_X1 U5692 ( .A(n6234), .ZN(n5292) );
  AOI21_X1 U5693 ( .B1(n6383), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n4636), 
        .ZN(n4637) );
  OAI21_X1 U5694 ( .B1(n5296), .B2(n6391), .A(n4637), .ZN(n4638) );
  AOI21_X1 U5695 ( .B1(n5292), .B2(n6379), .A(n4638), .ZN(n4639) );
  OAI21_X1 U5696 ( .B1(n4640), .B2(n6357), .A(n4639), .ZN(U2983) );
  OAI22_X1 U5697 ( .A1(n6233), .A2(n4641), .B1(n6238), .B2(n3205), .ZN(n4642)
         );
  AOI21_X1 U5698 ( .B1(n6386), .B2(n4383), .A(n4642), .ZN(n4643) );
  INV_X1 U5699 ( .A(n4643), .ZN(U2858) );
  OR2_X1 U5700 ( .A1(n4645), .A2(n4644), .ZN(n4647) );
  NAND2_X1 U5701 ( .A1(n4647), .A2(n4646), .ZN(n6430) );
  INV_X1 U5702 ( .A(EBX_REG_2__SCAN_IN), .ZN(n6193) );
  OAI22_X1 U5703 ( .A1(n6430), .A2(n6233), .B1(n6238), .B2(n6193), .ZN(n4648)
         );
  AOI21_X1 U5704 ( .B1(n6378), .B2(n4383), .A(n4648), .ZN(n4649) );
  INV_X1 U5705 ( .A(n4649), .ZN(U2857) );
  OAI222_X1 U5706 ( .A1(n6175), .A2(n6233), .B1(n6230), .B2(n4158), .C1(n4759), 
        .C2(n6226), .ZN(U2855) );
  NAND2_X1 U5707 ( .A1(n4587), .A2(n4652), .ZN(n4653) );
  NOR3_X1 U5708 ( .A1(n4924), .A2(n4659), .A3(n6519), .ZN(n4654) );
  INV_X1 U5709 ( .A(n5914), .ZN(n6463) );
  NAND2_X1 U5710 ( .A1(n6458), .A2(n3256), .ZN(n4660) );
  OAI21_X1 U5711 ( .B1(n4654), .B2(n6463), .A(n4660), .ZN(n4658) );
  NAND3_X1 U5712 ( .A1(n6594), .A2(n6590), .A3(n6586), .ZN(n4904) );
  NOR2_X1 U5713 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4904), .ZN(n4689)
         );
  INV_X1 U5714 ( .A(n4689), .ZN(n4656) );
  AND2_X1 U5715 ( .A1(n4661), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6456) );
  INV_X1 U5716 ( .A(n4812), .ZN(n4655) );
  NOR2_X1 U5717 ( .A1(n4655), .A2(n5065), .ZN(n4782) );
  OAI21_X1 U5718 ( .B1(n4782), .B2(n4969), .A(n5023), .ZN(n4776) );
  AOI211_X1 U5719 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4656), .A(n6456), .B(
        n4776), .ZN(n4657) );
  NAND2_X1 U5720 ( .A1(n4658), .A2(n4657), .ZN(n4685) );
  NAND2_X1 U5721 ( .A1(n4685), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4666) );
  INV_X1 U5722 ( .A(n4660), .ZN(n4900) );
  NAND2_X1 U5723 ( .A1(n4900), .A2(n5154), .ZN(n4663) );
  NOR2_X1 U5724 ( .A1(n4661), .A2(n4969), .ZN(n5157) );
  NAND2_X1 U5725 ( .A1(n4782), .A2(n5157), .ZN(n4662) );
  OAI22_X1 U5726 ( .A1(n4687), .A2(n6529), .B1(n4686), .B2(n5932), .ZN(n4664)
         );
  AOI21_X1 U5727 ( .B1(n6512), .B2(n4689), .A(n4664), .ZN(n4665) );
  OAI211_X1 U5728 ( .C1(n4692), .C2(n6472), .A(n4666), .B(n4665), .ZN(U3020)
         );
  NAND2_X1 U5729 ( .A1(n4685), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4669) );
  INV_X1 U5730 ( .A(n6537), .ZN(n5090) );
  OAI22_X1 U5731 ( .A1(n4687), .A2(n5090), .B1(n4686), .B2(n5169), .ZN(n4667)
         );
  AOI21_X1 U5732 ( .B1(n6536), .B2(n4689), .A(n4667), .ZN(n4668) );
  OAI211_X1 U5733 ( .C1(n4692), .C2(n6543), .A(n4669), .B(n4668), .ZN(U3022)
         );
  NAND2_X1 U5734 ( .A1(n4685), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4672) );
  OAI22_X1 U5735 ( .A1(n4687), .A2(n6567), .B1(n4686), .B2(n5194), .ZN(n4670)
         );
  AOI21_X1 U5736 ( .B1(n6562), .B2(n4689), .A(n4670), .ZN(n4671) );
  OAI211_X1 U5737 ( .C1(n4692), .C2(n6494), .A(n4672), .B(n4671), .ZN(U3026)
         );
  NAND2_X1 U5738 ( .A1(n4685), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4675) );
  OAI22_X1 U5739 ( .A1(n4687), .A2(n6561), .B1(n4686), .B2(n5179), .ZN(n4673)
         );
  AOI21_X1 U5740 ( .B1(n6556), .B2(n4689), .A(n4673), .ZN(n4674) );
  OAI211_X1 U5741 ( .C1(n4692), .C2(n6490), .A(n4675), .B(n4674), .ZN(U3025)
         );
  NAND2_X1 U5742 ( .A1(n4685), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4678) );
  OAI22_X1 U5743 ( .A1(n4687), .A2(n6555), .B1(n4686), .B2(n5174), .ZN(n4676)
         );
  AOI21_X1 U5744 ( .B1(n6550), .B2(n4689), .A(n4676), .ZN(n4677) );
  OAI211_X1 U5745 ( .C1(n4692), .C2(n6486), .A(n4678), .B(n4677), .ZN(U3024)
         );
  NAND2_X1 U5746 ( .A1(n4685), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4681) );
  OAI22_X1 U5747 ( .A1(n4687), .A2(n6549), .B1(n4686), .B2(n5206), .ZN(n4679)
         );
  AOI21_X1 U5748 ( .B1(n6544), .B2(n4689), .A(n4679), .ZN(n4680) );
  OAI211_X1 U5749 ( .C1(n4692), .C2(n6482), .A(n4681), .B(n4680), .ZN(U3023)
         );
  NAND2_X1 U5750 ( .A1(n4685), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4684) );
  OAI22_X1 U5751 ( .A1(n4687), .A2(n6578), .B1(n4686), .B2(n5184), .ZN(n4682)
         );
  AOI21_X1 U5752 ( .B1(n6569), .B2(n4689), .A(n4682), .ZN(n4683) );
  OAI211_X1 U5753 ( .C1(n4692), .C2(n6502), .A(n4684), .B(n4683), .ZN(U3027)
         );
  NAND2_X1 U5754 ( .A1(n4685), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4691) );
  OAI22_X1 U5755 ( .A1(n4687), .A2(n6535), .B1(n4686), .B2(n5189), .ZN(n4688)
         );
  AOI21_X1 U5756 ( .B1(n6530), .B2(n4689), .A(n4688), .ZN(n4690) );
  OAI211_X1 U5757 ( .C1(n4692), .C2(n6476), .A(n4691), .B(n4690), .ZN(U3021)
         );
  OR2_X1 U5758 ( .A1(n4587), .A2(n3577), .ZN(n4735) );
  AOI21_X1 U5759 ( .B1(n4697), .B2(STATEBS16_REG_SCAN_IN), .A(n6519), .ZN(
        n4778) );
  INV_X1 U5760 ( .A(n3170), .ZN(n6214) );
  AND2_X1 U5761 ( .A1(n4547), .A2(n6214), .ZN(n4928) );
  NAND2_X1 U5762 ( .A1(n4928), .A2(n4693), .ZN(n4777) );
  OR2_X1 U5763 ( .A1(n4777), .A2(n5233), .ZN(n4694) );
  NAND2_X1 U5764 ( .A1(n6586), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4929) );
  OR2_X1 U5765 ( .A1(n4929), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4775)
         );
  OR2_X1 U5766 ( .A1(n6580), .A2(n4775), .ZN(n4722) );
  NAND2_X1 U5767 ( .A1(n4694), .A2(n4722), .ZN(n4700) );
  INV_X1 U5768 ( .A(n4775), .ZN(n4695) );
  AOI22_X1 U5769 ( .A1(n4778), .A2(n4700), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4695), .ZN(n4728) );
  INV_X1 U5770 ( .A(n4697), .ZN(n4696) );
  NOR2_X2 U5771 ( .A1(n4696), .A2(n4962), .ZN(n4808) );
  INV_X1 U5772 ( .A(n6550), .ZN(n5170) );
  OAI22_X1 U5773 ( .A1(n4723), .A2(n6486), .B1(n5170), .B2(n4722), .ZN(n4698)
         );
  AOI21_X1 U5774 ( .B1(n6483), .B2(n4808), .A(n4698), .ZN(n4703) );
  INV_X1 U5775 ( .A(n4778), .ZN(n4701) );
  INV_X1 U5776 ( .A(n6521), .ZN(n5103) );
  AOI21_X1 U5777 ( .B1(n6519), .B2(n4775), .A(n5103), .ZN(n4699) );
  NAND2_X1 U5778 ( .A1(n4725), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4702) );
  OAI211_X1 U5779 ( .C1(n4728), .C2(n5174), .A(n4703), .B(n4702), .ZN(U3064)
         );
  OAI22_X1 U5780 ( .A1(n4723), .A2(n6543), .B1(n5165), .B2(n4722), .ZN(n4704)
         );
  AOI21_X1 U5781 ( .B1(n6537), .B2(n4808), .A(n4704), .ZN(n4706) );
  NAND2_X1 U5782 ( .A1(n4725), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4705) );
  OAI211_X1 U5783 ( .C1(n4728), .C2(n5169), .A(n4706), .B(n4705), .ZN(U3062)
         );
  OAI22_X1 U5784 ( .A1(n4723), .A2(n6482), .B1(n5201), .B2(n4722), .ZN(n4707)
         );
  AOI21_X1 U5785 ( .B1(n6479), .B2(n4808), .A(n4707), .ZN(n4709) );
  NAND2_X1 U5786 ( .A1(n4725), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4708) );
  OAI211_X1 U5787 ( .C1(n4728), .C2(n5206), .A(n4709), .B(n4708), .ZN(U3063)
         );
  INV_X1 U5788 ( .A(n6562), .ZN(n5190) );
  OAI22_X1 U5789 ( .A1(n4723), .A2(n6494), .B1(n5190), .B2(n4722), .ZN(n4710)
         );
  AOI21_X1 U5790 ( .B1(n6491), .B2(n4808), .A(n4710), .ZN(n4712) );
  NAND2_X1 U5791 ( .A1(n4725), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4711) );
  OAI211_X1 U5792 ( .C1(n4728), .C2(n5194), .A(n4712), .B(n4711), .ZN(U3066)
         );
  OAI22_X1 U5793 ( .A1(n4723), .A2(n6472), .B1(n5195), .B2(n4722), .ZN(n4713)
         );
  AOI21_X1 U5794 ( .B1(n6469), .B2(n4808), .A(n4713), .ZN(n4715) );
  NAND2_X1 U5795 ( .A1(n4725), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4714) );
  OAI211_X1 U5796 ( .C1(n4728), .C2(n5932), .A(n4715), .B(n4714), .ZN(U3060)
         );
  OAI22_X1 U5797 ( .A1(n4723), .A2(n6502), .B1(n5180), .B2(n4722), .ZN(n4716)
         );
  AOI21_X1 U5798 ( .B1(n6498), .B2(n4808), .A(n4716), .ZN(n4718) );
  NAND2_X1 U5799 ( .A1(n4725), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4717) );
  OAI211_X1 U5800 ( .C1(n4728), .C2(n5184), .A(n4718), .B(n4717), .ZN(U3067)
         );
  INV_X1 U5801 ( .A(n6530), .ZN(n5185) );
  OAI22_X1 U5802 ( .A1(n4723), .A2(n6476), .B1(n5185), .B2(n4722), .ZN(n4719)
         );
  AOI21_X1 U5803 ( .B1(n6473), .B2(n4808), .A(n4719), .ZN(n4721) );
  NAND2_X1 U5804 ( .A1(n4725), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4720) );
  OAI211_X1 U5805 ( .C1(n4728), .C2(n5189), .A(n4721), .B(n4720), .ZN(U3061)
         );
  INV_X1 U5806 ( .A(n6556), .ZN(n5175) );
  OAI22_X1 U5807 ( .A1(n4723), .A2(n6490), .B1(n5175), .B2(n4722), .ZN(n4724)
         );
  AOI21_X1 U5808 ( .B1(n6487), .B2(n4808), .A(n4724), .ZN(n4727) );
  NAND2_X1 U5809 ( .A1(n4725), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4726) );
  OAI211_X1 U5810 ( .C1(n4728), .C2(n5179), .A(n4727), .B(n4726), .ZN(U3065)
         );
  NAND2_X1 U5811 ( .A1(n5902), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5905) );
  INV_X1 U5812 ( .A(n5905), .ZN(n5909) );
  NOR2_X1 U5813 ( .A1(n5909), .A2(n6519), .ZN(n6515) );
  AOI21_X1 U5814 ( .B1(n5154), .B2(n4735), .A(n6515), .ZN(n4731) );
  OR2_X1 U5815 ( .A1(n5064), .A2(n4852), .ZN(n6462) );
  INV_X1 U5816 ( .A(n6462), .ZN(n4729) );
  INV_X1 U5817 ( .A(n4754), .ZN(n6504) );
  AOI21_X1 U5818 ( .B1(n4729), .B2(n3491), .A(n6504), .ZN(n4732) );
  INV_X1 U5819 ( .A(n6455), .ZN(n4730) );
  OAI22_X1 U5820 ( .A1(n4731), .A2(n4732), .B1(n4730), .B2(n4969), .ZN(n6506)
         );
  INV_X1 U5821 ( .A(n4731), .ZN(n4733) );
  NAND2_X1 U5822 ( .A1(n4733), .A2(n4732), .ZN(n4734) );
  OAI211_X1 U5823 ( .C1(n6455), .C2(n5154), .A(n4734), .B(n6521), .ZN(n6507)
         );
  NOR2_X1 U5824 ( .A1(n5165), .A2(n4754), .ZN(n4737) );
  INV_X1 U5825 ( .A(n5153), .ZN(n5019) );
  OAI22_X1 U5826 ( .A1(n5090), .A2(n6510), .B1(n6503), .B2(n6543), .ZN(n4736)
         );
  AOI211_X1 U5827 ( .C1(n6507), .C2(INSTQUEUE_REG_7__2__SCAN_IN), .A(n4737), 
        .B(n4736), .ZN(n4738) );
  OAI21_X1 U5828 ( .B1(n4758), .B2(n5169), .A(n4738), .ZN(U3078) );
  NOR2_X1 U5829 ( .A1(n5195), .A2(n4754), .ZN(n4740) );
  OAI22_X1 U5830 ( .A1(n6529), .A2(n6510), .B1(n6503), .B2(n6472), .ZN(n4739)
         );
  AOI211_X1 U5831 ( .C1(n6507), .C2(INSTQUEUE_REG_7__0__SCAN_IN), .A(n4740), 
        .B(n4739), .ZN(n4741) );
  OAI21_X1 U5832 ( .B1(n4758), .B2(n5932), .A(n4741), .ZN(U3076) );
  NOR2_X1 U5833 ( .A1(n5185), .A2(n4754), .ZN(n4743) );
  OAI22_X1 U5834 ( .A1(n6535), .A2(n6510), .B1(n6503), .B2(n6476), .ZN(n4742)
         );
  AOI211_X1 U5835 ( .C1(n6507), .C2(INSTQUEUE_REG_7__1__SCAN_IN), .A(n4743), 
        .B(n4742), .ZN(n4744) );
  OAI21_X1 U5836 ( .B1(n4758), .B2(n5189), .A(n4744), .ZN(U3077) );
  NOR2_X1 U5837 ( .A1(n5190), .A2(n4754), .ZN(n4746) );
  OAI22_X1 U5838 ( .A1(n6567), .A2(n6510), .B1(n6503), .B2(n6494), .ZN(n4745)
         );
  AOI211_X1 U5839 ( .C1(n6507), .C2(INSTQUEUE_REG_7__6__SCAN_IN), .A(n4746), 
        .B(n4745), .ZN(n4747) );
  OAI21_X1 U5840 ( .B1(n4758), .B2(n5194), .A(n4747), .ZN(U3082) );
  NOR2_X1 U5841 ( .A1(n5180), .A2(n4754), .ZN(n4749) );
  OAI22_X1 U5842 ( .A1(n6578), .A2(n6510), .B1(n6503), .B2(n6502), .ZN(n4748)
         );
  AOI211_X1 U5843 ( .C1(n6507), .C2(INSTQUEUE_REG_7__7__SCAN_IN), .A(n4749), 
        .B(n4748), .ZN(n4750) );
  OAI21_X1 U5844 ( .B1(n4758), .B2(n5184), .A(n4750), .ZN(U3083) );
  NOR2_X1 U5845 ( .A1(n5201), .A2(n4754), .ZN(n4752) );
  OAI22_X1 U5846 ( .A1(n6549), .A2(n6510), .B1(n6503), .B2(n6482), .ZN(n4751)
         );
  AOI211_X1 U5847 ( .C1(n6507), .C2(INSTQUEUE_REG_7__3__SCAN_IN), .A(n4752), 
        .B(n4751), .ZN(n4753) );
  OAI21_X1 U5848 ( .B1(n4758), .B2(n5206), .A(n4753), .ZN(U3079) );
  NOR2_X1 U5849 ( .A1(n5170), .A2(n4754), .ZN(n4756) );
  OAI22_X1 U5850 ( .A1(n6555), .A2(n6510), .B1(n6503), .B2(n6486), .ZN(n4755)
         );
  AOI211_X1 U5851 ( .C1(n6507), .C2(INSTQUEUE_REG_7__4__SCAN_IN), .A(n4756), 
        .B(n4755), .ZN(n4757) );
  OAI21_X1 U5852 ( .B1(n4758), .B2(n5174), .A(n4757), .ZN(U3080) );
  INV_X1 U5853 ( .A(n4759), .ZN(n6186) );
  AOI21_X1 U5854 ( .B1(n6383), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n4760), 
        .ZN(n4761) );
  OAI21_X1 U5855 ( .B1(n6189), .B2(n6391), .A(n4761), .ZN(n4762) );
  AOI21_X1 U5856 ( .B1(n6186), .B2(n6379), .A(n4762), .ZN(n4763) );
  OAI21_X1 U5857 ( .B1(n6357), .B2(n4764), .A(n4763), .ZN(U2982) );
  NAND2_X1 U5858 ( .A1(n4584), .A2(n4766), .ZN(n4767) );
  AND2_X1 U5859 ( .A1(n4765), .A2(n4767), .ZN(n6368) );
  INV_X1 U5860 ( .A(n6368), .ZN(n4772) );
  OAI222_X1 U5861 ( .A1(n4772), .A2(n5983), .B1(n5360), .B2(n6941), .C1(n5449), 
        .C2(n3618), .ZN(U2886) );
  INV_X1 U5862 ( .A(EBX_REG_5__SCAN_IN), .ZN(n6167) );
  INV_X1 U5863 ( .A(n4768), .ZN(n4769) );
  XNOR2_X1 U5864 ( .A(n4770), .B(n4769), .ZN(n6172) );
  INV_X1 U5865 ( .A(n6172), .ZN(n4771) );
  OAI222_X1 U5866 ( .A1(n6226), .A2(n4772), .B1(n6230), .B2(n6167), .C1(n6233), 
        .C2(n4771), .ZN(U2854) );
  NAND2_X1 U5867 ( .A1(n4587), .A2(n4773), .ZN(n4774) );
  OR2_X1 U5868 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4775), .ZN(n4806)
         );
  AOI211_X1 U5869 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4806), .A(n5157), .B(
        n4776), .ZN(n4780) );
  OAI211_X1 U5870 ( .C1(n6463), .C2(n5128), .A(n4778), .B(n4777), .ZN(n4779)
         );
  NAND2_X1 U5871 ( .A1(n4780), .A2(n4779), .ZN(n4804) );
  NAND2_X1 U5872 ( .A1(n4804), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4785) );
  INV_X1 U5873 ( .A(n4928), .ZN(n4781) );
  NOR2_X1 U5874 ( .A1(n4781), .A2(n6519), .ZN(n4860) );
  AOI22_X1 U5875 ( .A1(n4860), .A2(n6458), .B1(n6456), .B2(n4782), .ZN(n4805)
         );
  OAI22_X1 U5876 ( .A1(n5190), .A2(n4806), .B1(n4805), .B2(n5194), .ZN(n4783)
         );
  AOI21_X1 U5877 ( .B1(n6563), .B2(n4808), .A(n4783), .ZN(n4784) );
  OAI211_X1 U5878 ( .C1(n5128), .C2(n6567), .A(n4785), .B(n4784), .ZN(U3058)
         );
  NAND2_X1 U5879 ( .A1(n4804), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4788) );
  OAI22_X1 U5880 ( .A1(n5175), .A2(n4806), .B1(n4805), .B2(n5179), .ZN(n4786)
         );
  AOI21_X1 U5881 ( .B1(n6557), .B2(n4808), .A(n4786), .ZN(n4787) );
  OAI211_X1 U5882 ( .C1(n5128), .C2(n6561), .A(n4788), .B(n4787), .ZN(U3057)
         );
  NAND2_X1 U5883 ( .A1(n4804), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4791) );
  OAI22_X1 U5884 ( .A1(n5165), .A2(n4806), .B1(n4805), .B2(n5169), .ZN(n4789)
         );
  AOI21_X1 U5885 ( .B1(n5053), .B2(n4808), .A(n4789), .ZN(n4790) );
  OAI211_X1 U5886 ( .C1(n5128), .C2(n5090), .A(n4791), .B(n4790), .ZN(U3054)
         );
  NAND2_X1 U5887 ( .A1(n4804), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4794) );
  OAI22_X1 U5888 ( .A1(n5185), .A2(n4806), .B1(n4805), .B2(n5189), .ZN(n4792)
         );
  AOI21_X1 U5889 ( .B1(n6531), .B2(n4808), .A(n4792), .ZN(n4793) );
  OAI211_X1 U5890 ( .C1(n5128), .C2(n6535), .A(n4794), .B(n4793), .ZN(U3053)
         );
  NAND2_X1 U5891 ( .A1(n4804), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4797) );
  OAI22_X1 U5892 ( .A1(n5180), .A2(n4806), .B1(n4805), .B2(n5184), .ZN(n4795)
         );
  AOI21_X1 U5893 ( .B1(n6570), .B2(n4808), .A(n4795), .ZN(n4796) );
  OAI211_X1 U5894 ( .C1(n5128), .C2(n6578), .A(n4797), .B(n4796), .ZN(U3059)
         );
  NAND2_X1 U5895 ( .A1(n4804), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4800) );
  OAI22_X1 U5896 ( .A1(n5170), .A2(n4806), .B1(n4805), .B2(n5174), .ZN(n4798)
         );
  AOI21_X1 U5897 ( .B1(n6551), .B2(n4808), .A(n4798), .ZN(n4799) );
  OAI211_X1 U5898 ( .C1(n5128), .C2(n6555), .A(n4800), .B(n4799), .ZN(U3056)
         );
  NAND2_X1 U5899 ( .A1(n4804), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4803) );
  OAI22_X1 U5900 ( .A1(n5201), .A2(n4806), .B1(n4805), .B2(n5206), .ZN(n4801)
         );
  AOI21_X1 U5901 ( .B1(n6545), .B2(n4808), .A(n4801), .ZN(n4802) );
  OAI211_X1 U5902 ( .C1(n5128), .C2(n6549), .A(n4803), .B(n4802), .ZN(U3055)
         );
  NAND2_X1 U5903 ( .A1(n4804), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4810) );
  OAI22_X1 U5904 ( .A1(n5195), .A2(n4806), .B1(n4805), .B2(n5932), .ZN(n4807)
         );
  AOI21_X1 U5905 ( .B1(n6513), .B2(n4808), .A(n4807), .ZN(n4809) );
  OAI211_X1 U5906 ( .C1(n5128), .C2(n6529), .A(n4810), .B(n4809), .ZN(U3052)
         );
  NAND3_X1 U5907 ( .A1(n4972), .A2(n5154), .A3(n6503), .ZN(n4811) );
  AND2_X1 U5908 ( .A1(n3256), .A2(n3171), .ZN(n4817) );
  AOI21_X1 U5909 ( .B1(n4811), .B2(n5914), .A(n4817), .ZN(n4816) );
  NAND3_X1 U5910 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6590), .A3(n6586), .ZN(n4968) );
  NOR2_X1 U5911 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4968), .ZN(n4845)
         );
  INV_X1 U5912 ( .A(n6456), .ZN(n4814) );
  OR2_X1 U5913 ( .A1(n5065), .A2(n4812), .ZN(n4818) );
  AOI21_X1 U5914 ( .B1(n4818), .B2(STATE2_REG_2__SCAN_IN), .A(n4813), .ZN(
        n4853) );
  OAI211_X1 U5915 ( .C1(n6683), .C2(n4845), .A(n4814), .B(n4853), .ZN(n4815)
         );
  NAND2_X1 U5916 ( .A1(n4842), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4823) );
  NAND2_X1 U5917 ( .A1(n4817), .A2(n5154), .ZN(n4820) );
  INV_X1 U5918 ( .A(n4818), .ZN(n4859) );
  NAND2_X1 U5919 ( .A1(n5157), .A2(n4859), .ZN(n4819) );
  AND2_X1 U5920 ( .A1(n4820), .A2(n4819), .ZN(n4843) );
  OAI22_X1 U5921 ( .A1(n6503), .A2(n6555), .B1(n4843), .B2(n5174), .ZN(n4821)
         );
  AOI21_X1 U5922 ( .B1(n6550), .B2(n4845), .A(n4821), .ZN(n4822) );
  OAI211_X1 U5923 ( .C1(n6486), .C2(n4972), .A(n4823), .B(n4822), .ZN(U3088)
         );
  NAND2_X1 U5924 ( .A1(n4842), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4826) );
  OAI22_X1 U5925 ( .A1(n6503), .A2(n6549), .B1(n4843), .B2(n5206), .ZN(n4824)
         );
  AOI21_X1 U5926 ( .B1(n6544), .B2(n4845), .A(n4824), .ZN(n4825) );
  OAI211_X1 U5927 ( .C1(n6482), .C2(n4972), .A(n4826), .B(n4825), .ZN(U3087)
         );
  NAND2_X1 U5928 ( .A1(n4842), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4829) );
  OAI22_X1 U5929 ( .A1(n6503), .A2(n6578), .B1(n4843), .B2(n5184), .ZN(n4827)
         );
  AOI21_X1 U5930 ( .B1(n6569), .B2(n4845), .A(n4827), .ZN(n4828) );
  OAI211_X1 U5931 ( .C1(n6502), .C2(n4972), .A(n4829), .B(n4828), .ZN(U3091)
         );
  NAND2_X1 U5932 ( .A1(n4842), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4832) );
  OAI22_X1 U5933 ( .A1(n6503), .A2(n6567), .B1(n4843), .B2(n5194), .ZN(n4830)
         );
  AOI21_X1 U5934 ( .B1(n6562), .B2(n4845), .A(n4830), .ZN(n4831) );
  OAI211_X1 U5935 ( .C1(n6494), .C2(n4972), .A(n4832), .B(n4831), .ZN(U3090)
         );
  NAND2_X1 U5936 ( .A1(n4842), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4835) );
  OAI22_X1 U5937 ( .A1(n6503), .A2(n6561), .B1(n4843), .B2(n5179), .ZN(n4833)
         );
  AOI21_X1 U5938 ( .B1(n6556), .B2(n4845), .A(n4833), .ZN(n4834) );
  OAI211_X1 U5939 ( .C1(n6490), .C2(n4972), .A(n4835), .B(n4834), .ZN(U3089)
         );
  NAND2_X1 U5940 ( .A1(n4842), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4838) );
  OAI22_X1 U5941 ( .A1(n6503), .A2(n5090), .B1(n4843), .B2(n5169), .ZN(n4836)
         );
  AOI21_X1 U5942 ( .B1(n6536), .B2(n4845), .A(n4836), .ZN(n4837) );
  OAI211_X1 U5943 ( .C1(n6543), .C2(n4972), .A(n4838), .B(n4837), .ZN(U3086)
         );
  NAND2_X1 U5944 ( .A1(n4842), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4841) );
  OAI22_X1 U5945 ( .A1(n6503), .A2(n6535), .B1(n4843), .B2(n5189), .ZN(n4839)
         );
  AOI21_X1 U5946 ( .B1(n6530), .B2(n4845), .A(n4839), .ZN(n4840) );
  OAI211_X1 U5947 ( .C1(n6476), .C2(n4972), .A(n4841), .B(n4840), .ZN(U3085)
         );
  NAND2_X1 U5948 ( .A1(n4842), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4847) );
  OAI22_X1 U5949 ( .A1(n6503), .A2(n6529), .B1(n4843), .B2(n5932), .ZN(n4844)
         );
  AOI21_X1 U5950 ( .B1(n6512), .B2(n4845), .A(n4844), .ZN(n4846) );
  OAI211_X1 U5951 ( .C1(n4972), .C2(n6472), .A(n4847), .B(n4846), .ZN(U3084)
         );
  NAND2_X1 U5952 ( .A1(n4931), .A2(n4850), .ZN(n4857) );
  AOI21_X1 U5953 ( .B1(n4857), .B2(n6542), .A(n6786), .ZN(n4851) );
  AOI211_X1 U5954 ( .C1(n4928), .C2(n4852), .A(n6519), .B(n4851), .ZN(n4856)
         );
  NOR2_X1 U5955 ( .A1(n6594), .A2(n4929), .ZN(n4933) );
  AND2_X1 U5956 ( .A1(n6580), .A2(n4933), .ZN(n4858) );
  INV_X1 U5957 ( .A(n5157), .ZN(n4854) );
  OAI211_X1 U5958 ( .C1(n6683), .C2(n4858), .A(n4854), .B(n4853), .ZN(n4855)
         );
  NAND2_X1 U5959 ( .A1(n4882), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4863)
         );
  INV_X1 U5960 ( .A(n4858), .ZN(n4884) );
  AOI22_X1 U5961 ( .A1(n4860), .A2(n3171), .B1(n6456), .B2(n4859), .ZN(n4883)
         );
  OAI22_X1 U5962 ( .A1(n5201), .A2(n4884), .B1(n4883), .B2(n5206), .ZN(n4861)
         );
  AOI21_X1 U5963 ( .B1(n6545), .B2(n4951), .A(n4861), .ZN(n4862) );
  OAI211_X1 U5964 ( .C1(n6542), .C2(n6549), .A(n4863), .B(n4862), .ZN(U3119)
         );
  NAND2_X1 U5965 ( .A1(n4882), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4866)
         );
  OAI22_X1 U5966 ( .A1(n5170), .A2(n4884), .B1(n4883), .B2(n5174), .ZN(n4864)
         );
  AOI21_X1 U5967 ( .B1(n6551), .B2(n4951), .A(n4864), .ZN(n4865) );
  OAI211_X1 U5968 ( .C1(n6542), .C2(n6555), .A(n4866), .B(n4865), .ZN(U3120)
         );
  NAND2_X1 U5969 ( .A1(n4882), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4869)
         );
  OAI22_X1 U5970 ( .A1(n5180), .A2(n4884), .B1(n4883), .B2(n5184), .ZN(n4867)
         );
  AOI21_X1 U5971 ( .B1(n6570), .B2(n4951), .A(n4867), .ZN(n4868) );
  OAI211_X1 U5972 ( .C1(n6542), .C2(n6578), .A(n4869), .B(n4868), .ZN(U3123)
         );
  NAND2_X1 U5973 ( .A1(n4882), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4872)
         );
  OAI22_X1 U5974 ( .A1(n5190), .A2(n4884), .B1(n4883), .B2(n5194), .ZN(n4870)
         );
  AOI21_X1 U5975 ( .B1(n6563), .B2(n4951), .A(n4870), .ZN(n4871) );
  OAI211_X1 U5976 ( .C1(n6542), .C2(n6567), .A(n4872), .B(n4871), .ZN(U3122)
         );
  NAND2_X1 U5977 ( .A1(n4882), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4875)
         );
  OAI22_X1 U5978 ( .A1(n5175), .A2(n4884), .B1(n4883), .B2(n5179), .ZN(n4873)
         );
  AOI21_X1 U5979 ( .B1(n6557), .B2(n4951), .A(n4873), .ZN(n4874) );
  OAI211_X1 U5980 ( .C1(n6542), .C2(n6561), .A(n4875), .B(n4874), .ZN(U3121)
         );
  NAND2_X1 U5981 ( .A1(n4882), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4878)
         );
  OAI22_X1 U5982 ( .A1(n5165), .A2(n4884), .B1(n4883), .B2(n5169), .ZN(n4876)
         );
  AOI21_X1 U5983 ( .B1(n5053), .B2(n4951), .A(n4876), .ZN(n4877) );
  OAI211_X1 U5984 ( .C1(n6542), .C2(n5090), .A(n4878), .B(n4877), .ZN(U3118)
         );
  NAND2_X1 U5985 ( .A1(n4882), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4881)
         );
  OAI22_X1 U5986 ( .A1(n5185), .A2(n4884), .B1(n4883), .B2(n5189), .ZN(n4879)
         );
  AOI21_X1 U5987 ( .B1(n6531), .B2(n4951), .A(n4879), .ZN(n4880) );
  OAI211_X1 U5988 ( .C1(n6542), .C2(n6535), .A(n4881), .B(n4880), .ZN(U3117)
         );
  NAND2_X1 U5989 ( .A1(n4882), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4887)
         );
  OAI22_X1 U5990 ( .A1(n5195), .A2(n4884), .B1(n4883), .B2(n5932), .ZN(n4885)
         );
  AOI21_X1 U5991 ( .B1(n6513), .B2(n4951), .A(n4885), .ZN(n4886) );
  OAI211_X1 U5992 ( .C1(n6542), .C2(n6529), .A(n4887), .B(n4886), .ZN(U3116)
         );
  XNOR2_X1 U5993 ( .A(n4889), .B(n4888), .ZN(n5140) );
  INV_X1 U5994 ( .A(n4890), .ZN(n4891) );
  XNOR2_X1 U5995 ( .A(n4892), .B(n4891), .ZN(n6154) );
  INV_X1 U5996 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6652) );
  NOR2_X1 U5997 ( .A1(n6392), .A2(n6652), .ZN(n5135) );
  NOR2_X1 U5999 ( .A1(n4893), .A2(n4993), .ZN(n5143) );
  NAND2_X1 U6000 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n5143), .ZN(n4895)
         );
  INV_X1 U6001 ( .A(n6437), .ZN(n4894) );
  AOI21_X1 U6002 ( .B1(n4895), .B2(n6403), .A(n4894), .ZN(n5003) );
  OAI33_X1 U6003 ( .A1(1'b0), .A2(n5003), .A3(n4297), .B1(
        INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n5144), .B3(n4895), .ZN(n4897) );
  AOI211_X1 U6004 ( .C1(n6445), .C2(n6154), .A(n5135), .B(n4897), .ZN(n4898)
         );
  OAI21_X1 U6005 ( .B1(n6394), .B2(n5140), .A(n4898), .ZN(U3012) );
  NOR2_X1 U6006 ( .A1(n6580), .A2(n4904), .ZN(n4923) );
  AOI21_X1 U6007 ( .B1(n4900), .B2(n3491), .A(n4923), .ZN(n4905) );
  AOI21_X1 U6008 ( .B1(n4901), .B2(STATEBS16_REG_SCAN_IN), .A(n6519), .ZN(
        n4903) );
  AOI22_X1 U6009 ( .A1(n4905), .A2(n4903), .B1(n6519), .B2(n4904), .ZN(n4902)
         );
  NAND2_X1 U6010 ( .A1(n6521), .A2(n4902), .ZN(n4922) );
  INV_X1 U6011 ( .A(n4903), .ZN(n4906) );
  OAI22_X1 U6012 ( .A1(n4906), .A2(n4905), .B1(n4969), .B2(n4904), .ZN(n4921)
         );
  AOI22_X1 U6013 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4922), .B1(n6546), 
        .B2(n4921), .ZN(n4908) );
  AOI22_X1 U6014 ( .A1(n4924), .A2(n6479), .B1(n6544), .B2(n4923), .ZN(n4907)
         );
  OAI211_X1 U6015 ( .C1(n6482), .C2(n5056), .A(n4908), .B(n4907), .ZN(U3031)
         );
  AOI22_X1 U6016 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4922), .B1(n6552), 
        .B2(n4921), .ZN(n4910) );
  AOI22_X1 U6017 ( .A1(n4924), .A2(n6483), .B1(n6550), .B2(n4923), .ZN(n4909)
         );
  OAI211_X1 U6018 ( .C1(n6486), .C2(n5056), .A(n4910), .B(n4909), .ZN(U3032)
         );
  AOI22_X1 U6019 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4922), .B1(n6526), 
        .B2(n4921), .ZN(n4912) );
  AOI22_X1 U6020 ( .A1(n4924), .A2(n6469), .B1(n6512), .B2(n4923), .ZN(n4911)
         );
  OAI211_X1 U6021 ( .C1(n6472), .C2(n5056), .A(n4912), .B(n4911), .ZN(U3028)
         );
  AOI22_X1 U6022 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4922), .B1(n6573), 
        .B2(n4921), .ZN(n4914) );
  AOI22_X1 U6023 ( .A1(n4924), .A2(n6498), .B1(n6569), .B2(n4923), .ZN(n4913)
         );
  OAI211_X1 U6024 ( .C1(n6502), .C2(n5056), .A(n4914), .B(n4913), .ZN(U3035)
         );
  AOI22_X1 U6025 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4922), .B1(n6539), 
        .B2(n4921), .ZN(n4916) );
  AOI22_X1 U6026 ( .A1(n4924), .A2(n6537), .B1(n6536), .B2(n4923), .ZN(n4915)
         );
  OAI211_X1 U6027 ( .C1(n6543), .C2(n5056), .A(n4916), .B(n4915), .ZN(U3030)
         );
  AOI22_X1 U6028 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4922), .B1(n6564), 
        .B2(n4921), .ZN(n4918) );
  AOI22_X1 U6029 ( .A1(n4924), .A2(n6491), .B1(n6562), .B2(n4923), .ZN(n4917)
         );
  OAI211_X1 U6030 ( .C1(n6494), .C2(n5056), .A(n4918), .B(n4917), .ZN(U3034)
         );
  AOI22_X1 U6031 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4922), .B1(n6532), 
        .B2(n4921), .ZN(n4920) );
  AOI22_X1 U6032 ( .A1(n4924), .A2(n6473), .B1(n6530), .B2(n4923), .ZN(n4919)
         );
  OAI211_X1 U6033 ( .C1(n6476), .C2(n5056), .A(n4920), .B(n4919), .ZN(U3029)
         );
  AOI22_X1 U6034 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4922), .B1(n6558), 
        .B2(n4921), .ZN(n4926) );
  AOI22_X1 U6035 ( .A1(n4924), .A2(n6487), .B1(n6556), .B2(n4923), .ZN(n4925)
         );
  OAI211_X1 U6036 ( .C1(n6490), .C2(n5056), .A(n4926), .B(n4925), .ZN(U3033)
         );
  AND2_X1 U6037 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4933), .ZN(n4927)
         );
  INV_X1 U6038 ( .A(n4927), .ZN(n4956) );
  AOI22_X1 U6039 ( .A1(n4951), .A2(n6537), .B1(n5936), .B2(n5053), .ZN(n4938)
         );
  AOI21_X1 U6040 ( .B1(n4964), .B2(n4928), .A(n4927), .ZN(n4932) );
  NAND2_X1 U6041 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4930) );
  OAI22_X1 U6042 ( .A1(n4932), .A2(n6519), .B1(n4930), .B2(n4929), .ZN(n4953)
         );
  NAND2_X1 U6043 ( .A1(n4931), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5095) );
  NAND2_X1 U6044 ( .A1(n4932), .A2(n5095), .ZN(n4936) );
  INV_X1 U6045 ( .A(n4933), .ZN(n4934) );
  NAND2_X1 U6046 ( .A1(n6519), .A2(n4934), .ZN(n4935) );
  OAI211_X1 U6047 ( .C1(n6519), .C2(n4936), .A(n6521), .B(n4935), .ZN(n4952)
         );
  AOI22_X1 U6048 ( .A1(n4953), .A2(n6539), .B1(INSTQUEUE_REG_13__2__SCAN_IN), 
        .B2(n4952), .ZN(n4937) );
  OAI211_X1 U6049 ( .C1(n5165), .C2(n4956), .A(n4938), .B(n4937), .ZN(U3126)
         );
  AOI22_X1 U6050 ( .A1(n4951), .A2(n6473), .B1(n5936), .B2(n6531), .ZN(n4940)
         );
  AOI22_X1 U6051 ( .A1(n4953), .A2(n6532), .B1(INSTQUEUE_REG_13__1__SCAN_IN), 
        .B2(n4952), .ZN(n4939) );
  OAI211_X1 U6052 ( .C1(n5185), .C2(n4956), .A(n4940), .B(n4939), .ZN(U3125)
         );
  AOI22_X1 U6053 ( .A1(n4951), .A2(n6483), .B1(n5936), .B2(n6551), .ZN(n4942)
         );
  AOI22_X1 U6054 ( .A1(n4953), .A2(n6552), .B1(INSTQUEUE_REG_13__4__SCAN_IN), 
        .B2(n4952), .ZN(n4941) );
  OAI211_X1 U6055 ( .C1(n5170), .C2(n4956), .A(n4942), .B(n4941), .ZN(U3128)
         );
  AOI22_X1 U6056 ( .A1(n4951), .A2(n6479), .B1(n5936), .B2(n6545), .ZN(n4944)
         );
  AOI22_X1 U6057 ( .A1(n4953), .A2(n6546), .B1(INSTQUEUE_REG_13__3__SCAN_IN), 
        .B2(n4952), .ZN(n4943) );
  OAI211_X1 U6058 ( .C1(n5201), .C2(n4956), .A(n4944), .B(n4943), .ZN(U3127)
         );
  AOI22_X1 U6059 ( .A1(n4951), .A2(n6498), .B1(n5936), .B2(n6570), .ZN(n4946)
         );
  AOI22_X1 U6060 ( .A1(n4953), .A2(n6573), .B1(INSTQUEUE_REG_13__7__SCAN_IN), 
        .B2(n4952), .ZN(n4945) );
  OAI211_X1 U6061 ( .C1(n5180), .C2(n4956), .A(n4946), .B(n4945), .ZN(U3131)
         );
  AOI22_X1 U6062 ( .A1(n4951), .A2(n6469), .B1(n5936), .B2(n6513), .ZN(n4948)
         );
  AOI22_X1 U6063 ( .A1(n4953), .A2(n6526), .B1(INSTQUEUE_REG_13__0__SCAN_IN), 
        .B2(n4952), .ZN(n4947) );
  OAI211_X1 U6064 ( .C1(n5195), .C2(n4956), .A(n4948), .B(n4947), .ZN(U3124)
         );
  AOI22_X1 U6065 ( .A1(n4951), .A2(n6487), .B1(n5936), .B2(n6557), .ZN(n4950)
         );
  AOI22_X1 U6066 ( .A1(n4953), .A2(n6558), .B1(INSTQUEUE_REG_13__5__SCAN_IN), 
        .B2(n4952), .ZN(n4949) );
  OAI211_X1 U6067 ( .C1(n5175), .C2(n4956), .A(n4950), .B(n4949), .ZN(U3129)
         );
  AOI22_X1 U6068 ( .A1(n4951), .A2(n6491), .B1(n5936), .B2(n6563), .ZN(n4955)
         );
  AOI22_X1 U6069 ( .A1(n4953), .A2(n6564), .B1(INSTQUEUE_REG_13__6__SCAN_IN), 
        .B2(n4952), .ZN(n4954) );
  OAI211_X1 U6070 ( .C1(n5190), .C2(n4956), .A(n4955), .B(n4954), .ZN(U3130)
         );
  INV_X1 U6071 ( .A(EAX_REG_24__SCAN_IN), .ZN(n6290) );
  AOI22_X1 U6072 ( .A1(n6267), .A2(UWORD_REG_8__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4957) );
  OAI21_X1 U6073 ( .B1(n6290), .B2(n5012), .A(n4957), .ZN(U2899) );
  INV_X1 U6074 ( .A(EAX_REG_28__SCAN_IN), .ZN(n6296) );
  AOI22_X1 U6075 ( .A1(n6267), .A2(UWORD_REG_12__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4958) );
  OAI21_X1 U6076 ( .B1(n6296), .B2(n5012), .A(n4958), .ZN(U2895) );
  INV_X1 U6077 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6299) );
  AOI22_X1 U6078 ( .A1(n6267), .A2(UWORD_REG_14__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4959) );
  OAI21_X1 U6079 ( .B1(n6299), .B2(n5012), .A(n4959), .ZN(U2893) );
  INV_X1 U6080 ( .A(EAX_REG_26__SCAN_IN), .ZN(n6293) );
  AOI22_X1 U6081 ( .A1(n6267), .A2(UWORD_REG_10__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4960) );
  OAI21_X1 U6082 ( .B1(n6293), .B2(n5012), .A(n4960), .ZN(U2897) );
  INV_X1 U6083 ( .A(n4961), .ZN(n4963) );
  NOR2_X1 U6084 ( .A1(n6580), .A2(n4968), .ZN(n4989) );
  AOI21_X1 U6085 ( .B1(n4964), .B2(n3256), .A(n4989), .ZN(n4971) );
  OR3_X1 U6086 ( .A1(n6514), .A2(n5902), .A3(n6786), .ZN(n4965) );
  AOI22_X1 U6087 ( .A1(n4971), .A2(n4967), .B1(n6519), .B2(n4968), .ZN(n4966)
         );
  NAND2_X1 U6088 ( .A1(n6521), .A2(n4966), .ZN(n4988) );
  INV_X1 U6089 ( .A(n4967), .ZN(n4970) );
  OAI22_X1 U6090 ( .A1(n4971), .A2(n4970), .B1(n4969), .B2(n4968), .ZN(n4987)
         );
  AOI22_X1 U6091 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4988), .B1(n6526), 
        .B2(n4987), .ZN(n4974) );
  AOI22_X1 U6092 ( .A1(n4990), .A2(n6469), .B1(n6512), .B2(n4989), .ZN(n4973)
         );
  OAI211_X1 U6093 ( .C1(n5152), .C2(n6472), .A(n4974), .B(n4973), .ZN(U3092)
         );
  AOI22_X1 U6094 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4988), .B1(n6532), 
        .B2(n4987), .ZN(n4976) );
  AOI22_X1 U6095 ( .A1(n4990), .A2(n6473), .B1(n4989), .B2(n6530), .ZN(n4975)
         );
  OAI211_X1 U6096 ( .C1(n5152), .C2(n6476), .A(n4976), .B(n4975), .ZN(U3093)
         );
  AOI22_X1 U6097 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4988), .B1(n6546), 
        .B2(n4987), .ZN(n4978) );
  AOI22_X1 U6098 ( .A1(n4990), .A2(n6479), .B1(n4989), .B2(n6544), .ZN(n4977)
         );
  OAI211_X1 U6099 ( .C1(n5152), .C2(n6482), .A(n4978), .B(n4977), .ZN(U3095)
         );
  AOI22_X1 U6100 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4988), .B1(n6539), 
        .B2(n4987), .ZN(n4980) );
  AOI22_X1 U6101 ( .A1(n4990), .A2(n6537), .B1(n4989), .B2(n6536), .ZN(n4979)
         );
  OAI211_X1 U6102 ( .C1(n5152), .C2(n6543), .A(n4980), .B(n4979), .ZN(U3094)
         );
  AOI22_X1 U6103 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4988), .B1(n6564), 
        .B2(n4987), .ZN(n4982) );
  AOI22_X1 U6104 ( .A1(n4990), .A2(n6491), .B1(n4989), .B2(n6562), .ZN(n4981)
         );
  OAI211_X1 U6105 ( .C1(n5152), .C2(n6494), .A(n4982), .B(n4981), .ZN(U3098)
         );
  AOI22_X1 U6106 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4988), .B1(n6573), 
        .B2(n4987), .ZN(n4984) );
  AOI22_X1 U6107 ( .A1(n4990), .A2(n6498), .B1(n4989), .B2(n6569), .ZN(n4983)
         );
  OAI211_X1 U6108 ( .C1(n5152), .C2(n6502), .A(n4984), .B(n4983), .ZN(U3099)
         );
  AOI22_X1 U6109 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4988), .B1(n6558), 
        .B2(n4987), .ZN(n4986) );
  AOI22_X1 U6110 ( .A1(n4990), .A2(n6487), .B1(n4989), .B2(n6556), .ZN(n4985)
         );
  OAI211_X1 U6111 ( .C1(n5152), .C2(n6490), .A(n4986), .B(n4985), .ZN(U3097)
         );
  AOI22_X1 U6112 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4988), .B1(n6552), 
        .B2(n4987), .ZN(n4992) );
  AOI22_X1 U6113 ( .A1(n4990), .A2(n6483), .B1(n4989), .B2(n6550), .ZN(n4991)
         );
  OAI211_X1 U6114 ( .C1(n5152), .C2(n6486), .A(n4992), .B(n4991), .ZN(U3096)
         );
  AOI21_X1 U6115 ( .B1(n6425), .B2(n5143), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n5002) );
  NOR2_X1 U6116 ( .A1(n4994), .A2(n4993), .ZN(n5145) );
  NOR2_X1 U6117 ( .A1(n5385), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4995)
         );
  NAND2_X1 U6118 ( .A1(n5145), .A2(n4995), .ZN(n4996) );
  NAND2_X1 U6119 ( .A1(n6427), .A2(REIP_REG_5__SCAN_IN), .ZN(n6370) );
  NAND2_X1 U6120 ( .A1(n4996), .A2(n6370), .ZN(n4997) );
  AOI21_X1 U6121 ( .B1(n6445), .B2(n6172), .A(n4997), .ZN(n5001) );
  XOR2_X1 U6122 ( .A(n3162), .B(n4999), .Z(n6369) );
  NAND2_X1 U6123 ( .A1(n6369), .A2(n6439), .ZN(n5000) );
  OAI211_X1 U6124 ( .C1(n5003), .C2(n5002), .A(n5001), .B(n5000), .ZN(U3013)
         );
  INV_X1 U6125 ( .A(EAX_REG_19__SCAN_IN), .ZN(n6280) );
  INV_X2 U6126 ( .A(n6606), .ZN(n6267) );
  AOI22_X1 U6127 ( .A1(n6267), .A2(UWORD_REG_3__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n5004) );
  OAI21_X1 U6128 ( .B1(n6280), .B2(n5012), .A(n5004), .ZN(U2904) );
  INV_X1 U6129 ( .A(EAX_REG_17__SCAN_IN), .ZN(n6276) );
  AOI22_X1 U6130 ( .A1(n6267), .A2(UWORD_REG_1__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n5005) );
  OAI21_X1 U6131 ( .B1(n6276), .B2(n5012), .A(n5005), .ZN(U2906) );
  INV_X1 U6132 ( .A(EAX_REG_18__SCAN_IN), .ZN(n6278) );
  AOI22_X1 U6133 ( .A1(n6267), .A2(UWORD_REG_2__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n5006) );
  OAI21_X1 U6134 ( .B1(n6278), .B2(n5012), .A(n5006), .ZN(U2905) );
  INV_X1 U6135 ( .A(EAX_REG_22__SCAN_IN), .ZN(n6287) );
  AOI22_X1 U6136 ( .A1(n6267), .A2(UWORD_REG_6__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n5007) );
  OAI21_X1 U6137 ( .B1(n6287), .B2(n5012), .A(n5007), .ZN(U2901) );
  INV_X1 U6138 ( .A(EAX_REG_21__SCAN_IN), .ZN(n6285) );
  AOI22_X1 U6139 ( .A1(n6267), .A2(UWORD_REG_5__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n5008) );
  OAI21_X1 U6140 ( .B1(n6285), .B2(n5012), .A(n5008), .ZN(U2902) );
  AOI22_X1 U6141 ( .A1(n6267), .A2(UWORD_REG_7__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n5009) );
  OAI21_X1 U6142 ( .B1(n3905), .B2(n5012), .A(n5009), .ZN(U2900) );
  INV_X1 U6143 ( .A(EAX_REG_20__SCAN_IN), .ZN(n6282) );
  AOI22_X1 U6144 ( .A1(n6267), .A2(UWORD_REG_4__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n5010) );
  OAI21_X1 U6145 ( .B1(n6282), .B2(n5012), .A(n5010), .ZN(U2903) );
  INV_X1 U6146 ( .A(EAX_REG_16__SCAN_IN), .ZN(n6274) );
  AOI22_X1 U6147 ( .A1(n6267), .A2(UWORD_REG_0__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n5011) );
  OAI21_X1 U6148 ( .B1(n6274), .B2(n5012), .A(n5011), .ZN(U2907) );
  AND2_X1 U6149 ( .A1(n5013), .A2(n4765), .ZN(n5015) );
  OR2_X1 U6150 ( .A1(n5015), .A2(n5014), .ZN(n6161) );
  OAI222_X1 U6151 ( .A1(n6161), .A2(n5983), .B1(n5360), .B2(n5016), .C1(n6319), 
        .C2(n5449), .ZN(U2885) );
  INV_X1 U6152 ( .A(n6154), .ZN(n5017) );
  OAI222_X1 U6153 ( .A1(n6161), .A2(n6226), .B1(n5018), .B2(n6238), .C1(n6233), 
        .C2(n5017), .ZN(U2853) );
  INV_X1 U6154 ( .A(n5056), .ZN(n5021) );
  NAND2_X1 U6155 ( .A1(n5019), .A2(n4587), .ZN(n5020) );
  OAI21_X1 U6156 ( .B1(n5021), .B2(n3257), .A(n5914), .ZN(n5022) );
  NOR2_X1 U6157 ( .A1(n4547), .A2(n6214), .ZN(n5156) );
  NAND2_X1 U6158 ( .A1(n6458), .A2(n5156), .ZN(n5097) );
  AOI21_X1 U6159 ( .B1(n5022), .B2(n5097), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n5024) );
  NAND3_X1 U6160 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6594), .A3(n6590), .ZN(n5104) );
  NOR2_X1 U6161 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5104), .ZN(n5025)
         );
  OAI21_X1 U6162 ( .B1(n5065), .B2(n4969), .A(n5023), .ZN(n5058) );
  NOR2_X1 U6163 ( .A1(n6456), .A2(n5058), .ZN(n5162) );
  NAND2_X1 U6164 ( .A1(n5049), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5030) );
  INV_X1 U6165 ( .A(n5025), .ZN(n5051) );
  INV_X1 U6166 ( .A(n5097), .ZN(n5027) );
  INV_X1 U6167 ( .A(n5065), .ZN(n5026) );
  NOR2_X1 U6168 ( .A1(n5026), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6457)
         );
  AOI22_X1 U6169 ( .A1(n5027), .A2(n5154), .B1(n5157), .B2(n6457), .ZN(n5050)
         );
  OAI22_X1 U6170 ( .A1(n5201), .A2(n5051), .B1(n5050), .B2(n5206), .ZN(n5028)
         );
  AOI21_X1 U6171 ( .B1(n6545), .B2(n3257), .A(n5028), .ZN(n5029) );
  OAI211_X1 U6172 ( .C1(n5056), .C2(n6549), .A(n5030), .B(n5029), .ZN(U3039)
         );
  NAND2_X1 U6173 ( .A1(n5049), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5033) );
  OAI22_X1 U6174 ( .A1(n5185), .A2(n5051), .B1(n5050), .B2(n5189), .ZN(n5031)
         );
  AOI21_X1 U6175 ( .B1(n6531), .B2(n3257), .A(n5031), .ZN(n5032) );
  OAI211_X1 U6176 ( .C1(n5056), .C2(n6535), .A(n5033), .B(n5032), .ZN(U3037)
         );
  NAND2_X1 U6177 ( .A1(n5049), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5036) );
  OAI22_X1 U6178 ( .A1(n5195), .A2(n5051), .B1(n5050), .B2(n5932), .ZN(n5034)
         );
  AOI21_X1 U6179 ( .B1(n6513), .B2(n3257), .A(n5034), .ZN(n5035) );
  OAI211_X1 U6180 ( .C1(n5056), .C2(n6529), .A(n5036), .B(n5035), .ZN(U3036)
         );
  NAND2_X1 U6181 ( .A1(n5049), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5039) );
  OAI22_X1 U6182 ( .A1(n5175), .A2(n5051), .B1(n5050), .B2(n5179), .ZN(n5037)
         );
  AOI21_X1 U6183 ( .B1(n6557), .B2(n3257), .A(n5037), .ZN(n5038) );
  OAI211_X1 U6184 ( .C1(n5056), .C2(n6561), .A(n5039), .B(n5038), .ZN(U3041)
         );
  NAND2_X1 U6185 ( .A1(n5049), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5042) );
  OAI22_X1 U6186 ( .A1(n5170), .A2(n5051), .B1(n5050), .B2(n5174), .ZN(n5040)
         );
  AOI21_X1 U6187 ( .B1(n6551), .B2(n3257), .A(n5040), .ZN(n5041) );
  OAI211_X1 U6188 ( .C1(n5056), .C2(n6555), .A(n5042), .B(n5041), .ZN(U3040)
         );
  NAND2_X1 U6189 ( .A1(n5049), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5045) );
  OAI22_X1 U6190 ( .A1(n5180), .A2(n5051), .B1(n5050), .B2(n5184), .ZN(n5043)
         );
  AOI21_X1 U6191 ( .B1(n6570), .B2(n3257), .A(n5043), .ZN(n5044) );
  OAI211_X1 U6192 ( .C1(n5056), .C2(n6578), .A(n5045), .B(n5044), .ZN(U3043)
         );
  NAND2_X1 U6193 ( .A1(n5049), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5048) );
  OAI22_X1 U6194 ( .A1(n5190), .A2(n5051), .B1(n5050), .B2(n5194), .ZN(n5046)
         );
  AOI21_X1 U6195 ( .B1(n6563), .B2(n3257), .A(n5046), .ZN(n5047) );
  OAI211_X1 U6196 ( .C1(n5056), .C2(n6567), .A(n5048), .B(n5047), .ZN(U3042)
         );
  NAND2_X1 U6197 ( .A1(n5049), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5055) );
  OAI22_X1 U6198 ( .A1(n5165), .A2(n5051), .B1(n5050), .B2(n5169), .ZN(n5052)
         );
  AOI21_X1 U6199 ( .B1(n5053), .B2(n3257), .A(n5052), .ZN(n5054) );
  OAI211_X1 U6200 ( .C1(n5056), .C2(n5090), .A(n5055), .B(n5054), .ZN(U3038)
         );
  NOR3_X1 U6201 ( .A1(n5936), .A2(n5935), .A3(n6519), .ZN(n5057) );
  OAI21_X1 U6202 ( .B1(n5057), .B2(n6463), .A(n5064), .ZN(n5063) );
  NOR2_X1 U6203 ( .A1(n5157), .A2(n5058), .ZN(n6467) );
  INV_X1 U6204 ( .A(n5059), .ZN(n5060) );
  NOR2_X1 U6205 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5060), .ZN(n5937)
         );
  INV_X1 U6206 ( .A(n5937), .ZN(n5061) );
  AOI21_X1 U6207 ( .B1(n5061), .B2(STATE2_REG_3__SCAN_IN), .A(n6594), .ZN(
        n5062) );
  NAND3_X1 U6208 ( .A1(n5063), .A2(n6467), .A3(n5062), .ZN(n5931) );
  NAND2_X1 U6209 ( .A1(n5931), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5070)
         );
  INV_X1 U6210 ( .A(n5935), .ZN(n5086) );
  NOR2_X1 U6211 ( .A1(n5064), .A2(n6519), .ZN(n6459) );
  NAND2_X1 U6212 ( .A1(n6459), .A2(n3171), .ZN(n5067) );
  AND2_X1 U6213 ( .A1(n5065), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5158)
         );
  NAND2_X1 U6214 ( .A1(n6456), .A2(n5158), .ZN(n5066) );
  OAI22_X1 U6215 ( .A1(n5086), .A2(n6490), .B1(n5933), .B2(n5179), .ZN(n5068)
         );
  AOI21_X1 U6216 ( .B1(n6556), .B2(n5937), .A(n5068), .ZN(n5069) );
  OAI211_X1 U6217 ( .C1(n5091), .C2(n6561), .A(n5070), .B(n5069), .ZN(U3137)
         );
  NAND2_X1 U6218 ( .A1(n5931), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5073)
         );
  OAI22_X1 U6219 ( .A1(n5086), .A2(n6486), .B1(n5933), .B2(n5174), .ZN(n5071)
         );
  AOI21_X1 U6220 ( .B1(n6550), .B2(n5937), .A(n5071), .ZN(n5072) );
  OAI211_X1 U6221 ( .C1(n5091), .C2(n6555), .A(n5073), .B(n5072), .ZN(U3136)
         );
  NAND2_X1 U6222 ( .A1(n5931), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5076)
         );
  OAI22_X1 U6223 ( .A1(n5086), .A2(n6476), .B1(n5933), .B2(n5189), .ZN(n5074)
         );
  AOI21_X1 U6224 ( .B1(n6530), .B2(n5937), .A(n5074), .ZN(n5075) );
  OAI211_X1 U6225 ( .C1(n5091), .C2(n6535), .A(n5076), .B(n5075), .ZN(U3133)
         );
  NAND2_X1 U6226 ( .A1(n5931), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5079)
         );
  OAI22_X1 U6227 ( .A1(n5086), .A2(n6502), .B1(n5933), .B2(n5184), .ZN(n5077)
         );
  AOI21_X1 U6228 ( .B1(n6569), .B2(n5937), .A(n5077), .ZN(n5078) );
  OAI211_X1 U6229 ( .C1(n5091), .C2(n6578), .A(n5079), .B(n5078), .ZN(U3139)
         );
  NAND2_X1 U6230 ( .A1(n5931), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5082)
         );
  OAI22_X1 U6231 ( .A1(n5086), .A2(n6494), .B1(n5933), .B2(n5194), .ZN(n5080)
         );
  AOI21_X1 U6232 ( .B1(n6562), .B2(n5937), .A(n5080), .ZN(n5081) );
  OAI211_X1 U6233 ( .C1(n5091), .C2(n6567), .A(n5082), .B(n5081), .ZN(U3138)
         );
  NAND2_X1 U6234 ( .A1(n5931), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5085)
         );
  OAI22_X1 U6235 ( .A1(n5086), .A2(n6482), .B1(n5933), .B2(n5206), .ZN(n5083)
         );
  AOI21_X1 U6236 ( .B1(n6544), .B2(n5937), .A(n5083), .ZN(n5084) );
  OAI211_X1 U6237 ( .C1(n5091), .C2(n6549), .A(n5085), .B(n5084), .ZN(U3135)
         );
  NAND2_X1 U6238 ( .A1(n5931), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5089)
         );
  OAI22_X1 U6239 ( .A1(n5086), .A2(n6543), .B1(n5933), .B2(n5169), .ZN(n5087)
         );
  AOI21_X1 U6240 ( .B1(n6536), .B2(n5937), .A(n5087), .ZN(n5088) );
  OAI211_X1 U6241 ( .C1(n5091), .C2(n5090), .A(n5089), .B(n5088), .ZN(U3134)
         );
  NOR2_X1 U6242 ( .A1(n5014), .A2(n5093), .ZN(n5094) );
  OR2_X1 U6243 ( .A1(n5092), .A2(n5094), .ZN(n6360) );
  OAI222_X1 U6244 ( .A1(n6360), .A2(n5983), .B1(n5360), .B2(n6950), .C1(n5449), 
        .C2(n3655), .ZN(U2884) );
  NAND2_X1 U6245 ( .A1(n5095), .A2(n6514), .ZN(n5908) );
  NOR3_X1 U6246 ( .A1(n5908), .A2(n4586), .A3(n5905), .ZN(n5096) );
  NOR2_X1 U6247 ( .A1(n5096), .A2(n6519), .ZN(n5102) );
  OR2_X1 U6248 ( .A1(n5097), .A2(n5233), .ZN(n5099) );
  INV_X1 U6249 ( .A(n6511), .ZN(n5098) );
  NAND2_X1 U6250 ( .A1(n5098), .A2(n6594), .ZN(n5129) );
  NAND2_X1 U6251 ( .A1(n5099), .A2(n5129), .ZN(n5106) );
  INV_X1 U6252 ( .A(n5104), .ZN(n5100) );
  AOI22_X1 U6253 ( .A1(n5102), .A2(n5106), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5100), .ZN(n5134) );
  OAI22_X1 U6254 ( .A1(n5170), .A2(n5129), .B1(n6486), .B2(n5128), .ZN(n5101)
         );
  AOI21_X1 U6255 ( .B1(n6483), .B2(n3257), .A(n5101), .ZN(n5109) );
  INV_X1 U6256 ( .A(n5102), .ZN(n5107) );
  AOI21_X1 U6257 ( .B1(n6519), .B2(n5104), .A(n5103), .ZN(n5105) );
  NAND2_X1 U6258 ( .A1(n5131), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n5108) );
  OAI211_X1 U6259 ( .C1(n5134), .C2(n5174), .A(n5109), .B(n5108), .ZN(U3048)
         );
  OAI22_X1 U6260 ( .A1(n5195), .A2(n5129), .B1(n6472), .B2(n5128), .ZN(n5110)
         );
  AOI21_X1 U6261 ( .B1(n6469), .B2(n3257), .A(n5110), .ZN(n5112) );
  NAND2_X1 U6262 ( .A1(n5131), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n5111) );
  OAI211_X1 U6263 ( .C1(n5134), .C2(n5932), .A(n5112), .B(n5111), .ZN(U3044)
         );
  OAI22_X1 U6264 ( .A1(n5201), .A2(n5129), .B1(n6482), .B2(n5128), .ZN(n5113)
         );
  AOI21_X1 U6265 ( .B1(n6479), .B2(n3257), .A(n5113), .ZN(n5115) );
  NAND2_X1 U6266 ( .A1(n5131), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n5114) );
  OAI211_X1 U6267 ( .C1(n5134), .C2(n5206), .A(n5115), .B(n5114), .ZN(U3047)
         );
  OAI22_X1 U6268 ( .A1(n5190), .A2(n5129), .B1(n6494), .B2(n5128), .ZN(n5116)
         );
  AOI21_X1 U6269 ( .B1(n6491), .B2(n3257), .A(n5116), .ZN(n5118) );
  NAND2_X1 U6270 ( .A1(n5131), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n5117) );
  OAI211_X1 U6271 ( .C1(n5134), .C2(n5194), .A(n5118), .B(n5117), .ZN(U3050)
         );
  OAI22_X1 U6272 ( .A1(n5185), .A2(n5129), .B1(n6476), .B2(n5128), .ZN(n5119)
         );
  AOI21_X1 U6273 ( .B1(n6473), .B2(n3257), .A(n5119), .ZN(n5121) );
  NAND2_X1 U6274 ( .A1(n5131), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n5120) );
  OAI211_X1 U6275 ( .C1(n5134), .C2(n5189), .A(n5121), .B(n5120), .ZN(U3045)
         );
  OAI22_X1 U6276 ( .A1(n5180), .A2(n5129), .B1(n6502), .B2(n5128), .ZN(n5122)
         );
  AOI21_X1 U6277 ( .B1(n6498), .B2(n3257), .A(n5122), .ZN(n5124) );
  NAND2_X1 U6278 ( .A1(n5131), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5123) );
  OAI211_X1 U6279 ( .C1(n5134), .C2(n5184), .A(n5124), .B(n5123), .ZN(U3051)
         );
  OAI22_X1 U6280 ( .A1(n5165), .A2(n5129), .B1(n6543), .B2(n5128), .ZN(n5125)
         );
  AOI21_X1 U6281 ( .B1(n6537), .B2(n3257), .A(n5125), .ZN(n5127) );
  NAND2_X1 U6282 ( .A1(n5131), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n5126) );
  OAI211_X1 U6283 ( .C1(n5134), .C2(n5169), .A(n5127), .B(n5126), .ZN(U3046)
         );
  OAI22_X1 U6284 ( .A1(n5175), .A2(n5129), .B1(n6490), .B2(n5128), .ZN(n5130)
         );
  AOI21_X1 U6285 ( .B1(n6487), .B2(n3257), .A(n5130), .ZN(n5133) );
  NAND2_X1 U6286 ( .A1(n5131), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n5132) );
  OAI211_X1 U6287 ( .C1(n5134), .C2(n5179), .A(n5133), .B(n5132), .ZN(U3049)
         );
  INV_X1 U6288 ( .A(n6161), .ZN(n5138) );
  AOI21_X1 U6289 ( .B1(n6383), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n5135), 
        .ZN(n5136) );
  OAI21_X1 U6290 ( .B1(n6165), .B2(n6391), .A(n5136), .ZN(n5137) );
  AOI21_X1 U6291 ( .B1(n5138), .B2(n6379), .A(n5137), .ZN(n5139) );
  OAI21_X1 U6292 ( .B1(n6357), .B2(n5140), .A(n5139), .ZN(U2980) );
  XNOR2_X1 U6293 ( .A(n3161), .B(n5142), .ZN(n5255) );
  NAND3_X1 U6294 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n5143), .ZN(n5312) );
  NOR2_X1 U6295 ( .A1(n5312), .A2(n5144), .ZN(n6406) );
  NAND2_X1 U6296 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6404) );
  OAI211_X1 U6297 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6406), .B(n6404), .ZN(n5151) );
  NAND3_X1 U6298 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n5145), .ZN(n5311) );
  AOI22_X1 U6299 ( .A1(n6425), .A2(n5312), .B1(n5858), .B2(n5311), .ZN(n5146)
         );
  NAND2_X1 U6300 ( .A1(n5381), .A2(n5146), .ZN(n6402) );
  OAI21_X1 U6301 ( .B1(n5148), .B2(n5147), .A(n5259), .ZN(n6130) );
  INV_X1 U6302 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6656) );
  OAI22_X1 U6303 ( .A1(n6431), .A2(n6130), .B1(n6656), .B2(n6392), .ZN(n5149)
         );
  AOI21_X1 U6304 ( .B1(n6402), .B2(INSTADDRPOINTER_REG_8__SCAN_IN), .A(n5149), 
        .ZN(n5150) );
  OAI211_X1 U6305 ( .C1(n5255), .C2(n6394), .A(n5151), .B(n5150), .ZN(U3010)
         );
  INV_X1 U6306 ( .A(n6577), .ZN(n6538) );
  OAI21_X1 U6307 ( .B1(n5203), .B2(n6538), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5155) );
  NAND2_X1 U6308 ( .A1(n5155), .A2(n5154), .ZN(n5163) );
  INV_X1 U6309 ( .A(n5163), .ZN(n5159) );
  AND2_X1 U6310 ( .A1(n5156), .A2(n3171), .ZN(n6518) );
  NAND3_X1 U6311 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6590), .ZN(n6523) );
  NOR2_X1 U6312 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6523), .ZN(n5164)
         );
  OAI22_X1 U6313 ( .A1(n4969), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B1(n6683), .B2(n5164), .ZN(n5160) );
  INV_X1 U6314 ( .A(n5160), .ZN(n5161) );
  NAND2_X1 U6315 ( .A1(n5199), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5168)
         );
  INV_X1 U6316 ( .A(n5164), .ZN(n5200) );
  OAI22_X1 U6317 ( .A1(n5165), .A2(n5200), .B1(n6543), .B2(n6577), .ZN(n5166)
         );
  AOI21_X1 U6318 ( .B1(n5203), .B2(n6537), .A(n5166), .ZN(n5167) );
  OAI211_X1 U6319 ( .C1(n5207), .C2(n5169), .A(n5168), .B(n5167), .ZN(U3102)
         );
  NAND2_X1 U6320 ( .A1(n5199), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5173)
         );
  OAI22_X1 U6321 ( .A1(n5170), .A2(n5200), .B1(n6486), .B2(n6577), .ZN(n5171)
         );
  AOI21_X1 U6322 ( .B1(n5203), .B2(n6483), .A(n5171), .ZN(n5172) );
  OAI211_X1 U6323 ( .C1(n5207), .C2(n5174), .A(n5173), .B(n5172), .ZN(U3104)
         );
  NAND2_X1 U6324 ( .A1(n5199), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n5178)
         );
  OAI22_X1 U6325 ( .A1(n5175), .A2(n5200), .B1(n6490), .B2(n6577), .ZN(n5176)
         );
  AOI21_X1 U6326 ( .B1(n5203), .B2(n6487), .A(n5176), .ZN(n5177) );
  OAI211_X1 U6327 ( .C1(n5207), .C2(n5179), .A(n5178), .B(n5177), .ZN(U3105)
         );
  NAND2_X1 U6328 ( .A1(n5199), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5183)
         );
  OAI22_X1 U6329 ( .A1(n5180), .A2(n5200), .B1(n6502), .B2(n6577), .ZN(n5181)
         );
  AOI21_X1 U6330 ( .B1(n5203), .B2(n6498), .A(n5181), .ZN(n5182) );
  OAI211_X1 U6331 ( .C1(n5207), .C2(n5184), .A(n5183), .B(n5182), .ZN(U3107)
         );
  NAND2_X1 U6332 ( .A1(n5199), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5188)
         );
  OAI22_X1 U6333 ( .A1(n5185), .A2(n5200), .B1(n6476), .B2(n6577), .ZN(n5186)
         );
  AOI21_X1 U6334 ( .B1(n5203), .B2(n6473), .A(n5186), .ZN(n5187) );
  OAI211_X1 U6335 ( .C1(n5207), .C2(n5189), .A(n5188), .B(n5187), .ZN(U3101)
         );
  NAND2_X1 U6336 ( .A1(n5199), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5193)
         );
  OAI22_X1 U6337 ( .A1(n5190), .A2(n5200), .B1(n6494), .B2(n6577), .ZN(n5191)
         );
  AOI21_X1 U6338 ( .B1(n5203), .B2(n6491), .A(n5191), .ZN(n5192) );
  OAI211_X1 U6339 ( .C1(n5207), .C2(n5194), .A(n5193), .B(n5192), .ZN(U3106)
         );
  NAND2_X1 U6340 ( .A1(n5199), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n5198)
         );
  OAI22_X1 U6341 ( .A1(n5195), .A2(n5200), .B1(n6472), .B2(n6577), .ZN(n5196)
         );
  AOI21_X1 U6342 ( .B1(n5203), .B2(n6469), .A(n5196), .ZN(n5197) );
  OAI211_X1 U6343 ( .C1(n5207), .C2(n5932), .A(n5198), .B(n5197), .ZN(U3100)
         );
  NAND2_X1 U6344 ( .A1(n5199), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5205)
         );
  OAI22_X1 U6345 ( .A1(n5201), .A2(n5200), .B1(n6482), .B2(n6577), .ZN(n5202)
         );
  AOI21_X1 U6346 ( .B1(n5203), .B2(n6479), .A(n5202), .ZN(n5204) );
  OAI211_X1 U6347 ( .C1(n5207), .C2(n5206), .A(n5205), .B(n5204), .ZN(U3103)
         );
  OAI21_X1 U6348 ( .B1(n5092), .B2(n5210), .A(n5209), .ZN(n5249) );
  INV_X1 U6349 ( .A(DATAI_8_), .ZN(n7050) );
  INV_X1 U6350 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6324) );
  OAI222_X1 U6351 ( .A1(n5249), .A2(n5983), .B1(n5360), .B2(n7050), .C1(n5449), 
        .C2(n6324), .ZN(U2883) );
  INV_X1 U6352 ( .A(n6406), .ZN(n5219) );
  XOR2_X1 U6353 ( .A(n5211), .B(n5212), .Z(n6362) );
  NAND2_X1 U6354 ( .A1(n6362), .A2(n6439), .ZN(n5218) );
  INV_X1 U6355 ( .A(n5213), .ZN(n5214) );
  XNOR2_X1 U6356 ( .A(n5215), .B(n5214), .ZN(n6145) );
  INV_X1 U6357 ( .A(n6145), .ZN(n5221) );
  NAND2_X1 U6358 ( .A1(n6427), .A2(REIP_REG_7__SCAN_IN), .ZN(n6363) );
  OAI21_X1 U6359 ( .B1(n6431), .B2(n5221), .A(n6363), .ZN(n5216) );
  AOI21_X1 U6360 ( .B1(n6402), .B2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n5216), 
        .ZN(n5217) );
  OAI211_X1 U6361 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n5219), .A(n5218), 
        .B(n5217), .ZN(U3011) );
  INV_X1 U6362 ( .A(n6360), .ZN(n6149) );
  INV_X1 U6363 ( .A(EBX_REG_7__SCAN_IN), .ZN(n5220) );
  OAI22_X1 U6364 ( .A1(n6233), .A2(n5221), .B1(n6238), .B2(n5220), .ZN(n5222)
         );
  AOI21_X1 U6365 ( .B1(n6149), .B2(n4383), .A(n5222), .ZN(n5223) );
  INV_X1 U6366 ( .A(n5223), .ZN(U2852) );
  NOR3_X1 U6367 ( .A1(n6613), .A2(n6683), .A3(n6615), .ZN(n6611) );
  NOR3_X1 U6368 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n6626), .A3(n5454), .ZN(
        n6622) );
  OR2_X1 U6369 ( .A1(n5227), .A2(n5240), .ZN(n5228) );
  NAND2_X1 U6370 ( .A1(n6162), .A2(n5228), .ZN(n6221) );
  INV_X1 U6371 ( .A(n6221), .ZN(n5248) );
  NOR2_X1 U6372 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5239) );
  NAND2_X1 U6373 ( .A1(n6215), .A2(n6190), .ZN(n6062) );
  OR2_X1 U6374 ( .A1(n5232), .A2(n5240), .ZN(n6213) );
  NOR2_X1 U6375 ( .A1(n5233), .A2(n6213), .ZN(n5243) );
  NAND2_X1 U6376 ( .A1(n5234), .A2(n5239), .ZN(n6610) );
  NAND2_X1 U6377 ( .A1(n6271), .A2(n6610), .ZN(n5237) );
  NOR2_X1 U6378 ( .A1(EBX_REG_31__SCAN_IN), .A2(n5239), .ZN(n5235) );
  NAND2_X1 U6379 ( .A1(n3436), .A2(n5235), .ZN(n5236) );
  NAND2_X1 U6380 ( .A1(n5237), .A2(n5236), .ZN(n5238) );
  NOR2_X1 U6381 ( .A1(n5240), .A2(n5239), .ZN(n5241) );
  NAND2_X1 U6382 ( .A1(EBX_REG_31__SCAN_IN), .A2(n5241), .ZN(n6206) );
  OAI22_X1 U6383 ( .A1(n6224), .A2(n4144), .B1(n6202), .B2(n6441), .ZN(n5242)
         );
  AOI211_X1 U6384 ( .C1(n6062), .C2(REIP_REG_0__SCAN_IN), .A(n5243), .B(n5242), 
        .ZN(n5247) );
  OAI21_X1 U6385 ( .B1(n6212), .B2(n6211), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5246) );
  OAI211_X1 U6386 ( .C1(n5764), .C2(n5248), .A(n5247), .B(n5246), .ZN(U2827)
         );
  INV_X1 U6387 ( .A(n5249), .ZN(n6139) );
  INV_X1 U6388 ( .A(EBX_REG_8__SCAN_IN), .ZN(n6135) );
  OAI22_X1 U6389 ( .A1(n6233), .A2(n6130), .B1(n6238), .B2(n6135), .ZN(n5250)
         );
  AOI21_X1 U6390 ( .B1(n6139), .B2(n4383), .A(n5250), .ZN(n5251) );
  INV_X1 U6391 ( .A(n5251), .ZN(U2851) );
  AOI22_X1 U6392 ( .A1(n6383), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n6427), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n5252) );
  OAI21_X1 U6393 ( .B1(n6137), .B2(n6391), .A(n5252), .ZN(n5253) );
  AOI21_X1 U6394 ( .B1(n6139), .B2(n6379), .A(n5253), .ZN(n5254) );
  OAI21_X1 U6395 ( .B1(n5255), .B2(n6357), .A(n5254), .ZN(U2978) );
  NAND2_X1 U6396 ( .A1(n5209), .A2(n5257), .ZN(n5258) );
  AND2_X1 U6397 ( .A1(n5256), .A2(n5258), .ZN(n6125) );
  INV_X1 U6398 ( .A(n6125), .ZN(n5262) );
  AOI21_X1 U6399 ( .B1(n5260), .B2(n5259), .A(n5271), .ZN(n6416) );
  AOI22_X1 U6400 ( .A1(n5980), .A2(n6416), .B1(EBX_REG_9__SCAN_IN), .B2(n5605), 
        .ZN(n5261) );
  OAI21_X1 U6401 ( .B1(n5262), .B2(n6226), .A(n5261), .ZN(U2850) );
  INV_X1 U6402 ( .A(DATAI_9_), .ZN(n7017) );
  INV_X1 U6403 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6327) );
  OAI222_X1 U6404 ( .A1(n5262), .A2(n5983), .B1(n5360), .B2(n7017), .C1(n5449), 
        .C2(n6327), .ZN(U2882) );
  XNOR2_X1 U6405 ( .A(n5733), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5264)
         );
  XNOR2_X1 U6406 ( .A(n5263), .B(n5264), .ZN(n6415) );
  AOI22_X1 U6407 ( .A1(n6383), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .B1(n6427), 
        .B2(REIP_REG_9__SCAN_IN), .ZN(n5265) );
  OAI21_X1 U6408 ( .B1(n6391), .B2(n5266), .A(n5265), .ZN(n5267) );
  AOI21_X1 U6409 ( .B1(n6125), .B2(n6379), .A(n5267), .ZN(n5268) );
  OAI21_X1 U6410 ( .B1(n6415), .B2(n6357), .A(n5268), .ZN(U2977) );
  OR2_X1 U6411 ( .A1(n5256), .A2(n5270), .ZN(n5303) );
  INV_X1 U6412 ( .A(n5303), .ZN(n5269) );
  AOI21_X1 U6413 ( .B1(n5270), .B2(n5256), .A(n5269), .ZN(n5288) );
  INV_X1 U6414 ( .A(n5288), .ZN(n5291) );
  INV_X1 U6415 ( .A(n5286), .ZN(n5278) );
  OAI21_X1 U6416 ( .B1(n5272), .B2(n5271), .A(n6111), .ZN(n6410) );
  AOI22_X1 U6417 ( .A1(EBX_REG_10__SCAN_IN), .A2(n6156), .B1(
        PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n6212), .ZN(n5274) );
  NAND2_X1 U6418 ( .A1(n5273), .A2(n6215), .ZN(n6181) );
  OAI211_X1 U6419 ( .C1(n6202), .C2(n6410), .A(n5274), .B(n6181), .ZN(n5277)
         );
  INV_X1 U6420 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6659) );
  INV_X1 U6421 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6654) );
  INV_X1 U6422 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6651) );
  INV_X1 U6423 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6684) );
  INV_X1 U6424 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6648) );
  INV_X1 U6425 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6647) );
  NOR3_X1 U6426 ( .A1(n6684), .A2(n6648), .A3(n6647), .ZN(n6179) );
  NAND2_X1 U6427 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6179), .ZN(n6166) );
  NOR2_X1 U6428 ( .A1(n6651), .A2(n6166), .ZN(n6151) );
  NAND2_X1 U6429 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6151), .ZN(n6143) );
  NOR2_X1 U6430 ( .A1(n6654), .A2(n6143), .ZN(n6133) );
  NAND2_X1 U6431 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6133), .ZN(n5275) );
  NAND2_X1 U6432 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6123), .ZN(n5411) );
  INV_X1 U6433 ( .A(n6215), .ZN(n6191) );
  NOR2_X1 U6434 ( .A1(n6191), .A2(n5275), .ZN(n6121) );
  NAND3_X1 U6435 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .A3(
        n6121), .ZN(n5403) );
  NAND2_X1 U6436 ( .A1(n6062), .A2(n5403), .ZN(n6114) );
  AOI21_X1 U6437 ( .B1(n6659), .B2(n5411), .A(n6114), .ZN(n5276) );
  AOI211_X1 U6438 ( .C1(n6211), .C2(n5278), .A(n5277), .B(n5276), .ZN(n5279)
         );
  OAI21_X1 U6439 ( .B1(n5291), .B2(n6162), .A(n5279), .ZN(U2817) );
  INV_X1 U6440 ( .A(n5281), .ZN(n5283) );
  NAND2_X1 U6441 ( .A1(n5283), .A2(n5282), .ZN(n5284) );
  XNOR2_X1 U6442 ( .A(n5280), .B(n5284), .ZN(n6405) );
  AOI22_X1 U6443 ( .A1(n6383), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6427), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5285) );
  OAI21_X1 U6444 ( .B1(n5286), .B2(n6391), .A(n5285), .ZN(n5287) );
  AOI21_X1 U6445 ( .B1(n5288), .B2(n6379), .A(n5287), .ZN(n5289) );
  OAI21_X1 U6446 ( .B1(n6357), .B2(n6405), .A(n5289), .ZN(U2976) );
  INV_X1 U6447 ( .A(DATAI_10_), .ZN(n7039) );
  INV_X1 U6448 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6330) );
  OAI222_X1 U6449 ( .A1(n5291), .A2(n5983), .B1(n5360), .B2(n7039), .C1(n5449), 
        .C2(n6330), .ZN(U2881) );
  INV_X1 U6450 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5290) );
  OAI222_X1 U6451 ( .A1(n5291), .A2(n6226), .B1(n6230), .B2(n5290), .C1(n6410), 
        .C2(n6233), .ZN(U2849) );
  NAND2_X1 U6452 ( .A1(n5292), .A2(n6221), .ZN(n5301) );
  OAI21_X1 U6453 ( .B1(n6179), .B2(n6190), .A(n6215), .ZN(n6176) );
  AOI22_X1 U6454 ( .A1(n6231), .A2(n6178), .B1(n6156), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n5295) );
  INV_X1 U6455 ( .A(n6190), .ZN(n6192) );
  INV_X1 U6456 ( .A(n6179), .ZN(n5293) );
  NAND4_X1 U6457 ( .A1(n6192), .A2(REIP_REG_2__SCAN_IN), .A3(n5293), .A4(
        REIP_REG_1__SCAN_IN), .ZN(n5294) );
  NAND2_X1 U6458 ( .A1(n5295), .A2(n5294), .ZN(n5299) );
  OAI22_X1 U6459 ( .A1(n5297), .A2(n6198), .B1(n6205), .B2(n5296), .ZN(n5298)
         );
  AOI211_X1 U6460 ( .C1(REIP_REG_3__SCAN_IN), .C2(n6176), .A(n5299), .B(n5298), 
        .ZN(n5300) );
  OAI211_X1 U6461 ( .C1(n6458), .C2(n6213), .A(n5301), .B(n5300), .ZN(U2824)
         );
  AND2_X1 U6462 ( .A1(n5303), .A2(n5302), .ZN(n5304) );
  OR2_X1 U6463 ( .A1(n5304), .A2(n5307), .ZN(n6353) );
  INV_X1 U6464 ( .A(DATAI_11_), .ZN(n5305) );
  INV_X1 U6465 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6333) );
  OAI222_X1 U6466 ( .A1(n6353), .A2(n5983), .B1(n5360), .B2(n5305), .C1(n5449), 
        .C2(n6333), .ZN(U2880) );
  XOR2_X1 U6467 ( .A(n5307), .B(n5306), .Z(n6106) );
  INV_X1 U6468 ( .A(n6106), .ZN(n5325) );
  INV_X1 U6469 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6336) );
  INV_X1 U6470 ( .A(DATAI_12_), .ZN(n6854) );
  OAI222_X1 U6471 ( .A1(n5983), .A2(n5325), .B1(n5449), .B2(n6336), .C1(n6854), 
        .C2(n5360), .ZN(U2879) );
  NOR2_X1 U6472 ( .A1(n5309), .A2(n3192), .ZN(n5310) );
  XNOR2_X1 U6473 ( .A(n5308), .B(n5310), .ZN(n5324) );
  NAND2_X1 U6474 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5333) );
  INV_X1 U6475 ( .A(n5333), .ZN(n5336) );
  INV_X1 U6476 ( .A(n6404), .ZN(n6407) );
  NAND3_X1 U6477 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n6407), .ZN(n5313) );
  NOR2_X1 U6478 ( .A1(n5311), .A2(n5313), .ZN(n5375) );
  NAND2_X1 U6479 ( .A1(n5375), .A2(n6424), .ZN(n5859) );
  AOI21_X1 U6480 ( .B1(n5313), .B2(n6403), .A(n6402), .ZN(n6401) );
  OAI221_X1 U6481 ( .B1(n5336), .B2(n5853), .C1(n5336), .C2(n5859), .A(n6401), 
        .ZN(n5317) );
  NOR2_X1 U6482 ( .A1(n5313), .A2(n5312), .ZN(n5376) );
  NAND2_X1 U6483 ( .A1(n6425), .A2(n5376), .ZN(n5363) );
  NAND2_X1 U6484 ( .A1(n5859), .A2(n5363), .ZN(n6398) );
  INV_X1 U6485 ( .A(n6398), .ZN(n6018) );
  OAI21_X1 U6486 ( .B1(n6018), .B2(n6400), .A(n4324), .ZN(n5316) );
  OAI21_X1 U6487 ( .B1(n5314), .B2(n6110), .A(n5337), .ZN(n6103) );
  NAND2_X1 U6488 ( .A1(n6427), .A2(REIP_REG_12__SCAN_IN), .ZN(n5320) );
  OAI21_X1 U6489 ( .B1(n6431), .B2(n6103), .A(n5320), .ZN(n5315) );
  AOI21_X1 U6490 ( .B1(n5317), .B2(n5316), .A(n5315), .ZN(n5318) );
  OAI21_X1 U6491 ( .B1(n5324), .B2(n6394), .A(n5318), .ZN(U3006) );
  INV_X1 U6492 ( .A(n6105), .ZN(n5321) );
  NAND2_X1 U6493 ( .A1(n6383), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5319)
         );
  OAI211_X1 U6494 ( .C1(n6391), .C2(n5321), .A(n5320), .B(n5319), .ZN(n5322)
         );
  AOI21_X1 U6495 ( .B1(n6106), .B2(n6379), .A(n5322), .ZN(n5323) );
  OAI21_X1 U6496 ( .B1(n5324), .B2(n6357), .A(n5323), .ZN(U2974) );
  OAI222_X1 U6497 ( .A1(n6233), .A2(n6103), .B1(n6230), .B2(n4180), .C1(n6226), 
        .C2(n5325), .ZN(U2847) );
  OAI21_X1 U6498 ( .B1(n5326), .B2(n5328), .A(n5327), .ZN(n5997) );
  INV_X1 U6499 ( .A(DATAI_13_), .ZN(n6851) );
  INV_X1 U6500 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6339) );
  OAI222_X1 U6501 ( .A1(n5997), .A2(n5983), .B1(n5360), .B2(n6851), .C1(n5449), 
        .C2(n6339), .ZN(U2878) );
  OAI21_X1 U6502 ( .B1(n5331), .B2(n5330), .A(n5329), .ZN(n5999) );
  INV_X1 U6503 ( .A(n5999), .ZN(n5344) );
  NOR2_X1 U6504 ( .A1(n5335), .A2(n5333), .ZN(n5374) );
  NAND2_X1 U6505 ( .A1(n5333), .A2(n5332), .ZN(n5334) );
  OAI211_X1 U6506 ( .C1(n5374), .C2(n6450), .A(n6401), .B(n5334), .ZN(n5366)
         );
  NAND2_X1 U6507 ( .A1(n5336), .A2(n5335), .ZN(n5341) );
  XNOR2_X1 U6508 ( .A(n5338), .B(n5337), .ZN(n6091) );
  INV_X1 U6509 ( .A(n6091), .ZN(n5339) );
  NAND2_X1 U6510 ( .A1(n6445), .A2(n5339), .ZN(n5340) );
  NAND2_X1 U6511 ( .A1(n6427), .A2(REIP_REG_13__SCAN_IN), .ZN(n6000) );
  OAI211_X1 U6512 ( .C1(n6018), .C2(n5341), .A(n5340), .B(n6000), .ZN(n5342)
         );
  AOI21_X1 U6513 ( .B1(n5366), .B2(INSTADDRPOINTER_REG_13__SCAN_IN), .A(n5342), 
        .ZN(n5343) );
  OAI21_X1 U6514 ( .B1(n5344), .B2(n6394), .A(n5343), .ZN(U3005) );
  INV_X1 U6515 ( .A(n5997), .ZN(n6097) );
  INV_X1 U6516 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6092) );
  OAI22_X1 U6517 ( .A1(n6233), .A2(n6091), .B1(n6238), .B2(n6092), .ZN(n5345)
         );
  AOI21_X1 U6518 ( .B1(n6097), .B2(n4383), .A(n5345), .ZN(n5346) );
  INV_X1 U6519 ( .A(n5346), .ZN(U2846) );
  OR2_X1 U6520 ( .A1(n5348), .A2(n5347), .ZN(n5350) );
  NAND2_X1 U6521 ( .A1(n5350), .A2(n5349), .ZN(n6083) );
  INV_X1 U6522 ( .A(DATAI_14_), .ZN(n6953) );
  INV_X1 U6523 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6342) );
  OAI222_X1 U6524 ( .A1(n6083), .A2(n5983), .B1(n5360), .B2(n6953), .C1(n5449), 
        .C2(n6342), .ZN(U2877) );
  OAI21_X1 U6525 ( .B1(n5352), .B2(n5351), .A(n5357), .ZN(n6080) );
  OAI222_X1 U6526 ( .A1(n6083), .A2(n6226), .B1(n5353), .B2(n6230), .C1(n6080), 
        .C2(n6233), .ZN(U2845) );
  NAND2_X1 U6527 ( .A1(n5349), .A2(n5355), .ZN(n5356) );
  NAND2_X1 U6528 ( .A1(n5354), .A2(n5356), .ZN(n6072) );
  AOI21_X1 U6529 ( .B1(n5358), .B2(n5357), .A(n5629), .ZN(n6070) );
  AOI22_X1 U6530 ( .A1(n5980), .A2(n6070), .B1(EBX_REG_15__SCAN_IN), .B2(n5605), .ZN(n5359) );
  OAI21_X1 U6531 ( .B1(n6072), .B2(n6226), .A(n5359), .ZN(U2844) );
  INV_X1 U6532 ( .A(DATAI_15_), .ZN(n6949) );
  INV_X1 U6533 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6347) );
  OAI222_X1 U6534 ( .A1(n6072), .A2(n5983), .B1(n6949), .B2(n5360), .C1(n5449), 
        .C2(n6347), .ZN(U2876) );
  XNOR2_X1 U6535 ( .A(n5733), .B(n5367), .ZN(n5362) );
  XNOR2_X1 U6536 ( .A(n5361), .B(n5362), .ZN(n5763) );
  AOI21_X1 U6537 ( .B1(n5364), .B2(n5363), .A(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5365) );
  OAI21_X1 U6538 ( .B1(n5366), .B2(n5365), .A(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n5371) );
  NAND3_X1 U6539 ( .A1(n5374), .A2(n5367), .A3(n6398), .ZN(n5370) );
  INV_X1 U6540 ( .A(n6080), .ZN(n5368) );
  AOI22_X1 U6541 ( .A1(n6445), .A2(n5368), .B1(n6427), .B2(
        REIP_REG_14__SCAN_IN), .ZN(n5369) );
  AND3_X1 U6542 ( .A1(n5371), .A2(n5370), .A3(n5369), .ZN(n5372) );
  OAI21_X1 U6543 ( .B1(n5763), .B2(n6394), .A(n5372), .ZN(U3004) );
  INV_X1 U6544 ( .A(n5532), .ZN(n5373) );
  XNOR2_X1 U6545 ( .A(n5593), .B(n5373), .ZN(n5541) );
  NAND2_X1 U6546 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5374), .ZN(n5862) );
  NAND2_X1 U6547 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5894) );
  NOR2_X1 U6548 ( .A1(n5862), .A2(n5894), .ZN(n5851) );
  NAND2_X1 U6549 ( .A1(n5375), .A2(n5851), .ZN(n5857) );
  NAND4_X1 U6550 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A3(INSTADDRPOINTER_REG_19__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5377) );
  NOR2_X1 U6551 ( .A1(n5857), .A2(n5377), .ZN(n5378) );
  NAND2_X1 U6552 ( .A1(n5851), .A2(n5376), .ZN(n5852) );
  NOR2_X1 U6553 ( .A1(n5377), .A2(n5852), .ZN(n5382) );
  AOI22_X1 U6554 ( .A1(n5378), .A2(n6424), .B1(n6425), .B2(n5382), .ZN(n5835)
         );
  INV_X1 U6555 ( .A(n5835), .ZN(n5843) );
  NAND3_X1 U6556 ( .A1(n5836), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n5843), .ZN(n5389) );
  INV_X1 U6557 ( .A(n5378), .ZN(n5379) );
  NAND2_X1 U6558 ( .A1(n5858), .A2(n5379), .ZN(n5380) );
  OAI211_X1 U6559 ( .C1(n5382), .C2(n5853), .A(n5381), .B(n5380), .ZN(n5848)
         );
  INV_X1 U6560 ( .A(n5836), .ZN(n5383) );
  AND2_X1 U6561 ( .A1(n6403), .A2(n5383), .ZN(n5384) );
  NOR2_X1 U6562 ( .A1(n5848), .A2(n5384), .ZN(n5824) );
  NAND2_X1 U6563 ( .A1(n5385), .A2(n5853), .ZN(n5387) );
  INV_X1 U6564 ( .A(n5435), .ZN(n5386) );
  NAND2_X1 U6565 ( .A1(n5387), .A2(n5386), .ZN(n5388) );
  AOI21_X1 U6566 ( .B1(n5390), .B2(n5389), .A(n6002), .ZN(n5391) );
  AOI211_X1 U6567 ( .C1(n6445), .C2(n5541), .A(n5392), .B(n5391), .ZN(n5393)
         );
  OAI21_X1 U6568 ( .B1(n5394), .B2(n6394), .A(n5393), .ZN(U2994) );
  INV_X1 U6569 ( .A(n5395), .ZN(n5400) );
  AOI22_X1 U6570 ( .A1(n5397), .A2(n6027), .B1(n5396), .B2(n5927), .ZN(n5399)
         );
  INV_X1 U6571 ( .A(n4545), .ZN(n5917) );
  AOI21_X1 U6572 ( .B1(n5927), .B2(n5917), .A(n5460), .ZN(n5459) );
  OAI222_X1 U6573 ( .A1(n6614), .A2(n5400), .B1(n5460), .B2(n5399), .C1(n5398), 
        .C2(n5459), .ZN(U3456) );
  AOI22_X1 U6574 ( .A1(n6242), .A2(DATAI_30_), .B1(n6245), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5402) );
  NAND2_X1 U6575 ( .A1(n6246), .A2(DATAI_14_), .ZN(n5401) );
  OAI211_X1 U6576 ( .C1(n4356), .C2(n5983), .A(n5402), .B(n5401), .ZN(U2861)
         );
  INV_X1 U6577 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6660) );
  NOR2_X1 U6578 ( .A1(n6660), .A2(n5403), .ZN(n6090) );
  NAND4_X1 U6579 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6090), .A3(
        REIP_REG_13__SCAN_IN), .A4(REIP_REG_12__SCAN_IN), .ZN(n6061) );
  NAND3_X1 U6580 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .ZN(n5412) );
  NOR2_X1 U6581 ( .A1(n6061), .A2(n5412), .ZN(n5570) );
  INV_X1 U6582 ( .A(REIP_REG_20__SCAN_IN), .ZN(n7018) );
  NAND2_X1 U6583 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5976) );
  NOR2_X1 U6584 ( .A1(n7018), .A2(n5976), .ZN(n5404) );
  NAND2_X1 U6585 ( .A1(n5570), .A2(n5404), .ZN(n5405) );
  NAND3_X1 U6586 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n5413) );
  AND2_X1 U6587 ( .A1(n6062), .A2(n5413), .ZN(n5406) );
  AND2_X1 U6588 ( .A1(REIP_REG_26__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n5414) );
  NAND2_X1 U6589 ( .A1(n5414), .A2(REIP_REG_24__SCAN_IN), .ZN(n5407) );
  AND2_X1 U6590 ( .A1(n6062), .A2(n5407), .ZN(n5408) );
  NOR2_X1 U6591 ( .A1(n5529), .A2(n5408), .ZN(n5523) );
  NAND2_X1 U6592 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n5409) );
  NAND2_X1 U6593 ( .A1(n6192), .A2(n5409), .ZN(n5410) );
  NAND2_X1 U6594 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .ZN(
        n6095) );
  NAND2_X1 U6595 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6113), .ZN(n6109) );
  NAND4_X1 U6596 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .A4(n6056), .ZN(n5955) );
  NOR2_X1 U6597 ( .A1(n5955), .A2(n5413), .ZN(n5530) );
  NAND2_X1 U6598 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5530), .ZN(n5535) );
  INV_X1 U6599 ( .A(n5414), .ZN(n5415) );
  NOR2_X1 U6600 ( .A1(n5535), .A2(n5415), .ZN(n5505) );
  AND2_X1 U6601 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n5416) );
  NAND2_X1 U6602 ( .A1(n5505), .A2(n5416), .ZN(n5470) );
  OR2_X1 U6603 ( .A1(n5470), .A2(REIP_REG_29__SCAN_IN), .ZN(n5477) );
  AND2_X1 U6604 ( .A1(n5488), .A2(n5477), .ZN(n5463) );
  INV_X1 U6605 ( .A(n5463), .ZN(n5424) );
  NOR2_X1 U6606 ( .A1(n5790), .A2(n6202), .ZN(n5423) );
  INV_X1 U6607 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6946) );
  NOR3_X1 U6608 ( .A1(n5470), .A2(REIP_REG_30__SCAN_IN), .A3(n6946), .ZN(n5419) );
  NOR2_X1 U6609 ( .A1(n6224), .A2(n5417), .ZN(n5418) );
  AOI211_X1 U6610 ( .C1(n6212), .C2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5419), 
        .B(n5418), .ZN(n5420) );
  OAI21_X1 U6611 ( .B1(n5421), .B2(n6205), .A(n5420), .ZN(n5422) );
  OAI21_X1 U6612 ( .B1(n4356), .B2(n6162), .A(n5425), .ZN(U2797) );
  INV_X1 U6613 ( .A(n5429), .ZN(n5431) );
  INV_X1 U6614 ( .A(n5426), .ZN(n5430) );
  INV_X1 U6615 ( .A(n5427), .ZN(n5428) );
  INV_X1 U6616 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5438) );
  INV_X1 U6617 ( .A(n5432), .ZN(n5448) );
  AND2_X1 U6618 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5436) );
  INV_X1 U6619 ( .A(n5436), .ZN(n5816) );
  NAND2_X1 U6620 ( .A1(n6403), .A2(n5816), .ZN(n5433) );
  NAND2_X1 U6621 ( .A1(n6002), .A2(n5433), .ZN(n5810) );
  AND2_X1 U6622 ( .A1(n6403), .A2(n5437), .ZN(n5434) );
  NOR2_X1 U6623 ( .A1(n5810), .A2(n5434), .ZN(n5774) );
  INV_X1 U6624 ( .A(n5774), .ZN(n5441) );
  NAND2_X1 U6625 ( .A1(n6427), .A2(REIP_REG_29__SCAN_IN), .ZN(n5443) );
  NAND2_X1 U6626 ( .A1(n5826), .A2(n5435), .ZN(n6009) );
  INV_X1 U6627 ( .A(n6009), .ZN(n5817) );
  NAND2_X1 U6628 ( .A1(n5817), .A2(n5436), .ZN(n5807) );
  NOR2_X1 U6629 ( .A1(n5807), .A2(n5437), .ZN(n5787) );
  NAND2_X1 U6630 ( .A1(n5787), .A2(n5438), .ZN(n5439) );
  OAI211_X1 U6631 ( .C1(n5480), .C2(n6431), .A(n5443), .B(n5439), .ZN(n5440)
         );
  AOI21_X1 U6632 ( .B1(n5441), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5440), 
        .ZN(n5442) );
  OAI21_X1 U6633 ( .B1(n5448), .B2(n6394), .A(n5442), .ZN(U2989) );
  NAND2_X1 U6634 ( .A1(n6366), .A2(n5483), .ZN(n5444) );
  OAI211_X1 U6635 ( .C1(n5445), .C2(n6372), .A(n5444), .B(n5443), .ZN(n5446)
         );
  AOI21_X1 U6636 ( .B1(n5634), .B2(n6379), .A(n5446), .ZN(n5447) );
  OAI21_X1 U6637 ( .B1(n5448), .B2(n6357), .A(n5447), .ZN(U2957) );
  NAND3_X1 U6638 ( .A1(n5462), .A2(n5450), .A3(n5449), .ZN(n5452) );
  AOI22_X1 U6639 ( .A1(n6242), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6245), .ZN(n5451) );
  NAND2_X1 U6640 ( .A1(n5452), .A2(n5451), .ZN(U2860) );
  AOI22_X1 U6641 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5773), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n5453), .ZN(n5925) );
  INV_X1 U6642 ( .A(n5925), .ZN(n5457) );
  NOR2_X1 U6643 ( .A1(n5454), .A2(n6452), .ZN(n5924) );
  NOR2_X1 U6644 ( .A1(n6614), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5456)
         );
  AOI222_X1 U6645 ( .A1(n5457), .A2(n5924), .B1(n4545), .B2(n5456), .C1(n5455), 
        .C2(n6027), .ZN(n5461) );
  OAI22_X1 U6646 ( .A1(n5461), .A2(n5460), .B1(n5459), .B2(n3168), .ZN(U3459)
         );
  INV_X1 U6647 ( .A(n5462), .ZN(n5476) );
  OAI21_X1 U6648 ( .B1(REIP_REG_30__SCAN_IN), .B2(n6190), .A(n5463), .ZN(n5475) );
  OAI22_X1 U6649 ( .A1(n5464), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4159), .ZN(n5469) );
  NOR4_X1 U6650 ( .A1(n5470), .A2(REIP_REG_31__SCAN_IN), .A3(n6900), .A4(n6946), .ZN(n5473) );
  AND4_X1 U6651 ( .A1(n6271), .A2(EBX_REG_31__SCAN_IN), .A3(n6610), .A4(n5471), 
        .ZN(n5472) );
  AOI211_X1 U6652 ( .C1(n6212), .C2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5473), 
        .B(n5472), .ZN(n5474) );
  NAND2_X1 U6653 ( .A1(n5634), .A2(n6150), .ZN(n5485) );
  NAND2_X1 U6654 ( .A1(n6212), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5478)
         );
  OAI211_X1 U6655 ( .C1(n6224), .C2(n5479), .A(n5478), .B(n5477), .ZN(n5482)
         );
  NOR2_X1 U6656 ( .A1(n5480), .A2(n6202), .ZN(n5481) );
  AOI211_X1 U6657 ( .C1(n6211), .C2(n5483), .A(n5482), .B(n5481), .ZN(n5484)
         );
  OAI211_X1 U6658 ( .C1(n5488), .C2(n6946), .A(n5485), .B(n5484), .ZN(U2798)
         );
  INV_X1 U6659 ( .A(n5488), .ZN(n5497) );
  OR2_X1 U6660 ( .A1(n3186), .A2(n5489), .ZN(n5490) );
  NAND2_X1 U6661 ( .A1(n5491), .A2(n5490), .ZN(n5801) );
  INV_X1 U6662 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6673) );
  NOR2_X1 U6663 ( .A1(n6673), .A2(REIP_REG_28__SCAN_IN), .ZN(n5492) );
  AOI22_X1 U6664 ( .A1(n6156), .A2(EBX_REG_28__SCAN_IN), .B1(n5505), .B2(n5492), .ZN(n5493) );
  OAI21_X1 U6665 ( .B1(n5801), .B2(n6202), .A(n5493), .ZN(n5494) );
  AOI21_X1 U6666 ( .B1(PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6212), .A(n5494), 
        .ZN(n5495) );
  OAI21_X1 U6667 ( .B1(n5657), .B2(n6205), .A(n5495), .ZN(n5496) );
  AOI21_X1 U6668 ( .B1(n5497), .B2(REIP_REG_28__SCAN_IN), .A(n5496), .ZN(n5498) );
  OAI21_X1 U6669 ( .B1(n5667), .B2(n6162), .A(n5498), .ZN(U2799) );
  AOI21_X1 U6670 ( .B1(n5502), .B2(n5500), .A(n5501), .ZN(n5675) );
  INV_X1 U6671 ( .A(n5675), .ZN(n5642) );
  AND2_X1 U6672 ( .A1(n5517), .A2(n5503), .ZN(n5504) );
  OR2_X1 U6673 ( .A1(n3186), .A2(n5504), .ZN(n5805) );
  NAND2_X1 U6674 ( .A1(n6212), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5507)
         );
  AOI22_X1 U6675 ( .A1(n6156), .A2(EBX_REG_27__SCAN_IN), .B1(n5505), .B2(n6673), .ZN(n5506) );
  OAI211_X1 U6676 ( .C1(n6202), .C2(n5805), .A(n5507), .B(n5506), .ZN(n5509)
         );
  NOR2_X1 U6677 ( .A1(n5523), .A2(n6673), .ZN(n5508) );
  AOI211_X1 U6678 ( .C1(n6211), .C2(n5671), .A(n5509), .B(n5508), .ZN(n5510)
         );
  OAI21_X1 U6679 ( .B1(n5642), .B2(n6162), .A(n5510), .ZN(U2800) );
  OAI21_X1 U6680 ( .B1(n5511), .B2(n5512), .A(n5500), .ZN(n5683) );
  INV_X1 U6681 ( .A(n5535), .ZN(n5513) );
  AOI21_X1 U6682 ( .B1(n5513), .B2(REIP_REG_25__SCAN_IN), .A(
        REIP_REG_26__SCAN_IN), .ZN(n5522) );
  INV_X1 U6683 ( .A(n5677), .ZN(n5519) );
  OR2_X1 U6684 ( .A1(n5514), .A2(n5515), .ZN(n5516) );
  NAND2_X1 U6685 ( .A1(n5517), .A2(n5516), .ZN(n5814) );
  INV_X1 U6686 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5582) );
  OAI22_X1 U6687 ( .A1(n5814), .A2(n6202), .B1(n6224), .B2(n5582), .ZN(n5518)
         );
  AOI21_X1 U6688 ( .B1(n6211), .B2(n5519), .A(n5518), .ZN(n5521) );
  NAND2_X1 U6689 ( .A1(n6212), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5520)
         );
  OAI211_X1 U6690 ( .C1(n5523), .C2(n5522), .A(n5521), .B(n5520), .ZN(n5524)
         );
  INV_X1 U6691 ( .A(n5524), .ZN(n5525) );
  OAI21_X1 U6692 ( .B1(n5683), .B2(n6162), .A(n5525), .ZN(U2801) );
  AOI21_X1 U6693 ( .B1(n5527), .B2(n5526), .A(n5511), .ZN(n5528) );
  INV_X1 U6694 ( .A(n5528), .ZN(n5691) );
  INV_X1 U6695 ( .A(n5529), .ZN(n5945) );
  NAND2_X1 U6696 ( .A1(n6922), .A2(n5530), .ZN(n5542) );
  INV_X1 U6697 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6920) );
  AOI21_X1 U6698 ( .B1(n5945), .B2(n5542), .A(n6920), .ZN(n5539) );
  AOI21_X1 U6699 ( .B1(n5593), .B2(n5532), .A(n5531), .ZN(n5533) );
  OR2_X1 U6700 ( .A1(n5514), .A2(n5533), .ZN(n6004) );
  NOR2_X1 U6701 ( .A1(n6004), .A2(n6202), .ZN(n5538) );
  INV_X1 U6702 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5583) );
  OAI22_X1 U6703 ( .A1(n5583), .A2(n6224), .B1(n5684), .B2(n6198), .ZN(n5537)
         );
  OAI22_X1 U6704 ( .A1(REIP_REG_25__SCAN_IN), .A2(n5535), .B1(n5534), .B2(
        n6205), .ZN(n5536) );
  NOR4_X1 U6705 ( .A1(n5539), .A2(n5538), .A3(n5537), .A4(n5536), .ZN(n5540)
         );
  OAI21_X1 U6706 ( .B1(n5691), .B2(n6162), .A(n5540), .ZN(U2802) );
  NAND2_X1 U6707 ( .A1(n5586), .A2(n6150), .ZN(n5549) );
  INV_X1 U6708 ( .A(n5541), .ZN(n5588) );
  NAND2_X1 U6709 ( .A1(n6156), .A2(EBX_REG_24__SCAN_IN), .ZN(n5543) );
  OAI211_X1 U6710 ( .C1(n5588), .C2(n6202), .A(n5543), .B(n5542), .ZN(n5546)
         );
  NOR2_X1 U6711 ( .A1(n6198), .A2(n5544), .ZN(n5545) );
  AOI211_X1 U6712 ( .C1(n6211), .C2(n5547), .A(n5546), .B(n5545), .ZN(n5548)
         );
  OAI211_X1 U6713 ( .C1(n5945), .C2(n6922), .A(n5549), .B(n5548), .ZN(U2803)
         );
  NAND2_X1 U6714 ( .A1(n5551), .A2(n5552), .ZN(n5553) );
  INV_X1 U6715 ( .A(n5990), .ZN(n5607) );
  INV_X1 U6716 ( .A(n6056), .ZN(n5554) );
  OAI21_X1 U6717 ( .B1(n5976), .B2(n5554), .A(n7018), .ZN(n5564) );
  INV_X1 U6718 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5555) );
  OAI22_X1 U6719 ( .A1(n5555), .A2(n6198), .B1(n5720), .B2(n6205), .ZN(n5563)
         );
  MUX2_X1 U6720 ( .A(n5557), .B(n5611), .S(n5556), .Z(n5559) );
  XNOR2_X1 U6721 ( .A(n5559), .B(n5558), .ZN(n5868) );
  INV_X1 U6722 ( .A(n5868), .ZN(n5561) );
  INV_X1 U6723 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5560) );
  OAI22_X1 U6724 ( .A1(n5561), .A2(n6202), .B1(n5560), .B2(n6224), .ZN(n5562)
         );
  AOI211_X1 U6725 ( .C1(n5564), .C2(n5960), .A(n5563), .B(n5562), .ZN(n5565)
         );
  OAI21_X1 U6726 ( .B1(n5607), .B2(n6162), .A(n5565), .ZN(U2807) );
  INV_X1 U6727 ( .A(n5568), .ZN(n5569) );
  AOI21_X1 U6728 ( .B1(n3228), .B2(n3227), .A(n5569), .ZN(n5743) );
  INV_X1 U6729 ( .A(n5743), .ZN(n5656) );
  NAND2_X1 U6730 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n6060) );
  INV_X1 U6731 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6916) );
  OAI21_X1 U6732 ( .B1(n6060), .B2(n6078), .A(n6916), .ZN(n5577) );
  INV_X1 U6733 ( .A(n6062), .ZN(n6122) );
  NOR2_X1 U6734 ( .A1(n6122), .A2(n5570), .ZN(n6052) );
  AND2_X1 U6735 ( .A1(n5571), .A2(n5628), .ZN(n5572) );
  NOR2_X1 U6736 ( .A1(n5617), .A2(n5572), .ZN(n6013) );
  INV_X1 U6737 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5624) );
  OAI22_X1 U6738 ( .A1(n5624), .A2(n6224), .B1(n5573), .B2(n6198), .ZN(n5574)
         );
  AOI211_X1 U6739 ( .C1(n6013), .C2(n6178), .A(n6169), .B(n5574), .ZN(n5575)
         );
  OAI21_X1 U6740 ( .B1(n6205), .B2(n5741), .A(n5575), .ZN(n5576) );
  AOI21_X1 U6741 ( .B1(n5577), .B2(n6052), .A(n5576), .ZN(n5578) );
  OAI21_X1 U6742 ( .B1(n5656), .B2(n6162), .A(n5578), .ZN(U2810) );
  INV_X1 U6743 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5579) );
  OAI22_X1 U6744 ( .A1(n5772), .A2(n6233), .B1(n6238), .B2(n5579), .ZN(U2828)
         );
  INV_X1 U6745 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5580) );
  OAI222_X1 U6746 ( .A1(n6226), .A2(n5667), .B1(n5580), .B2(n6230), .C1(n5801), 
        .C2(n6233), .ZN(U2831) );
  OAI222_X1 U6747 ( .A1(n6226), .A2(n5642), .B1(n5581), .B2(n6230), .C1(n5805), 
        .C2(n6233), .ZN(U2832) );
  OAI222_X1 U6748 ( .A1(n6226), .A2(n5683), .B1(n5582), .B2(n6230), .C1(n5814), 
        .C2(n6233), .ZN(U2833) );
  OAI22_X1 U6749 ( .A1(n6233), .A2(n6004), .B1(n5583), .B2(n6238), .ZN(n5584)
         );
  INV_X1 U6750 ( .A(n5584), .ZN(n5585) );
  OAI21_X1 U6751 ( .B1(n5691), .B2(n6226), .A(n5585), .ZN(U2834) );
  INV_X1 U6752 ( .A(n5586), .ZN(n5649) );
  OAI222_X1 U6753 ( .A1(n6233), .A2(n5588), .B1(n6226), .B2(n5649), .C1(n5587), 
        .C2(n6238), .ZN(U2835) );
  AOI21_X1 U6754 ( .B1(n5590), .B2(n5589), .A(n4372), .ZN(n5699) );
  INV_X1 U6755 ( .A(n5699), .ZN(n5946) );
  INV_X1 U6756 ( .A(n5834), .ZN(n5592) );
  AOI21_X1 U6757 ( .B1(n5592), .B2(n5833), .A(n5591), .ZN(n5594) );
  OR2_X1 U6758 ( .A1(n5594), .A2(n5593), .ZN(n5943) );
  INV_X1 U6759 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5951) );
  OAI22_X1 U6760 ( .A1(n6233), .A2(n5943), .B1(n5951), .B2(n6238), .ZN(n5595)
         );
  INV_X1 U6761 ( .A(n5595), .ZN(n5596) );
  OAI21_X1 U6762 ( .B1(n5946), .B2(n6226), .A(n5596), .ZN(U2836) );
  AND2_X1 U6763 ( .A1(n5550), .A2(n5598), .ZN(n5599) );
  NOR2_X1 U6764 ( .A1(n5597), .A2(n5599), .ZN(n5987) );
  INV_X1 U6765 ( .A(n5987), .ZN(n5604) );
  NAND2_X1 U6766 ( .A1(n5601), .A2(n5600), .ZN(n5602) );
  NAND2_X1 U6767 ( .A1(n5834), .A2(n5602), .ZN(n5962) );
  OAI222_X1 U6768 ( .A1(n6226), .A2(n5604), .B1(n5603), .B2(n6230), .C1(n5962), 
        .C2(n6233), .ZN(U2838) );
  AOI22_X1 U6769 ( .A1(n5980), .A2(n5868), .B1(EBX_REG_20__SCAN_IN), .B2(n5605), .ZN(n5606) );
  OAI21_X1 U6770 ( .B1(n5607), .B2(n6226), .A(n5606), .ZN(U2839) );
  OR2_X1 U6771 ( .A1(n5608), .A2(n5609), .ZN(n5610) );
  NAND2_X1 U6772 ( .A1(n5551), .A2(n5610), .ZN(n5973) );
  INV_X1 U6773 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5616) );
  NAND2_X1 U6774 ( .A1(n5611), .A2(n4150), .ZN(n5614) );
  OR2_X1 U6775 ( .A1(n5612), .A2(n4150), .ZN(n5613) );
  NAND2_X1 U6776 ( .A1(n5614), .A2(n5613), .ZN(n5618) );
  NAND2_X1 U6777 ( .A1(n5618), .A2(n5617), .ZN(n5619) );
  XNOR2_X1 U6778 ( .A(n5619), .B(n5615), .ZN(n5877) );
  INV_X1 U6779 ( .A(n5877), .ZN(n5972) );
  OAI222_X1 U6780 ( .A1(n5973), .A2(n6226), .B1(n6230), .B2(n5616), .C1(n6233), 
        .C2(n5972), .ZN(U2840) );
  OR2_X1 U6781 ( .A1(n5618), .A2(n5617), .ZN(n5620) );
  NAND2_X1 U6782 ( .A1(n5620), .A2(n5619), .ZN(n6059) );
  NOR2_X1 U6783 ( .A1(n5569), .A2(n5621), .ZN(n5622) );
  OR2_X1 U6784 ( .A1(n5608), .A2(n5622), .ZN(n5993) );
  OAI222_X1 U6785 ( .A1(n6233), .A2(n6059), .B1(n5623), .B2(n6230), .C1(n5993), 
        .C2(n6226), .ZN(U2841) );
  INV_X1 U6786 ( .A(n6013), .ZN(n5625) );
  OAI22_X1 U6787 ( .A1(n6233), .A2(n5625), .B1(n5624), .B2(n6238), .ZN(n5626)
         );
  AOI21_X1 U6788 ( .B1(n5743), .B2(n4383), .A(n5626), .ZN(n5627) );
  INV_X1 U6789 ( .A(n5627), .ZN(U2842) );
  OAI21_X1 U6790 ( .B1(n5630), .B2(n5629), .A(n5628), .ZN(n6064) );
  AOI21_X1 U6791 ( .B1(n5631), .B2(n5354), .A(n5567), .ZN(n6244) );
  INV_X1 U6792 ( .A(n6244), .ZN(n5632) );
  OAI222_X1 U6793 ( .A1(n6064), .A2(n6233), .B1(n5633), .B2(n6230), .C1(n5632), 
        .C2(n6226), .ZN(U2843) );
  INV_X1 U6794 ( .A(n5634), .ZN(n5637) );
  AOI22_X1 U6795 ( .A1(n6242), .A2(DATAI_29_), .B1(n6245), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5636) );
  NAND2_X1 U6796 ( .A1(n6246), .A2(DATAI_13_), .ZN(n5635) );
  OAI211_X1 U6797 ( .C1(n5637), .C2(n5983), .A(n5636), .B(n5635), .ZN(U2862)
         );
  AOI22_X1 U6798 ( .A1(n6242), .A2(DATAI_28_), .B1(n6245), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5639) );
  NAND2_X1 U6799 ( .A1(n6246), .A2(DATAI_12_), .ZN(n5638) );
  OAI211_X1 U6800 ( .C1(n5667), .C2(n5983), .A(n5639), .B(n5638), .ZN(U2863)
         );
  AOI22_X1 U6801 ( .A1(n6242), .A2(DATAI_27_), .B1(n6245), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5641) );
  NAND2_X1 U6802 ( .A1(n6246), .A2(DATAI_11_), .ZN(n5640) );
  OAI211_X1 U6803 ( .C1(n5642), .C2(n5983), .A(n5641), .B(n5640), .ZN(U2864)
         );
  AOI22_X1 U6804 ( .A1(n6242), .A2(DATAI_26_), .B1(n6245), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5644) );
  NAND2_X1 U6805 ( .A1(n6246), .A2(DATAI_10_), .ZN(n5643) );
  OAI211_X1 U6806 ( .C1(n5683), .C2(n5983), .A(n5644), .B(n5643), .ZN(U2865)
         );
  AOI22_X1 U6807 ( .A1(n6242), .A2(DATAI_25_), .B1(n6245), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5646) );
  NAND2_X1 U6808 ( .A1(n6246), .A2(DATAI_9_), .ZN(n5645) );
  OAI211_X1 U6809 ( .C1(n5691), .C2(n5983), .A(n5646), .B(n5645), .ZN(U2866)
         );
  AOI22_X1 U6810 ( .A1(n6242), .A2(DATAI_24_), .B1(n6245), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5648) );
  NAND2_X1 U6811 ( .A1(n6246), .A2(DATAI_8_), .ZN(n5647) );
  OAI211_X1 U6812 ( .C1(n5649), .C2(n5983), .A(n5648), .B(n5647), .ZN(U2867)
         );
  AOI22_X1 U6813 ( .A1(n6246), .A2(DATAI_7_), .B1(n6245), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5651) );
  NAND2_X1 U6814 ( .A1(n6242), .A2(DATAI_23_), .ZN(n5650) );
  OAI211_X1 U6815 ( .C1(n5946), .C2(n5983), .A(n5651), .B(n5650), .ZN(U2868)
         );
  AOI22_X1 U6816 ( .A1(n6246), .A2(DATAI_3_), .B1(n6245), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5653) );
  NAND2_X1 U6817 ( .A1(n6242), .A2(DATAI_19_), .ZN(n5652) );
  OAI211_X1 U6818 ( .C1(n5973), .C2(n5983), .A(n5653), .B(n5652), .ZN(U2872)
         );
  AOI22_X1 U6819 ( .A1(n6242), .A2(DATAI_17_), .B1(n6245), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5655) );
  NAND2_X1 U6820 ( .A1(n6246), .A2(DATAI_1_), .ZN(n5654) );
  OAI211_X1 U6821 ( .C1(n5656), .C2(n5983), .A(n5655), .B(n5654), .ZN(U2874)
         );
  AND2_X1 U6822 ( .A1(n6427), .A2(REIP_REG_28__SCAN_IN), .ZN(n5797) );
  NOR2_X1 U6823 ( .A1(n6391), .A2(n5657), .ZN(n5658) );
  AOI211_X1 U6824 ( .C1(PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n6383), .A(n5797), 
        .B(n5658), .ZN(n5666) );
  INV_X1 U6825 ( .A(n5680), .ZN(n5659) );
  NAND3_X1 U6826 ( .A1(n5659), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5729), .ZN(n5663) );
  CLKBUF_X1 U6827 ( .A(n5660), .Z(n5688) );
  NAND2_X1 U6828 ( .A1(n5661), .A2(n5823), .ZN(n5815) );
  NOR2_X1 U6829 ( .A1(n5729), .A2(n5815), .ZN(n5662) );
  NAND2_X1 U6830 ( .A1(n5688), .A2(n5662), .ZN(n5668) );
  AOI22_X1 U6831 ( .A1(n5663), .A2(n5668), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5823), .ZN(n5664) );
  XNOR2_X1 U6832 ( .A(n5664), .B(n5796), .ZN(n5795) );
  NAND2_X1 U6833 ( .A1(n5795), .A2(n6387), .ZN(n5665) );
  OAI211_X1 U6834 ( .C1(n5667), .C2(n6359), .A(n5666), .B(n5665), .ZN(U2958)
         );
  NAND2_X1 U6835 ( .A1(n5669), .A2(n5668), .ZN(n5670) );
  XNOR2_X1 U6836 ( .A(n5670), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5812)
         );
  NAND2_X1 U6837 ( .A1(n6366), .A2(n5671), .ZN(n5672) );
  NAND2_X1 U6838 ( .A1(n6427), .A2(REIP_REG_27__SCAN_IN), .ZN(n5806) );
  OAI211_X1 U6839 ( .C1(n5673), .C2(n6372), .A(n5672), .B(n5806), .ZN(n5674)
         );
  AOI21_X1 U6840 ( .B1(n5675), .B2(n6379), .A(n5674), .ZN(n5676) );
  OAI21_X1 U6841 ( .B1(n5812), .B2(n6357), .A(n5676), .ZN(U2959) );
  INV_X1 U6842 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6947) );
  NOR2_X1 U6843 ( .A1(n6392), .A2(n6947), .ZN(n5819) );
  NOR2_X1 U6844 ( .A1(n6391), .A2(n5677), .ZN(n5678) );
  AOI211_X1 U6845 ( .C1(PHYADDRPOINTER_REG_26__SCAN_IN), .C2(n6383), .A(n5819), 
        .B(n5678), .ZN(n5682) );
  XNOR2_X1 U6846 ( .A(n5733), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5679)
         );
  XNOR2_X1 U6847 ( .A(n5680), .B(n5679), .ZN(n5813) );
  NAND2_X1 U6848 ( .A1(n5813), .A2(n6387), .ZN(n5681) );
  OAI211_X1 U6849 ( .C1(n5683), .C2(n6359), .A(n5682), .B(n5681), .ZN(U2960)
         );
  OAI22_X1 U6850 ( .A1(n6372), .A2(n5684), .B1(n6392), .B2(n6920), .ZN(n5685)
         );
  AOI21_X1 U6851 ( .B1(n6366), .B2(n5686), .A(n5685), .ZN(n5690) );
  OAI21_X1 U6852 ( .B1(n5688), .B2(n5687), .A(n4394), .ZN(n6006) );
  NAND2_X1 U6853 ( .A1(n6006), .A2(n6387), .ZN(n5689) );
  OAI211_X1 U6854 ( .C1(n5691), .C2(n6359), .A(n5690), .B(n5689), .ZN(U2961)
         );
  NAND2_X1 U6855 ( .A1(n5836), .A2(n5864), .ZN(n5694) );
  OAI21_X1 U6856 ( .B1(n5692), .B2(n5694), .A(n5693), .ZN(n5695) );
  XNOR2_X1 U6857 ( .A(n5695), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5832)
         );
  NAND2_X1 U6858 ( .A1(n6366), .A2(n5942), .ZN(n5696) );
  NAND2_X1 U6859 ( .A1(n6427), .A2(REIP_REG_23__SCAN_IN), .ZN(n5828) );
  OAI211_X1 U6860 ( .C1(n6372), .C2(n5697), .A(n5696), .B(n5828), .ZN(n5698)
         );
  AOI21_X1 U6861 ( .B1(n5699), .B2(n6379), .A(n5698), .ZN(n5700) );
  OAI21_X1 U6862 ( .B1(n5832), .B2(n6357), .A(n5700), .ZN(U2963) );
  AOI21_X1 U6863 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5733), .A(n5702), 
        .ZN(n5703) );
  XNOR2_X1 U6864 ( .A(n5701), .B(n5703), .ZN(n5842) );
  OAI21_X1 U6865 ( .B1(n5597), .B2(n5704), .A(n5589), .ZN(n5705) );
  NOR2_X1 U6866 ( .A1(n6392), .A2(n6913), .ZN(n5839) );
  AOI21_X1 U6867 ( .B1(n6383), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5839), 
        .ZN(n5706) );
  OAI21_X1 U6868 ( .B1(n5952), .B2(n6391), .A(n5706), .ZN(n5707) );
  AOI21_X1 U6869 ( .B1(n5984), .B2(n6379), .A(n5707), .ZN(n5708) );
  OAI21_X1 U6870 ( .B1(n5842), .B2(n6357), .A(n5708), .ZN(U2964) );
  AOI21_X1 U6871 ( .B1(n5711), .B2(n5710), .A(n5709), .ZN(n5850) );
  INV_X1 U6872 ( .A(n5961), .ZN(n5713) );
  NAND2_X1 U6873 ( .A1(n6383), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5712)
         );
  NAND2_X1 U6874 ( .A1(n6427), .A2(REIP_REG_21__SCAN_IN), .ZN(n5846) );
  OAI211_X1 U6875 ( .C1(n6391), .C2(n5713), .A(n5712), .B(n5846), .ZN(n5714)
         );
  AOI21_X1 U6876 ( .B1(n5987), .B2(n6379), .A(n5714), .ZN(n5715) );
  OAI21_X1 U6877 ( .B1(n5850), .B2(n6357), .A(n5715), .ZN(U2965) );
  NAND2_X1 U6878 ( .A1(n5717), .A2(n5716), .ZN(n5718) );
  NAND2_X1 U6879 ( .A1(n5692), .A2(n5718), .ZN(n5871) );
  AOI22_X1 U6880 ( .A1(n6383), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .B1(n6427), 
        .B2(REIP_REG_20__SCAN_IN), .ZN(n5719) );
  OAI21_X1 U6881 ( .B1(n5720), .B2(n6391), .A(n5719), .ZN(n5721) );
  AOI21_X1 U6882 ( .B1(n5990), .B2(n6379), .A(n5721), .ZN(n5722) );
  OAI21_X1 U6883 ( .B1(n5871), .B2(n6357), .A(n5722), .ZN(U2966) );
  OAI21_X1 U6884 ( .B1(n5724), .B2(n5874), .A(n5723), .ZN(n5725) );
  XNOR2_X1 U6885 ( .A(n5725), .B(n5733), .ZN(n5879) );
  OAI22_X1 U6886 ( .A1(n6372), .A2(n5971), .B1(n6392), .B2(n6667), .ZN(n5727)
         );
  NOR2_X1 U6887 ( .A1(n5973), .A2(n6359), .ZN(n5726) );
  AOI211_X1 U6888 ( .C1(n6366), .C2(n5969), .A(n5727), .B(n5726), .ZN(n5728)
         );
  OAI21_X1 U6889 ( .B1(n5879), .B2(n6357), .A(n5728), .ZN(U2967) );
  NAND2_X1 U6890 ( .A1(n5729), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5881) );
  INV_X1 U6891 ( .A(n5881), .ZN(n5739) );
  INV_X1 U6893 ( .A(n5732), .ZN(n5735) );
  NOR2_X1 U6894 ( .A1(n5733), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5736)
         );
  NAND3_X1 U6895 ( .A1(n5735), .A2(n5736), .A3(n5734), .ZN(n5880) );
  INV_X1 U6896 ( .A(n5880), .ZN(n5738) );
  AOI211_X1 U6897 ( .C1(n5731), .C2(n5745), .A(n5736), .B(n5739), .ZN(n5737)
         );
  AOI211_X1 U6898 ( .C1(n5739), .C2(n5731), .A(n5738), .B(n5737), .ZN(n6012)
         );
  AOI22_X1 U6899 ( .A1(n6383), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .B1(n6427), 
        .B2(REIP_REG_17__SCAN_IN), .ZN(n5740) );
  OAI21_X1 U6900 ( .B1(n5741), .B2(n6391), .A(n5740), .ZN(n5742) );
  AOI21_X1 U6901 ( .B1(n5743), .B2(n6379), .A(n5742), .ZN(n5744) );
  OAI21_X1 U6902 ( .B1(n6012), .B2(n6357), .A(n5744), .ZN(U2969) );
  INV_X1 U6903 ( .A(n5745), .ZN(n5749) );
  OAI21_X1 U6904 ( .B1(n5747), .B2(n5749), .A(n5746), .ZN(n5748) );
  OAI21_X1 U6905 ( .B1(n5731), .B2(n5749), .A(n5748), .ZN(n5901) );
  NAND2_X1 U6906 ( .A1(n6427), .A2(REIP_REG_16__SCAN_IN), .ZN(n5897) );
  NAND2_X1 U6907 ( .A1(n6383), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5750)
         );
  OAI211_X1 U6908 ( .C1(n6391), .C2(n6065), .A(n5897), .B(n5750), .ZN(n5751)
         );
  AOI21_X1 U6909 ( .B1(n6244), .B2(n6379), .A(n5751), .ZN(n5752) );
  OAI21_X1 U6910 ( .B1(n5901), .B2(n6357), .A(n5752), .ZN(U2970) );
  OAI21_X1 U6911 ( .B1(n3167), .B2(n5753), .A(n5732), .ZN(n6022) );
  NAND2_X1 U6912 ( .A1(n6022), .A2(n6387), .ZN(n5758) );
  NAND2_X1 U6913 ( .A1(n6427), .A2(REIP_REG_15__SCAN_IN), .ZN(n6019) );
  OAI21_X1 U6914 ( .B1(n6372), .B2(n5755), .A(n6019), .ZN(n5756) );
  AOI21_X1 U6915 ( .B1(n6366), .B2(n6071), .A(n5756), .ZN(n5757) );
  OAI211_X1 U6916 ( .C1(n6359), .C2(n6072), .A(n5758), .B(n5757), .ZN(U2971)
         );
  INV_X1 U6917 ( .A(REIP_REG_14__SCAN_IN), .ZN(n5759) );
  OAI22_X1 U6918 ( .A1(n6372), .A2(n6081), .B1(n6392), .B2(n5759), .ZN(n5761)
         );
  NOR2_X1 U6919 ( .A1(n6083), .A2(n6359), .ZN(n5760) );
  AOI211_X1 U6920 ( .C1(n6366), .C2(n6084), .A(n5761), .B(n5760), .ZN(n5762)
         );
  OAI21_X1 U6921 ( .B1(n6357), .B2(n5763), .A(n5762), .ZN(U2972) );
  INV_X1 U6922 ( .A(n5764), .ZN(n5765) );
  NAND2_X1 U6923 ( .A1(n5765), .A2(n6379), .ZN(n5771) );
  OR2_X1 U6924 ( .A1(n5767), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6440)
         );
  NAND3_X1 U6925 ( .A1(n5766), .A2(n6440), .A3(n6387), .ZN(n5770) );
  NAND2_X1 U6926 ( .A1(n6427), .A2(REIP_REG_0__SCAN_IN), .ZN(n6442) );
  OAI21_X1 U6927 ( .B1(n6383), .B2(n5768), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5769) );
  NAND4_X1 U6928 ( .A1(n5771), .A2(n5770), .A3(n6442), .A4(n5769), .ZN(U2986)
         );
  INV_X1 U6929 ( .A(n5772), .ZN(n5781) );
  NAND3_X1 U6930 ( .A1(n5787), .A2(n5775), .A3(n5773), .ZN(n5779) );
  INV_X1 U6931 ( .A(n6403), .ZN(n5893) );
  OAI21_X1 U6932 ( .B1(n5893), .B2(n5775), .A(n5774), .ZN(n5792) );
  INV_X1 U6933 ( .A(n5776), .ZN(n5777) );
  OAI21_X1 U6934 ( .B1(n5783), .B2(n6394), .A(n5782), .ZN(U2987) );
  INV_X1 U6935 ( .A(n5784), .ZN(n5794) );
  INV_X1 U6936 ( .A(n5785), .ZN(n5789) );
  INV_X1 U6937 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5786) );
  NAND3_X1 U6938 ( .A1(n5787), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5786), .ZN(n5788) );
  OAI211_X1 U6939 ( .C1(n5790), .C2(n6431), .A(n5789), .B(n5788), .ZN(n5791)
         );
  AOI21_X1 U6940 ( .B1(n5792), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5791), 
        .ZN(n5793) );
  OAI21_X1 U6941 ( .B1(n5794), .B2(n6394), .A(n5793), .ZN(U2988) );
  INV_X1 U6942 ( .A(n5795), .ZN(n5804) );
  INV_X1 U6943 ( .A(n5807), .ZN(n5799) );
  XNOR2_X1 U6944 ( .A(n5796), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5798)
         );
  AOI21_X1 U6945 ( .B1(n5799), .B2(n5798), .A(n5797), .ZN(n5800) );
  OAI21_X1 U6946 ( .B1(n5801), .B2(n6431), .A(n5800), .ZN(n5802) );
  AOI21_X1 U6947 ( .B1(n5810), .B2(INSTADDRPOINTER_REG_28__SCAN_IN), .A(n5802), 
        .ZN(n5803) );
  OAI21_X1 U6948 ( .B1(n5804), .B2(n6394), .A(n5803), .ZN(U2990) );
  NOR2_X1 U6949 ( .A1(n5805), .A2(n6431), .ZN(n5809) );
  OAI21_X1 U6950 ( .B1(n5807), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5806), 
        .ZN(n5808) );
  AOI211_X1 U6951 ( .C1(n5810), .C2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5809), .B(n5808), .ZN(n5811) );
  OAI21_X1 U6952 ( .B1(n5812), .B2(n6394), .A(n5811), .ZN(U2991) );
  NAND2_X1 U6953 ( .A1(n5813), .A2(n6439), .ZN(n5822) );
  INV_X1 U6954 ( .A(n5814), .ZN(n5820) );
  AND3_X1 U6955 ( .A1(n5817), .A2(n5816), .A3(n5815), .ZN(n5818) );
  AOI211_X1 U6956 ( .C1(n5820), .C2(n6445), .A(n5819), .B(n5818), .ZN(n5821)
         );
  OAI211_X1 U6957 ( .C1(n6002), .C2(n5823), .A(n5822), .B(n5821), .ZN(U2992)
         );
  INV_X1 U6958 ( .A(n5824), .ZN(n5830) );
  NAND2_X1 U6959 ( .A1(n5826), .A2(n5825), .ZN(n5827) );
  OAI211_X1 U6960 ( .C1(n6431), .C2(n5943), .A(n5828), .B(n5827), .ZN(n5829)
         );
  AOI21_X1 U6961 ( .B1(n5830), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n5829), 
        .ZN(n5831) );
  OAI21_X1 U6962 ( .B1(n5832), .B2(n6394), .A(n5831), .ZN(U2995) );
  XNOR2_X1 U6963 ( .A(n5834), .B(n5833), .ZN(n5979) );
  NOR3_X1 U6964 ( .A1(n5837), .A2(n5836), .A3(n5835), .ZN(n5838) );
  AOI211_X1 U6965 ( .C1(n6445), .C2(n5979), .A(n5839), .B(n5838), .ZN(n5841)
         );
  NAND2_X1 U6966 ( .A1(n5848), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5840) );
  OAI211_X1 U6967 ( .C1(n5842), .C2(n6394), .A(n5841), .B(n5840), .ZN(U2996)
         );
  NAND2_X1 U6968 ( .A1(n5844), .A2(n5843), .ZN(n5845) );
  OAI211_X1 U6969 ( .C1(n6431), .C2(n5962), .A(n5846), .B(n5845), .ZN(n5847)
         );
  AOI21_X1 U6970 ( .B1(n5848), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5847), 
        .ZN(n5849) );
  OAI21_X1 U6971 ( .B1(n5850), .B2(n6394), .A(n5849), .ZN(U2997) );
  INV_X1 U6972 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5860) );
  INV_X1 U6973 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5886) );
  NAND2_X1 U6974 ( .A1(n5851), .A2(n5886), .ZN(n6017) );
  INV_X1 U6975 ( .A(n5852), .ZN(n5854) );
  AOI21_X1 U6976 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5854), .A(n5853), 
        .ZN(n5856) );
  AOI211_X1 U6977 ( .C1(n5858), .C2(n5857), .A(n5856), .B(n5855), .ZN(n6010)
         );
  OAI21_X1 U6978 ( .B1(n5859), .B2(n6017), .A(n6010), .ZN(n5885) );
  AOI21_X1 U6979 ( .B1(n5860), .B2(n6403), .A(n5885), .ZN(n5873) );
  NOR2_X1 U6980 ( .A1(n5861), .A2(n5873), .ZN(n5867) );
  INV_X1 U6981 ( .A(n5862), .ZN(n5892) );
  NAND2_X1 U6982 ( .A1(n5892), .A2(n6398), .ZN(n6025) );
  NOR2_X1 U6983 ( .A1(n5894), .A2(n6025), .ZN(n5888) );
  NAND2_X1 U6984 ( .A1(n5863), .A2(n5888), .ZN(n5875) );
  NOR3_X1 U6985 ( .A1(n5865), .A2(n5864), .A3(n5875), .ZN(n5866) );
  AOI211_X1 U6986 ( .C1(n6427), .C2(REIP_REG_20__SCAN_IN), .A(n5867), .B(n5866), .ZN(n5870) );
  NAND2_X1 U6987 ( .A1(n6445), .A2(n5868), .ZN(n5869) );
  OAI211_X1 U6988 ( .C1(n5871), .C2(n6394), .A(n5870), .B(n5869), .ZN(U2998)
         );
  NAND2_X1 U6989 ( .A1(n6384), .A2(REIP_REG_19__SCAN_IN), .ZN(n5872) );
  OAI221_X1 U6990 ( .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n5875), .C1(
        n5874), .C2(n5873), .A(n5872), .ZN(n5876) );
  AOI21_X1 U6991 ( .B1(n6445), .B2(n5877), .A(n5876), .ZN(n5878) );
  OAI21_X1 U6992 ( .B1(n5879), .B2(n6394), .A(n5878), .ZN(U2999) );
  OAI21_X1 U6993 ( .B1(n5731), .B2(n5881), .A(n5880), .ZN(n5882) );
  XOR2_X1 U6994 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .B(n5882), .Z(n5994) );
  INV_X1 U6995 ( .A(n5994), .ZN(n5891) );
  INV_X1 U6996 ( .A(REIP_REG_18__SCAN_IN), .ZN(n5883) );
  OAI22_X1 U6997 ( .A1(n6431), .A2(n6059), .B1(n6392), .B2(n5883), .ZN(n5884)
         );
  AOI21_X1 U6998 ( .B1(n5885), .B2(INSTADDRPOINTER_REG_18__SCAN_IN), .A(n5884), 
        .ZN(n5890) );
  NOR2_X1 U6999 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n5886), .ZN(n5887)
         );
  NAND2_X1 U7000 ( .A1(n5888), .A2(n5887), .ZN(n5889) );
  OAI211_X1 U7001 ( .C1(n5891), .C2(n6394), .A(n5890), .B(n5889), .ZN(U3000)
         );
  OAI21_X1 U7002 ( .B1(n5893), .B2(n5892), .A(n6401), .ZN(n6021) );
  OAI21_X1 U7003 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A(n5894), .ZN(n5898) );
  INV_X1 U7004 ( .A(n6064), .ZN(n5895) );
  NAND2_X1 U7005 ( .A1(n6445), .A2(n5895), .ZN(n5896) );
  OAI211_X1 U7006 ( .C1(n6025), .C2(n5898), .A(n5897), .B(n5896), .ZN(n5899)
         );
  AOI21_X1 U7007 ( .B1(n6021), .B2(INSTADDRPOINTER_REG_16__SCAN_IN), .A(n5899), 
        .ZN(n5900) );
  OAI21_X1 U7008 ( .B1(n5901), .B2(n6394), .A(n5900), .ZN(U3002) );
  OAI21_X1 U7009 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n5902), .A(n6515), .ZN(
        n5903) );
  OAI21_X1 U7010 ( .B1(n5911), .B2(n6214), .A(n5903), .ZN(n5904) );
  MUX2_X1 U7011 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5904), .S(n6453), 
        .Z(U3464) );
  XNOR2_X1 U7012 ( .A(n4587), .B(n5905), .ZN(n5906) );
  OAI22_X1 U7013 ( .A1(n5906), .A2(n6519), .B1(n6196), .B2(n5911), .ZN(n5907)
         );
  MUX2_X1 U7014 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5907), .S(n6453), 
        .Z(U3463) );
  INV_X1 U7015 ( .A(n4651), .ZN(n5913) );
  AOI21_X1 U7016 ( .B1(n5910), .B2(n5909), .A(n5908), .ZN(n5912) );
  OAI222_X1 U7017 ( .A1(n5914), .A2(n5913), .B1(n6519), .B2(n5912), .C1(n5911), 
        .C2(n6458), .ZN(n5915) );
  MUX2_X1 U7018 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n5915), .S(n6453), 
        .Z(U3462) );
  INV_X1 U7019 ( .A(n5916), .ZN(n5922) );
  NAND2_X1 U7020 ( .A1(n5918), .A2(n5917), .ZN(n5923) );
  OAI22_X1 U7021 ( .A1(n5920), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(n5923), .B2(n5919), .ZN(n5921) );
  AOI21_X1 U7022 ( .B1(n3170), .B2(n5922), .A(n5921), .ZN(n6582) );
  INV_X1 U7023 ( .A(n6027), .ZN(n5929) );
  INV_X1 U7024 ( .A(n5923), .ZN(n5926) );
  AOI22_X1 U7025 ( .A1(n5927), .A2(n5926), .B1(n5925), .B2(n5924), .ZN(n5928)
         );
  OAI21_X1 U7026 ( .B1(n6582), .B2(n5929), .A(n5928), .ZN(n5930) );
  MUX2_X1 U7027 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n5930), .S(n6032), 
        .Z(U3460) );
  NAND2_X1 U7028 ( .A1(n5931), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5941)
         );
  NOR2_X1 U7029 ( .A1(n5933), .A2(n5932), .ZN(n5934) );
  AOI21_X1 U7030 ( .B1(n5935), .B2(n6513), .A(n5934), .ZN(n5940) );
  NAND2_X1 U7031 ( .A1(n5936), .A2(n6469), .ZN(n5939) );
  NAND2_X1 U7032 ( .A1(n6512), .A2(n5937), .ZN(n5938) );
  NAND4_X1 U7033 ( .A1(n5941), .A2(n5940), .A3(n5939), .A4(n5938), .ZN(U3132)
         );
  AND2_X1 U7034 ( .A1(n6266), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI22_X1 U7035 ( .A1(PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n6212), .B1(n5942), 
        .B2(n6211), .ZN(n5950) );
  INV_X1 U7036 ( .A(n5943), .ZN(n5948) );
  INV_X1 U7037 ( .A(REIP_REG_21__SCAN_IN), .ZN(n7024) );
  NOR2_X1 U7038 ( .A1(n7024), .A2(n5955), .ZN(n5954) );
  AOI21_X1 U7039 ( .B1(REIP_REG_22__SCAN_IN), .B2(n5954), .A(
        REIP_REG_23__SCAN_IN), .ZN(n5944) );
  OAI22_X1 U7040 ( .A1(n5946), .A2(n6162), .B1(n5945), .B2(n5944), .ZN(n5947)
         );
  AOI21_X1 U7041 ( .B1(n5948), .B2(n6178), .A(n5947), .ZN(n5949) );
  OAI211_X1 U7042 ( .C1(n5951), .C2(n6224), .A(n5950), .B(n5949), .ZN(U2804)
         );
  AOI22_X1 U7043 ( .A1(EBX_REG_22__SCAN_IN), .A2(n6156), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6212), .ZN(n5959) );
  INV_X1 U7044 ( .A(n5952), .ZN(n5953) );
  AOI22_X1 U7045 ( .A1(n5953), .A2(n6211), .B1(n5979), .B2(n6178), .ZN(n5958)
         );
  INV_X1 U7046 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6913) );
  AOI22_X1 U7047 ( .A1(n5984), .A2(n6150), .B1(n6913), .B2(n5954), .ZN(n5957)
         );
  NOR2_X1 U7048 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5955), .ZN(n5964) );
  OAI21_X1 U7049 ( .B1(n5960), .B2(n5964), .A(REIP_REG_22__SCAN_IN), .ZN(n5956) );
  NAND4_X1 U7050 ( .A1(n5959), .A2(n5958), .A3(n5957), .A4(n5956), .ZN(U2805)
         );
  AOI22_X1 U7051 ( .A1(EBX_REG_21__SCAN_IN), .A2(n6156), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6212), .ZN(n5968) );
  AOI22_X1 U7052 ( .A1(n5961), .A2(n6211), .B1(REIP_REG_21__SCAN_IN), .B2(
        n5960), .ZN(n5967) );
  NOR2_X1 U7053 ( .A1(n5962), .A2(n6202), .ZN(n5963) );
  AOI21_X1 U7054 ( .B1(n5987), .B2(n6150), .A(n5963), .ZN(n5966) );
  INV_X1 U7055 ( .A(n5964), .ZN(n5965) );
  NAND4_X1 U7056 ( .A1(n5968), .A2(n5967), .A3(n5966), .A4(n5965), .ZN(U2806)
         );
  AOI22_X1 U7057 ( .A1(n5969), .A2(n6211), .B1(REIP_REG_19__SCAN_IN), .B2(
        n6052), .ZN(n5970) );
  OAI211_X1 U7058 ( .C1(n6198), .C2(n5971), .A(n5970), .B(n6181), .ZN(n5975)
         );
  OAI22_X1 U7059 ( .A1(n5973), .A2(n6162), .B1(n5972), .B2(n6202), .ZN(n5974)
         );
  AOI211_X1 U7060 ( .C1(EBX_REG_19__SCAN_IN), .C2(n6156), .A(n5975), .B(n5974), 
        .ZN(n5978) );
  OAI211_X1 U7061 ( .C1(REIP_REG_19__SCAN_IN), .C2(REIP_REG_18__SCAN_IN), .A(
        n6056), .B(n5976), .ZN(n5977) );
  NAND2_X1 U7062 ( .A1(n5978), .A2(n5977), .ZN(U2808) );
  AOI22_X1 U7063 ( .A1(n5984), .A2(n4383), .B1(n5980), .B2(n5979), .ZN(n5981)
         );
  OAI21_X1 U7064 ( .B1(n6230), .B2(n5982), .A(n5981), .ZN(U2837) );
  INV_X1 U7065 ( .A(n5983), .ZN(n6243) );
  AOI22_X1 U7066 ( .A1(n5984), .A2(n6243), .B1(n6242), .B2(DATAI_22_), .ZN(
        n5986) );
  AOI22_X1 U7067 ( .A1(n6246), .A2(DATAI_6_), .B1(n6245), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5985) );
  NAND2_X1 U7068 ( .A1(n5986), .A2(n5985), .ZN(U2869) );
  AOI22_X1 U7069 ( .A1(n5987), .A2(n6243), .B1(n6242), .B2(DATAI_21_), .ZN(
        n5989) );
  AOI22_X1 U7070 ( .A1(n6246), .A2(DATAI_5_), .B1(n6245), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5988) );
  NAND2_X1 U7071 ( .A1(n5989), .A2(n5988), .ZN(U2870) );
  AOI22_X1 U7072 ( .A1(n5990), .A2(n6243), .B1(n6242), .B2(DATAI_20_), .ZN(
        n5992) );
  AOI22_X1 U7073 ( .A1(n6246), .A2(DATAI_4_), .B1(n6245), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5991) );
  NAND2_X1 U7074 ( .A1(n5992), .A2(n5991), .ZN(U2871) );
  AOI22_X1 U7075 ( .A1(n6384), .A2(REIP_REG_18__SCAN_IN), .B1(n6383), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5996) );
  AOI22_X1 U7076 ( .A1(n5994), .A2(n6387), .B1(n6379), .B2(n6239), .ZN(n5995)
         );
  OAI211_X1 U7077 ( .C1(n6391), .C2(n6054), .A(n5996), .B(n5995), .ZN(U2968)
         );
  OAI22_X1 U7078 ( .A1(n5997), .A2(n6359), .B1(n6100), .B2(n6391), .ZN(n5998)
         );
  AOI21_X1 U7079 ( .B1(n6387), .B2(n5999), .A(n5998), .ZN(n6001) );
  OAI211_X1 U7080 ( .C1(n3725), .C2(n6372), .A(n6001), .B(n6000), .ZN(U2973)
         );
  INV_X1 U7081 ( .A(n6002), .ZN(n6003) );
  AOI22_X1 U7082 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n6003), .B1(n6384), .B2(REIP_REG_25__SCAN_IN), .ZN(n6008) );
  INV_X1 U7083 ( .A(n6004), .ZN(n6005) );
  AOI22_X1 U7084 ( .A1(n6006), .A2(n6439), .B1(n6445), .B2(n6005), .ZN(n6007)
         );
  OAI211_X1 U7085 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n6009), .A(n6008), .B(n6007), .ZN(U2993) );
  INV_X1 U7086 ( .A(n6010), .ZN(n6011) );
  AOI22_X1 U7087 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n6011), .B1(n6384), .B2(REIP_REG_17__SCAN_IN), .ZN(n6016) );
  INV_X1 U7088 ( .A(n6012), .ZN(n6014) );
  AOI22_X1 U7089 ( .A1(n6014), .A2(n6439), .B1(n6445), .B2(n6013), .ZN(n6015)
         );
  OAI211_X1 U7090 ( .C1(n6018), .C2(n6017), .A(n6016), .B(n6015), .ZN(U3001)
         );
  INV_X1 U7091 ( .A(n6019), .ZN(n6020) );
  AOI21_X1 U7092 ( .B1(n6445), .B2(n6070), .A(n6020), .ZN(n6024) );
  AOI22_X1 U7093 ( .A1(n6022), .A2(n6439), .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n6021), .ZN(n6023) );
  OAI211_X1 U7094 ( .C1(INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n6025), .A(n6024), .B(n6023), .ZN(U3003) );
  INV_X1 U7095 ( .A(n6184), .ZN(n6029) );
  NAND4_X1 U7096 ( .A1(n6029), .A2(n6028), .A3(n6027), .A4(n6026), .ZN(n6030)
         );
  OAI21_X1 U7097 ( .B1(n6032), .B2(n6031), .A(n6030), .ZN(U3455) );
  NAND2_X1 U7098 ( .A1(n6961), .A2(STATE_REG_1__SCAN_IN), .ZN(n7093) );
  INV_X2 U7099 ( .A(n7093), .ZN(n7094) );
  INV_X1 U7100 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6923) );
  INV_X1 U7101 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6936) );
  OAI221_X2 U7102 ( .B1(n6936), .B2(n6961), .C1(STATE_REG_1__SCAN_IN), .C2(
        n6961), .A(n7093), .ZN(n6629) );
  OAI21_X1 U7103 ( .B1(n7094), .B2(n6923), .A(n6629), .ZN(U2789) );
  OAI21_X1 U7104 ( .B1(n6033), .B2(n6620), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6034) );
  OAI21_X1 U7105 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6621), .A(n6034), .ZN(
        U2790) );
  INV_X1 U7106 ( .A(D_C_N_REG_SCAN_IN), .ZN(n6958) );
  NOR2_X1 U7107 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6036) );
  NOR2_X1 U7108 ( .A1(n7094), .A2(n6036), .ZN(n6035) );
  AOI22_X1 U7109 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(n7094), .B1(n6958), .B2(
        n6035), .ZN(U2791) );
  INV_X1 U7110 ( .A(n6629), .ZN(n6679) );
  OAI21_X1 U7111 ( .B1(BS16_N), .B2(n6036), .A(n6679), .ZN(n6678) );
  OAI21_X1 U7112 ( .B1(n6679), .B2(n6786), .A(n6678), .ZN(U2792) );
  OAI21_X1 U7113 ( .B1(n6037), .B2(n7063), .A(n6357), .ZN(U2793) );
  NOR4_X1 U7114 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(
        DATAWIDTH_REG_14__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(
        DATAWIDTH_REG_7__SCAN_IN), .ZN(n6041) );
  NOR4_X1 U7115 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(
        DATAWIDTH_REG_10__SCAN_IN), .A3(DATAWIDTH_REG_23__SCAN_IN), .A4(
        DATAWIDTH_REG_3__SCAN_IN), .ZN(n6040) );
  NOR4_X1 U7116 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6039) );
  NOR4_X1 U7117 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n6038) );
  NAND4_X1 U7118 ( .A1(n6041), .A2(n6040), .A3(n6039), .A4(n6038), .ZN(n6047)
         );
  NOR4_X1 U7119 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(DATAWIDTH_REG_6__SCAN_IN), .A3(DATAWIDTH_REG_5__SCAN_IN), .A4(DATAWIDTH_REG_20__SCAN_IN), .ZN(n6045) );
  AOI211_X1 U7120 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_11__SCAN_IN), .B(
        DATAWIDTH_REG_2__SCAN_IN), .ZN(n6044) );
  NOR4_X1 U7121 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_17__SCAN_IN), .A4(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n6043) );
  NOR4_X1 U7122 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(DATAWIDTH_REG_16__SCAN_IN), .A3(DATAWIDTH_REG_9__SCAN_IN), .A4(DATAWIDTH_REG_8__SCAN_IN), .ZN(n6042) );
  NAND4_X1 U7123 ( .A1(n6045), .A2(n6044), .A3(n6043), .A4(n6042), .ZN(n6046)
         );
  NOR2_X1 U7124 ( .A1(n6047), .A2(n6046), .ZN(n6689) );
  INV_X1 U7125 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6675) );
  NOR3_X1 U7126 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6049) );
  OAI21_X1 U7127 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6049), .A(n6689), .ZN(n6048)
         );
  OAI21_X1 U7128 ( .B1(n6689), .B2(n6675), .A(n6048), .ZN(U2794) );
  INV_X1 U7129 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6831) );
  AOI21_X1 U7130 ( .B1(n6684), .B2(n6831), .A(n6049), .ZN(n6051) );
  INV_X1 U7131 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6050) );
  INV_X1 U7132 ( .A(n6689), .ZN(n6686) );
  AOI22_X1 U7133 ( .A1(n6689), .A2(n6051), .B1(n6050), .B2(n6686), .ZN(U2795)
         );
  AOI22_X1 U7134 ( .A1(EBX_REG_18__SCAN_IN), .A2(n6156), .B1(
        REIP_REG_18__SCAN_IN), .B2(n6052), .ZN(n6053) );
  OAI21_X1 U7135 ( .B1(n6054), .B2(n6205), .A(n6053), .ZN(n6055) );
  AOI211_X1 U7136 ( .C1(n6212), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6169), 
        .B(n6055), .ZN(n6058) );
  AOI22_X1 U7137 ( .A1(n6239), .A2(n6150), .B1(n5883), .B2(n6056), .ZN(n6057)
         );
  OAI211_X1 U7138 ( .C1(n6202), .C2(n6059), .A(n6058), .B(n6057), .ZN(U2809)
         );
  OAI21_X1 U7139 ( .B1(REIP_REG_16__SCAN_IN), .B2(REIP_REG_15__SCAN_IN), .A(
        n6060), .ZN(n6069) );
  INV_X1 U7140 ( .A(REIP_REG_16__SCAN_IN), .ZN(n7036) );
  NAND2_X1 U7141 ( .A1(n6062), .A2(n6061), .ZN(n6088) );
  AOI22_X1 U7142 ( .A1(EBX_REG_16__SCAN_IN), .A2(n6156), .B1(
        PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n6212), .ZN(n6063) );
  OAI211_X1 U7143 ( .C1(n7036), .C2(n6088), .A(n6063), .B(n6181), .ZN(n6067)
         );
  OAI22_X1 U7144 ( .A1(n6205), .A2(n6065), .B1(n6202), .B2(n6064), .ZN(n6066)
         );
  AOI211_X1 U7145 ( .C1(n6244), .C2(n6150), .A(n6067), .B(n6066), .ZN(n6068)
         );
  OAI21_X1 U7146 ( .B1(n6078), .B2(n6069), .A(n6068), .ZN(U2811) );
  AOI22_X1 U7147 ( .A1(n6071), .A2(n6211), .B1(n6178), .B2(n6070), .ZN(n6077)
         );
  INV_X1 U7148 ( .A(n6072), .ZN(n6075) );
  INV_X1 U7149 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6665) );
  AOI22_X1 U7150 ( .A1(EBX_REG_15__SCAN_IN), .A2(n6156), .B1(
        PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n6212), .ZN(n6073) );
  OAI211_X1 U7151 ( .C1(n6665), .C2(n6088), .A(n6073), .B(n6181), .ZN(n6074)
         );
  AOI21_X1 U7152 ( .B1(n6075), .B2(n6150), .A(n6074), .ZN(n6076) );
  OAI211_X1 U7153 ( .C1(REIP_REG_15__SCAN_IN), .C2(n6078), .A(n6077), .B(n6076), .ZN(U2812) );
  NOR2_X1 U7154 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6079), .ZN(n6089) );
  OAI22_X1 U7155 ( .A1(n6081), .A2(n6198), .B1(n6202), .B2(n6080), .ZN(n6082)
         );
  AOI211_X1 U7156 ( .C1(n6156), .C2(EBX_REG_14__SCAN_IN), .A(n6169), .B(n6082), 
        .ZN(n6087) );
  INV_X1 U7157 ( .A(n6083), .ZN(n6085) );
  AOI22_X1 U7158 ( .A1(n6085), .A2(n6150), .B1(n6211), .B2(n6084), .ZN(n6086)
         );
  OAI211_X1 U7159 ( .C1(n6089), .C2(n6088), .A(n6087), .B(n6086), .ZN(U2813)
         );
  NOR2_X1 U7160 ( .A1(n6122), .A2(n6090), .ZN(n6101) );
  OAI21_X1 U7161 ( .B1(n6198), .B2(n3725), .A(n6181), .ZN(n6094) );
  OAI22_X1 U7162 ( .A1(n6092), .A2(n6224), .B1(n6202), .B2(n6091), .ZN(n6093)
         );
  AOI211_X1 U7163 ( .C1(REIP_REG_13__SCAN_IN), .C2(n6101), .A(n6094), .B(n6093), .ZN(n6099) );
  INV_X1 U7164 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6662) );
  INV_X1 U7165 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6661) );
  AOI21_X1 U7166 ( .B1(n6662), .B2(n6661), .A(n6109), .ZN(n6096) );
  AOI22_X1 U7167 ( .A1(n6097), .A2(n6150), .B1(n6096), .B2(n6095), .ZN(n6098)
         );
  OAI211_X1 U7168 ( .C1(n6100), .C2(n6205), .A(n6099), .B(n6098), .ZN(U2814)
         );
  AOI22_X1 U7169 ( .A1(EBX_REG_12__SCAN_IN), .A2(n6156), .B1(
        REIP_REG_12__SCAN_IN), .B2(n6101), .ZN(n6102) );
  OAI21_X1 U7170 ( .B1(n6202), .B2(n6103), .A(n6102), .ZN(n6104) );
  AOI211_X1 U7171 ( .C1(n6212), .C2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n6169), 
        .B(n6104), .ZN(n6108) );
  AOI22_X1 U7172 ( .A1(n6106), .A2(n6150), .B1(n6105), .B2(n6211), .ZN(n6107)
         );
  OAI211_X1 U7173 ( .C1(REIP_REG_12__SCAN_IN), .C2(n6109), .A(n6108), .B(n6107), .ZN(U2815) );
  AOI21_X1 U7174 ( .B1(n6112), .B2(n6111), .A(n6110), .ZN(n6225) );
  AOI22_X1 U7175 ( .A1(n6178), .A2(n6225), .B1(n6113), .B2(n6660), .ZN(n6120)
         );
  OAI22_X1 U7176 ( .A1(n6115), .A2(n6198), .B1(n6660), .B2(n6114), .ZN(n6116)
         );
  AOI211_X1 U7177 ( .C1(n6156), .C2(EBX_REG_11__SCAN_IN), .A(n6169), .B(n6116), 
        .ZN(n6119) );
  OAI22_X1 U7178 ( .A1(n6353), .A2(n6162), .B1(n6205), .B2(n6352), .ZN(n6117)
         );
  INV_X1 U7179 ( .A(n6117), .ZN(n6118) );
  NAND3_X1 U7180 ( .A1(n6120), .A2(n6119), .A3(n6118), .ZN(U2816) );
  NOR2_X1 U7181 ( .A1(n6122), .A2(n6121), .ZN(n6131) );
  AOI22_X1 U7182 ( .A1(n6178), .A2(n6416), .B1(REIP_REG_9__SCAN_IN), .B2(n6131), .ZN(n6129) );
  AOI22_X1 U7183 ( .A1(EBX_REG_9__SCAN_IN), .A2(n6156), .B1(
        PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n6212), .ZN(n6128) );
  INV_X1 U7184 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6657) );
  AOI21_X1 U7185 ( .B1(n6123), .B2(n6657), .A(n6169), .ZN(n6127) );
  AOI22_X1 U7186 ( .A1(n6125), .A2(n6150), .B1(n6211), .B2(n6124), .ZN(n6126)
         );
  NAND4_X1 U7187 ( .A1(n6129), .A2(n6128), .A3(n6127), .A4(n6126), .ZN(U2818)
         );
  INV_X1 U7188 ( .A(n6130), .ZN(n6132) );
  AOI22_X1 U7189 ( .A1(n6178), .A2(n6132), .B1(REIP_REG_8__SCAN_IN), .B2(n6131), .ZN(n6142) );
  NAND3_X1 U7190 ( .A1(n6192), .A2(n6133), .A3(n6656), .ZN(n6134) );
  OAI211_X1 U7191 ( .C1(n6224), .C2(n6135), .A(n6181), .B(n6134), .ZN(n6136)
         );
  AOI21_X1 U7192 ( .B1(PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n6212), .A(n6136), 
        .ZN(n6141) );
  INV_X1 U7193 ( .A(n6137), .ZN(n6138) );
  AOI22_X1 U7194 ( .A1(n6139), .A2(n6150), .B1(n6138), .B2(n6211), .ZN(n6140)
         );
  NAND3_X1 U7195 ( .A1(n6142), .A2(n6141), .A3(n6140), .ZN(U2819) );
  OR3_X1 U7196 ( .A1(n6190), .A2(n6143), .A3(REIP_REG_7__SCAN_IN), .ZN(n6144)
         );
  OAI211_X1 U7197 ( .C1(n6198), .C2(n3650), .A(n6181), .B(n6144), .ZN(n6148)
         );
  AOI22_X1 U7198 ( .A1(EBX_REG_7__SCAN_IN), .A2(n6156), .B1(n6178), .B2(n6145), 
        .ZN(n6146) );
  INV_X1 U7199 ( .A(n6146), .ZN(n6147) );
  AOI211_X1 U7200 ( .C1(n6150), .C2(n6149), .A(n6148), .B(n6147), .ZN(n6153)
         );
  OAI21_X1 U7201 ( .B1(n6151), .B2(n6190), .A(n6215), .ZN(n6171) );
  AND3_X1 U7202 ( .A1(n6192), .A2(n6652), .A3(n6151), .ZN(n6155) );
  OAI21_X1 U7203 ( .B1(n6171), .B2(n6155), .A(REIP_REG_7__SCAN_IN), .ZN(n6152)
         );
  OAI211_X1 U7204 ( .C1(n6205), .C2(n6358), .A(n6153), .B(n6152), .ZN(U2820)
         );
  AOI22_X1 U7205 ( .A1(n6178), .A2(n6154), .B1(REIP_REG_6__SCAN_IN), .B2(n6171), .ZN(n6160) );
  AOI211_X1 U7206 ( .C1(n6156), .C2(EBX_REG_6__SCAN_IN), .A(n6169), .B(n6155), 
        .ZN(n6157) );
  INV_X1 U7207 ( .A(n6157), .ZN(n6158) );
  AOI21_X1 U7208 ( .B1(n6212), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6158), 
        .ZN(n6159) );
  OAI211_X1 U7209 ( .C1(n6162), .C2(n6161), .A(n6160), .B(n6159), .ZN(n6163)
         );
  INV_X1 U7210 ( .A(n6163), .ZN(n6164) );
  OAI21_X1 U7211 ( .B1(n6165), .B2(n6205), .A(n6164), .ZN(U2821) );
  OAI21_X1 U7212 ( .B1(n6190), .B2(n6166), .A(n6651), .ZN(n6170) );
  INV_X1 U7213 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6373) );
  OAI22_X1 U7214 ( .A1(n6167), .A2(n6224), .B1(n6373), .B2(n6198), .ZN(n6168)
         );
  AOI211_X1 U7215 ( .C1(n6171), .C2(n6170), .A(n6169), .B(n6168), .ZN(n6174)
         );
  AOI22_X1 U7216 ( .A1(n6368), .A2(n6221), .B1(n6178), .B2(n6172), .ZN(n6173)
         );
  OAI211_X1 U7217 ( .C1(n6365), .C2(n6205), .A(n6174), .B(n6173), .ZN(U2822)
         );
  INV_X1 U7218 ( .A(n6175), .ZN(n6177) );
  AOI22_X1 U7219 ( .A1(n6178), .A2(n6177), .B1(REIP_REG_4__SCAN_IN), .B2(n6176), .ZN(n6188) );
  NAND3_X1 U7220 ( .A1(n6192), .A2(n6179), .A3(n6649), .ZN(n6180) );
  OAI211_X1 U7221 ( .C1(n6224), .C2(n4158), .A(n6181), .B(n6180), .ZN(n6182)
         );
  AOI21_X1 U7222 ( .B1(n6212), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6182), 
        .ZN(n6183) );
  OAI21_X1 U7223 ( .B1(n6184), .B2(n6213), .A(n6183), .ZN(n6185) );
  AOI21_X1 U7224 ( .B1(n6186), .B2(n6221), .A(n6185), .ZN(n6187) );
  OAI211_X1 U7225 ( .C1(n6189), .C2(n6205), .A(n6188), .B(n6187), .ZN(U2823)
         );
  NOR2_X1 U7226 ( .A1(n6190), .A2(REIP_REG_1__SCAN_IN), .ZN(n6207) );
  NOR3_X1 U7227 ( .A1(n6191), .A2(n6647), .A3(n6207), .ZN(n6195) );
  AOI21_X1 U7228 ( .B1(n6192), .B2(REIP_REG_1__SCAN_IN), .A(
        REIP_REG_2__SCAN_IN), .ZN(n6194) );
  OAI22_X1 U7229 ( .A1(n6195), .A2(n6194), .B1(n6193), .B2(n6224), .ZN(n6200)
         );
  OAI22_X1 U7230 ( .A1(n6198), .A2(n6197), .B1(n6196), .B2(n6213), .ZN(n6199)
         );
  NOR2_X1 U7231 ( .A1(n6200), .A2(n6199), .ZN(n6201) );
  OAI21_X1 U7232 ( .B1(n6202), .B2(n6430), .A(n6201), .ZN(n6203) );
  AOI21_X1 U7233 ( .B1(n6378), .B2(n6221), .A(n6203), .ZN(n6204) );
  OAI21_X1 U7234 ( .B1(n6382), .B2(n6205), .A(n6204), .ZN(U2825) );
  INV_X1 U7235 ( .A(n6206), .ZN(n6208) );
  AOI21_X1 U7236 ( .B1(n6209), .B2(n6208), .A(n6207), .ZN(n6223) );
  INV_X1 U7237 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6210) );
  NAND2_X1 U7238 ( .A1(n6211), .A2(n6210), .ZN(n6219) );
  NAND2_X1 U7239 ( .A1(n6212), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6218)
         );
  OAI22_X1 U7240 ( .A1(n6215), .A2(n6684), .B1(n6214), .B2(n6213), .ZN(n6216)
         );
  INV_X1 U7241 ( .A(n6216), .ZN(n6217) );
  NAND3_X1 U7242 ( .A1(n6219), .A2(n6218), .A3(n6217), .ZN(n6220) );
  AOI21_X1 U7243 ( .B1(n6386), .B2(n6221), .A(n6220), .ZN(n6222) );
  OAI211_X1 U7244 ( .C1(n3205), .C2(n6224), .A(n6223), .B(n6222), .ZN(U2826)
         );
  INV_X1 U7245 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6229) );
  INV_X1 U7246 ( .A(n6225), .ZN(n6393) );
  OAI22_X1 U7247 ( .A1(n6353), .A2(n6226), .B1(n6233), .B2(n6393), .ZN(n6227)
         );
  INV_X1 U7248 ( .A(n6227), .ZN(n6228) );
  OAI21_X1 U7249 ( .B1(n6230), .B2(n6229), .A(n6228), .ZN(U2848) );
  INV_X1 U7250 ( .A(EBX_REG_3__SCAN_IN), .ZN(n6237) );
  INV_X1 U7251 ( .A(n6231), .ZN(n6232) );
  OAI22_X1 U7252 ( .A1(n6234), .A2(n6226), .B1(n6233), .B2(n6232), .ZN(n6235)
         );
  INV_X1 U7253 ( .A(n6235), .ZN(n6236) );
  OAI21_X1 U7254 ( .B1(n6238), .B2(n6237), .A(n6236), .ZN(U2856) );
  AOI22_X1 U7255 ( .A1(n6239), .A2(n6243), .B1(n6242), .B2(DATAI_18_), .ZN(
        n6241) );
  AOI22_X1 U7256 ( .A1(n6246), .A2(DATAI_2_), .B1(n6245), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6240) );
  NAND2_X1 U7257 ( .A1(n6241), .A2(n6240), .ZN(U2873) );
  AOI22_X1 U7258 ( .A1(n6244), .A2(n6243), .B1(n6242), .B2(DATAI_16_), .ZN(
        n6248) );
  AOI22_X1 U7259 ( .A1(n6246), .A2(DATAI_0_), .B1(n6245), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6247) );
  NAND2_X1 U7260 ( .A1(n6248), .A2(n6247), .ZN(U2875) );
  AOI22_X1 U7261 ( .A1(n6267), .A2(LWORD_REG_15__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6250) );
  OAI21_X1 U7262 ( .B1(n6347), .B2(n6269), .A(n6250), .ZN(U2908) );
  AOI22_X1 U7263 ( .A1(n6267), .A2(LWORD_REG_14__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6251) );
  OAI21_X1 U7264 ( .B1(n6342), .B2(n6269), .A(n6251), .ZN(U2909) );
  AOI22_X1 U7265 ( .A1(n6267), .A2(LWORD_REG_13__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6252) );
  OAI21_X1 U7266 ( .B1(n6339), .B2(n6269), .A(n6252), .ZN(U2910) );
  AOI22_X1 U7267 ( .A1(n6267), .A2(LWORD_REG_12__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6253) );
  OAI21_X1 U7268 ( .B1(n6336), .B2(n6269), .A(n6253), .ZN(U2911) );
  AOI22_X1 U7269 ( .A1(n6267), .A2(LWORD_REG_11__SCAN_IN), .B1(n6261), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6254) );
  OAI21_X1 U7270 ( .B1(n6333), .B2(n6269), .A(n6254), .ZN(U2912) );
  AOI22_X1 U7271 ( .A1(n6267), .A2(LWORD_REG_10__SCAN_IN), .B1(n6261), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6255) );
  OAI21_X1 U7272 ( .B1(n6330), .B2(n6269), .A(n6255), .ZN(U2913) );
  AOI22_X1 U7273 ( .A1(n6267), .A2(LWORD_REG_9__SCAN_IN), .B1(n6261), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6256) );
  OAI21_X1 U7274 ( .B1(n6327), .B2(n6269), .A(n6256), .ZN(U2914) );
  AOI22_X1 U7275 ( .A1(n6267), .A2(LWORD_REG_8__SCAN_IN), .B1(n6261), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6257) );
  OAI21_X1 U7276 ( .B1(n6324), .B2(n6269), .A(n6257), .ZN(U2915) );
  AOI22_X1 U7277 ( .A1(n6267), .A2(LWORD_REG_7__SCAN_IN), .B1(n6261), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6258) );
  OAI21_X1 U7278 ( .B1(n3655), .B2(n6269), .A(n6258), .ZN(U2916) );
  AOI22_X1 U7279 ( .A1(n6267), .A2(LWORD_REG_6__SCAN_IN), .B1(n6261), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6259) );
  OAI21_X1 U7280 ( .B1(n6319), .B2(n6269), .A(n6259), .ZN(U2917) );
  AOI22_X1 U7281 ( .A1(n6267), .A2(LWORD_REG_5__SCAN_IN), .B1(n6261), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6260) );
  OAI21_X1 U7282 ( .B1(n3618), .B2(n6269), .A(n6260), .ZN(U2918) );
  AOI22_X1 U7283 ( .A1(n6267), .A2(LWORD_REG_4__SCAN_IN), .B1(n6261), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6262) );
  OAI21_X1 U7284 ( .B1(n6314), .B2(n6269), .A(n6262), .ZN(U2919) );
  AOI22_X1 U7285 ( .A1(n6267), .A2(LWORD_REG_3__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6263) );
  OAI21_X1 U7286 ( .B1(n6311), .B2(n6269), .A(n6263), .ZN(U2920) );
  AOI22_X1 U7287 ( .A1(n6267), .A2(LWORD_REG_2__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6264) );
  OAI21_X1 U7288 ( .B1(n6308), .B2(n6269), .A(n6264), .ZN(U2921) );
  AOI22_X1 U7289 ( .A1(n6267), .A2(LWORD_REG_1__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6265) );
  OAI21_X1 U7290 ( .B1(n6305), .B2(n6269), .A(n6265), .ZN(U2922) );
  AOI22_X1 U7291 ( .A1(n6267), .A2(LWORD_REG_0__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6268) );
  OAI21_X1 U7292 ( .B1(n6302), .B2(n6269), .A(n6268), .ZN(U2923) );
  AND2_X1 U7293 ( .A1(n6343), .A2(DATAI_0_), .ZN(n6300) );
  AOI21_X1 U7294 ( .B1(UWORD_REG_0__SCAN_IN), .B2(n6283), .A(n6300), .ZN(n6273) );
  OAI21_X1 U7295 ( .B1(n6274), .B2(n6346), .A(n6273), .ZN(U2924) );
  AND2_X1 U7296 ( .A1(n6343), .A2(DATAI_1_), .ZN(n6303) );
  AOI21_X1 U7297 ( .B1(UWORD_REG_1__SCAN_IN), .B2(n6283), .A(n6303), .ZN(n6275) );
  OAI21_X1 U7298 ( .B1(n6276), .B2(n6346), .A(n6275), .ZN(U2925) );
  AND2_X1 U7299 ( .A1(n6343), .A2(DATAI_2_), .ZN(n6306) );
  AOI21_X1 U7300 ( .B1(UWORD_REG_2__SCAN_IN), .B2(n6283), .A(n6306), .ZN(n6277) );
  OAI21_X1 U7301 ( .B1(n6278), .B2(n6346), .A(n6277), .ZN(U2926) );
  AND2_X1 U7302 ( .A1(n6343), .A2(DATAI_3_), .ZN(n6309) );
  AOI21_X1 U7303 ( .B1(UWORD_REG_3__SCAN_IN), .B2(n6283), .A(n6309), .ZN(n6279) );
  OAI21_X1 U7304 ( .B1(n6280), .B2(n6346), .A(n6279), .ZN(U2927) );
  AND2_X1 U7305 ( .A1(n6343), .A2(DATAI_4_), .ZN(n6312) );
  AOI21_X1 U7306 ( .B1(UWORD_REG_4__SCAN_IN), .B2(n6344), .A(n6312), .ZN(n6281) );
  OAI21_X1 U7307 ( .B1(n6282), .B2(n6346), .A(n6281), .ZN(U2928) );
  AND2_X1 U7308 ( .A1(n6343), .A2(DATAI_5_), .ZN(n6315) );
  AOI21_X1 U7309 ( .B1(UWORD_REG_5__SCAN_IN), .B2(n6283), .A(n6315), .ZN(n6284) );
  OAI21_X1 U7310 ( .B1(n6285), .B2(n6346), .A(n6284), .ZN(U2929) );
  AND2_X1 U7311 ( .A1(n6343), .A2(DATAI_6_), .ZN(n6317) );
  AOI21_X1 U7312 ( .B1(UWORD_REG_6__SCAN_IN), .B2(n6344), .A(n6317), .ZN(n6286) );
  OAI21_X1 U7313 ( .B1(n6287), .B2(n6346), .A(n6286), .ZN(U2930) );
  AND2_X1 U7314 ( .A1(n6343), .A2(DATAI_7_), .ZN(n6320) );
  AOI21_X1 U7315 ( .B1(UWORD_REG_7__SCAN_IN), .B2(n6344), .A(n6320), .ZN(n6288) );
  OAI21_X1 U7316 ( .B1(n3905), .B2(n6346), .A(n6288), .ZN(U2931) );
  AND2_X1 U7317 ( .A1(n6343), .A2(DATAI_8_), .ZN(n6322) );
  AOI21_X1 U7318 ( .B1(UWORD_REG_8__SCAN_IN), .B2(n6344), .A(n6322), .ZN(n6289) );
  OAI21_X1 U7319 ( .B1(n6290), .B2(n6346), .A(n6289), .ZN(U2932) );
  AND2_X1 U7320 ( .A1(n6343), .A2(DATAI_9_), .ZN(n6325) );
  AOI21_X1 U7321 ( .B1(UWORD_REG_9__SCAN_IN), .B2(n6344), .A(n6325), .ZN(n6291) );
  OAI21_X1 U7322 ( .B1(n3940), .B2(n6346), .A(n6291), .ZN(U2933) );
  AND2_X1 U7323 ( .A1(n6343), .A2(DATAI_10_), .ZN(n6328) );
  AOI21_X1 U7324 ( .B1(UWORD_REG_10__SCAN_IN), .B2(n6344), .A(n6328), .ZN(
        n6292) );
  OAI21_X1 U7325 ( .B1(n6293), .B2(n6346), .A(n6292), .ZN(U2934) );
  AND2_X1 U7326 ( .A1(n6343), .A2(DATAI_11_), .ZN(n6331) );
  AOI21_X1 U7327 ( .B1(UWORD_REG_11__SCAN_IN), .B2(n6344), .A(n6331), .ZN(
        n6294) );
  OAI21_X1 U7328 ( .B1(n3978), .B2(n6346), .A(n6294), .ZN(U2935) );
  AND2_X1 U7329 ( .A1(n6343), .A2(DATAI_12_), .ZN(n6334) );
  AOI21_X1 U7330 ( .B1(UWORD_REG_12__SCAN_IN), .B2(n6344), .A(n6334), .ZN(
        n6295) );
  OAI21_X1 U7331 ( .B1(n6296), .B2(n6346), .A(n6295), .ZN(U2936) );
  AND2_X1 U7332 ( .A1(n6343), .A2(DATAI_13_), .ZN(n6337) );
  AOI21_X1 U7333 ( .B1(UWORD_REG_13__SCAN_IN), .B2(n6344), .A(n6337), .ZN(
        n6297) );
  OAI21_X1 U7334 ( .B1(n4019), .B2(n6346), .A(n6297), .ZN(U2937) );
  AND2_X1 U7335 ( .A1(n6343), .A2(DATAI_14_), .ZN(n6340) );
  AOI21_X1 U7336 ( .B1(UWORD_REG_14__SCAN_IN), .B2(n6344), .A(n6340), .ZN(
        n6298) );
  OAI21_X1 U7337 ( .B1(n6299), .B2(n6346), .A(n6298), .ZN(U2938) );
  AOI21_X1 U7338 ( .B1(LWORD_REG_0__SCAN_IN), .B2(n6344), .A(n6300), .ZN(n6301) );
  OAI21_X1 U7339 ( .B1(n6302), .B2(n6346), .A(n6301), .ZN(U2939) );
  AOI21_X1 U7340 ( .B1(LWORD_REG_1__SCAN_IN), .B2(n6344), .A(n6303), .ZN(n6304) );
  OAI21_X1 U7341 ( .B1(n6305), .B2(n6346), .A(n6304), .ZN(U2940) );
  AOI21_X1 U7342 ( .B1(LWORD_REG_2__SCAN_IN), .B2(n6344), .A(n6306), .ZN(n6307) );
  OAI21_X1 U7343 ( .B1(n6308), .B2(n6346), .A(n6307), .ZN(U2941) );
  AOI21_X1 U7344 ( .B1(LWORD_REG_3__SCAN_IN), .B2(n6344), .A(n6309), .ZN(n6310) );
  OAI21_X1 U7345 ( .B1(n6311), .B2(n6346), .A(n6310), .ZN(U2942) );
  AOI21_X1 U7346 ( .B1(LWORD_REG_4__SCAN_IN), .B2(n6344), .A(n6312), .ZN(n6313) );
  OAI21_X1 U7347 ( .B1(n6314), .B2(n6346), .A(n6313), .ZN(U2943) );
  AOI21_X1 U7348 ( .B1(LWORD_REG_5__SCAN_IN), .B2(n6344), .A(n6315), .ZN(n6316) );
  OAI21_X1 U7349 ( .B1(n3618), .B2(n6346), .A(n6316), .ZN(U2944) );
  AOI21_X1 U7350 ( .B1(LWORD_REG_6__SCAN_IN), .B2(n6344), .A(n6317), .ZN(n6318) );
  OAI21_X1 U7351 ( .B1(n6319), .B2(n6346), .A(n6318), .ZN(U2945) );
  AOI21_X1 U7352 ( .B1(LWORD_REG_7__SCAN_IN), .B2(n6344), .A(n6320), .ZN(n6321) );
  OAI21_X1 U7353 ( .B1(n3655), .B2(n6346), .A(n6321), .ZN(U2946) );
  AOI21_X1 U7354 ( .B1(LWORD_REG_8__SCAN_IN), .B2(n6344), .A(n6322), .ZN(n6323) );
  OAI21_X1 U7355 ( .B1(n6324), .B2(n6346), .A(n6323), .ZN(U2947) );
  AOI21_X1 U7356 ( .B1(LWORD_REG_9__SCAN_IN), .B2(n6344), .A(n6325), .ZN(n6326) );
  OAI21_X1 U7357 ( .B1(n6327), .B2(n6346), .A(n6326), .ZN(U2948) );
  AOI21_X1 U7358 ( .B1(LWORD_REG_10__SCAN_IN), .B2(n6344), .A(n6328), .ZN(
        n6329) );
  OAI21_X1 U7359 ( .B1(n6330), .B2(n6346), .A(n6329), .ZN(U2949) );
  AOI21_X1 U7360 ( .B1(LWORD_REG_11__SCAN_IN), .B2(n6344), .A(n6331), .ZN(
        n6332) );
  OAI21_X1 U7361 ( .B1(n6333), .B2(n6346), .A(n6332), .ZN(U2950) );
  AOI21_X1 U7362 ( .B1(LWORD_REG_12__SCAN_IN), .B2(n6344), .A(n6334), .ZN(
        n6335) );
  OAI21_X1 U7363 ( .B1(n6336), .B2(n6346), .A(n6335), .ZN(U2951) );
  AOI21_X1 U7364 ( .B1(LWORD_REG_13__SCAN_IN), .B2(n6344), .A(n6337), .ZN(
        n6338) );
  OAI21_X1 U7365 ( .B1(n6339), .B2(n6346), .A(n6338), .ZN(U2952) );
  AOI21_X1 U7366 ( .B1(LWORD_REG_14__SCAN_IN), .B2(n6344), .A(n6340), .ZN(
        n6341) );
  OAI21_X1 U7367 ( .B1(n6342), .B2(n6346), .A(n6341), .ZN(U2953) );
  AOI22_X1 U7368 ( .A1(n6344), .A2(LWORD_REG_15__SCAN_IN), .B1(n6343), .B2(
        DATAI_15_), .ZN(n6345) );
  OAI21_X1 U7369 ( .B1(n6347), .B2(n6346), .A(n6345), .ZN(U2954) );
  NAND2_X1 U7370 ( .A1(n6349), .A2(n6348), .ZN(n6351) );
  XOR2_X1 U7371 ( .A(n6351), .B(n6350), .Z(n6395) );
  AOI22_X1 U7372 ( .A1(n6384), .A2(REIP_REG_11__SCAN_IN), .B1(n6383), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6356) );
  OAI22_X1 U7373 ( .A1(n6353), .A2(n6359), .B1(n6391), .B2(n6352), .ZN(n6354)
         );
  INV_X1 U7374 ( .A(n6354), .ZN(n6355) );
  OAI211_X1 U7375 ( .C1(n6395), .C2(n6357), .A(n6356), .B(n6355), .ZN(U2975)
         );
  OAI22_X1 U7376 ( .A1(n6360), .A2(n6359), .B1(n6358), .B2(n6391), .ZN(n6361)
         );
  AOI21_X1 U7377 ( .B1(n6362), .B2(n6387), .A(n6361), .ZN(n6364) );
  OAI211_X1 U7378 ( .C1(n3650), .C2(n6372), .A(n6364), .B(n6363), .ZN(U2979)
         );
  INV_X1 U7379 ( .A(n6365), .ZN(n6367) );
  AOI222_X1 U7380 ( .A1(n6369), .A2(n6387), .B1(n6379), .B2(n6368), .C1(n6367), 
        .C2(n6366), .ZN(n6371) );
  OAI211_X1 U7381 ( .C1(n6373), .C2(n6372), .A(n6371), .B(n6370), .ZN(U2981)
         );
  AOI22_X1 U7382 ( .A1(n6384), .A2(REIP_REG_2__SCAN_IN), .B1(n6383), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6381) );
  NAND2_X1 U7383 ( .A1(n6376), .A2(n3159), .ZN(n6377) );
  XOR2_X1 U7384 ( .A(n6374), .B(n6377), .Z(n6435) );
  AOI22_X1 U7385 ( .A1(n6435), .A2(n6387), .B1(n6379), .B2(n6378), .ZN(n6380)
         );
  OAI211_X1 U7386 ( .C1(n6391), .C2(n6382), .A(n6381), .B(n6380), .ZN(U2984)
         );
  AOI22_X1 U7387 ( .A1(n6384), .A2(REIP_REG_1__SCAN_IN), .B1(n6383), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6390) );
  INV_X1 U7388 ( .A(n6385), .ZN(n6388) );
  AOI22_X1 U7389 ( .A1(n6388), .A2(n6387), .B1(n6386), .B2(n6379), .ZN(n6389)
         );
  OAI211_X1 U7390 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n6391), .A(n6390), 
        .B(n6389), .ZN(U2985) );
  OAI22_X1 U7391 ( .A1(n6431), .A2(n6393), .B1(n6660), .B2(n6392), .ZN(n6397)
         );
  NOR2_X1 U7392 ( .A1(n6395), .A2(n6394), .ZN(n6396) );
  AOI211_X1 U7393 ( .C1(n6400), .C2(n6398), .A(n6397), .B(n6396), .ZN(n6399)
         );
  OAI21_X1 U7394 ( .B1(n6401), .B2(n6400), .A(n6399), .ZN(U3007) );
  AOI21_X1 U7395 ( .B1(n6404), .B2(n6403), .A(n6402), .ZN(n6423) );
  INV_X1 U7396 ( .A(n6405), .ZN(n6412) );
  NAND2_X1 U7397 ( .A1(n6407), .A2(n6406), .ZN(n6418) );
  AOI221_X1 U7398 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .C1(n6422), .C2(n6414), .A(n6418), 
        .ZN(n6408) );
  AOI21_X1 U7399 ( .B1(n6427), .B2(REIP_REG_10__SCAN_IN), .A(n6408), .ZN(n6409) );
  OAI21_X1 U7400 ( .B1(n6431), .B2(n6410), .A(n6409), .ZN(n6411) );
  AOI21_X1 U7401 ( .B1(n6412), .B2(n6439), .A(n6411), .ZN(n6413) );
  OAI21_X1 U7402 ( .B1(n6423), .B2(n6414), .A(n6413), .ZN(U3008) );
  INV_X1 U7403 ( .A(n6415), .ZN(n6420) );
  AOI22_X1 U7404 ( .A1(n6445), .A2(n6416), .B1(n6427), .B2(REIP_REG_9__SCAN_IN), .ZN(n6417) );
  OAI21_X1 U7405 ( .B1(n6418), .B2(INSTADDRPOINTER_REG_9__SCAN_IN), .A(n6417), 
        .ZN(n6419) );
  AOI21_X1 U7406 ( .B1(n6420), .B2(n6439), .A(n6419), .ZN(n6421) );
  OAI21_X1 U7407 ( .B1(n6423), .B2(n6422), .A(n6421), .ZN(U3009) );
  NAND2_X1 U7408 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6424), .ZN(n6438)
         );
  NAND3_X1 U7409 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n6426), .A3(n6425), 
        .ZN(n6429) );
  NAND2_X1 U7410 ( .A1(n6427), .A2(REIP_REG_2__SCAN_IN), .ZN(n6428) );
  OAI211_X1 U7411 ( .C1(n6431), .C2(n6430), .A(n6429), .B(n6428), .ZN(n6434)
         );
  INV_X1 U7412 ( .A(n6432), .ZN(n6433) );
  AOI211_X1 U7413 ( .C1(n6435), .C2(n6439), .A(n6434), .B(n6433), .ZN(n6436)
         );
  OAI221_X1 U7414 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6438), .C1(n4258), .C2(n6437), .A(n6436), .ZN(U3016) );
  NAND3_X1 U7415 ( .A1(n6440), .A2(n5766), .A3(n6439), .ZN(n6448) );
  INV_X1 U7416 ( .A(n6441), .ZN(n6444) );
  INV_X1 U7417 ( .A(n6442), .ZN(n6443) );
  AOI21_X1 U7418 ( .B1(n6445), .B2(n6444), .A(n6443), .ZN(n6447) );
  AND3_X1 U7419 ( .A1(n6448), .A2(n6447), .A3(n6446), .ZN(n6449) );
  OAI221_X1 U7420 ( .B1(n6452), .B2(n6451), .C1(n6452), .C2(n6450), .A(n6449), 
        .ZN(U3018) );
  NOR2_X1 U7421 ( .A1(n6454), .A2(n6453), .ZN(U3019) );
  NAND2_X1 U7422 ( .A1(n6580), .A2(n6455), .ZN(n6465) );
  INV_X1 U7423 ( .A(n6465), .ZN(n6496) );
  AOI22_X1 U7424 ( .A1(n6459), .A2(n6458), .B1(n6457), .B2(n6456), .ZN(n6460)
         );
  AOI22_X1 U7425 ( .A1(n6512), .A2(n6496), .B1(n6526), .B2(n6495), .ZN(n6471)
         );
  INV_X1 U7426 ( .A(n6510), .ZN(n6461) );
  NOR3_X1 U7427 ( .A1(n6497), .A2(n6461), .A3(n6519), .ZN(n6464) );
  OAI21_X1 U7428 ( .B1(n6464), .B2(n6463), .A(n6462), .ZN(n6468) );
  AOI21_X1 U7429 ( .B1(n6465), .B2(STATE2_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6466) );
  NAND3_X1 U7430 ( .A1(n6468), .A2(n6467), .A3(n6466), .ZN(n6499) );
  AOI22_X1 U7431 ( .A1(n6499), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6469), 
        .B2(n6497), .ZN(n6470) );
  OAI211_X1 U7432 ( .C1(n6472), .C2(n6510), .A(n6471), .B(n6470), .ZN(U3068)
         );
  AOI22_X1 U7433 ( .A1(n6530), .A2(n6496), .B1(n6532), .B2(n6495), .ZN(n6475)
         );
  AOI22_X1 U7434 ( .A1(n6499), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6473), 
        .B2(n6497), .ZN(n6474) );
  OAI211_X1 U7435 ( .C1(n6476), .C2(n6510), .A(n6475), .B(n6474), .ZN(U3069)
         );
  AOI22_X1 U7436 ( .A1(n6536), .A2(n6496), .B1(n6539), .B2(n6495), .ZN(n6478)
         );
  AOI22_X1 U7437 ( .A1(n6499), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6537), 
        .B2(n6497), .ZN(n6477) );
  OAI211_X1 U7438 ( .C1(n6543), .C2(n6510), .A(n6478), .B(n6477), .ZN(U3070)
         );
  AOI22_X1 U7439 ( .A1(n6544), .A2(n6496), .B1(n6546), .B2(n6495), .ZN(n6481)
         );
  AOI22_X1 U7440 ( .A1(n6499), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6479), 
        .B2(n6497), .ZN(n6480) );
  OAI211_X1 U7441 ( .C1(n6482), .C2(n6510), .A(n6481), .B(n6480), .ZN(U3071)
         );
  AOI22_X1 U7442 ( .A1(n6550), .A2(n6496), .B1(n6552), .B2(n6495), .ZN(n6485)
         );
  AOI22_X1 U7443 ( .A1(n6499), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6483), 
        .B2(n6497), .ZN(n6484) );
  OAI211_X1 U7444 ( .C1(n6486), .C2(n6510), .A(n6485), .B(n6484), .ZN(U3072)
         );
  AOI22_X1 U7445 ( .A1(n6556), .A2(n6496), .B1(n6558), .B2(n6495), .ZN(n6489)
         );
  AOI22_X1 U7446 ( .A1(n6499), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6487), 
        .B2(n6497), .ZN(n6488) );
  OAI211_X1 U7447 ( .C1(n6490), .C2(n6510), .A(n6489), .B(n6488), .ZN(U3073)
         );
  AOI22_X1 U7448 ( .A1(n6562), .A2(n6496), .B1(n6564), .B2(n6495), .ZN(n6493)
         );
  AOI22_X1 U7449 ( .A1(n6499), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6491), 
        .B2(n6497), .ZN(n6492) );
  OAI211_X1 U7450 ( .C1(n6494), .C2(n6510), .A(n6493), .B(n6492), .ZN(U3074)
         );
  AOI22_X1 U7451 ( .A1(n6569), .A2(n6496), .B1(n6573), .B2(n6495), .ZN(n6501)
         );
  AOI22_X1 U7452 ( .A1(n6499), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6498), 
        .B2(n6497), .ZN(n6500) );
  OAI211_X1 U7453 ( .C1(n6502), .C2(n6510), .A(n6501), .B(n6500), .ZN(U3075)
         );
  INV_X1 U7454 ( .A(n6503), .ZN(n6505) );
  AOI22_X1 U7455 ( .A1(n6557), .A2(n6505), .B1(n6556), .B2(n6504), .ZN(n6509)
         );
  AOI22_X1 U7456 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6507), .B1(n6558), 
        .B2(n6506), .ZN(n6508) );
  OAI211_X1 U7457 ( .C1(n6561), .C2(n6510), .A(n6509), .B(n6508), .ZN(U3081)
         );
  NOR2_X1 U7458 ( .A1(n6511), .A2(n6594), .ZN(n6568) );
  AOI22_X1 U7459 ( .A1(n6571), .A2(n6513), .B1(n6512), .B2(n6568), .ZN(n6528)
         );
  INV_X1 U7460 ( .A(n6514), .ZN(n6517) );
  INV_X1 U7461 ( .A(n6515), .ZN(n6516) );
  OAI21_X1 U7462 ( .B1(n6517), .B2(n6519), .A(n6516), .ZN(n6522) );
  AOI21_X1 U7463 ( .B1(n6518), .B2(n3491), .A(n6568), .ZN(n6524) );
  AOI22_X1 U7464 ( .A1(n6522), .A2(n6524), .B1(n6523), .B2(n6519), .ZN(n6520)
         );
  NAND2_X1 U7465 ( .A1(n6521), .A2(n6520), .ZN(n6574) );
  INV_X1 U7466 ( .A(n6522), .ZN(n6525) );
  OAI22_X1 U7467 ( .A1(n6525), .A2(n6524), .B1(n6523), .B2(n4969), .ZN(n6572)
         );
  AOI22_X1 U7468 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6574), .B1(n6526), 
        .B2(n6572), .ZN(n6527) );
  OAI211_X1 U7469 ( .C1(n6529), .C2(n6577), .A(n6528), .B(n6527), .ZN(U3108)
         );
  AOI22_X1 U7470 ( .A1(n6571), .A2(n6531), .B1(n6530), .B2(n6568), .ZN(n6534)
         );
  AOI22_X1 U7471 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6574), .B1(n6532), 
        .B2(n6572), .ZN(n6533) );
  OAI211_X1 U7472 ( .C1(n6535), .C2(n6577), .A(n6534), .B(n6533), .ZN(U3109)
         );
  AOI22_X1 U7473 ( .A1(n6538), .A2(n6537), .B1(n6536), .B2(n6568), .ZN(n6541)
         );
  AOI22_X1 U7474 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6574), .B1(n6539), 
        .B2(n6572), .ZN(n6540) );
  OAI211_X1 U7475 ( .C1(n6543), .C2(n6542), .A(n6541), .B(n6540), .ZN(U3110)
         );
  AOI22_X1 U7476 ( .A1(n6571), .A2(n6545), .B1(n6544), .B2(n6568), .ZN(n6548)
         );
  AOI22_X1 U7477 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6574), .B1(n6546), 
        .B2(n6572), .ZN(n6547) );
  OAI211_X1 U7478 ( .C1(n6549), .C2(n6577), .A(n6548), .B(n6547), .ZN(U3111)
         );
  AOI22_X1 U7479 ( .A1(n6571), .A2(n6551), .B1(n6550), .B2(n6568), .ZN(n6554)
         );
  AOI22_X1 U7480 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6574), .B1(n6552), 
        .B2(n6572), .ZN(n6553) );
  OAI211_X1 U7481 ( .C1(n6555), .C2(n6577), .A(n6554), .B(n6553), .ZN(U3112)
         );
  AOI22_X1 U7482 ( .A1(n6571), .A2(n6557), .B1(n6556), .B2(n6568), .ZN(n6560)
         );
  AOI22_X1 U7483 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6574), .B1(n6558), 
        .B2(n6572), .ZN(n6559) );
  OAI211_X1 U7484 ( .C1(n6561), .C2(n6577), .A(n6560), .B(n6559), .ZN(U3113)
         );
  AOI22_X1 U7485 ( .A1(n6571), .A2(n6563), .B1(n6562), .B2(n6568), .ZN(n6566)
         );
  AOI22_X1 U7486 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6574), .B1(n6564), 
        .B2(n6572), .ZN(n6565) );
  OAI211_X1 U7487 ( .C1(n6567), .C2(n6577), .A(n6566), .B(n6565), .ZN(U3114)
         );
  AOI22_X1 U7488 ( .A1(n6571), .A2(n6570), .B1(n6569), .B2(n6568), .ZN(n6576)
         );
  AOI22_X1 U7489 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6574), .B1(n6573), 
        .B2(n6572), .ZN(n6575) );
  OAI211_X1 U7490 ( .C1(n6578), .C2(n6577), .A(n6576), .B(n6575), .ZN(U3115)
         );
  AOI211_X1 U7491 ( .C1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n6581), .A(n6580), .B(n6579), .ZN(n6588) );
  INV_X1 U7492 ( .A(n6588), .ZN(n6585) );
  INV_X1 U7493 ( .A(n6582), .ZN(n6584) );
  OAI211_X1 U7494 ( .C1(n6586), .C2(n6585), .A(n6584), .B(n6583), .ZN(n6587)
         );
  OAI21_X1 U7495 ( .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n6588), .A(n6587), 
        .ZN(n6589) );
  AOI222_X1 U7496 ( .A1(n6591), .A2(n6590), .B1(n6591), .B2(n6589), .C1(n6590), 
        .C2(n6589), .ZN(n6596) );
  INV_X1 U7497 ( .A(n6596), .ZN(n6593) );
  AOI21_X1 U7498 ( .B1(n6594), .B2(n6593), .A(n6592), .ZN(n6595) );
  AOI211_X1 U7499 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6596), .A(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B(n6595), .ZN(n6605) );
  INV_X1 U7500 ( .A(n6597), .ZN(n6600) );
  OAI21_X1 U7501 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6598), 
        .ZN(n6599) );
  NAND4_X1 U7502 ( .A1(n6602), .A2(n6601), .A3(n6600), .A4(n6599), .ZN(n6603)
         );
  NOR3_X1 U7503 ( .A1(n6605), .A2(n6604), .A3(n6603), .ZN(n6618) );
  INV_X1 U7504 ( .A(n6618), .ZN(n6607) );
  OAI22_X1 U7505 ( .A1(n6607), .A2(n6620), .B1(n7066), .B2(n6606), .ZN(n6608)
         );
  OAI21_X1 U7506 ( .B1(n6610), .B2(n6609), .A(n6608), .ZN(n6682) );
  OAI21_X1 U7507 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n7066), .A(n6682), .ZN(
        n6619) );
  AOI221_X1 U7508 ( .B1(n6612), .B2(STATE2_REG_0__SCAN_IN), .C1(n6619), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6611), .ZN(n6617) );
  OAI211_X1 U7509 ( .C1(n6615), .C2(n6614), .A(n6613), .B(n6682), .ZN(n6616)
         );
  OAI211_X1 U7510 ( .C1(n6618), .C2(n6620), .A(n6617), .B(n6616), .ZN(U3148)
         );
  NAND3_X1 U7511 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6626), .A3(n6619), .ZN(
        n6625) );
  OAI21_X1 U7512 ( .B1(READY_N), .B2(n6621), .A(n6620), .ZN(n6623) );
  AOI21_X1 U7513 ( .B1(n6623), .B2(n6682), .A(n6622), .ZN(n6624) );
  NAND2_X1 U7514 ( .A1(n6625), .A2(n6624), .ZN(U3149) );
  OAI211_X1 U7515 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n7066), .A(n6680), .B(
        n6626), .ZN(n6628) );
  OAI21_X1 U7516 ( .B1(n6694), .B2(n6628), .A(n6627), .ZN(U3150) );
  AND2_X1 U7517 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6629), .ZN(U3151) );
  AND2_X1 U7518 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6629), .ZN(U3152) );
  AND2_X1 U7519 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6629), .ZN(U3153) );
  AND2_X1 U7520 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6629), .ZN(U3154) );
  AND2_X1 U7521 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6629), .ZN(U3155) );
  AND2_X1 U7522 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6629), .ZN(U3156) );
  AND2_X1 U7523 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6629), .ZN(U3157) );
  AND2_X1 U7524 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6629), .ZN(U3158) );
  INV_X1 U7525 ( .A(DATAWIDTH_REG_23__SCAN_IN), .ZN(n6934) );
  NOR2_X1 U7526 ( .A1(n6679), .A2(n6934), .ZN(U3159) );
  AND2_X1 U7527 ( .A1(n6629), .A2(DATAWIDTH_REG_22__SCAN_IN), .ZN(U3160) );
  INV_X1 U7528 ( .A(DATAWIDTH_REG_21__SCAN_IN), .ZN(n6852) );
  NOR2_X1 U7529 ( .A1(n6679), .A2(n6852), .ZN(U3161) );
  AND2_X1 U7530 ( .A1(n6629), .A2(DATAWIDTH_REG_20__SCAN_IN), .ZN(U3162) );
  AND2_X1 U7531 ( .A1(n6629), .A2(DATAWIDTH_REG_19__SCAN_IN), .ZN(U3163) );
  INV_X1 U7532 ( .A(DATAWIDTH_REG_18__SCAN_IN), .ZN(n6944) );
  NOR2_X1 U7533 ( .A1(n6679), .A2(n6944), .ZN(U3164) );
  INV_X1 U7534 ( .A(DATAWIDTH_REG_17__SCAN_IN), .ZN(n6903) );
  NOR2_X1 U7535 ( .A1(n6679), .A2(n6903), .ZN(U3165) );
  INV_X1 U7536 ( .A(DATAWIDTH_REG_16__SCAN_IN), .ZN(n6774) );
  NOR2_X1 U7537 ( .A1(n6679), .A2(n6774), .ZN(U3166) );
  INV_X1 U7538 ( .A(DATAWIDTH_REG_15__SCAN_IN), .ZN(n6844) );
  NOR2_X1 U7539 ( .A1(n6679), .A2(n6844), .ZN(U3167) );
  INV_X1 U7540 ( .A(DATAWIDTH_REG_14__SCAN_IN), .ZN(n7047) );
  NOR2_X1 U7541 ( .A1(n6679), .A2(n7047), .ZN(U3168) );
  AND2_X1 U7542 ( .A1(n6629), .A2(DATAWIDTH_REG_13__SCAN_IN), .ZN(U3169) );
  AND2_X1 U7543 ( .A1(n6629), .A2(DATAWIDTH_REG_12__SCAN_IN), .ZN(U3170) );
  INV_X1 U7544 ( .A(DATAWIDTH_REG_11__SCAN_IN), .ZN(n6857) );
  NOR2_X1 U7545 ( .A1(n6679), .A2(n6857), .ZN(U3171) );
  AND2_X1 U7546 ( .A1(n6629), .A2(DATAWIDTH_REG_10__SCAN_IN), .ZN(U3172) );
  AND2_X1 U7547 ( .A1(n6629), .A2(DATAWIDTH_REG_9__SCAN_IN), .ZN(U3173) );
  INV_X1 U7548 ( .A(DATAWIDTH_REG_8__SCAN_IN), .ZN(n6856) );
  NOR2_X1 U7549 ( .A1(n6679), .A2(n6856), .ZN(U3174) );
  AND2_X1 U7550 ( .A1(n6629), .A2(DATAWIDTH_REG_7__SCAN_IN), .ZN(U3175) );
  INV_X1 U7551 ( .A(DATAWIDTH_REG_6__SCAN_IN), .ZN(n6807) );
  NOR2_X1 U7552 ( .A1(n6679), .A2(n6807), .ZN(U3176) );
  INV_X1 U7553 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n6800) );
  NOR2_X1 U7554 ( .A1(n6679), .A2(n6800), .ZN(U3177) );
  INV_X1 U7555 ( .A(DATAWIDTH_REG_4__SCAN_IN), .ZN(n6806) );
  NOR2_X1 U7556 ( .A1(n6679), .A2(n6806), .ZN(U3178) );
  INV_X1 U7557 ( .A(DATAWIDTH_REG_3__SCAN_IN), .ZN(n7014) );
  NOR2_X1 U7558 ( .A1(n6679), .A2(n7014), .ZN(U3179) );
  AND2_X1 U7559 ( .A1(n6629), .A2(DATAWIDTH_REG_2__SCAN_IN), .ZN(U3180) );
  NAND2_X1 U7560 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6634) );
  NAND2_X1 U7561 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6635) );
  NAND2_X1 U7562 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .ZN(n6641) );
  NAND2_X1 U7563 ( .A1(n6635), .A2(n6641), .ZN(n6631) );
  INV_X1 U7564 ( .A(NA_N), .ZN(n6630) );
  AOI221_X1 U7565 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6630), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6645) );
  AOI21_X1 U7566 ( .B1(n6632), .B2(n6631), .A(n6645), .ZN(n6633) );
  OAI221_X1 U7567 ( .B1(n7094), .B2(REQUESTPENDING_REG_SCAN_IN), .C1(n7094), 
        .C2(n6634), .A(n6633), .ZN(U3181) );
  INV_X1 U7568 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6642) );
  NOR2_X1 U7569 ( .A1(n6961), .A2(n6642), .ZN(n6637) );
  INV_X1 U7570 ( .A(n6634), .ZN(n6636) );
  OAI21_X1 U7571 ( .B1(n6637), .B2(n6636), .A(n6635), .ZN(n6638) );
  NAND3_X1 U7572 ( .A1(n6639), .A2(n6641), .A3(n6638), .ZN(U3182) );
  AOI221_X1 U7573 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n7066), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6640) );
  AOI221_X1 U7574 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6640), .C2(HOLD), .A(n6961), .ZN(n6646) );
  OR4_X1 U7575 ( .A1(n6642), .A2(n6961), .A3(n6641), .A4(NA_N), .ZN(n6644) );
  NAND3_X1 U7576 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .A3(
        STATE_REG_2__SCAN_IN), .ZN(n6643) );
  OAI211_X1 U7577 ( .C1(n6646), .C2(n6645), .A(n6644), .B(n6643), .ZN(U3183)
         );
  NAND2_X1 U7578 ( .A1(n7094), .A2(n6936), .ZN(n6663) );
  INV_X1 U7579 ( .A(ADDRESS_REG_0__SCAN_IN), .ZN(n6992) );
  OAI222_X1 U7580 ( .A1(n6663), .A2(n6647), .B1(n6992), .B2(n7094), .C1(n6684), 
        .C2(n6671), .ZN(U3184) );
  INV_X1 U7581 ( .A(ADDRESS_REG_1__SCAN_IN), .ZN(n6914) );
  CLKBUF_X1 U7582 ( .A(n6663), .Z(n6674) );
  OAI222_X1 U7583 ( .A1(n6671), .A2(n6647), .B1(n6914), .B2(n7094), .C1(n6648), 
        .C2(n6674), .ZN(U3185) );
  INV_X1 U7584 ( .A(ADDRESS_REG_2__SCAN_IN), .ZN(n7033) );
  OAI222_X1 U7585 ( .A1(n6671), .A2(n6648), .B1(n7033), .B2(n7094), .C1(n6649), 
        .C2(n6674), .ZN(U3186) );
  INV_X1 U7586 ( .A(ADDRESS_REG_3__SCAN_IN), .ZN(n7065) );
  OAI222_X1 U7587 ( .A1(n6671), .A2(n6649), .B1(n7065), .B2(n7094), .C1(n6651), 
        .C2(n6663), .ZN(U3187) );
  INV_X1 U7588 ( .A(ADDRESS_REG_4__SCAN_IN), .ZN(n6650) );
  OAI222_X1 U7589 ( .A1(n6671), .A2(n6651), .B1(n6650), .B2(n7094), .C1(n6652), 
        .C2(n6674), .ZN(U3188) );
  INV_X1 U7590 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n7046) );
  OAI222_X1 U7591 ( .A1(n6671), .A2(n6652), .B1(n7046), .B2(n7094), .C1(n6654), 
        .C2(n6674), .ZN(U3189) );
  INV_X1 U7592 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n6653) );
  OAI222_X1 U7593 ( .A1(n6671), .A2(n6654), .B1(n6653), .B2(n7094), .C1(n6656), 
        .C2(n6663), .ZN(U3190) );
  INV_X1 U7594 ( .A(ADDRESS_REG_7__SCAN_IN), .ZN(n6655) );
  OAI222_X1 U7595 ( .A1(n6671), .A2(n6656), .B1(n6655), .B2(n7094), .C1(n6657), 
        .C2(n6674), .ZN(U3191) );
  INV_X1 U7596 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n7052) );
  OAI222_X1 U7597 ( .A1(n6671), .A2(n6657), .B1(n7052), .B2(n7094), .C1(n6659), 
        .C2(n6663), .ZN(U3192) );
  INV_X1 U7598 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n6658) );
  OAI222_X1 U7599 ( .A1(n6671), .A2(n6659), .B1(n6658), .B2(n7094), .C1(n6660), 
        .C2(n6663), .ZN(U3193) );
  INV_X1 U7600 ( .A(ADDRESS_REG_10__SCAN_IN), .ZN(n6929) );
  OAI222_X1 U7601 ( .A1(n6663), .A2(n6661), .B1(n6929), .B2(n7094), .C1(n6660), 
        .C2(n6671), .ZN(U3194) );
  INV_X1 U7602 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n6809) );
  OAI222_X1 U7603 ( .A1(n6671), .A2(n6661), .B1(n6809), .B2(n7094), .C1(n6662), 
        .C2(n6663), .ZN(U3195) );
  INV_X1 U7604 ( .A(ADDRESS_REG_12__SCAN_IN), .ZN(n7030) );
  OAI222_X1 U7605 ( .A1(n6671), .A2(n6662), .B1(n7030), .B2(n7094), .C1(n5759), 
        .C2(n6663), .ZN(U3196) );
  INV_X1 U7606 ( .A(ADDRESS_REG_13__SCAN_IN), .ZN(n6781) );
  OAI222_X1 U7607 ( .A1(n6663), .A2(n6665), .B1(n6781), .B2(n7094), .C1(n5759), 
        .C2(n6671), .ZN(U3197) );
  INV_X1 U7608 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n6664) );
  OAI222_X1 U7609 ( .A1(n6671), .A2(n6665), .B1(n6664), .B2(n7094), .C1(n7036), 
        .C2(n6663), .ZN(U3198) );
  INV_X1 U7610 ( .A(ADDRESS_REG_15__SCAN_IN), .ZN(n6666) );
  OAI222_X1 U7611 ( .A1(n6671), .A2(n7036), .B1(n6666), .B2(n7094), .C1(n6916), 
        .C2(n6674), .ZN(U3199) );
  INV_X1 U7612 ( .A(ADDRESS_REG_16__SCAN_IN), .ZN(n6783) );
  OAI222_X1 U7613 ( .A1(n6674), .A2(n5883), .B1(n6783), .B2(n7094), .C1(n6916), 
        .C2(n6671), .ZN(U3200) );
  INV_X1 U7614 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n7060) );
  INV_X1 U7615 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6667) );
  OAI222_X1 U7616 ( .A1(n6671), .A2(n5883), .B1(n7060), .B2(n7094), .C1(n6667), 
        .C2(n6674), .ZN(U3201) );
  INV_X1 U7617 ( .A(ADDRESS_REG_18__SCAN_IN), .ZN(n6835) );
  OAI222_X1 U7618 ( .A1(n6671), .A2(n6667), .B1(n6835), .B2(n7094), .C1(n7018), 
        .C2(n6674), .ZN(U3202) );
  INV_X1 U7619 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n6668) );
  OAI222_X1 U7620 ( .A1(n6671), .A2(n7018), .B1(n6668), .B2(n7094), .C1(n7024), 
        .C2(n6674), .ZN(U3203) );
  INV_X1 U7621 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n6930) );
  OAI222_X1 U7622 ( .A1(n6671), .A2(n7024), .B1(n6930), .B2(n7094), .C1(n6913), 
        .C2(n6674), .ZN(U3204) );
  INV_X1 U7623 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n6669) );
  INV_X1 U7624 ( .A(REIP_REG_23__SCAN_IN), .ZN(n7015) );
  OAI222_X1 U7625 ( .A1(n6671), .A2(n6913), .B1(n6669), .B2(n7094), .C1(n7015), 
        .C2(n6674), .ZN(U3205) );
  INV_X1 U7626 ( .A(ADDRESS_REG_22__SCAN_IN), .ZN(n7037) );
  OAI222_X1 U7627 ( .A1(n6671), .A2(n7015), .B1(n7037), .B2(n7094), .C1(n6922), 
        .C2(n6674), .ZN(U3206) );
  INV_X1 U7628 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n7049) );
  OAI222_X1 U7629 ( .A1(n6674), .A2(n6920), .B1(n7049), .B2(n7094), .C1(n6922), 
        .C2(n6671), .ZN(U3207) );
  INV_X1 U7630 ( .A(ADDRESS_REG_24__SCAN_IN), .ZN(n6670) );
  OAI222_X1 U7631 ( .A1(n6671), .A2(n6920), .B1(n6670), .B2(n7094), .C1(n6947), 
        .C2(n6674), .ZN(U3208) );
  INV_X1 U7632 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n7053) );
  OAI222_X1 U7633 ( .A1(n6671), .A2(n6947), .B1(n7053), .B2(n7094), .C1(n6673), 
        .C2(n6674), .ZN(U3209) );
  INV_X1 U7634 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n6672) );
  INV_X1 U7635 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6780) );
  OAI222_X1 U7636 ( .A1(n6671), .A2(n6673), .B1(n6672), .B2(n7094), .C1(n6780), 
        .C2(n6674), .ZN(U3210) );
  INV_X1 U7637 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n6799) );
  OAI222_X1 U7638 ( .A1(n6671), .A2(n6780), .B1(n6799), .B2(n7094), .C1(n6946), 
        .C2(n6674), .ZN(U3211) );
  INV_X1 U7639 ( .A(ADDRESS_REG_28__SCAN_IN), .ZN(n6794) );
  OAI222_X1 U7640 ( .A1(n6671), .A2(n6946), .B1(n6794), .B2(n7094), .C1(n6900), 
        .C2(n6674), .ZN(U3212) );
  INV_X1 U7641 ( .A(REIP_REG_31__SCAN_IN), .ZN(n7062) );
  INV_X1 U7642 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n6902) );
  OAI222_X1 U7643 ( .A1(n6674), .A2(n7062), .B1(n6902), .B2(n7094), .C1(n6900), 
        .C2(n6671), .ZN(U3213) );
  INV_X1 U7644 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6932) );
  INV_X1 U7645 ( .A(BE_N_REG_2__SCAN_IN), .ZN(n6833) );
  AOI22_X1 U7646 ( .A1(n7094), .A2(n6932), .B1(n6833), .B2(n7093), .ZN(U3446)
         );
  INV_X1 U7647 ( .A(BE_N_REG_1__SCAN_IN), .ZN(n6825) );
  AOI22_X1 U7648 ( .A1(n7094), .A2(n6675), .B1(n6825), .B2(n7093), .ZN(U3447)
         );
  OAI22_X1 U7649 ( .A1(n7093), .A2(BYTEENABLE_REG_0__SCAN_IN), .B1(
        BE_N_REG_0__SCAN_IN), .B2(n7094), .ZN(n6676) );
  INV_X1 U7650 ( .A(n6676), .ZN(U3448) );
  OAI21_X1 U7651 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6679), .A(n6678), .ZN(
        n6677) );
  INV_X1 U7652 ( .A(n6677), .ZN(U3451) );
  OAI21_X1 U7653 ( .B1(n6679), .B2(n6831), .A(n6678), .ZN(U3452) );
  OAI211_X1 U7654 ( .C1(n6683), .C2(n6682), .A(n6681), .B(n6680), .ZN(U3453)
         );
  AOI21_X1 U7655 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6685) );
  AOI22_X1 U7656 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6685), .B2(n6684), .ZN(n6687) );
  AOI22_X1 U7657 ( .A1(n6689), .A2(n6687), .B1(n6932), .B2(n6686), .ZN(U3468)
         );
  INV_X1 U7658 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6959) );
  OAI21_X1 U7659 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6689), .ZN(n6688) );
  OAI21_X1 U7660 ( .B1(n6689), .B2(n6959), .A(n6688), .ZN(U3469) );
  INV_X1 U7661 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6964) );
  AOI22_X1 U7662 ( .A1(n7094), .A2(READREQUEST_REG_SCAN_IN), .B1(n6964), .B2(
        n7093), .ZN(U3470) );
  AOI211_X1 U7663 ( .C1(n6267), .C2(n7066), .A(n6691), .B(n6690), .ZN(n6698)
         );
  OAI211_X1 U7664 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6693), .A(n6692), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6695) );
  AOI21_X1 U7665 ( .B1(n6695), .B2(STATE2_REG_0__SCAN_IN), .A(n6694), .ZN(
        n6697) );
  NAND2_X1 U7666 ( .A1(n6698), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6696) );
  OAI21_X1 U7667 ( .B1(n6698), .B2(n6697), .A(n6696), .ZN(U3472) );
  INV_X1 U7668 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n7069) );
  INV_X1 U7669 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n6943) );
  AOI22_X1 U7670 ( .A1(n7094), .A2(n7069), .B1(n6943), .B2(n7093), .ZN(U3473)
         );
  OAI22_X1 U7671 ( .A1(STATE_REG_0__SCAN_IN), .A2(keyinput_g103), .B1(
        DATAI_17_), .B2(keyinput_g14), .ZN(n6699) );
  AOI221_X1 U7672 ( .B1(STATE_REG_0__SCAN_IN), .B2(keyinput_g103), .C1(
        keyinput_g14), .C2(DATAI_17_), .A(n6699), .ZN(n6706) );
  OAI22_X1 U7673 ( .A1(READREQUEST_REG_SCAN_IN), .A2(keyinput_g37), .B1(
        keyinput_g126), .B2(DATAWIDTH_REG_22__SCAN_IN), .ZN(n6700) );
  AOI221_X1 U7674 ( .B1(READREQUEST_REG_SCAN_IN), .B2(keyinput_g37), .C1(
        DATAWIDTH_REG_22__SCAN_IN), .C2(keyinput_g126), .A(n6700), .ZN(n6705)
         );
  OAI22_X1 U7675 ( .A1(REIP_REG_29__SCAN_IN), .A2(keyinput_g53), .B1(DATAI_11_), .B2(keyinput_g20), .ZN(n6701) );
  AOI221_X1 U7676 ( .B1(REIP_REG_29__SCAN_IN), .B2(keyinput_g53), .C1(
        keyinput_g20), .C2(DATAI_11_), .A(n6701), .ZN(n6704) );
  OAI22_X1 U7677 ( .A1(REIP_REG_26__SCAN_IN), .A2(keyinput_g56), .B1(
        keyinput_g96), .B2(ADDRESS_REG_4__SCAN_IN), .ZN(n6702) );
  AOI221_X1 U7678 ( .B1(REIP_REG_26__SCAN_IN), .B2(keyinput_g56), .C1(
        ADDRESS_REG_4__SCAN_IN), .C2(keyinput_g96), .A(n6702), .ZN(n6703) );
  NAND4_X1 U7679 ( .A1(n6706), .A2(n6705), .A3(n6704), .A4(n6703), .ZN(n6734)
         );
  OAI22_X1 U7680 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(keyinput_g121), .B1(
        DATAWIDTH_REG_14__SCAN_IN), .B2(keyinput_g118), .ZN(n6707) );
  AOI221_X1 U7681 ( .B1(DATAWIDTH_REG_17__SCAN_IN), .B2(keyinput_g121), .C1(
        keyinput_g118), .C2(DATAWIDTH_REG_14__SCAN_IN), .A(n6707), .ZN(n6714)
         );
  OAI22_X1 U7682 ( .A1(ADDRESS_REG_0__SCAN_IN), .A2(keyinput_g100), .B1(
        keyinput_g76), .B2(ADDRESS_REG_24__SCAN_IN), .ZN(n6708) );
  AOI221_X1 U7683 ( .B1(ADDRESS_REG_0__SCAN_IN), .B2(keyinput_g100), .C1(
        ADDRESS_REG_24__SCAN_IN), .C2(keyinput_g76), .A(n6708), .ZN(n6713) );
  OAI22_X1 U7684 ( .A1(DATAI_19_), .A2(keyinput_g12), .B1(keyinput_g111), .B2(
        DATAWIDTH_REG_7__SCAN_IN), .ZN(n6709) );
  AOI221_X1 U7685 ( .B1(DATAI_19_), .B2(keyinput_g12), .C1(
        DATAWIDTH_REG_7__SCAN_IN), .C2(keyinput_g111), .A(n6709), .ZN(n6712)
         );
  OAI22_X1 U7686 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(keyinput_g104), .B1(
        keyinput_g117), .B2(DATAWIDTH_REG_13__SCAN_IN), .ZN(n6710) );
  AOI221_X1 U7687 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(keyinput_g104), .C1(
        DATAWIDTH_REG_13__SCAN_IN), .C2(keyinput_g117), .A(n6710), .ZN(n6711)
         );
  NAND4_X1 U7688 ( .A1(n6714), .A2(n6713), .A3(n6712), .A4(n6711), .ZN(n6733)
         );
  OAI22_X1 U7689 ( .A1(DATAI_22_), .A2(keyinput_g9), .B1(
        DATAWIDTH_REG_10__SCAN_IN), .B2(keyinput_g114), .ZN(n6715) );
  AOI221_X1 U7690 ( .B1(DATAI_22_), .B2(keyinput_g9), .C1(keyinput_g114), .C2(
        DATAWIDTH_REG_10__SCAN_IN), .A(n6715), .ZN(n6722) );
  OAI22_X1 U7691 ( .A1(REIP_REG_27__SCAN_IN), .A2(keyinput_g55), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(keyinput_g75), .ZN(n6716) );
  AOI221_X1 U7692 ( .B1(REIP_REG_27__SCAN_IN), .B2(keyinput_g55), .C1(
        keyinput_g75), .C2(ADDRESS_REG_25__SCAN_IN), .A(n6716), .ZN(n6721) );
  OAI22_X1 U7693 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(keyinput_g113), .B1(
        ADS_N_REG_SCAN_IN), .B2(keyinput_g38), .ZN(n6717) );
  AOI221_X1 U7694 ( .B1(DATAWIDTH_REG_9__SCAN_IN), .B2(keyinput_g113), .C1(
        keyinput_g38), .C2(ADS_N_REG_SCAN_IN), .A(n6717), .ZN(n6720) );
  OAI22_X1 U7695 ( .A1(DATAI_1_), .A2(keyinput_g30), .B1(
        DATAWIDTH_REG_19__SCAN_IN), .B2(keyinput_g123), .ZN(n6718) );
  AOI221_X1 U7696 ( .B1(DATAI_1_), .B2(keyinput_g30), .C1(keyinput_g123), .C2(
        DATAWIDTH_REG_19__SCAN_IN), .A(n6718), .ZN(n6719) );
  NAND4_X1 U7697 ( .A1(n6722), .A2(n6721), .A3(n6720), .A4(n6719), .ZN(n6732)
         );
  OAI22_X1 U7698 ( .A1(DATAI_28_), .A2(keyinput_g3), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(keyinput_g79), .ZN(n6723) );
  AOI221_X1 U7699 ( .B1(DATAI_28_), .B2(keyinput_g3), .C1(keyinput_g79), .C2(
        ADDRESS_REG_21__SCAN_IN), .A(n6723), .ZN(n6730) );
  OAI22_X1 U7700 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(keyinput_g106), .B1(
        DATAWIDTH_REG_18__SCAN_IN), .B2(keyinput_g122), .ZN(n6724) );
  AOI221_X1 U7701 ( .B1(DATAWIDTH_REG_2__SCAN_IN), .B2(keyinput_g106), .C1(
        keyinput_g122), .C2(DATAWIDTH_REG_18__SCAN_IN), .A(n6724), .ZN(n6729)
         );
  OAI22_X1 U7702 ( .A1(DATAI_20_), .A2(keyinput_g11), .B1(DATAI_18_), .B2(
        keyinput_g13), .ZN(n6725) );
  AOI221_X1 U7703 ( .B1(DATAI_20_), .B2(keyinput_g11), .C1(keyinput_g13), .C2(
        DATAI_18_), .A(n6725), .ZN(n6728) );
  OAI22_X1 U7704 ( .A1(DATAI_16_), .A2(keyinput_g15), .B1(keyinput_g50), .B2(
        BYTEENABLE_REG_3__SCAN_IN), .ZN(n6726) );
  AOI221_X1 U7705 ( .B1(DATAI_16_), .B2(keyinput_g15), .C1(
        BYTEENABLE_REG_3__SCAN_IN), .C2(keyinput_g50), .A(n6726), .ZN(n6727)
         );
  NAND4_X1 U7706 ( .A1(n6730), .A2(n6729), .A3(n6728), .A4(n6727), .ZN(n6731)
         );
  NOR4_X1 U7707 ( .A1(n6734), .A2(n6733), .A3(n6732), .A4(n6731), .ZN(n7092)
         );
  OAI22_X1 U7708 ( .A1(M_IO_N_REG_SCAN_IN), .A2(keyinput_g40), .B1(
        keyinput_g116), .B2(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6735) );
  AOI221_X1 U7709 ( .B1(M_IO_N_REG_SCAN_IN), .B2(keyinput_g40), .C1(
        DATAWIDTH_REG_12__SCAN_IN), .C2(keyinput_g116), .A(n6735), .ZN(n6742)
         );
  OAI22_X1 U7710 ( .A1(ADDRESS_REG_6__SCAN_IN), .A2(keyinput_g94), .B1(
        BE_N_REG_0__SCAN_IN), .B2(keyinput_g70), .ZN(n6736) );
  AOI221_X1 U7711 ( .B1(ADDRESS_REG_6__SCAN_IN), .B2(keyinput_g94), .C1(
        keyinput_g70), .C2(BE_N_REG_0__SCAN_IN), .A(n6736), .ZN(n6741) );
  OAI22_X1 U7712 ( .A1(REIP_REG_25__SCAN_IN), .A2(keyinput_g57), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(keyinput_g93), .ZN(n6737) );
  AOI221_X1 U7713 ( .B1(REIP_REG_25__SCAN_IN), .B2(keyinput_g57), .C1(
        keyinput_g93), .C2(ADDRESS_REG_7__SCAN_IN), .A(n6737), .ZN(n6740) );
  OAI22_X1 U7714 ( .A1(MORE_REG_SCAN_IN), .A2(keyinput_g44), .B1(
        BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_g48), .ZN(n6738) );
  AOI221_X1 U7715 ( .B1(MORE_REG_SCAN_IN), .B2(keyinput_g44), .C1(keyinput_g48), .C2(BYTEENABLE_REG_1__SCAN_IN), .A(n6738), .ZN(n6739) );
  NAND4_X1 U7716 ( .A1(n6742), .A2(n6741), .A3(n6740), .A4(n6739), .ZN(n6870)
         );
  OAI22_X1 U7717 ( .A1(STATE_REG_2__SCAN_IN), .A2(keyinput_g101), .B1(
        keyinput_g25), .B2(DATAI_6_), .ZN(n6743) );
  AOI221_X1 U7718 ( .B1(STATE_REG_2__SCAN_IN), .B2(keyinput_g101), .C1(
        DATAI_6_), .C2(keyinput_g25), .A(n6743), .ZN(n6769) );
  INV_X1 U7719 ( .A(DATAI_24_), .ZN(n6749) );
  OAI22_X1 U7720 ( .A1(W_R_N_REG_SCAN_IN), .A2(keyinput_g46), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(keyinput_g92), .ZN(n6744) );
  AOI221_X1 U7721 ( .B1(W_R_N_REG_SCAN_IN), .B2(keyinput_g46), .C1(
        keyinput_g92), .C2(ADDRESS_REG_8__SCAN_IN), .A(n6744), .ZN(n6747) );
  OAI22_X1 U7722 ( .A1(HOLD), .A2(keyinput_g36), .B1(ADDRESS_REG_19__SCAN_IN), 
        .B2(keyinput_g81), .ZN(n6745) );
  AOI221_X1 U7723 ( .B1(HOLD), .B2(keyinput_g36), .C1(keyinput_g81), .C2(
        ADDRESS_REG_19__SCAN_IN), .A(n6745), .ZN(n6746) );
  OAI211_X1 U7724 ( .C1(n6749), .C2(keyinput_g7), .A(n6747), .B(n6746), .ZN(
        n6748) );
  AOI21_X1 U7725 ( .B1(n6749), .B2(keyinput_g7), .A(n6748), .ZN(n6768) );
  AOI22_X1 U7726 ( .A1(DATAI_9_), .A2(keyinput_g22), .B1(DATAI_31_), .B2(
        keyinput_g0), .ZN(n6750) );
  OAI221_X1 U7727 ( .B1(DATAI_9_), .B2(keyinput_g22), .C1(DATAI_31_), .C2(
        keyinput_g0), .A(n6750), .ZN(n6757) );
  AOI22_X1 U7728 ( .A1(DATAI_15_), .A2(keyinput_g16), .B1(DATAI_3_), .B2(
        keyinput_g28), .ZN(n6751) );
  OAI221_X1 U7729 ( .B1(DATAI_15_), .B2(keyinput_g16), .C1(DATAI_3_), .C2(
        keyinput_g28), .A(n6751), .ZN(n6756) );
  AOI22_X1 U7730 ( .A1(BYTEENABLE_REG_2__SCAN_IN), .A2(keyinput_g49), .B1(
        REIP_REG_21__SCAN_IN), .B2(keyinput_g61), .ZN(n6752) );
  OAI221_X1 U7731 ( .B1(BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_g49), .C1(
        REIP_REG_21__SCAN_IN), .C2(keyinput_g61), .A(n6752), .ZN(n6755) );
  AOI22_X1 U7732 ( .A1(ADDRESS_REG_1__SCAN_IN), .A2(keyinput_g99), .B1(
        DATAWIDTH_REG_20__SCAN_IN), .B2(keyinput_g124), .ZN(n6753) );
  OAI221_X1 U7733 ( .B1(ADDRESS_REG_1__SCAN_IN), .B2(keyinput_g99), .C1(
        DATAWIDTH_REG_20__SCAN_IN), .C2(keyinput_g124), .A(n6753), .ZN(n6754)
         );
  NOR4_X1 U7734 ( .A1(n6757), .A2(n6756), .A3(n6755), .A4(n6754), .ZN(n6767)
         );
  AOI22_X1 U7735 ( .A1(ADDRESS_REG_15__SCAN_IN), .A2(keyinput_g85), .B1(
        DATAI_29_), .B2(keyinput_g2), .ZN(n6758) );
  OAI221_X1 U7736 ( .B1(ADDRESS_REG_15__SCAN_IN), .B2(keyinput_g85), .C1(
        DATAI_29_), .C2(keyinput_g2), .A(n6758), .ZN(n6765) );
  AOI22_X1 U7737 ( .A1(ADDRESS_REG_14__SCAN_IN), .A2(keyinput_g86), .B1(
        MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_g32), .ZN(n6759) );
  OAI221_X1 U7738 ( .B1(ADDRESS_REG_14__SCAN_IN), .B2(keyinput_g86), .C1(
        MEMORYFETCH_REG_SCAN_IN), .C2(keyinput_g32), .A(n6759), .ZN(n6764) );
  AOI22_X1 U7739 ( .A1(ADDRESS_REG_26__SCAN_IN), .A2(keyinput_g74), .B1(
        DATAI_2_), .B2(keyinput_g29), .ZN(n6760) );
  OAI221_X1 U7740 ( .B1(ADDRESS_REG_26__SCAN_IN), .B2(keyinput_g74), .C1(
        DATAI_2_), .C2(keyinput_g29), .A(n6760), .ZN(n6763) );
  AOI22_X1 U7741 ( .A1(BE_N_REG_3__SCAN_IN), .A2(keyinput_g67), .B1(
        REIP_REG_22__SCAN_IN), .B2(keyinput_g60), .ZN(n6761) );
  OAI221_X1 U7742 ( .B1(BE_N_REG_3__SCAN_IN), .B2(keyinput_g67), .C1(
        REIP_REG_22__SCAN_IN), .C2(keyinput_g60), .A(n6761), .ZN(n6762) );
  NOR4_X1 U7743 ( .A1(n6765), .A2(n6764), .A3(n6763), .A4(n6762), .ZN(n6766)
         );
  NAND4_X1 U7744 ( .A1(n6769), .A2(n6768), .A3(n6767), .A4(n6766), .ZN(n6869)
         );
  AOI22_X1 U7745 ( .A1(ADDRESS_REG_9__SCAN_IN), .A2(keyinput_g91), .B1(
        REIP_REG_17__SCAN_IN), .B2(keyinput_g65), .ZN(n6770) );
  OAI221_X1 U7746 ( .B1(ADDRESS_REG_9__SCAN_IN), .B2(keyinput_g91), .C1(
        REIP_REG_17__SCAN_IN), .C2(keyinput_g65), .A(n6770), .ZN(n6778) );
  AOI22_X1 U7747 ( .A1(ADDRESS_REG_29__SCAN_IN), .A2(keyinput_g71), .B1(
        REIP_REG_24__SCAN_IN), .B2(keyinput_g58), .ZN(n6771) );
  OAI221_X1 U7748 ( .B1(ADDRESS_REG_29__SCAN_IN), .B2(keyinput_g71), .C1(
        REIP_REG_24__SCAN_IN), .C2(keyinput_g58), .A(n6771), .ZN(n6777) );
  AOI22_X1 U7749 ( .A1(NA_N), .A2(keyinput_g33), .B1(REIP_REG_19__SCAN_IN), 
        .B2(keyinput_g63), .ZN(n6772) );
  OAI221_X1 U7750 ( .B1(NA_N), .B2(keyinput_g33), .C1(REIP_REG_19__SCAN_IN), 
        .C2(keyinput_g63), .A(n6772), .ZN(n6776) );
  AOI22_X1 U7751 ( .A1(n6897), .A2(keyinput_g31), .B1(keyinput_g120), .B2(
        n6774), .ZN(n6773) );
  OAI221_X1 U7752 ( .B1(n6897), .B2(keyinput_g31), .C1(n6774), .C2(
        keyinput_g120), .A(n6773), .ZN(n6775) );
  NOR4_X1 U7753 ( .A1(n6778), .A2(n6777), .A3(n6776), .A4(n6775), .ZN(n6819)
         );
  AOI22_X1 U7754 ( .A1(n6781), .A2(keyinput_g87), .B1(n6780), .B2(keyinput_g54), .ZN(n6779) );
  OAI221_X1 U7755 ( .B1(n6781), .B2(keyinput_g87), .C1(n6780), .C2(
        keyinput_g54), .A(n6779), .ZN(n6791) );
  INV_X1 U7756 ( .A(BS16_N), .ZN(n6784) );
  AOI22_X1 U7757 ( .A1(n6784), .A2(keyinput_g34), .B1(n6783), .B2(keyinput_g84), .ZN(n6782) );
  OAI221_X1 U7758 ( .B1(n6784), .B2(keyinput_g34), .C1(n6783), .C2(
        keyinput_g84), .A(n6782), .ZN(n6790) );
  AOI22_X1 U7759 ( .A1(n6786), .A2(keyinput_g43), .B1(keyinput_g78), .B2(n7037), .ZN(n6785) );
  OAI221_X1 U7760 ( .B1(n6786), .B2(keyinput_g43), .C1(n7037), .C2(
        keyinput_g78), .A(n6785), .ZN(n6789) );
  AOI22_X1 U7761 ( .A1(n7014), .A2(keyinput_g107), .B1(n7033), .B2(
        keyinput_g98), .ZN(n6787) );
  OAI221_X1 U7762 ( .B1(n7014), .B2(keyinput_g107), .C1(n7033), .C2(
        keyinput_g98), .A(n6787), .ZN(n6788) );
  NOR4_X1 U7763 ( .A1(n6791), .A2(n6790), .A3(n6789), .A4(n6788), .ZN(n6818)
         );
  INV_X1 U7764 ( .A(DATAI_30_), .ZN(n6793) );
  AOI22_X1 U7765 ( .A1(n6794), .A2(keyinput_g72), .B1(n6793), .B2(keyinput_g1), 
        .ZN(n6792) );
  OAI221_X1 U7766 ( .B1(n6794), .B2(keyinput_g72), .C1(n6793), .C2(keyinput_g1), .A(n6792), .ZN(n6804) );
  INV_X1 U7767 ( .A(DATAI_27_), .ZN(n6796) );
  AOI22_X1 U7768 ( .A1(n6796), .A2(keyinput_g4), .B1(n5883), .B2(keyinput_g64), 
        .ZN(n6795) );
  OAI221_X1 U7769 ( .B1(n6796), .B2(keyinput_g4), .C1(n5883), .C2(keyinput_g64), .A(n6795), .ZN(n6803) );
  INV_X1 U7770 ( .A(DATAI_25_), .ZN(n7023) );
  AOI22_X1 U7771 ( .A1(n6950), .A2(keyinput_g24), .B1(n7023), .B2(keyinput_g6), 
        .ZN(n6797) );
  OAI221_X1 U7772 ( .B1(n6950), .B2(keyinput_g24), .C1(n7023), .C2(keyinput_g6), .A(n6797), .ZN(n6802) );
  AOI22_X1 U7773 ( .A1(n6800), .A2(keyinput_g109), .B1(keyinput_g73), .B2(
        n6799), .ZN(n6798) );
  OAI221_X1 U7774 ( .B1(n6800), .B2(keyinput_g109), .C1(n6799), .C2(
        keyinput_g73), .A(n6798), .ZN(n6801) );
  NOR4_X1 U7775 ( .A1(n6804), .A2(n6803), .A3(n6802), .A4(n6801), .ZN(n6817)
         );
  AOI22_X1 U7776 ( .A1(n6807), .A2(keyinput_g110), .B1(keyinput_g108), .B2(
        n6806), .ZN(n6805) );
  OAI221_X1 U7777 ( .B1(n6807), .B2(keyinput_g110), .C1(n6806), .C2(
        keyinput_g108), .A(n6805), .ZN(n6815) );
  AOI22_X1 U7778 ( .A1(n7066), .A2(keyinput_g35), .B1(keyinput_g89), .B2(n6809), .ZN(n6808) );
  OAI221_X1 U7779 ( .B1(n7066), .B2(keyinput_g35), .C1(n6809), .C2(
        keyinput_g89), .A(n6808), .ZN(n6814) );
  INV_X1 U7780 ( .A(STATE_REG_1__SCAN_IN), .ZN(n7021) );
  AOI22_X1 U7781 ( .A1(n7021), .A2(keyinput_g102), .B1(keyinput_g23), .B2(
        n7050), .ZN(n6810) );
  OAI221_X1 U7782 ( .B1(n7021), .B2(keyinput_g102), .C1(n7050), .C2(
        keyinput_g23), .A(n6810), .ZN(n6813) );
  AOI22_X1 U7783 ( .A1(n7030), .A2(keyinput_g88), .B1(n6929), .B2(keyinput_g90), .ZN(n6811) );
  OAI221_X1 U7784 ( .B1(n7030), .B2(keyinput_g88), .C1(n6929), .C2(
        keyinput_g90), .A(n6811), .ZN(n6812) );
  NOR4_X1 U7785 ( .A1(n6815), .A2(n6814), .A3(n6813), .A4(n6812), .ZN(n6816)
         );
  NAND4_X1 U7786 ( .A1(n6819), .A2(n6818), .A3(n6817), .A4(n6816), .ZN(n6868)
         );
  AOI22_X1 U7787 ( .A1(n6900), .A2(keyinput_g52), .B1(keyinput_g83), .B2(n7060), .ZN(n6820) );
  OAI221_X1 U7788 ( .B1(n6900), .B2(keyinput_g52), .C1(n7060), .C2(
        keyinput_g83), .A(n6820), .ZN(n6829) );
  AOI22_X1 U7789 ( .A1(n7063), .A2(keyinput_g45), .B1(n6941), .B2(keyinput_g26), .ZN(n6821) );
  OAI221_X1 U7790 ( .B1(n7063), .B2(keyinput_g45), .C1(n6941), .C2(
        keyinput_g26), .A(n6821), .ZN(n6828) );
  INV_X1 U7791 ( .A(DATAI_21_), .ZN(n6823) );
  AOI22_X1 U7792 ( .A1(n6823), .A2(keyinput_g10), .B1(n7039), .B2(keyinput_g21), .ZN(n6822) );
  OAI221_X1 U7793 ( .B1(n6823), .B2(keyinput_g10), .C1(n7039), .C2(
        keyinput_g21), .A(n6822), .ZN(n6827) );
  AOI22_X1 U7794 ( .A1(n6958), .A2(keyinput_g41), .B1(n6825), .B2(keyinput_g69), .ZN(n6824) );
  OAI221_X1 U7795 ( .B1(n6958), .B2(keyinput_g41), .C1(n6825), .C2(
        keyinput_g69), .A(n6824), .ZN(n6826) );
  NOR4_X1 U7796 ( .A1(n6829), .A2(n6828), .A3(n6827), .A4(n6826), .ZN(n6866)
         );
  AOI22_X1 U7797 ( .A1(n6831), .A2(keyinput_g105), .B1(n6965), .B2(keyinput_g5), .ZN(n6830) );
  OAI221_X1 U7798 ( .B1(n6831), .B2(keyinput_g105), .C1(n6965), .C2(
        keyinput_g5), .A(n6830), .ZN(n6840) );
  INV_X1 U7799 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6937) );
  AOI22_X1 U7800 ( .A1(n6937), .A2(keyinput_g39), .B1(keyinput_g68), .B2(n6833), .ZN(n6832) );
  OAI221_X1 U7801 ( .B1(n6937), .B2(keyinput_g39), .C1(n6833), .C2(
        keyinput_g68), .A(n6832), .ZN(n6839) );
  AOI22_X1 U7802 ( .A1(n6835), .A2(keyinput_g82), .B1(n7062), .B2(keyinput_g51), .ZN(n6834) );
  OAI221_X1 U7803 ( .B1(n6835), .B2(keyinput_g82), .C1(n7062), .C2(
        keyinput_g51), .A(n6834), .ZN(n6838) );
  AOI22_X1 U7804 ( .A1(n7018), .A2(keyinput_g62), .B1(n7036), .B2(keyinput_g66), .ZN(n6836) );
  OAI221_X1 U7805 ( .B1(n7018), .B2(keyinput_g62), .C1(n7036), .C2(
        keyinput_g66), .A(n6836), .ZN(n6837) );
  NOR4_X1 U7806 ( .A1(n6840), .A2(n6839), .A3(n6838), .A4(n6837), .ZN(n6865)
         );
  AOI22_X1 U7807 ( .A1(n7015), .A2(keyinput_g59), .B1(keyinput_g95), .B2(n7046), .ZN(n6841) );
  OAI221_X1 U7808 ( .B1(n7015), .B2(keyinput_g59), .C1(n7046), .C2(
        keyinput_g95), .A(n6841), .ZN(n6849) );
  INV_X1 U7809 ( .A(DATAI_23_), .ZN(n6952) );
  AOI22_X1 U7810 ( .A1(n6952), .A2(keyinput_g8), .B1(keyinput_g97), .B2(n7065), 
        .ZN(n6842) );
  OAI221_X1 U7811 ( .B1(n6952), .B2(keyinput_g8), .C1(n7065), .C2(keyinput_g97), .A(n6842), .ZN(n6848) );
  AOI22_X1 U7812 ( .A1(n6899), .A2(keyinput_g27), .B1(keyinput_g119), .B2(
        n6844), .ZN(n6843) );
  OAI221_X1 U7813 ( .B1(n6899), .B2(keyinput_g27), .C1(n6844), .C2(
        keyinput_g119), .A(n6843), .ZN(n6847) );
  AOI22_X1 U7814 ( .A1(n6930), .A2(keyinput_g80), .B1(n6953), .B2(keyinput_g17), .ZN(n6845) );
  OAI221_X1 U7815 ( .B1(n6930), .B2(keyinput_g80), .C1(n6953), .C2(
        keyinput_g17), .A(n6845), .ZN(n6846) );
  NOR4_X1 U7816 ( .A1(n6849), .A2(n6848), .A3(n6847), .A4(n6846), .ZN(n6864)
         );
  AOI22_X1 U7817 ( .A1(n6852), .A2(keyinput_g125), .B1(n6851), .B2(
        keyinput_g18), .ZN(n6850) );
  OAI221_X1 U7818 ( .B1(n6852), .B2(keyinput_g125), .C1(n6851), .C2(
        keyinput_g18), .A(n6850), .ZN(n6862) );
  AOI22_X1 U7819 ( .A1(n6959), .A2(keyinput_g47), .B1(n6854), .B2(keyinput_g19), .ZN(n6853) );
  OAI221_X1 U7820 ( .B1(n6959), .B2(keyinput_g47), .C1(n6854), .C2(
        keyinput_g19), .A(n6853), .ZN(n6861) );
  AOI22_X1 U7821 ( .A1(n6857), .A2(keyinput_g115), .B1(keyinput_g112), .B2(
        n6856), .ZN(n6855) );
  OAI221_X1 U7822 ( .B1(n6857), .B2(keyinput_g115), .C1(n6856), .C2(
        keyinput_g112), .A(n6855), .ZN(n6860) );
  AOI22_X1 U7823 ( .A1(n6934), .A2(keyinput_g127), .B1(keyinput_g77), .B2(
        n7049), .ZN(n6858) );
  OAI221_X1 U7824 ( .B1(n6934), .B2(keyinput_g127), .C1(n7049), .C2(
        keyinput_g77), .A(n6858), .ZN(n6859) );
  NOR4_X1 U7825 ( .A1(n6862), .A2(n6861), .A3(n6860), .A4(n6859), .ZN(n6863)
         );
  NAND4_X1 U7826 ( .A1(n6866), .A2(n6865), .A3(n6864), .A4(n6863), .ZN(n6867)
         );
  NOR4_X1 U7827 ( .A1(n6870), .A2(n6869), .A3(n6868), .A4(n6867), .ZN(n7091)
         );
  OAI22_X1 U7828 ( .A1(keyinput_f87), .A2(ADDRESS_REG_13__SCAN_IN), .B1(
        keyinput_f86), .B2(ADDRESS_REG_14__SCAN_IN), .ZN(n6871) );
  AOI221_X1 U7829 ( .B1(keyinput_f87), .B2(ADDRESS_REG_13__SCAN_IN), .C1(
        ADDRESS_REG_14__SCAN_IN), .C2(keyinput_f86), .A(n6871), .ZN(n6878) );
  OAI22_X1 U7830 ( .A1(keyinput_f120), .A2(DATAWIDTH_REG_16__SCAN_IN), .B1(
        keyinput_f72), .B2(ADDRESS_REG_28__SCAN_IN), .ZN(n6872) );
  AOI221_X1 U7831 ( .B1(keyinput_f120), .B2(DATAWIDTH_REG_16__SCAN_IN), .C1(
        ADDRESS_REG_28__SCAN_IN), .C2(keyinput_f72), .A(n6872), .ZN(n6877) );
  OAI22_X1 U7832 ( .A1(keyinput_f73), .A2(ADDRESS_REG_27__SCAN_IN), .B1(
        keyinput_f113), .B2(DATAWIDTH_REG_9__SCAN_IN), .ZN(n6873) );
  AOI221_X1 U7833 ( .B1(keyinput_f73), .B2(ADDRESS_REG_27__SCAN_IN), .C1(
        DATAWIDTH_REG_9__SCAN_IN), .C2(keyinput_f113), .A(n6873), .ZN(n6876)
         );
  OAI22_X1 U7834 ( .A1(DATAI_27_), .A2(keyinput_f4), .B1(keyinput_f33), .B2(
        NA_N), .ZN(n6874) );
  AOI221_X1 U7835 ( .B1(DATAI_27_), .B2(keyinput_f4), .C1(NA_N), .C2(
        keyinput_f33), .A(n6874), .ZN(n6875) );
  NAND4_X1 U7836 ( .A1(n6878), .A2(n6877), .A3(n6876), .A4(n6875), .ZN(n6911)
         );
  OAI22_X1 U7837 ( .A1(DATAI_13_), .A2(keyinput_f18), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(keyinput_f76), .ZN(n6879) );
  AOI221_X1 U7838 ( .B1(DATAI_13_), .B2(keyinput_f18), .C1(keyinput_f76), .C2(
        ADDRESS_REG_24__SCAN_IN), .A(n6879), .ZN(n6886) );
  OAI22_X1 U7839 ( .A1(keyinput_f70), .A2(BE_N_REG_0__SCAN_IN), .B1(
        keyinput_f93), .B2(ADDRESS_REG_7__SCAN_IN), .ZN(n6880) );
  AOI221_X1 U7840 ( .B1(keyinput_f70), .B2(BE_N_REG_0__SCAN_IN), .C1(
        ADDRESS_REG_7__SCAN_IN), .C2(keyinput_f93), .A(n6880), .ZN(n6885) );
  OAI22_X1 U7841 ( .A1(REIP_REG_28__SCAN_IN), .A2(keyinput_f54), .B1(
        keyinput_f64), .B2(REIP_REG_18__SCAN_IN), .ZN(n6881) );
  AOI221_X1 U7842 ( .B1(REIP_REG_28__SCAN_IN), .B2(keyinput_f54), .C1(
        REIP_REG_18__SCAN_IN), .C2(keyinput_f64), .A(n6881), .ZN(n6884) );
  OAI22_X1 U7843 ( .A1(DATAI_11_), .A2(keyinput_f20), .B1(keyinput_f30), .B2(
        DATAI_1_), .ZN(n6882) );
  AOI221_X1 U7844 ( .B1(DATAI_11_), .B2(keyinput_f20), .C1(DATAI_1_), .C2(
        keyinput_f30), .A(n6882), .ZN(n6883) );
  NAND4_X1 U7845 ( .A1(n6886), .A2(n6885), .A3(n6884), .A4(n6883), .ZN(n6910)
         );
  OAI22_X1 U7846 ( .A1(DATAI_12_), .A2(keyinput_f19), .B1(keyinput_f112), .B2(
        DATAWIDTH_REG_8__SCAN_IN), .ZN(n6887) );
  AOI221_X1 U7847 ( .B1(DATAI_12_), .B2(keyinput_f19), .C1(
        DATAWIDTH_REG_8__SCAN_IN), .C2(keyinput_f112), .A(n6887), .ZN(n6894)
         );
  OAI22_X1 U7848 ( .A1(keyinput_f119), .A2(DATAWIDTH_REG_15__SCAN_IN), .B1(
        keyinput_f36), .B2(HOLD), .ZN(n6888) );
  AOI221_X1 U7849 ( .B1(keyinput_f119), .B2(DATAWIDTH_REG_15__SCAN_IN), .C1(
        HOLD), .C2(keyinput_f36), .A(n6888), .ZN(n6893) );
  OAI22_X1 U7850 ( .A1(DATAI_24_), .A2(keyinput_f7), .B1(keyinput_f29), .B2(
        DATAI_2_), .ZN(n6889) );
  AOI221_X1 U7851 ( .B1(DATAI_24_), .B2(keyinput_f7), .C1(DATAI_2_), .C2(
        keyinput_f29), .A(n6889), .ZN(n6892) );
  OAI22_X1 U7852 ( .A1(keyinput_f117), .A2(DATAWIDTH_REG_13__SCAN_IN), .B1(
        keyinput_f48), .B2(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6890) );
  AOI221_X1 U7853 ( .B1(keyinput_f117), .B2(DATAWIDTH_REG_13__SCAN_IN), .C1(
        BYTEENABLE_REG_1__SCAN_IN), .C2(keyinput_f48), .A(n6890), .ZN(n6891)
         );
  NAND4_X1 U7854 ( .A1(n6894), .A2(n6893), .A3(n6892), .A4(n6891), .ZN(n6909)
         );
  OAI22_X1 U7855 ( .A1(keyinput_f81), .A2(ADDRESS_REG_19__SCAN_IN), .B1(
        keyinput_f68), .B2(BE_N_REG_2__SCAN_IN), .ZN(n6895) );
  AOI221_X1 U7856 ( .B1(keyinput_f81), .B2(ADDRESS_REG_19__SCAN_IN), .C1(
        BE_N_REG_2__SCAN_IN), .C2(keyinput_f68), .A(n6895), .ZN(n6907) );
  OAI22_X1 U7857 ( .A1(n6897), .A2(keyinput_f31), .B1(ADDRESS_REG_15__SCAN_IN), 
        .B2(keyinput_f85), .ZN(n6896) );
  AOI221_X1 U7858 ( .B1(n6897), .B2(keyinput_f31), .C1(keyinput_f85), .C2(
        ADDRESS_REG_15__SCAN_IN), .A(n6896), .ZN(n6906) );
  OAI22_X1 U7859 ( .A1(n6900), .A2(keyinput_f52), .B1(n6899), .B2(keyinput_f27), .ZN(n6898) );
  AOI221_X1 U7860 ( .B1(n6900), .B2(keyinput_f52), .C1(keyinput_f27), .C2(
        n6899), .A(n6898), .ZN(n6905) );
  OAI22_X1 U7861 ( .A1(keyinput_f121), .A2(n6903), .B1(n6902), .B2(
        keyinput_f71), .ZN(n6901) );
  AOI221_X1 U7862 ( .B1(n6903), .B2(keyinput_f121), .C1(n6902), .C2(
        keyinput_f71), .A(n6901), .ZN(n6904) );
  NAND4_X1 U7863 ( .A1(n6907), .A2(n6906), .A3(n6905), .A4(n6904), .ZN(n6908)
         );
  NOR4_X1 U7864 ( .A1(n6911), .A2(n6910), .A3(n6909), .A4(n6908), .ZN(n7085)
         );
  AOI22_X1 U7865 ( .A1(n6914), .A2(keyinput_f99), .B1(n6913), .B2(keyinput_f60), .ZN(n6912) );
  OAI221_X1 U7866 ( .B1(n6914), .B2(keyinput_f99), .C1(n6913), .C2(
        keyinput_f60), .A(n6912), .ZN(n6927) );
  INV_X1 U7867 ( .A(DATAI_17_), .ZN(n6917) );
  AOI22_X1 U7868 ( .A1(n6917), .A2(keyinput_f14), .B1(n6916), .B2(keyinput_f65), .ZN(n6915) );
  OAI221_X1 U7869 ( .B1(n6917), .B2(keyinput_f14), .C1(n6916), .C2(
        keyinput_f65), .A(n6915), .ZN(n6926) );
  INV_X1 U7870 ( .A(DATAI_16_), .ZN(n6919) );
  AOI22_X1 U7871 ( .A1(n6920), .A2(keyinput_f57), .B1(keyinput_f15), .B2(n6919), .ZN(n6918) );
  OAI221_X1 U7872 ( .B1(n6920), .B2(keyinput_f57), .C1(n6919), .C2(
        keyinput_f15), .A(n6918), .ZN(n6925) );
  AOI22_X1 U7873 ( .A1(n6923), .A2(keyinput_f38), .B1(n6922), .B2(keyinput_f58), .ZN(n6921) );
  OAI221_X1 U7874 ( .B1(n6923), .B2(keyinput_f38), .C1(n6922), .C2(
        keyinput_f58), .A(n6921), .ZN(n6924) );
  NOR4_X1 U7875 ( .A1(n6927), .A2(n6926), .A3(n6925), .A4(n6924), .ZN(n7084)
         );
  AOI22_X1 U7876 ( .A1(n6930), .A2(keyinput_f80), .B1(keyinput_f90), .B2(n6929), .ZN(n6928) );
  OAI221_X1 U7877 ( .B1(n6930), .B2(keyinput_f80), .C1(n6929), .C2(
        keyinput_f90), .A(n6928), .ZN(n6977) );
  INV_X1 U7878 ( .A(DATAI_29_), .ZN(n6933) );
  AOI22_X1 U7879 ( .A1(n6933), .A2(keyinput_f2), .B1(keyinput_f49), .B2(n6932), 
        .ZN(n6931) );
  OAI221_X1 U7880 ( .B1(n6933), .B2(keyinput_f2), .C1(n6932), .C2(keyinput_f49), .A(n6931), .ZN(n6976) );
  XNOR2_X1 U7881 ( .A(keyinput_f127), .B(n6934), .ZN(n6939) );
  AOI22_X1 U7882 ( .A1(n6937), .A2(keyinput_f39), .B1(n6936), .B2(
        keyinput_f101), .ZN(n6935) );
  OAI221_X1 U7883 ( .B1(n6937), .B2(keyinput_f39), .C1(n6936), .C2(
        keyinput_f101), .A(n6935), .ZN(n6938) );
  AOI211_X1 U7884 ( .C1(n6941), .C2(keyinput_f26), .A(n6939), .B(n6938), .ZN(
        n6940) );
  OAI21_X1 U7885 ( .B1(n6941), .B2(keyinput_f26), .A(n6940), .ZN(n6975) );
  OAI22_X1 U7886 ( .A1(keyinput_f122), .A2(n6944), .B1(n6943), .B2(
        keyinput_f40), .ZN(n6942) );
  AOI221_X1 U7887 ( .B1(n6944), .B2(keyinput_f122), .C1(n6943), .C2(
        keyinput_f40), .A(n6942), .ZN(n6973) );
  AOI22_X1 U7888 ( .A1(n6947), .A2(keyinput_f56), .B1(n6946), .B2(keyinput_f53), .ZN(n6945) );
  OAI221_X1 U7889 ( .B1(n6947), .B2(keyinput_f56), .C1(n6946), .C2(
        keyinput_f53), .A(n6945), .ZN(n6956) );
  AOI22_X1 U7890 ( .A1(n6950), .A2(keyinput_f24), .B1(keyinput_f16), .B2(n6949), .ZN(n6948) );
  OAI221_X1 U7891 ( .B1(n6950), .B2(keyinput_f24), .C1(n6949), .C2(
        keyinput_f16), .A(n6948), .ZN(n6955) );
  AOI22_X1 U7892 ( .A1(n6953), .A2(keyinput_f17), .B1(keyinput_f8), .B2(n6952), 
        .ZN(n6951) );
  OAI221_X1 U7893 ( .B1(n6953), .B2(keyinput_f17), .C1(n6952), .C2(keyinput_f8), .A(n6951), .ZN(n6954) );
  NOR3_X1 U7894 ( .A1(n6956), .A2(n6955), .A3(n6954), .ZN(n6972) );
  OAI22_X1 U7895 ( .A1(keyinput_f47), .A2(n6959), .B1(n6958), .B2(keyinput_f41), .ZN(n6957) );
  AOI221_X1 U7896 ( .B1(n6959), .B2(keyinput_f47), .C1(n6958), .C2(
        keyinput_f41), .A(n6957), .ZN(n6971) );
  XOR2_X1 U7897 ( .A(keyinput_f116), .B(DATAWIDTH_REG_12__SCAN_IN), .Z(n6969)
         );
  XOR2_X1 U7898 ( .A(keyinput_f114), .B(DATAWIDTH_REG_10__SCAN_IN), .Z(n6968)
         );
  INV_X1 U7899 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6962) );
  AOI22_X1 U7900 ( .A1(n6962), .A2(keyinput_f37), .B1(n6961), .B2(
        keyinput_f103), .ZN(n6960) );
  OAI221_X1 U7901 ( .B1(n6962), .B2(keyinput_f37), .C1(n6961), .C2(
        keyinput_f103), .A(n6960), .ZN(n6967) );
  AOI22_X1 U7902 ( .A1(n6965), .A2(keyinput_f5), .B1(keyinput_f46), .B2(n6964), 
        .ZN(n6963) );
  OAI221_X1 U7903 ( .B1(n6965), .B2(keyinput_f5), .C1(n6964), .C2(keyinput_f46), .A(n6963), .ZN(n6966) );
  NOR4_X1 U7904 ( .A1(n6969), .A2(n6968), .A3(n6967), .A4(n6966), .ZN(n6970)
         );
  NAND4_X1 U7905 ( .A1(n6973), .A2(n6972), .A3(n6971), .A4(n6970), .ZN(n6974)
         );
  NOR4_X1 U7906 ( .A1(n6977), .A2(n6976), .A3(n6975), .A4(n6974), .ZN(n7083)
         );
  OAI22_X1 U7907 ( .A1(keyinput_f106), .A2(DATAWIDTH_REG_2__SCAN_IN), .B1(
        keyinput_f115), .B2(DATAWIDTH_REG_11__SCAN_IN), .ZN(n6978) );
  AOI221_X1 U7908 ( .B1(keyinput_f106), .B2(DATAWIDTH_REG_2__SCAN_IN), .C1(
        DATAWIDTH_REG_11__SCAN_IN), .C2(keyinput_f115), .A(n6978), .ZN(n6985)
         );
  OAI22_X1 U7909 ( .A1(REIP_REG_27__SCAN_IN), .A2(keyinput_f55), .B1(
        BE_N_REG_1__SCAN_IN), .B2(keyinput_f69), .ZN(n6979) );
  AOI221_X1 U7910 ( .B1(REIP_REG_27__SCAN_IN), .B2(keyinput_f55), .C1(
        keyinput_f69), .C2(BE_N_REG_1__SCAN_IN), .A(n6979), .ZN(n6984) );
  OAI22_X1 U7911 ( .A1(keyinput_f104), .A2(DATAWIDTH_REG_0__SCAN_IN), .B1(
        keyinput_f91), .B2(ADDRESS_REG_9__SCAN_IN), .ZN(n6980) );
  AOI221_X1 U7912 ( .B1(keyinput_f104), .B2(DATAWIDTH_REG_0__SCAN_IN), .C1(
        ADDRESS_REG_9__SCAN_IN), .C2(keyinput_f91), .A(n6980), .ZN(n6983) );
  OAI22_X1 U7913 ( .A1(DATAI_21_), .A2(keyinput_f10), .B1(keyinput_f89), .B2(
        ADDRESS_REG_11__SCAN_IN), .ZN(n6981) );
  AOI221_X1 U7914 ( .B1(DATAI_21_), .B2(keyinput_f10), .C1(
        ADDRESS_REG_11__SCAN_IN), .C2(keyinput_f89), .A(n6981), .ZN(n6982) );
  NAND4_X1 U7915 ( .A1(n6985), .A2(n6984), .A3(n6983), .A4(n6982), .ZN(n7081)
         );
  OAI22_X1 U7916 ( .A1(keyinput_f84), .A2(ADDRESS_REG_16__SCAN_IN), .B1(
        keyinput_f34), .B2(BS16_N), .ZN(n6986) );
  AOI221_X1 U7917 ( .B1(keyinput_f84), .B2(ADDRESS_REG_16__SCAN_IN), .C1(
        BS16_N), .C2(keyinput_f34), .A(n6986), .ZN(n7012) );
  OAI22_X1 U7918 ( .A1(DATAI_28_), .A2(keyinput_f3), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(keyinput_f96), .ZN(n6987) );
  AOI221_X1 U7919 ( .B1(DATAI_28_), .B2(keyinput_f3), .C1(keyinput_f96), .C2(
        ADDRESS_REG_4__SCAN_IN), .A(n6987), .ZN(n6990) );
  OAI22_X1 U7920 ( .A1(DATAI_19_), .A2(keyinput_f12), .B1(
        DATAWIDTH_REG_1__SCAN_IN), .B2(keyinput_f105), .ZN(n6988) );
  AOI221_X1 U7921 ( .B1(DATAI_19_), .B2(keyinput_f12), .C1(keyinput_f105), 
        .C2(DATAWIDTH_REG_1__SCAN_IN), .A(n6988), .ZN(n6989) );
  OAI211_X1 U7922 ( .C1(n6992), .C2(keyinput_f100), .A(n6990), .B(n6989), .ZN(
        n6991) );
  AOI21_X1 U7923 ( .B1(n6992), .B2(keyinput_f100), .A(n6991), .ZN(n7011) );
  AOI22_X1 U7924 ( .A1(keyinput_f79), .A2(ADDRESS_REG_21__SCAN_IN), .B1(
        keyinput_f123), .B2(DATAWIDTH_REG_19__SCAN_IN), .ZN(n6993) );
  OAI221_X1 U7925 ( .B1(keyinput_f79), .B2(ADDRESS_REG_21__SCAN_IN), .C1(
        keyinput_f123), .C2(DATAWIDTH_REG_19__SCAN_IN), .A(n6993), .ZN(n7000)
         );
  AOI22_X1 U7926 ( .A1(keyinput_f50), .A2(BYTEENABLE_REG_3__SCAN_IN), .B1(
        REIP_REG_19__SCAN_IN), .B2(keyinput_f63), .ZN(n6994) );
  OAI221_X1 U7927 ( .B1(keyinput_f50), .B2(BYTEENABLE_REG_3__SCAN_IN), .C1(
        REIP_REG_19__SCAN_IN), .C2(keyinput_f63), .A(n6994), .ZN(n6999) );
  AOI22_X1 U7928 ( .A1(keyinput_f67), .A2(BE_N_REG_3__SCAN_IN), .B1(DATAI_6_), 
        .B2(keyinput_f25), .ZN(n6995) );
  OAI221_X1 U7929 ( .B1(keyinput_f67), .B2(BE_N_REG_3__SCAN_IN), .C1(DATAI_6_), 
        .C2(keyinput_f25), .A(n6995), .ZN(n6998) );
  AOI22_X1 U7930 ( .A1(keyinput_f94), .A2(ADDRESS_REG_6__SCAN_IN), .B1(
        keyinput_f110), .B2(DATAWIDTH_REG_6__SCAN_IN), .ZN(n6996) );
  OAI221_X1 U7931 ( .B1(keyinput_f94), .B2(ADDRESS_REG_6__SCAN_IN), .C1(
        keyinput_f110), .C2(DATAWIDTH_REG_6__SCAN_IN), .A(n6996), .ZN(n6997)
         );
  NOR4_X1 U7932 ( .A1(n7000), .A2(n6999), .A3(n6998), .A4(n6997), .ZN(n7010)
         );
  AOI22_X1 U7933 ( .A1(keyinput_f109), .A2(DATAWIDTH_REG_5__SCAN_IN), .B1(
        DATAI_30_), .B2(keyinput_f1), .ZN(n7001) );
  OAI221_X1 U7934 ( .B1(keyinput_f109), .B2(DATAWIDTH_REG_5__SCAN_IN), .C1(
        DATAI_30_), .C2(keyinput_f1), .A(n7001), .ZN(n7008) );
  AOI22_X1 U7935 ( .A1(keyinput_f124), .A2(DATAWIDTH_REG_20__SCAN_IN), .B1(
        MORE_REG_SCAN_IN), .B2(keyinput_f44), .ZN(n7002) );
  OAI221_X1 U7936 ( .B1(keyinput_f124), .B2(DATAWIDTH_REG_20__SCAN_IN), .C1(
        MORE_REG_SCAN_IN), .C2(keyinput_f44), .A(n7002), .ZN(n7007) );
  AOI22_X1 U7937 ( .A1(keyinput_f108), .A2(DATAWIDTH_REG_4__SCAN_IN), .B1(
        keyinput_f74), .B2(ADDRESS_REG_26__SCAN_IN), .ZN(n7003) );
  OAI221_X1 U7938 ( .B1(keyinput_f108), .B2(DATAWIDTH_REG_4__SCAN_IN), .C1(
        keyinput_f74), .C2(ADDRESS_REG_26__SCAN_IN), .A(n7003), .ZN(n7006) );
  AOI22_X1 U7939 ( .A1(keyinput_f82), .A2(ADDRESS_REG_18__SCAN_IN), .B1(
        STATEBS16_REG_SCAN_IN), .B2(keyinput_f43), .ZN(n7004) );
  OAI221_X1 U7940 ( .B1(keyinput_f82), .B2(ADDRESS_REG_18__SCAN_IN), .C1(
        STATEBS16_REG_SCAN_IN), .C2(keyinput_f43), .A(n7004), .ZN(n7005) );
  NOR4_X1 U7941 ( .A1(n7008), .A2(n7007), .A3(n7006), .A4(n7005), .ZN(n7009)
         );
  NAND4_X1 U7942 ( .A1(n7012), .A2(n7011), .A3(n7010), .A4(n7009), .ZN(n7080)
         );
  OAI22_X1 U7943 ( .A1(n7015), .A2(keyinput_f59), .B1(n7014), .B2(
        keyinput_f107), .ZN(n7013) );
  AOI221_X1 U7944 ( .B1(n7015), .B2(keyinput_f59), .C1(keyinput_f107), .C2(
        n7014), .A(n7013), .ZN(n7028) );
  OAI22_X1 U7945 ( .A1(n7018), .A2(keyinput_f62), .B1(n7017), .B2(keyinput_f22), .ZN(n7016) );
  AOI221_X1 U7946 ( .B1(n7018), .B2(keyinput_f62), .C1(keyinput_f22), .C2(
        n7017), .A(n7016), .ZN(n7027) );
  INV_X1 U7947 ( .A(keyinput_f125), .ZN(n7020) );
  OAI22_X1 U7948 ( .A1(n7021), .A2(keyinput_f102), .B1(n7020), .B2(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n7019) );
  AOI221_X1 U7949 ( .B1(n7021), .B2(keyinput_f102), .C1(
        DATAWIDTH_REG_21__SCAN_IN), .C2(n7020), .A(n7019), .ZN(n7026) );
  OAI22_X1 U7950 ( .A1(n7024), .A2(keyinput_f61), .B1(n7023), .B2(keyinput_f6), 
        .ZN(n7022) );
  AOI221_X1 U7951 ( .B1(n7024), .B2(keyinput_f61), .C1(keyinput_f6), .C2(n7023), .A(n7022), .ZN(n7025) );
  NAND4_X1 U7952 ( .A1(n7028), .A2(n7027), .A3(n7026), .A4(n7025), .ZN(n7079)
         );
  INV_X1 U7953 ( .A(DATAI_18_), .ZN(n7031) );
  AOI22_X1 U7954 ( .A1(n7031), .A2(keyinput_f13), .B1(keyinput_f88), .B2(n7030), .ZN(n7029) );
  OAI221_X1 U7955 ( .B1(n7031), .B2(keyinput_f13), .C1(n7030), .C2(
        keyinput_f88), .A(n7029), .ZN(n7044) );
  AOI22_X1 U7956 ( .A1(n7034), .A2(keyinput_f28), .B1(keyinput_f98), .B2(n7033), .ZN(n7032) );
  OAI221_X1 U7957 ( .B1(n7034), .B2(keyinput_f28), .C1(n7033), .C2(
        keyinput_f98), .A(n7032), .ZN(n7043) );
  AOI22_X1 U7958 ( .A1(n7037), .A2(keyinput_f78), .B1(n7036), .B2(keyinput_f66), .ZN(n7035) );
  OAI221_X1 U7959 ( .B1(n7037), .B2(keyinput_f78), .C1(n7036), .C2(
        keyinput_f66), .A(n7035), .ZN(n7042) );
  INV_X1 U7960 ( .A(DATAI_31_), .ZN(n7040) );
  AOI22_X1 U7961 ( .A1(n7040), .A2(keyinput_f0), .B1(keyinput_f21), .B2(n7039), 
        .ZN(n7038) );
  OAI221_X1 U7962 ( .B1(n7040), .B2(keyinput_f0), .C1(n7039), .C2(keyinput_f21), .A(n7038), .ZN(n7041) );
  NOR4_X1 U7963 ( .A1(n7044), .A2(n7043), .A3(n7042), .A4(n7041), .ZN(n7077)
         );
  OAI22_X1 U7964 ( .A1(keyinput_f118), .A2(n7047), .B1(n7046), .B2(
        keyinput_f95), .ZN(n7045) );
  AOI221_X1 U7965 ( .B1(n7047), .B2(keyinput_f118), .C1(n7046), .C2(
        keyinput_f95), .A(n7045), .ZN(n7076) );
  XOR2_X1 U7966 ( .A(keyinput_f126), .B(DATAWIDTH_REG_22__SCAN_IN), .Z(n7057)
         );
  XOR2_X1 U7967 ( .A(keyinput_f111), .B(DATAWIDTH_REG_7__SCAN_IN), .Z(n7056)
         );
  AOI22_X1 U7968 ( .A1(n7050), .A2(keyinput_f23), .B1(keyinput_f77), .B2(n7049), .ZN(n7048) );
  OAI221_X1 U7969 ( .B1(n7050), .B2(keyinput_f23), .C1(n7049), .C2(
        keyinput_f77), .A(n7048), .ZN(n7055) );
  AOI22_X1 U7970 ( .A1(n7053), .A2(keyinput_f75), .B1(keyinput_f92), .B2(n7052), .ZN(n7051) );
  OAI221_X1 U7971 ( .B1(n7053), .B2(keyinput_f75), .C1(n7052), .C2(
        keyinput_f92), .A(n7051), .ZN(n7054) );
  NOR4_X1 U7972 ( .A1(n7057), .A2(n7056), .A3(n7055), .A4(n7054), .ZN(n7075)
         );
  INV_X1 U7973 ( .A(DATAI_20_), .ZN(n7059) );
  AOI22_X1 U7974 ( .A1(n7060), .A2(keyinput_f83), .B1(n7059), .B2(keyinput_f11), .ZN(n7058) );
  OAI221_X1 U7975 ( .B1(n7060), .B2(keyinput_f83), .C1(n7059), .C2(
        keyinput_f11), .A(n7058), .ZN(n7073) );
  AOI22_X1 U7976 ( .A1(n7063), .A2(keyinput_f45), .B1(n7062), .B2(keyinput_f51), .ZN(n7061) );
  OAI221_X1 U7977 ( .B1(n7063), .B2(keyinput_f45), .C1(n7062), .C2(
        keyinput_f51), .A(n7061), .ZN(n7072) );
  AOI22_X1 U7978 ( .A1(n7066), .A2(keyinput_f35), .B1(keyinput_f97), .B2(n7065), .ZN(n7064) );
  OAI221_X1 U7979 ( .B1(n7066), .B2(keyinput_f35), .C1(n7065), .C2(
        keyinput_f97), .A(n7064), .ZN(n7071) );
  INV_X1 U7980 ( .A(DATAI_22_), .ZN(n7068) );
  AOI22_X1 U7981 ( .A1(n7069), .A2(keyinput_f32), .B1(n7068), .B2(keyinput_f9), 
        .ZN(n7067) );
  OAI221_X1 U7982 ( .B1(n7069), .B2(keyinput_f32), .C1(n7068), .C2(keyinput_f9), .A(n7067), .ZN(n7070) );
  NOR4_X1 U7983 ( .A1(n7073), .A2(n7072), .A3(n7071), .A4(n7070), .ZN(n7074)
         );
  NAND4_X1 U7984 ( .A1(n7077), .A2(n7076), .A3(n7075), .A4(n7074), .ZN(n7078)
         );
  NOR4_X1 U7985 ( .A1(n7081), .A2(n7080), .A3(n7079), .A4(n7078), .ZN(n7082)
         );
  NAND4_X1 U7986 ( .A1(n7085), .A2(n7084), .A3(n7083), .A4(n7082), .ZN(n7087)
         );
  AOI21_X1 U7987 ( .B1(keyinput_f42), .B2(n7087), .A(
        REQUESTPENDING_REG_SCAN_IN), .ZN(n7089) );
  INV_X1 U7988 ( .A(keyinput_f42), .ZN(n7086) );
  AOI21_X1 U7989 ( .B1(n7087), .B2(n7086), .A(keyinput_g42), .ZN(n7088) );
  AOI22_X1 U7990 ( .A1(keyinput_g42), .A2(n7089), .B1(
        REQUESTPENDING_REG_SCAN_IN), .B2(n7088), .ZN(n7090) );
  AOI21_X1 U7991 ( .B1(n7092), .B2(n7091), .A(n7090), .ZN(n7096) );
  AOI22_X1 U7992 ( .A1(n7094), .A2(BYTEENABLE_REG_3__SCAN_IN), .B1(
        BE_N_REG_3__SCAN_IN), .B2(n7093), .ZN(n7095) );
  XNOR2_X1 U7993 ( .A(n7096), .B(n7095), .ZN(U3445) );
  AND2_X2 U3733 ( .A1(n4542), .A2(n4545), .ZN(n3374) );
  CLKBUF_X2 U3607 ( .A(n3351), .Z(n3470) );
  INV_X2 U3605 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n4969) );
  AND2_X1 U3626 ( .A1(n4462), .A2(n4248), .ZN(n6374) );
  INV_X1 U3669 ( .A(n4314), .ZN(n5733) );
  CLKBUF_X1 U3620 ( .A(n3510), .Z(n3169) );
  NAND2_X1 U3624 ( .A1(n4264), .A2(n4263), .ZN(n4266) );
  CLKBUF_X1 U3636 ( .A(n4591), .Z(n3170) );
  CLKBUF_X1 U3752 ( .A(n4550), .Z(n3171) );
  CLKBUF_X1 U3987 ( .A(n5730), .Z(n5731) );
  CLKBUF_X1 U6892 ( .A(n4650), .Z(n4651) );
endmodule

