

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4260, n4262, n4263, n4264, n4265, n4266, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10171;

  INV_X4 U4764 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U4765 ( .A(P2_STATE_REG_SCAN_IN), .ZN(n10171) );
  INV_X1 U4766 ( .A(n6553), .ZN(n6660) );
  XNOR2_X1 U4767 ( .A(n4971), .B(n4973), .ZN(n5489) );
  INV_X1 U4768 ( .A(n10171), .ZN(n4260) );
  INV_X1 U4769 ( .A(n4260), .ZN(P2_U3152) );
  INV_X1 U4770 ( .A(n4260), .ZN(n4262) );
  INV_X1 U4771 ( .A(n5986), .ZN(n4264) );
  INV_X1 U4773 ( .A(n8115), .ZN(n5298) );
  AND2_X1 U4774 ( .A1(n4763), .A2(n4762), .ZN(n5139) );
  INV_X1 U4775 ( .A(n5968), .ZN(n5615) );
  INV_X2 U4776 ( .A(n5643), .ZN(n4266) );
  INV_X1 U4777 ( .A(n5929), .ZN(n6267) );
  INV_X4 U4778 ( .A(n4264), .ZN(n4265) );
  INV_X1 U4779 ( .A(n8405), .ZN(n8480) );
  AND3_X2 U4780 ( .A1(n5007), .A2(n4811), .A3(n4810), .ZN(n6556) );
  NAND2_X1 U4781 ( .A1(n5489), .A2(n7745), .ZN(n5088) );
  INV_X1 U4782 ( .A(n5049), .ZN(n5416) );
  INV_X2 U4783 ( .A(n5050), .ZN(n5074) );
  INV_X1 U4784 ( .A(n8063), .ZN(n8096) );
  NAND2_X1 U4785 ( .A1(n9632), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4993) );
  NAND2_X1 U4787 ( .A1(n4500), .A2(n4503), .ZN(n8438) );
  INV_X1 U4788 ( .A(n5088), .ZN(n6161) );
  NAND2_X1 U4789 ( .A1(n5188), .A2(n5187), .ZN(n8830) );
  NAND2_X1 U4790 ( .A1(n5175), .A2(n5174), .ZN(n8914) );
  NAND2_X1 U4791 ( .A1(n4440), .A2(n4859), .ZN(n5092) );
  AND2_X1 U4792 ( .A1(n4837), .A2(n4483), .ZN(n6052) );
  INV_X1 U4793 ( .A(n6933), .ZN(n9259) );
  NAND2_X2 U4794 ( .A1(n8484), .A2(n4505), .ZN(n8468) );
  MUX2_X2 U4795 ( .A(n8970), .B(n8969), .S(n9068), .Z(n8982) );
  XNOR2_X2 U4796 ( .A(n8438), .B(n8437), .ZN(n8701) );
  NAND2_X1 U4797 ( .A1(n5489), .A2(n7745), .ZN(n4263) );
  INV_X4 U4798 ( .A(n7794), .ZN(n5577) );
  AND2_X4 U4799 ( .A1(n4508), .A2(n4509), .ZN(n7794) );
  INV_X1 U4800 ( .A(n5648), .ZN(n5986) );
  OAI21_X2 U4801 ( .B1(n8567), .B2(n6111), .A(n6079), .ZN(n8541) );
  XNOR2_X2 U4802 ( .A(n5576), .B(n5549), .ZN(n6125) );
  OAI21_X1 U4803 ( .B1(n8065), .B2(n4278), .A(n4324), .ZN(n8859) );
  NAND2_X1 U4804 ( .A1(n6774), .A2(n7954), .ZN(n6773) );
  NAND2_X2 U4805 ( .A1(n7821), .A2(n7819), .ZN(n7948) );
  NAND2_X1 U4806 ( .A1(n9259), .A2(n7087), .ZN(n9192) );
  NAND2_X2 U4807 ( .A1(n6092), .A2(n6093), .ZN(n7092) );
  INV_X1 U4808 ( .A(n9255), .ZN(n7157) );
  INV_X2 U4809 ( .A(n6661), .ZN(n7263) );
  NAND2_X2 U4810 ( .A1(n6051), .A2(n7101), .ZN(n6092) );
  INV_X1 U4811 ( .A(n6568), .ZN(n6897) );
  CLKBUF_X2 U4812 ( .A(n5122), .Z(n8114) );
  INV_X1 U4814 ( .A(n5648), .ZN(n5603) );
  OR2_X1 U4815 ( .A1(n7798), .A2(n6199), .ZN(n5600) );
  NAND2_X4 U4816 ( .A1(n6034), .A2(n6125), .ZN(n5592) );
  NOR2_X1 U4817 ( .A1(n4310), .A2(n7986), .ZN(n7994) );
  NAND2_X1 U4818 ( .A1(n8808), .A2(n8059), .ZN(n8065) );
  AOI22_X1 U4819 ( .A1(n9180), .A2(n9117), .B1(n5464), .B2(n9177), .ZN(n9179)
         );
  AOI21_X1 U4820 ( .B1(n8670), .B2(n8130), .A(n8124), .ZN(n8125) );
  AOI21_X1 U4821 ( .B1(n8748), .B2(n8130), .A(n8129), .ZN(n8131) );
  MUX2_X1 U4822 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8128), .S(n10120), .Z(n8124) );
  MUX2_X1 U4823 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8128), .S(n10101), .Z(n8129) );
  NOR2_X1 U4824 ( .A1(n8505), .A2(n8506), .ZN(n8504) );
  NAND2_X1 U4825 ( .A1(n8841), .A2(n8014), .ZN(n8850) );
  NAND2_X1 U4826 ( .A1(n8470), .A2(n8471), .ZN(n8469) );
  NAND2_X1 U4827 ( .A1(n7747), .A2(n6077), .ZN(n8574) );
  AND2_X1 U4828 ( .A1(n7536), .A2(n7507), .ZN(n7506) );
  NAND3_X1 U4829 ( .A1(n7497), .A2(n7489), .A3(n7498), .ZN(n7536) );
  AND2_X1 U4830 ( .A1(n4617), .A2(n4616), .ZN(n4621) );
  AND2_X1 U4831 ( .A1(n4622), .A2(n8776), .ZN(n4279) );
  AND2_X1 U4832 ( .A1(n4602), .A2(n7258), .ZN(n7269) );
  AND2_X1 U4833 ( .A1(n7690), .A2(n8772), .ZN(n7677) );
  OR2_X1 U4834 ( .A1(n8566), .A2(n8549), .ZN(n8550) );
  OR2_X1 U4835 ( .A1(n7681), .A2(n8878), .ZN(n8772) );
  NAND2_X1 U4836 ( .A1(n7029), .A2(n7028), .ZN(n7258) );
  NOR2_X1 U4837 ( .A1(n8580), .A2(n8742), .ZN(n8581) );
  OR2_X1 U4838 ( .A1(n7757), .A2(n8747), .ZN(n8580) );
  OAI21_X1 U4839 ( .B1(n9969), .B2(n4582), .A(n4580), .ZN(n6104) );
  OR2_X1 U4840 ( .A1(n4271), .A2(n8143), .ZN(n7757) );
  OR2_X1 U4841 ( .A1(n6064), .A2(n6063), .ZN(n9951) );
  AND2_X1 U4842 ( .A1(n7845), .A2(n7844), .ZN(n7957) );
  AND2_X1 U4843 ( .A1(n7841), .A2(n7842), .ZN(n7956) );
  NAND2_X1 U4844 ( .A1(n5710), .A2(n5709), .ZN(n10070) );
  INV_X4 U4845 ( .A(n7263), .ZN(n4269) );
  XNOR2_X1 U4846 ( .A(n5171), .B(n5170), .ZN(n6238) );
  NAND2_X1 U4847 ( .A1(n5129), .A2(n5128), .ZN(n7540) );
  NAND2_X1 U4848 ( .A1(n5468), .A2(n5467), .ZN(n9198) );
  INV_X2 U4849 ( .A(n6660), .ZN(n8073) );
  AND4_X1 U4850 ( .A1(n5717), .A2(n5716), .A3(n5715), .A4(n5714), .ZN(n6969)
         );
  AND4_X1 U4851 ( .A1(n5701), .A2(n5700), .A3(n5699), .A4(n5698), .ZN(n7129)
         );
  INV_X1 U4852 ( .A(n10043), .ZN(n7079) );
  AND2_X1 U4853 ( .A1(n6416), .A2(n7259), .ZN(n6553) );
  INV_X2 U4854 ( .A(n8324), .ZN(n6051) );
  AND2_X1 U4855 ( .A1(n4301), .A2(n5609), .ZN(n7832) );
  INV_X2 U4856 ( .A(n8303), .ZN(P2_U3966) );
  AND2_X1 U4857 ( .A1(n5039), .A2(n5038), .ZN(n7087) );
  NAND2_X2 U4858 ( .A1(n5581), .A2(n5580), .ZN(n5968) );
  AND2_X2 U4859 ( .A1(n6554), .A2(n6417), .ZN(n8063) );
  AND2_X1 U4860 ( .A1(n6417), .A2(n6697), .ZN(n7259) );
  NAND4_X1 U4861 ( .A1(n5013), .A2(n5012), .A3(n5011), .A4(n5010), .ZN(n6568)
         );
  NAND2_X1 U4862 ( .A1(n7608), .A2(n5511), .ZN(n6697) );
  CLKBUF_X3 U4864 ( .A(n5051), .Z(n5492) );
  AOI21_X1 U4865 ( .B1(n6245), .B2(P1_REG2_REG_1__SCAN_IN), .A(n4809), .ZN(
        n4808) );
  AND3_X1 U4866 ( .A1(n5614), .A2(n5613), .A3(n5612), .ZN(n7247) );
  AND2_X1 U4867 ( .A1(n9637), .A2(n4996), .ZN(n5050) );
  AND2_X2 U4868 ( .A1(n4997), .A2(n9643), .ZN(n6245) );
  AND2_X1 U4869 ( .A1(n8764), .A2(n5558), .ZN(n5607) );
  AND2_X2 U4870 ( .A1(n8764), .A2(n8767), .ZN(n5918) );
  OAI211_X2 U4871 ( .C1(n5592), .C2(n6438), .A(n5601), .B(n5600), .ZN(n9991)
         );
  INV_X1 U4872 ( .A(n4996), .ZN(n9643) );
  NAND2_X4 U4873 ( .A1(n4997), .A2(n4996), .ZN(n5049) );
  INV_X1 U4874 ( .A(n7798), .ZN(n5862) );
  XNOR2_X1 U4875 ( .A(n5297), .B(n5453), .ZN(n9878) );
  NAND2_X1 U4876 ( .A1(n5556), .A2(n5555), .ZN(n8767) );
  NAND2_X1 U4877 ( .A1(n5555), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5551) );
  NAND2_X1 U4878 ( .A1(n5554), .A2(n5553), .ZN(n5556) );
  OAI21_X1 U4879 ( .B1(n5455), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5457) );
  NAND2_X1 U4880 ( .A1(n4881), .A2(n4870), .ZN(n5120) );
  OR2_X1 U4881 ( .A1(n5575), .A2(n6000), .ZN(n5576) );
  AND2_X1 U4882 ( .A1(n5512), .A2(n4970), .ZN(n5505) );
  AND2_X1 U4883 ( .A1(n4833), .A2(n4838), .ZN(n4831) );
  INV_X2 U4884 ( .A(n6576), .ZN(n4268) );
  AND3_X1 U4885 ( .A1(n4598), .A2(n4788), .A3(n4597), .ZN(n4596) );
  AND2_X1 U4886 ( .A1(n4604), .A2(n4337), .ZN(n4603) );
  INV_X1 U4887 ( .A(n4835), .ZN(n4599) );
  AND2_X1 U4888 ( .A1(n4963), .A2(n5089), .ZN(n5185) );
  AND2_X1 U4889 ( .A1(n4605), .A2(n5266), .ZN(n4604) );
  AND2_X1 U4890 ( .A1(n5539), .A2(n4836), .ZN(n4598) );
  NOR2_X1 U4891 ( .A1(n5250), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n4605) );
  AND2_X1 U4892 ( .A1(n5542), .A2(n4789), .ZN(n4788) );
  AND2_X1 U4893 ( .A1(n5540), .A2(n5541), .ZN(n4789) );
  NAND2_X1 U4894 ( .A1(n5563), .A2(n6279), .ZN(n5564) );
  AND2_X1 U4895 ( .A1(n5548), .A2(n4414), .ZN(n4597) );
  AND4_X1 U4896 ( .A1(n4962), .A2(n4961), .A3(n4960), .A4(n5104), .ZN(n4963)
         );
  NAND2_X1 U4897 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5550), .ZN(n5553) );
  NOR2_X1 U4898 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5535) );
  INV_X1 U4899 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5538) );
  NOR2_X1 U4900 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5536) );
  INV_X1 U4901 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4959) );
  INV_X1 U4902 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6389) );
  INV_X1 U4903 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6025) );
  NOR2_X1 U4904 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5565) );
  AND2_X1 U4905 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7448) );
  OAI21_X2 U4906 ( .B1(n5508), .B2(n4972), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n4971) );
  AND4_X2 U4907 ( .A1(n5045), .A2(n5044), .A3(n5043), .A4(n5042), .ZN(n6933)
         );
  NOR2_X2 U4908 ( .A1(n6417), .A2(n6420), .ZN(n6661) );
  OR2_X2 U4909 ( .A1(n5464), .A2(n9183), .ZN(n6417) );
  NOR2_X2 U4910 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5598) );
  NAND2_X1 U4911 ( .A1(n8486), .A2(n8485), .ZN(n8484) );
  AOI22_X2 U4912 ( .A1(n8527), .A2(n6080), .B1(n6117), .B2(n8533), .ZN(n8515)
         );
  AND2_X2 U4913 ( .A1(n7553), .A2(n6071), .ZN(n7576) );
  OR2_X2 U4914 ( .A1(n8454), .A2(n8456), .ZN(n4500) );
  OAI22_X2 U4915 ( .A1(n8515), .A2(n8517), .B1(n8302), .B2(n8647), .ZN(n8505)
         );
  AOI21_X1 U4916 ( .B1(n4664), .B2(n4666), .A(n4320), .ZN(n4662) );
  NAND2_X1 U4917 ( .A1(n5201), .A2(n4909), .ZN(n5214) );
  NAND2_X1 U4918 ( .A1(n4903), .A2(n4902), .ZN(n5183) );
  OR2_X1 U4919 ( .A1(n4883), .A2(n5140), .ZN(n4885) );
  AND2_X1 U4920 ( .A1(n4433), .A2(n7857), .ZN(n4431) );
  INV_X1 U4921 ( .A(n4435), .ZN(n4433) );
  NOR2_X1 U4922 ( .A1(n8143), .A2(n4444), .ZN(n4443) );
  OR2_X1 U4923 ( .A1(n7880), .A2(n7904), .ZN(n4444) );
  NOR2_X1 U4924 ( .A1(n7907), .A2(n4311), .ZN(n4424) );
  INV_X1 U4925 ( .A(n7905), .ZN(n4425) );
  INV_X1 U4926 ( .A(n8022), .ZN(n4615) );
  NAND2_X1 U4927 ( .A1(n4576), .A2(n8480), .ZN(n4573) );
  NAND2_X1 U4928 ( .A1(n8689), .A2(n8414), .ZN(n7939) );
  AOI21_X1 U4929 ( .B1(n4451), .B2(n4450), .A(n4449), .ZN(n4448) );
  AND2_X1 U4930 ( .A1(n7926), .A2(n7807), .ZN(n4450) );
  NOR2_X1 U4931 ( .A1(n7926), .A2(n7807), .ZN(n4449) );
  OAI21_X1 U4932 ( .B1(n7929), .B2(n8296), .A(n7925), .ZN(n4451) );
  INV_X1 U4933 ( .A(n8767), .ZN(n5558) );
  AND2_X1 U4934 ( .A1(n7862), .A2(n7863), .ZN(n7964) );
  AND2_X1 U4935 ( .A1(n7980), .A2(n7947), .ZN(n6090) );
  OR2_X1 U4936 ( .A1(n8130), .A2(n6782), .ZN(n7926) );
  AND2_X1 U4937 ( .A1(n4598), .A2(n4414), .ZN(n5739) );
  AND2_X1 U4938 ( .A1(n9329), .A2(n9080), .ZN(n4689) );
  OR2_X1 U4939 ( .A1(n9429), .A2(n9411), .ZN(n9149) );
  NOR2_X1 U4940 ( .A1(n4701), .A2(n5212), .ZN(n4699) );
  NOR2_X1 U4941 ( .A1(n4283), .A2(n4703), .ZN(n4702) );
  INV_X1 U4942 ( .A(n4704), .ZN(n4703) );
  NOR2_X1 U4943 ( .A1(n7038), .A2(n7264), .ZN(n4538) );
  NAND2_X1 U4944 ( .A1(n6947), .A2(n6849), .ZN(n9199) );
  NAND2_X1 U4945 ( .A1(n9258), .A2(n9912), .ZN(n9196) );
  NAND2_X1 U4946 ( .A1(n6824), .A2(n6933), .ZN(n9193) );
  NAND2_X1 U4947 ( .A1(n5392), .A2(n5391), .ZN(n5408) );
  AND2_X1 U4948 ( .A1(n5390), .A2(n5369), .ZN(n4757) );
  NAND2_X1 U4949 ( .A1(n5312), .A2(n5311), .ZN(n4944) );
  OAI21_X1 U4950 ( .B1(n5293), .B2(n5292), .A(n4938), .ZN(n5312) );
  OAI21_X1 U4951 ( .B1(n5265), .B2(n4929), .A(n4928), .ZN(n5279) );
  AND2_X1 U4952 ( .A1(n4924), .A2(n4923), .ZN(n5247) );
  NAND2_X1 U4953 ( .A1(n4895), .A2(SI_11_), .ZN(n4896) );
  NAND2_X1 U4954 ( .A1(n4386), .A2(n4384), .ZN(n8183) );
  AND2_X1 U4955 ( .A1(n5873), .A2(n4385), .ZN(n4384) );
  NAND2_X1 U4956 ( .A1(n7611), .A2(n5794), .ZN(n7620) );
  NAND2_X1 U4957 ( .A1(n6968), .A2(n6967), .ZN(n4781) );
  INV_X1 U4958 ( .A(n4769), .ZN(n4768) );
  OAI21_X1 U4959 ( .B1(n7296), .B2(n4770), .A(n7388), .ZN(n4769) );
  AND2_X1 U4960 ( .A1(n4523), .A2(n4522), .ZN(n6540) );
  NAND2_X1 U4961 ( .A1(n6538), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4522) );
  OR2_X1 U4962 ( .A1(n6540), .A2(n6539), .ZN(n4521) );
  NAND2_X1 U4963 ( .A1(n6072), .A2(n4517), .ZN(n4513) );
  AND2_X1 U4964 ( .A1(n6075), .A2(n6074), .ZN(n7967) );
  AND2_X1 U4965 ( .A1(n7966), .A2(n4515), .ZN(n4514) );
  NAND2_X1 U4966 ( .A1(n4516), .A2(n6072), .ZN(n4515) );
  AND2_X1 U4967 ( .A1(n4516), .A2(n6106), .ZN(n4583) );
  AND2_X1 U4968 ( .A1(n6070), .A2(n7554), .ZN(n4518) );
  AOI21_X1 U4969 ( .B1(n4499), .B2(n4495), .A(n4494), .ZN(n4493) );
  NOR2_X1 U4970 ( .A1(n8616), .A2(n8296), .ZN(n4494) );
  NOR2_X1 U4971 ( .A1(n4497), .A2(n8427), .ZN(n4495) );
  NOR2_X1 U4972 ( .A1(n8708), .A2(n8299), .ZN(n6081) );
  AND2_X1 U4973 ( .A1(n8155), .A2(n4331), .ZN(n4657) );
  OR2_X1 U4974 ( .A1(n4287), .A2(n7691), .ZN(n4627) );
  NOR2_X1 U4975 ( .A1(n8065), .A2(n4643), .ZN(n4641) );
  OR2_X1 U4976 ( .A1(n5097), .A2(n6222), .ZN(n4810) );
  OR2_X1 U4977 ( .A1(n5062), .A2(n6224), .ZN(n4811) );
  AOI21_X1 U4978 ( .B1(n9284), .B2(n9283), .A(n9863), .ZN(n9286) );
  AOI21_X1 U4979 ( .B1(n4667), .B2(n4665), .A(n4314), .ZN(n4664) );
  INV_X1 U4980 ( .A(n4291), .ZN(n4665) );
  OR2_X1 U4981 ( .A1(n9570), .A2(n9463), .ZN(n4671) );
  NAND2_X1 U4982 ( .A1(n4670), .A2(n4291), .ZN(n4669) );
  INV_X1 U4983 ( .A(n9438), .ZN(n4670) );
  AOI21_X1 U4984 ( .B1(n4677), .B2(n5277), .A(n4275), .ZN(n4675) );
  AND2_X1 U4985 ( .A1(n9095), .A2(n5080), .ZN(n4710) );
  XNOR2_X1 U4986 ( .A(n7797), .B(n7796), .ZN(n8758) );
  OAI21_X1 U4987 ( .B1(n7790), .B2(n4761), .A(n7793), .ZN(n7797) );
  NAND2_X1 U4988 ( .A1(n5352), .A2(n4958), .ZN(n5371) );
  NAND2_X1 U4989 ( .A1(n4743), .A2(n4741), .ZN(n5201) );
  AOI21_X1 U4990 ( .B1(n4744), .B2(n4284), .A(n4742), .ZN(n4741) );
  INV_X1 U4991 ( .A(n5198), .ZN(n4742) );
  OR2_X1 U4992 ( .A1(n8362), .A2(n8361), .ZN(n4531) );
  NAND2_X1 U4993 ( .A1(n7843), .A2(n7957), .ZN(n4435) );
  AND2_X1 U4994 ( .A1(n7956), .A2(n7838), .ZN(n4436) );
  AND2_X1 U4995 ( .A1(n4429), .A2(n4428), .ZN(n7866) );
  AND2_X1 U4996 ( .A1(n4442), .A2(n4441), .ZN(n7895) );
  NOR2_X1 U4997 ( .A1(n7885), .A2(n8558), .ZN(n4441) );
  OAI21_X1 U4998 ( .B1(n4445), .B2(n4443), .A(n7886), .ZN(n4442) );
  AND2_X1 U4999 ( .A1(n7908), .A2(n4339), .ZN(n4423) );
  NOR2_X1 U5000 ( .A1(n4274), .A2(n4322), .ZN(n4421) );
  NOR2_X1 U5001 ( .A1(n7936), .A2(n4360), .ZN(n4577) );
  NAND2_X1 U5002 ( .A1(n4481), .A2(n8446), .ZN(n4480) );
  NAND2_X1 U5003 ( .A1(n8509), .A2(n8533), .ZN(n4469) );
  INV_X1 U5004 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5541) );
  OR2_X1 U5005 ( .A1(n8977), .A2(n8976), .ZN(n9135) );
  OR2_X1 U5006 ( .A1(n7058), .A2(n6824), .ZN(n6823) );
  NAND2_X1 U5007 ( .A1(n4873), .A2(n4872), .ZN(n4884) );
  NAND2_X1 U5008 ( .A1(n4868), .A2(n4867), .ZN(n4881) );
  NOR2_X1 U5009 ( .A1(n5835), .A2(n8363), .ZN(n4373) );
  INV_X1 U5010 ( .A(n4588), .ZN(n4587) );
  NOR2_X1 U5011 ( .A1(n8514), .A2(n4589), .ZN(n4588) );
  INV_X1 U5012 ( .A(n7899), .ZN(n4589) );
  OR2_X1 U5013 ( .A1(n8549), .A2(n8197), .ZN(n7897) );
  OR2_X1 U5014 ( .A1(n5787), .A2(n7477), .ZN(n5820) );
  AND2_X1 U5015 ( .A1(n6098), .A2(n7809), .ZN(n4842) );
  NAND2_X1 U5016 ( .A1(n10043), .A2(n8320), .ZN(n7828) );
  INV_X1 U5017 ( .A(n7974), .ZN(n4488) );
  OR2_X1 U5018 ( .A1(n8626), .A2(n6082), .ZN(n7915) );
  INV_X1 U5019 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5540) );
  AND2_X1 U5020 ( .A1(n8892), .A2(n8066), .ZN(n4643) );
  OR2_X1 U5021 ( .A1(n8851), .A2(n4615), .ZN(n4614) );
  INV_X1 U5022 ( .A(n7685), .ZN(n4622) );
  OR2_X1 U5023 ( .A1(n4287), .A2(n4630), .ZN(n4629) );
  INV_X1 U5024 ( .A(n7688), .ZN(n4630) );
  OR2_X1 U5025 ( .A1(n9530), .A2(n9337), .ZN(n9167) );
  NOR2_X1 U5026 ( .A1(n9535), .A2(n9356), .ZN(n4692) );
  NOR2_X1 U5027 ( .A1(n9391), .A2(n4805), .ZN(n4804) );
  AND2_X1 U5028 ( .A1(n9155), .A2(n9033), .ZN(n9083) );
  OR2_X1 U5029 ( .A1(n9570), .A2(n5479), .ZN(n9085) );
  NOR2_X1 U5030 ( .A1(n9582), .A2(n9587), .ZN(n4547) );
  OAI21_X1 U5031 ( .B1(n7543), .B2(n9107), .A(n9135), .ZN(n7594) );
  INV_X1 U5032 ( .A(n4702), .ZN(n4696) );
  NOR2_X1 U5033 ( .A1(n4283), .A2(n5197), .ZN(n4701) );
  NOR2_X1 U5034 ( .A1(n9676), .A2(n4814), .ZN(n4813) );
  INV_X1 U5035 ( .A(n9129), .ZN(n4814) );
  INV_X1 U5036 ( .A(n8972), .ZN(n4816) );
  NAND2_X1 U5037 ( .A1(n5474), .A2(n9123), .ZN(n7105) );
  NOR2_X1 U5038 ( .A1(n5049), .A2(n6903), .ZN(n4809) );
  OR2_X1 U5039 ( .A1(n9430), .A2(n9560), .ZN(n9399) );
  OR2_X1 U5040 ( .A1(n4541), .A2(n8977), .ZN(n4540) );
  NOR2_X1 U5041 ( .A1(n6823), .A2(n6947), .ZN(n6940) );
  XNOR2_X1 U5042 ( .A(n7792), .B(n7791), .ZN(n7790) );
  NAND2_X1 U5043 ( .A1(n4723), .A2(n4722), .ZN(n7782) );
  AOI21_X1 U5044 ( .B1(n4725), .B2(n4727), .A(n4363), .ZN(n4722) );
  NAND2_X1 U5045 ( .A1(n5423), .A2(n4725), .ZN(n4723) );
  NAND2_X1 U5046 ( .A1(n5352), .A2(n4759), .ZN(n4758) );
  NOR2_X1 U5047 ( .A1(n5370), .A2(n4760), .ZN(n4759) );
  INV_X1 U5048 ( .A(n4958), .ZN(n4760) );
  NAND2_X1 U5049 ( .A1(n4933), .A2(n4932), .ZN(n5293) );
  NAND2_X1 U5050 ( .A1(n5279), .A2(n4930), .ZN(n4933) );
  AOI21_X1 U5051 ( .B1(n4732), .B2(n4735), .A(n4730), .ZN(n4729) );
  INV_X1 U5052 ( .A(n4924), .ZN(n4730) );
  NOR2_X1 U5053 ( .A1(n4897), .A2(n4749), .ZN(n4748) );
  INV_X1 U5054 ( .A(n4892), .ZN(n4749) );
  INV_X1 U5055 ( .A(n5170), .ZN(n4897) );
  XNOR2_X1 U5056 ( .A(n4894), .B(SI_11_), .ZN(n5170) );
  AND2_X1 U5057 ( .A1(n4892), .A2(n4891), .ZN(n5155) );
  INV_X1 U5058 ( .A(n4882), .ZN(n5140) );
  OAI21_X1 U5059 ( .B1(n5118), .B2(n5120), .A(n4881), .ZN(n4882) );
  NAND2_X1 U5060 ( .A1(n4764), .A2(n5095), .ZN(n4763) );
  INV_X1 U5061 ( .A(n5093), .ZN(n4764) );
  NAND2_X1 U5062 ( .A1(n4378), .A2(n4864), .ZN(n4861) );
  INV_X1 U5063 ( .A(n5060), .ZN(n4378) );
  OAI211_X1 U5064 ( .C1(n7794), .C2(P2_DATAO_REG_0__SCAN_IN), .A(SI_0_), .B(
        n4416), .ZN(n4849) );
  NAND2_X1 U5065 ( .A1(n7794), .A2(n4417), .ZN(n4416) );
  AND2_X1 U5066 ( .A1(n4844), .A2(n5633), .ZN(n4392) );
  AOI21_X1 U5067 ( .B1(n8246), .B2(n8245), .A(n5911), .ZN(n5935) );
  INV_X1 U5068 ( .A(n8321), .ZN(n6807) );
  NAND2_X1 U5069 ( .A1(n4771), .A2(n4775), .ZN(n6141) );
  INV_X1 U5070 ( .A(n4776), .ZN(n4775) );
  OAI21_X1 U5071 ( .B1(n4341), .B2(n4777), .A(n6140), .ZN(n4776) );
  INV_X1 U5072 ( .A(n5686), .ZN(n4394) );
  INV_X1 U5073 ( .A(n5685), .ZN(n4393) );
  OR2_X1 U5074 ( .A1(n8189), .A2(n5897), .ZN(n8191) );
  NAND2_X1 U5075 ( .A1(n8183), .A2(n4782), .ZN(n8192) );
  NOR2_X1 U5076 ( .A1(n4317), .A2(n4783), .ZN(n4782) );
  INV_X1 U5077 ( .A(n5877), .ZN(n4783) );
  AND2_X1 U5078 ( .A1(n5935), .A2(n5934), .ZN(n8222) );
  NAND2_X1 U5079 ( .A1(n5620), .A2(n4784), .ZN(n6794) );
  AND2_X1 U5080 ( .A1(n5632), .A2(n5619), .ZN(n4784) );
  INV_X1 U5081 ( .A(n6796), .ZN(n5632) );
  INV_X1 U5082 ( .A(n5753), .ZN(n4770) );
  INV_X1 U5083 ( .A(n7389), .ZN(n4766) );
  NAND2_X1 U5084 ( .A1(n4403), .A2(n5738), .ZN(n4402) );
  INV_X1 U5085 ( .A(n4405), .ZN(n4403) );
  NAND2_X1 U5086 ( .A1(n4296), .A2(n4404), .ZN(n4399) );
  INV_X1 U5087 ( .A(n5738), .ZN(n4404) );
  NAND2_X1 U5088 ( .A1(n4781), .A2(n4306), .ZN(n7125) );
  INV_X1 U5089 ( .A(n4388), .ZN(n4387) );
  OAI21_X1 U5090 ( .B1(n4785), .B2(n4389), .A(n8258), .ZN(n4388) );
  INV_X1 U5091 ( .A(n4571), .ZN(n4570) );
  NAND2_X1 U5092 ( .A1(n7991), .A2(n8480), .ZN(n7983) );
  AOI21_X1 U5093 ( .B1(n7938), .B2(n4448), .A(n7937), .ZN(n7943) );
  AOI21_X1 U5094 ( .B1(n8447), .B2(n6038), .A(n5971), .ZN(n8162) );
  AND4_X1 U5095 ( .A1(n5735), .A2(n5734), .A3(n5733), .A4(n5732), .ZN(n7286)
         );
  AND4_X1 U5096 ( .A1(n5642), .A2(n5641), .A3(n5640), .A4(n5639), .ZN(n6798)
         );
  OR2_X1 U5097 ( .A1(n6492), .A2(n6491), .ZN(n4527) );
  OR2_X1 U5098 ( .A1(n6479), .A2(n6478), .ZN(n4523) );
  NAND2_X1 U5099 ( .A1(n6738), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4520) );
  NOR2_X1 U5100 ( .A1(n7008), .A2(n4356), .ZN(n7013) );
  AND2_X1 U5101 ( .A1(n7324), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4525) );
  OR2_X1 U5102 ( .A1(n5983), .A2(n5982), .ZN(n6131) );
  NAND2_X1 U5103 ( .A1(n8455), .A2(n7916), .ZN(n8440) );
  NAND2_X1 U5104 ( .A1(n8469), .A2(n6121), .ZN(n8455) );
  NAND2_X1 U5105 ( .A1(n6110), .A2(n4309), .ZN(n4563) );
  NAND2_X1 U5106 ( .A1(n7708), .A2(n4564), .ZN(n4559) );
  NAND2_X1 U5107 ( .A1(n7967), .A2(n4517), .ZN(n4510) );
  NAND2_X1 U5108 ( .A1(n4512), .A2(n7967), .ZN(n4511) );
  INV_X1 U5109 ( .A(n4513), .ZN(n4512) );
  NAND2_X1 U5110 ( .A1(n7556), .A2(n7962), .ZN(n4584) );
  AND2_X1 U5111 ( .A1(n6069), .A2(n6068), .ZN(n4519) );
  NAND3_X1 U5112 ( .A1(n8598), .A2(n4307), .A3(n6061), .ZN(n9952) );
  NAND2_X1 U5113 ( .A1(n9969), .A2(n4292), .ZN(n7167) );
  NAND2_X1 U5114 ( .A1(n5592), .A2(n4482), .ZN(n4483) );
  OR2_X1 U5115 ( .A1(n6834), .A2(n6088), .ZN(n7095) );
  NAND2_X1 U5116 ( .A1(n4491), .A2(n7974), .ZN(n4490) );
  INV_X1 U5117 ( .A(n4496), .ZN(n4491) );
  NAND2_X1 U5118 ( .A1(n7926), .A2(n7925), .ZN(n7974) );
  NAND2_X1 U5119 ( .A1(n4493), .A2(n4486), .ZN(n4485) );
  NAND2_X1 U5120 ( .A1(n4496), .A2(n4488), .ZN(n4486) );
  NAND2_X1 U5121 ( .A1(n7743), .A2(n5706), .ZN(n5979) );
  NOR2_X1 U5122 ( .A1(n4312), .A2(n4498), .ZN(n4497) );
  INV_X1 U5123 ( .A(n4503), .ZN(n4498) );
  OR2_X1 U5124 ( .A1(n4501), .A2(n4312), .ZN(n4499) );
  AND2_X1 U5125 ( .A1(n8439), .A2(n4502), .ZN(n4501) );
  NAND2_X1 U5126 ( .A1(n8456), .A2(n4503), .ZN(n4502) );
  NAND2_X1 U5127 ( .A1(n6082), .A2(n4504), .ZN(n4503) );
  AND2_X1 U5128 ( .A1(n7915), .A2(n7916), .ZN(n8456) );
  NAND2_X1 U5129 ( .A1(n8226), .A2(n4506), .ZN(n4505) );
  NAND2_X1 U5130 ( .A1(n5771), .A2(n5770), .ZN(n8680) );
  AND2_X1 U5131 ( .A1(n6004), .A2(n7648), .ZN(n10012) );
  OR2_X1 U5132 ( .A1(n7572), .A2(n6003), .ZN(n6004) );
  XNOR2_X1 U5133 ( .A(n5566), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7980) );
  INV_X1 U5134 ( .A(n4410), .ZN(n4407) );
  OR2_X1 U5135 ( .A1(n5567), .A2(n6000), .ZN(n5572) );
  NOR3_X1 U5136 ( .A1(n5812), .A2(P2_IR_REG_16__SCAN_IN), .A3(n5564), .ZN(
        n5567) );
  INV_X1 U5137 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5571) );
  NAND2_X1 U5138 ( .A1(n5739), .A2(n4788), .ZN(n5812) );
  NAND2_X1 U5139 ( .A1(n7689), .A2(n4628), .ZN(n4620) );
  INV_X1 U5140 ( .A(n4629), .ZN(n4628) );
  AND2_X1 U5141 ( .A1(n4848), .A2(n8817), .ZN(n8771) );
  NAND2_X1 U5142 ( .A1(n7689), .A2(n7685), .ZN(n4626) );
  NAND2_X1 U5143 ( .A1(n4642), .A2(n4640), .ZN(n4639) );
  OAI22_X1 U5144 ( .A1(n7263), .A2(n6557), .B1(n6556), .B2(n6658), .ZN(n6558)
         );
  NAND2_X1 U5145 ( .A1(n4636), .A2(n8071), .ZN(n4635) );
  NAND2_X1 U5146 ( .A1(n4642), .A2(n4643), .ZN(n4636) );
  AOI21_X1 U5147 ( .B1(n4638), .B2(n4643), .A(n8789), .ZN(n4637) );
  INV_X1 U5148 ( .A(n4639), .ZN(n4638) );
  NAND2_X1 U5149 ( .A1(n4637), .A2(n4639), .ZN(n4632) );
  OR2_X1 U5150 ( .A1(n4635), .A2(n4642), .ZN(n4633) );
  NAND2_X1 U5151 ( .A1(n9069), .A2(n9065), .ZN(n9229) );
  NAND2_X1 U5152 ( .A1(n5488), .A2(n9878), .ZN(n6554) );
  OR2_X1 U5153 ( .A1(n9525), .A2(n9075), .ZN(n9230) );
  XNOR2_X1 U5154 ( .A(n6223), .B(n4463), .ZN(n6580) );
  INV_X1 U5155 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n4463) );
  NAND2_X1 U5156 ( .A1(n6641), .A2(n6605), .ZN(n6178) );
  NOR2_X1 U5157 ( .A1(n6611), .A2(n4315), .ZN(n9747) );
  NAND2_X1 U5158 ( .A1(n9747), .A2(n9748), .ZN(n9746) );
  NOR2_X1 U5159 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n4609) );
  NOR2_X1 U5160 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n4608) );
  AND2_X1 U5161 ( .A1(n4959), .A2(n4606), .ZN(n4607) );
  NAND2_X1 U5162 ( .A1(n6519), .A2(n6520), .ZN(n6518) );
  NAND2_X1 U5163 ( .A1(n6518), .A2(n4456), .ZN(n9776) );
  NAND2_X1 U5164 ( .A1(n6208), .A2(n4457), .ZN(n4456) );
  OAI21_X1 U5165 ( .B1(n9816), .B2(n4459), .A(n4458), .ZN(n9827) );
  NAND2_X1 U5166 ( .A1(n4462), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n4459) );
  NAND2_X1 U5167 ( .A1(n9267), .A2(n4462), .ZN(n4458) );
  INV_X1 U5168 ( .A(n9828), .ZN(n4462) );
  OR2_X1 U5169 ( .A1(n9816), .A2(n7599), .ZN(n4461) );
  NAND2_X1 U5170 ( .A1(n4551), .A2(n4550), .ZN(n9297) );
  INV_X1 U5171 ( .A(n9356), .ZN(n9320) );
  OR2_X1 U5172 ( .A1(n9535), .A2(n9320), .ZN(n9316) );
  AND2_X1 U5173 ( .A1(n9167), .A2(n9060), .ZN(n9317) );
  NOR2_X1 U5174 ( .A1(n9317), .A2(n4692), .ZN(n4691) );
  INV_X1 U5175 ( .A(n4692), .ZN(n4690) );
  OR2_X1 U5176 ( .A1(n9543), .A2(n9382), .ZN(n9351) );
  AND2_X1 U5177 ( .A1(n8946), .A2(n9378), .ZN(n9217) );
  AND2_X1 U5178 ( .A1(n9351), .A2(n9043), .ZN(n9370) );
  OR2_X1 U5179 ( .A1(n9555), .A2(n9412), .ZN(n9378) );
  NAND2_X1 U5180 ( .A1(n4718), .A2(n4347), .ZN(n9377) );
  NAND2_X1 U5181 ( .A1(n9390), .A2(n4343), .ZN(n4718) );
  NAND2_X1 U5182 ( .A1(n5480), .A2(n4804), .ZN(n9392) );
  INV_X1 U5183 ( .A(n9447), .ZN(n9411) );
  OR2_X1 U5184 ( .A1(n9439), .A2(n9429), .ZN(n9430) );
  INV_X1 U5185 ( .A(n4671), .ZN(n4668) );
  INV_X1 U5186 ( .A(n4675), .ZN(n4674) );
  AND2_X1 U5187 ( .A1(n9023), .A2(n9022), .ZN(n9457) );
  INV_X1 U5188 ( .A(n5276), .ZN(n4678) );
  NAND2_X1 U5189 ( .A1(n4681), .A2(n4680), .ZN(n4679) );
  INV_X1 U5190 ( .A(n9487), .ZN(n4681) );
  AND2_X1 U5191 ( .A1(n8951), .A2(n9458), .ZN(n9481) );
  NOR2_X1 U5192 ( .A1(n9508), .A2(n4823), .ZN(n4822) );
  INV_X1 U5193 ( .A(n9140), .ZN(n4823) );
  NAND2_X1 U5194 ( .A1(n7594), .A2(n9138), .ZN(n4824) );
  NOR2_X1 U5195 ( .A1(n4270), .A2(n9599), .ZN(n9515) );
  NAND2_X1 U5196 ( .A1(n9141), .A2(n9120), .ZN(n9508) );
  AND2_X1 U5197 ( .A1(n4332), .A2(n5168), .ZN(n4704) );
  AOI21_X1 U5198 ( .B1(n9098), .B2(n4708), .A(n4707), .ZN(n4706) );
  NOR2_X1 U5199 ( .A1(n7494), .A2(n9253), .ZN(n4707) );
  NOR2_X1 U5200 ( .A1(n7043), .A2(n7540), .ZN(n7110) );
  OR2_X1 U5201 ( .A1(n5116), .A2(n9098), .ZN(n7041) );
  NAND2_X1 U5202 ( .A1(n7152), .A2(n9200), .ZN(n4830) );
  AND2_X1 U5203 ( .A1(n5079), .A2(n6841), .ZN(n4713) );
  INV_X1 U5204 ( .A(n9094), .ZN(n4714) );
  NAND2_X1 U5205 ( .A1(n4793), .A2(n4791), .ZN(n4794) );
  NAND2_X1 U5206 ( .A1(n6818), .A2(n9089), .ZN(n6842) );
  INV_X1 U5207 ( .A(n9681), .ZN(n9499) );
  AND2_X1 U5208 ( .A1(n6892), .A2(n5016), .ZN(n7055) );
  INV_X1 U5209 ( .A(n9685), .ZN(n9510) );
  OR2_X1 U5210 ( .A1(n9079), .A2(n9736), .ZN(n9681) );
  INV_X1 U5211 ( .A(n5464), .ZN(n9186) );
  OAI21_X1 U5212 ( .B1(n4944), .B2(n4753), .A(n4751), .ZN(n5349) );
  INV_X1 U5213 ( .A(n4752), .ZN(n4751) );
  OAI21_X1 U5214 ( .B1(n4755), .B2(n4753), .A(n4952), .ZN(n4752) );
  NAND2_X1 U5215 ( .A1(n4754), .A2(n4947), .ZN(n4753) );
  NAND2_X1 U5216 ( .A1(n4750), .A2(n4947), .ZN(n5338) );
  NAND2_X1 U5217 ( .A1(n4944), .A2(n4755), .ZN(n4750) );
  NAND2_X1 U5218 ( .A1(n4944), .A2(n4943), .ZN(n5324) );
  NAND2_X1 U5219 ( .A1(n4731), .A2(n4736), .ZN(n5248) );
  NAND2_X1 U5220 ( .A1(n5214), .A2(n4738), .ZN(n4731) );
  OAI21_X1 U5221 ( .B1(n5214), .B2(n4740), .A(n4912), .ZN(n5230) );
  INV_X1 U5222 ( .A(P1_RD_REG_SCAN_IN), .ZN(n6391) );
  AND2_X1 U5223 ( .A1(n4909), .A2(n4908), .ZN(n5198) );
  NAND2_X1 U5224 ( .A1(n5156), .A2(n5155), .ZN(n4893) );
  INV_X1 U5225 ( .A(n4896), .ZN(n4746) );
  INV_X1 U5226 ( .A(n4745), .ZN(n4744) );
  OAI21_X1 U5227 ( .B1(n4748), .B2(n4284), .A(n4903), .ZN(n4745) );
  NOR2_X1 U5228 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5019) );
  OR2_X1 U5229 ( .A1(n5019), .A2(n9631), .ZN(n5021) );
  AND4_X1 U5230 ( .A1(n5777), .A2(n5776), .A3(n5775), .A4(n5774), .ZN(n7868)
         );
  AND2_X1 U5231 ( .A1(n8169), .A2(n8168), .ZN(n8223) );
  XNOR2_X1 U5232 ( .A(n5935), .B(n5914), .ZN(n8169) );
  INV_X1 U5233 ( .A(n5934), .ZN(n5914) );
  NAND2_X1 U5234 ( .A1(n5826), .A2(n8144), .ZN(n8149) );
  NAND2_X1 U5235 ( .A1(n7518), .A2(n7519), .ZN(n7611) );
  INV_X1 U5236 ( .A(n8273), .ZN(n8285) );
  NAND2_X1 U5237 ( .A1(n4774), .A2(n4778), .ZN(n6139) );
  NAND2_X1 U5238 ( .A1(n8205), .A2(n4341), .ZN(n4774) );
  AND2_X1 U5239 ( .A1(n8365), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4532) );
  INV_X1 U5240 ( .A(n4529), .ZN(n8391) );
  NOR2_X1 U5241 ( .A1(n8411), .A2(n10086), .ZN(n8607) );
  NAND2_X1 U5242 ( .A1(n7095), .A2(n8479), .ZN(n10009) );
  NAND2_X1 U5243 ( .A1(n5967), .A2(n5966), .ZN(n8699) );
  NAND2_X1 U5244 ( .A1(n7728), .A2(n5706), .ZN(n5967) );
  OAI21_X1 U5245 ( .B1(n4325), .B2(n4652), .A(n4647), .ZN(n4646) );
  NAND2_X1 U5246 ( .A1(n4286), .A2(n4648), .ZN(n4647) );
  NAND2_X1 U5247 ( .A1(n8150), .A2(n8151), .ZN(n4654) );
  AND4_X1 U5248 ( .A1(n5087), .A2(n5086), .A3(n5085), .A4(n5084), .ZN(n7262)
         );
  AND2_X1 U5249 ( .A1(n5066), .A2(n5065), .ZN(n4719) );
  OR2_X1 U5250 ( .A1(n5646), .A2(n5097), .ZN(n4720) );
  INV_X1 U5251 ( .A(n9355), .ZN(n9382) );
  NAND2_X1 U5252 ( .A1(n4978), .A2(n4977), .ZN(n9550) );
  NAND2_X1 U5253 ( .A1(n5204), .A2(n5203), .ZN(n9605) );
  NAND2_X1 U5254 ( .A1(n5406), .A2(n5405), .ZN(n9372) );
  NAND2_X1 U5255 ( .A1(n5003), .A2(n5002), .ZN(n9394) );
  INV_X1 U5256 ( .A(n7156), .ZN(n9257) );
  NAND2_X1 U5257 ( .A1(n9820), .A2(n9278), .ZN(n9834) );
  OR2_X1 U5258 ( .A1(n9291), .A2(n9288), .ZN(n4367) );
  NAND2_X1 U5259 ( .A1(n9292), .A2(n9878), .ZN(n4368) );
  OAI21_X1 U5260 ( .B1(n4685), .B2(n4684), .A(n4682), .ZN(n5452) );
  INV_X1 U5261 ( .A(n4688), .ZN(n4684) );
  AND2_X1 U5262 ( .A1(n4686), .A2(n4683), .ZN(n4682) );
  AND2_X1 U5263 ( .A1(n5037), .A2(n5036), .ZN(n5038) );
  OR2_X1 U5264 ( .A1(n4430), .A2(n7840), .ZN(n4429) );
  AOI21_X1 U5265 ( .B1(n4434), .B2(n7857), .A(n7856), .ZN(n4428) );
  OAI21_X1 U5266 ( .B1(n4435), .B2(n4436), .A(n4321), .ZN(n4434) );
  AOI211_X1 U5267 ( .C1(n4447), .C2(n4446), .A(n7879), .B(n7967), .ZN(n4445)
         );
  NOR2_X1 U5268 ( .A1(n7876), .A2(n7966), .ZN(n4446) );
  NAND2_X1 U5269 ( .A1(n7878), .A2(n7877), .ZN(n4447) );
  NAND2_X1 U5270 ( .A1(n7899), .A2(n7807), .ZN(n4426) );
  OAI21_X1 U5271 ( .B1(n7895), .B2(n8558), .A(n8545), .ZN(n7898) );
  NAND2_X1 U5272 ( .A1(n4422), .A2(n4424), .ZN(n4420) );
  NAND2_X1 U5273 ( .A1(n4330), .A2(n4575), .ZN(n4574) );
  INV_X1 U5274 ( .A(n4577), .ZN(n4575) );
  AOI21_X1 U5275 ( .B1(n4577), .B2(n7934), .A(n7941), .ZN(n4576) );
  OR2_X1 U5276 ( .A1(n7782), .A2(n7781), .ZN(n7786) );
  INV_X1 U5277 ( .A(n4726), .ZN(n4725) );
  OAI21_X1 U5278 ( .B1(n5424), .B2(n4727), .A(n5440), .ZN(n4726) );
  INV_X1 U5279 ( .A(n5425), .ZN(n4727) );
  AOI21_X1 U5280 ( .B1(n4736), .B2(n4734), .A(n4733), .ZN(n4732) );
  INV_X1 U5281 ( .A(n5247), .ZN(n4733) );
  INV_X1 U5282 ( .A(n4738), .ZN(n4734) );
  INV_X1 U5283 ( .A(n4736), .ZN(n4735) );
  NAND2_X1 U5284 ( .A1(n4387), .A2(n4389), .ZN(n4385) );
  NAND2_X1 U5285 ( .A1(n4778), .A2(n5965), .ZN(n4777) );
  NOR2_X1 U5286 ( .A1(n4777), .A2(n4773), .ZN(n4772) );
  INV_X1 U5287 ( .A(n4839), .ZN(n4773) );
  INV_X1 U5288 ( .A(n8157), .ZN(n4779) );
  AND2_X1 U5289 ( .A1(n4574), .A2(n8405), .ZN(n4572) );
  OAI22_X1 U5290 ( .A1(n4574), .A2(n4573), .B1(n4576), .B2(n8480), .ZN(n4571)
         );
  MUX2_X1 U5291 ( .A(n7936), .B(n7944), .S(n7807), .Z(n7937) );
  NAND2_X1 U5292 ( .A1(n8329), .A2(n4374), .ZN(n8348) );
  NAND2_X1 U5293 ( .A1(n8327), .A2(n4375), .ZN(n4374) );
  INV_X1 U5294 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n4375) );
  NOR2_X1 U5295 ( .A1(n8130), .A2(n4480), .ZN(n4479) );
  NOR2_X1 U5296 ( .A1(n5942), .A2(n8207), .ZN(n4371) );
  OR3_X1 U5297 ( .A1(n5916), .A2(n5915), .A3(n8254), .ZN(n5925) );
  NOR2_X1 U5298 ( .A1(n5880), .A2(n8240), .ZN(n4372) );
  OR2_X1 U5299 ( .A1(n7722), .A2(n4475), .ZN(n4474) );
  OR2_X1 U5300 ( .A1(n8680), .A2(n7416), .ZN(n4475) );
  INV_X1 U5301 ( .A(n7845), .ZN(n4582) );
  OR2_X1 U5302 ( .A1(n7189), .A2(n7286), .ZN(n7850) );
  INV_X1 U5303 ( .A(n10070), .ZN(n4467) );
  NAND2_X1 U5304 ( .A1(n4499), .A2(n8424), .ZN(n4496) );
  INV_X1 U5305 ( .A(n4480), .ZN(n4478) );
  OR2_X1 U5306 ( .A1(n8647), .A2(n8636), .ZN(n4468) );
  OR2_X1 U5307 ( .A1(n8636), .A2(n8226), .ZN(n7908) );
  NOR3_X1 U5308 ( .A1(n8550), .A2(n8647), .A3(n8728), .ZN(n8520) );
  NOR2_X1 U5309 ( .A1(n5564), .A2(n4411), .ZN(n4410) );
  INV_X1 U5310 ( .A(n5565), .ZN(n4411) );
  AND2_X1 U5311 ( .A1(n5739), .A2(n4789), .ZN(n5769) );
  NAND2_X1 U5312 ( .A1(n4613), .A2(n4303), .ZN(n4612) );
  NAND2_X1 U5313 ( .A1(n4295), .A2(n4615), .ZN(n4613) );
  AND2_X1 U5314 ( .A1(n9043), .A2(n9368), .ZN(n9219) );
  INV_X1 U5315 ( .A(n6697), .ZN(n6420) );
  NOR2_X1 U5316 ( .A1(n9802), .A2(n4355), .ZN(n9263) );
  OR2_X1 U5317 ( .A1(n9306), .A2(n9321), .ZN(n9168) );
  AND2_X1 U5318 ( .A1(n9041), .A2(n9351), .ZN(n9169) );
  INV_X1 U5319 ( .A(n9219), .ZN(n4801) );
  NOR2_X1 U5320 ( .A1(n9550), .A2(n9555), .ZN(n4556) );
  NOR2_X1 U5321 ( .A1(n9543), .A2(n4555), .ZN(n4554) );
  INV_X1 U5322 ( .A(n4556), .ZN(n4555) );
  OR2_X1 U5323 ( .A1(n9446), .A2(n9084), .ZN(n4798) );
  AOI21_X1 U5324 ( .B1(n4675), .B2(n4676), .A(n4313), .ZN(n4673) );
  NOR2_X1 U5325 ( .A1(n5288), .A2(n5287), .ZN(n5286) );
  NAND2_X1 U5326 ( .A1(n7461), .A2(n4542), .ZN(n4541) );
  OR2_X1 U5327 ( .A1(n9694), .A2(n7512), .ZN(n9130) );
  NOR2_X1 U5328 ( .A1(n5154), .A2(n4709), .ZN(n4708) );
  INV_X1 U5329 ( .A(n5137), .ZN(n4709) );
  INV_X1 U5330 ( .A(n9192), .ZN(n4792) );
  NAND2_X1 U5331 ( .A1(n9413), .A2(n9404), .ZN(n9397) );
  INV_X1 U5332 ( .A(n9399), .ZN(n9413) );
  NAND2_X1 U5333 ( .A1(n4817), .A2(n8972), .ZN(n9678) );
  NAND2_X1 U5334 ( .A1(n7105), .A2(n9129), .ZN(n4817) );
  NAND2_X1 U5335 ( .A1(n9678), .A2(n9679), .ZN(n9677) );
  NAND2_X1 U5336 ( .A1(n6414), .A2(n9434), .ZN(n9068) );
  INV_X1 U5337 ( .A(SI_30_), .ZN(n4761) );
  INV_X1 U5338 ( .A(n5337), .ZN(n4754) );
  NOR2_X1 U5339 ( .A1(n4948), .A2(n4756), .ZN(n4755) );
  INV_X1 U5340 ( .A(n4943), .ZN(n4756) );
  NOR2_X1 U5341 ( .A1(n5229), .A2(n4739), .ZN(n4738) );
  INV_X1 U5342 ( .A(n4912), .ZN(n4739) );
  AOI21_X1 U5343 ( .B1(n4740), .B2(n4738), .A(n4737), .ZN(n4736) );
  INV_X1 U5344 ( .A(n4917), .ZN(n4737) );
  INV_X1 U5345 ( .A(n5213), .ZN(n4740) );
  AND2_X1 U5346 ( .A1(n5117), .A2(n4871), .ZN(n5138) );
  AND2_X1 U5347 ( .A1(n4884), .A2(n4875), .ZN(n5142) );
  OR2_X1 U5348 ( .A1(n4880), .A2(n4879), .ZN(n5118) );
  XNOR2_X1 U5349 ( .A(n4878), .B(SI_7_), .ZN(n5102) );
  INV_X1 U5350 ( .A(SI_5_), .ZN(n6334) );
  NAND2_X1 U5351 ( .A1(n8222), .A2(n4413), .ZN(n5938) );
  OR2_X1 U5352 ( .A1(n5936), .A2(n5937), .ZN(n4413) );
  AND2_X1 U5353 ( .A1(n5845), .A2(n5830), .ZN(n4785) );
  INV_X1 U5354 ( .A(n8212), .ZN(n5845) );
  NAND2_X1 U5355 ( .A1(n5817), .A2(n5816), .ZN(n5835) );
  NAND2_X1 U5356 ( .A1(n8183), .A2(n5877), .ZN(n8237) );
  OR2_X1 U5357 ( .A1(n5866), .A2(n5865), .ZN(n5880) );
  INV_X1 U5358 ( .A(n4372), .ZN(n5893) );
  NAND2_X1 U5359 ( .A1(n8192), .A2(n5902), .ZN(n5910) );
  AND2_X1 U5360 ( .A1(n5724), .A2(n4406), .ZN(n4405) );
  INV_X1 U5361 ( .A(n7118), .ZN(n4406) );
  NAND2_X1 U5362 ( .A1(n5583), .A2(n5582), .ZN(n5593) );
  XNOR2_X1 U5363 ( .A(n5615), .B(n9991), .ZN(n4382) );
  INV_X1 U5364 ( .A(n5846), .ZN(n4389) );
  AND2_X1 U5365 ( .A1(n5872), .A2(n5861), .ZN(n8258) );
  NAND2_X1 U5366 ( .A1(n4373), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5866) );
  INV_X1 U5367 ( .A(n4373), .ZN(n5852) );
  NAND2_X1 U5368 ( .A1(n4779), .A2(n5950), .ZN(n4778) );
  NAND2_X1 U5369 ( .A1(n7620), .A2(n4346), .ZN(n8280) );
  AND4_X1 U5370 ( .A1(n5840), .A2(n5839), .A3(n5838), .A4(n5837), .ZN(n8268)
         );
  AND4_X1 U5371 ( .A1(n5792), .A2(n5791), .A3(n5790), .A4(n5789), .ZN(n7709)
         );
  AND4_X1 U5372 ( .A1(n5764), .A2(n5763), .A3(n5762), .A4(n5761), .ZN(n7520)
         );
  AND4_X1 U5373 ( .A1(n5749), .A2(n5748), .A3(n5747), .A4(n5746), .ZN(n7393)
         );
  AND4_X1 U5374 ( .A1(n5681), .A2(n5680), .A3(n5679), .A4(n5678), .ZN(n6970)
         );
  AND4_X1 U5375 ( .A1(n5657), .A2(n5656), .A3(n5655), .A4(n5654), .ZN(n6871)
         );
  NOR3_X1 U5376 ( .A1(n9946), .A2(n10008), .A3(n9652), .ZN(n9651) );
  NOR2_X1 U5377 ( .A1(n9665), .A2(n9664), .ZN(n9663) );
  NAND2_X1 U5378 ( .A1(n6457), .A2(n4536), .ZN(n4535) );
  NAND2_X1 U5379 ( .A1(n6458), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4536) );
  AND2_X1 U5380 ( .A1(n6914), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4528) );
  NOR2_X1 U5381 ( .A1(n6915), .A2(n6916), .ZN(n7008) );
  NAND2_X1 U5382 ( .A1(n7013), .A2(n7012), .ZN(n7211) );
  NAND2_X1 U5383 ( .A1(n7327), .A2(n7326), .ZN(n7473) );
  NAND2_X1 U5384 ( .A1(n7473), .A2(n4524), .ZN(n7475) );
  OR2_X1 U5385 ( .A1(n7474), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4524) );
  NAND2_X1 U5386 ( .A1(n7475), .A2(n7476), .ZN(n8329) );
  XNOR2_X1 U5387 ( .A(n4529), .B(n8396), .ZN(n8383) );
  NOR2_X1 U5388 ( .A1(n5812), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5847) );
  NAND2_X1 U5389 ( .A1(n4531), .A2(n4530), .ZN(n4529) );
  NAND2_X1 U5390 ( .A1(n8381), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4530) );
  AND2_X1 U5391 ( .A1(n8463), .A2(n4476), .ZN(n8418) );
  NOR2_X1 U5392 ( .A1(n8420), .A2(n4477), .ZN(n4476) );
  INV_X1 U5393 ( .A(n4479), .ZN(n4477) );
  AOI21_X1 U5394 ( .B1(n4594), .B2(n4593), .A(n4592), .ZN(n4591) );
  INV_X1 U5395 ( .A(n7921), .ZN(n4592) );
  INV_X1 U5396 ( .A(n6121), .ZN(n4593) );
  INV_X1 U5397 ( .A(n8699), .ZN(n8446) );
  AND2_X1 U5398 ( .A1(n4504), .A2(n8475), .ZN(n8463) );
  NAND2_X1 U5399 ( .A1(n4371), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5983) );
  INV_X1 U5400 ( .A(n4371), .ZN(n5954) );
  OR2_X1 U5401 ( .A1(n8708), .A2(n8158), .ZN(n8457) );
  NOR2_X1 U5402 ( .A1(n8493), .A2(n8708), .ZN(n8475) );
  NAND2_X1 U5403 ( .A1(n4586), .A2(n6118), .ZN(n4585) );
  NAND2_X1 U5404 ( .A1(n4587), .A2(n6119), .ZN(n4586) );
  OR2_X1 U5405 ( .A1(n8647), .A2(n8196), .ZN(n8499) );
  AND2_X1 U5406 ( .A1(n8499), .A2(n7890), .ZN(n8517) );
  NAND2_X1 U5407 ( .A1(n6116), .A2(n6115), .ZN(n4590) );
  NAND2_X1 U5408 ( .A1(n4590), .A2(n4588), .ZN(n8516) );
  NAND2_X1 U5409 ( .A1(n4372), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5916) );
  INV_X1 U5410 ( .A(n4563), .ZN(n4562) );
  AOI21_X1 U5411 ( .B1(n4565), .B2(n4563), .A(n4561), .ZN(n4560) );
  AND2_X1 U5412 ( .A1(n4566), .A2(n6107), .ZN(n7767) );
  NAND2_X1 U5413 ( .A1(n7708), .A2(n7803), .ZN(n4566) );
  NOR2_X1 U5414 ( .A1(n7412), .A2(n4474), .ZN(n7714) );
  NOR2_X1 U5415 ( .A1(n7412), .A2(n4475), .ZN(n7585) );
  NAND2_X1 U5416 ( .A1(n7290), .A2(n10085), .ZN(n7412) );
  AND3_X1 U5417 ( .A1(n9979), .A2(n4280), .A3(n10078), .ZN(n7290) );
  OR2_X1 U5418 ( .A1(n5712), .A2(n5711), .ZN(n5730) );
  NAND2_X1 U5419 ( .A1(n9979), .A2(n4272), .ZN(n9960) );
  OR2_X1 U5420 ( .A1(n5696), .A2(n5695), .ZN(n5712) );
  NAND2_X1 U5421 ( .A1(n9979), .A2(n10057), .ZN(n9978) );
  INV_X1 U5422 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5675) );
  OR2_X1 U5423 ( .A1(n5676), .A2(n5675), .ZN(n5696) );
  AND2_X1 U5424 ( .A1(n9965), .A2(n7837), .ZN(n8600) );
  NOR2_X1 U5425 ( .A1(n7954), .A2(n7829), .ZN(n6100) );
  OR2_X1 U5426 ( .A1(n7075), .A2(n7079), .ZN(n8601) );
  NOR2_X1 U5427 ( .A1(n10034), .A2(n9991), .ZN(n6775) );
  NOR2_X1 U5428 ( .A1(n8504), .A2(n4507), .ZN(n8486) );
  NOR2_X1 U5429 ( .A1(n8250), .A2(n8509), .ZN(n4507) );
  AND2_X1 U5430 ( .A1(n7906), .A2(n6118), .ZN(n8506) );
  INV_X1 U5431 ( .A(n8517), .ZN(n8514) );
  NAND2_X1 U5432 ( .A1(n5879), .A2(n5878), .ZN(n8549) );
  NAND2_X1 U5433 ( .A1(n7576), .A2(n7946), .ZN(n7577) );
  NAND2_X1 U5434 ( .A1(n7947), .A2(n4415), .ZN(n10086) );
  OAI211_X1 U5435 ( .C1(n5592), .C2(n6512), .A(n5661), .B(n5660), .ZN(n10048)
         );
  AND2_X1 U5436 ( .A1(n4455), .A2(n4452), .ZN(n10043) );
  OR2_X1 U5437 ( .A1(n5646), .A2(n5610), .ZN(n4455) );
  AND2_X1 U5438 ( .A1(n5647), .A2(n4453), .ZN(n4452) );
  NAND2_X1 U5439 ( .A1(n4454), .A2(n6480), .ZN(n4453) );
  OR2_X1 U5440 ( .A1(n7101), .A2(n7096), .ZN(n10034) );
  AND2_X1 U5441 ( .A1(n5549), .A2(n5573), .ZN(n4567) );
  NAND2_X1 U5442 ( .A1(n4471), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5574) );
  NOR2_X1 U5443 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n4472) );
  OAI21_X1 U5444 ( .B1(n5812), .B2(n4408), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5995) );
  NAND2_X1 U5445 ( .A1(n4410), .A2(n4409), .ZN(n4408) );
  NOR2_X1 U5446 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n4409) );
  AND2_X1 U5447 ( .A1(n5739), .A2(n5540), .ZN(n5754) );
  INV_X1 U5448 ( .A(n4598), .ZN(n5725) );
  NOR2_X1 U5449 ( .A1(n4659), .A2(n4652), .ZN(n4648) );
  AND2_X1 U5450 ( .A1(n4657), .A2(n4653), .ZN(n4652) );
  OR2_X1 U5451 ( .A1(n5148), .A2(n5147), .ZN(n5162) );
  OR2_X1 U5452 ( .A1(n4600), .A2(n8063), .ZN(n4847) );
  NAND2_X1 U5453 ( .A1(n4985), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5270) );
  INV_X1 U5454 ( .A(n5256), .ZN(n4985) );
  NAND2_X1 U5455 ( .A1(n8850), .A2(n8851), .ZN(n8849) );
  NAND2_X1 U5456 ( .A1(n4377), .A2(n4376), .ZN(n8879) );
  INV_X1 U5457 ( .A(n7680), .ZN(n4376) );
  NAND2_X1 U5458 ( .A1(n8819), .A2(n7676), .ZN(n4377) );
  NOR2_X1 U5459 ( .A1(n4644), .A2(n8067), .ZN(n8893) );
  INV_X1 U5460 ( .A(n8065), .ZN(n4644) );
  NAND2_X1 U5461 ( .A1(n4982), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5189) );
  INV_X1 U5462 ( .A(n5177), .ZN(n4982) );
  AND3_X1 U5463 ( .A1(n5024), .A2(n5023), .A3(n5022), .ZN(n6673) );
  NAND2_X1 U5464 ( .A1(n8849), .A2(n8022), .ZN(n8799) );
  NOR2_X1 U5465 ( .A1(n4624), .A2(n4627), .ZN(n4623) );
  NAND2_X1 U5466 ( .A1(n4629), .A2(n4627), .ZN(n4617) );
  NAND2_X1 U5467 ( .A1(n4279), .A2(n7683), .ZN(n4616) );
  OR2_X1 U5468 ( .A1(n5041), .A2(n5025), .ZN(n5027) );
  OR2_X1 U5469 ( .A1(n5049), .A2(n7062), .ZN(n5026) );
  NAND2_X1 U5470 ( .A1(n6174), .A2(n6175), .ZN(n6641) );
  NAND2_X1 U5471 ( .A1(n9746), .A2(n4348), .ZN(n9763) );
  NAND2_X1 U5472 ( .A1(n9763), .A2(n9762), .ZN(n9761) );
  NOR2_X1 U5473 ( .A1(n6596), .A2(n4342), .ZN(n6519) );
  OR2_X1 U5474 ( .A1(n5123), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5124) );
  AOI21_X1 U5475 ( .B1(n9776), .B2(n9775), .A(n6166), .ZN(n6170) );
  NOR2_X1 U5476 ( .A1(n6628), .A2(n4466), .ZN(n6631) );
  AND2_X1 U5477 ( .A1(n6629), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4466) );
  NOR2_X1 U5478 ( .A1(n6631), .A2(n6630), .ZN(n6683) );
  NOR2_X1 U5479 ( .A1(n6683), .A2(n4465), .ZN(n6687) );
  AND2_X1 U5480 ( .A1(n6684), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4465) );
  NAND2_X1 U5481 ( .A1(n6687), .A2(n6686), .ZN(n7363) );
  NOR2_X1 U5482 ( .A1(n9787), .A2(n4354), .ZN(n9803) );
  NOR2_X1 U5483 ( .A1(n9803), .A2(n9804), .ZN(n9802) );
  XNOR2_X1 U5484 ( .A(n9263), .B(n9275), .ZN(n7368) );
  NAND2_X1 U5485 ( .A1(n8117), .A2(n8116), .ZN(n9298) );
  NOR2_X1 U5486 ( .A1(n9297), .A2(n9298), .ZN(n9296) );
  NAND2_X1 U5487 ( .A1(n4688), .A2(n9082), .ZN(n4683) );
  NAND2_X1 U5488 ( .A1(n4687), .A2(n4294), .ZN(n4686) );
  INV_X1 U5489 ( .A(n4691), .ZN(n4687) );
  AND2_X1 U5490 ( .A1(n4689), .A2(n4294), .ZN(n4688) );
  OR2_X1 U5491 ( .A1(n9331), .A2(n9329), .ZN(n9332) );
  OAI21_X1 U5492 ( .B1(n5480), .B2(n4803), .A(n4800), .ZN(n9352) );
  INV_X1 U5493 ( .A(n9217), .ZN(n4803) );
  AOI21_X1 U5494 ( .B1(n9217), .B2(n4802), .A(n4801), .ZN(n4800) );
  INV_X1 U5495 ( .A(n4804), .ZN(n4802) );
  AND2_X1 U5496 ( .A1(n9413), .A2(n4552), .ZN(n9348) );
  AND2_X1 U5497 ( .A1(n4554), .A2(n4553), .ZN(n4552) );
  OR2_X1 U5498 ( .A1(n9082), .A2(n9081), .ZN(n9354) );
  NAND2_X1 U5499 ( .A1(n9413), .A2(n4554), .ZN(n9362) );
  INV_X1 U5500 ( .A(n4715), .ZN(n9361) );
  OAI21_X1 U5501 ( .B1(n9377), .B2(n4717), .A(n4716), .ZN(n4715) );
  AND2_X1 U5502 ( .A1(n9550), .A2(n9394), .ZN(n4717) );
  NAND2_X1 U5503 ( .A1(n9387), .A2(n5481), .ZN(n4716) );
  NAND2_X1 U5504 ( .A1(n4987), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5359) );
  OR2_X1 U5505 ( .A1(n5359), .A2(n4988), .ZN(n5380) );
  INV_X1 U5506 ( .A(n4664), .ZN(n4663) );
  NAND2_X1 U5507 ( .A1(n4986), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5357) );
  INV_X1 U5508 ( .A(n5341), .ZN(n4986) );
  INV_X1 U5509 ( .A(n9246), .ZN(n9412) );
  NAND2_X1 U5510 ( .A1(n4797), .A2(n4795), .ZN(n9409) );
  AOI21_X1 U5511 ( .B1(n4285), .B2(n9084), .A(n4796), .ZN(n4795) );
  INV_X1 U5512 ( .A(n9031), .ZN(n4796) );
  AND2_X1 U5513 ( .A1(n4798), .A2(n9085), .ZN(n9423) );
  NAND2_X1 U5514 ( .A1(n4798), .A2(n4285), .ZN(n9422) );
  NOR2_X1 U5515 ( .A1(n9570), .A2(n4545), .ZN(n4543) );
  OR2_X1 U5516 ( .A1(n5270), .A2(n5269), .ZN(n5288) );
  NAND2_X1 U5517 ( .A1(n9516), .A2(n4547), .ZN(n9474) );
  AOI21_X1 U5518 ( .B1(n4822), .B2(n4820), .A(n4819), .ZN(n4818) );
  INV_X1 U5519 ( .A(n4822), .ZN(n4821) );
  INV_X1 U5520 ( .A(n9138), .ZN(n4820) );
  NAND2_X1 U5521 ( .A1(n9516), .A2(n9494), .ZN(n9488) );
  AND2_X1 U5522 ( .A1(n9515), .A2(n9520), .ZN(n9516) );
  NAND2_X1 U5523 ( .A1(n4984), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5238) );
  INV_X1 U5524 ( .A(n5221), .ZN(n4984) );
  OAI21_X1 U5525 ( .B1(n5169), .B2(n4697), .A(n4695), .ZN(n7546) );
  AOI21_X1 U5526 ( .B1(n4699), .B2(n4696), .A(n4319), .ZN(n4695) );
  INV_X1 U5527 ( .A(n4699), .ZN(n4697) );
  NAND2_X1 U5528 ( .A1(n4983), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5206) );
  INV_X1 U5529 ( .A(n5189), .ZN(n4983) );
  OR2_X1 U5530 ( .A1(n5206), .A2(n5205), .ZN(n5221) );
  INV_X1 U5531 ( .A(n9250), .ZN(n8885) );
  NAND2_X1 U5532 ( .A1(n4700), .A2(n4698), .ZN(n7451) );
  INV_X1 U5533 ( .A(n4701), .ZN(n4698) );
  NAND2_X1 U5534 ( .A1(n5169), .A2(n4702), .ZN(n4700) );
  NOR3_X1 U5535 ( .A1(n9695), .A2(n8830), .A3(n8914), .ZN(n7459) );
  AOI21_X1 U5536 ( .B1(n9679), .B2(n4816), .A(n4351), .ZN(n4815) );
  NOR2_X1 U5537 ( .A1(n9695), .A2(n8914), .ZN(n7312) );
  OR2_X1 U5538 ( .A1(n7111), .A2(n9694), .ZN(n9695) );
  OAI21_X1 U5539 ( .B1(n7152), .B2(n4828), .A(n4825), .ZN(n7048) );
  INV_X1 U5540 ( .A(n4826), .ZN(n4825) );
  OAI21_X1 U5541 ( .B1(n4828), .B2(n9200), .A(n9122), .ZN(n4826) );
  NAND2_X1 U5542 ( .A1(n4981), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5148) );
  INV_X1 U5543 ( .A(n5130), .ZN(n4981) );
  NAND2_X1 U5544 ( .A1(n6940), .A2(n4277), .ZN(n7043) );
  NAND2_X1 U5545 ( .A1(n4979), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5109) );
  NAND2_X1 U5546 ( .A1(n7145), .A2(n5100), .ZN(n6990) );
  NAND2_X1 U5547 ( .A1(n6940), .A2(n4538), .ZN(n7149) );
  NAND2_X1 U5548 ( .A1(n6940), .A2(n9874), .ZN(n7147) );
  NAND2_X1 U5549 ( .A1(n9199), .A2(n9196), .ZN(n9094) );
  AND4_X1 U5550 ( .A1(n5078), .A2(n5077), .A3(n5076), .A4(n5075), .ZN(n6849)
         );
  INV_X1 U5551 ( .A(n6673), .ZN(n7059) );
  OR2_X1 U5552 ( .A1(n7056), .A2(n7059), .ZN(n7058) );
  NAND2_X1 U5553 ( .A1(n5015), .A2(n5014), .ZN(n6892) );
  NAND2_X1 U5554 ( .A1(n5050), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4807) );
  NAND2_X1 U5555 ( .A1(n5051), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n4806) );
  NAND2_X1 U5556 ( .A1(n5415), .A2(n5414), .ZN(n9535) );
  NAND2_X1 U5557 ( .A1(n7607), .A2(n8114), .ZN(n5398) );
  AND3_X1 U5558 ( .A1(n5073), .A2(n5072), .A3(n5071), .ZN(n9912) );
  INV_X1 U5559 ( .A(n9921), .ZN(n9713) );
  XNOR2_X1 U5560 ( .A(n7790), .B(SI_30_), .ZN(n8763) );
  XNOR2_X1 U5561 ( .A(n7782), .B(n5444), .ZN(n8766) );
  XNOR2_X1 U5562 ( .A(n5408), .B(n5407), .ZN(n7607) );
  NAND2_X1 U5563 ( .A1(n4758), .A2(n5369), .ZN(n5388) );
  NAND2_X1 U5564 ( .A1(n5349), .A2(n4957), .ZN(n5352) );
  NAND2_X1 U5565 ( .A1(n5217), .A2(n4604), .ZN(n5295) );
  NAND2_X1 U5566 ( .A1(n4893), .A2(n4748), .ZN(n4747) );
  NAND2_X1 U5567 ( .A1(n4893), .A2(n4892), .ZN(n5171) );
  NAND2_X1 U5568 ( .A1(n4329), .A2(n4861), .ZN(n5093) );
  XNOR2_X1 U5569 ( .A(n4860), .B(n6334), .ZN(n5060) );
  AND2_X1 U5570 ( .A1(n5034), .A2(n5020), .ZN(n4790) );
  AND2_X1 U5571 ( .A1(n4959), .A2(n5020), .ZN(n4610) );
  NAND2_X1 U5572 ( .A1(n4856), .A2(n4855), .ZN(n5032) );
  NAND2_X1 U5573 ( .A1(n7448), .A2(n4721), .ZN(n4508) );
  NAND2_X1 U5574 ( .A1(n7447), .A2(n6391), .ZN(n4509) );
  INV_X1 U5575 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4721) );
  INV_X1 U5576 ( .A(n5674), .ZN(n4396) );
  NAND2_X1 U5577 ( .A1(n6794), .A2(n4392), .ZN(n4397) );
  NAND2_X1 U5578 ( .A1(n7125), .A2(n5724), .ZN(n7119) );
  OAI21_X1 U5579 ( .B1(n6724), .B2(n6723), .A(n4379), .ZN(n6730) );
  NAND2_X1 U5580 ( .A1(n4381), .A2(n4380), .ZN(n4379) );
  INV_X1 U5581 ( .A(n4382), .ZN(n4380) );
  INV_X1 U5582 ( .A(n5602), .ZN(n4381) );
  OR2_X1 U5583 ( .A1(n6021), .A2(n6020), .ZN(n6022) );
  NAND2_X1 U5584 ( .A1(n4391), .A2(n4390), .ZN(n6968) );
  AOI21_X1 U5585 ( .B1(n5674), .B2(n4395), .A(n4327), .ZN(n4390) );
  NAND2_X1 U5586 ( .A1(n4767), .A2(n5753), .ZN(n7390) );
  NAND2_X1 U5587 ( .A1(n7297), .A2(n7296), .ZN(n4767) );
  NAND2_X1 U5588 ( .A1(n5939), .A2(n4412), .ZN(n8205) );
  AND2_X1 U5589 ( .A1(n5938), .A2(n4839), .ZN(n4412) );
  NAND2_X1 U5590 ( .A1(n8205), .A2(n8204), .ZN(n8156) );
  NAND2_X1 U5591 ( .A1(n5815), .A2(n5814), .ZN(n8143) );
  NAND2_X1 U5592 ( .A1(n6794), .A2(n5633), .ZN(n6952) );
  NAND2_X1 U5593 ( .A1(n8149), .A2(n4785), .ZN(n8261) );
  NAND2_X1 U5594 ( .A1(n8149), .A2(n5830), .ZN(n8213) );
  NOR2_X1 U5595 ( .A1(n8223), .A2(n8222), .ZN(n8225) );
  NAND2_X1 U5596 ( .A1(n5620), .A2(n5619), .ZN(n6797) );
  NAND2_X1 U5597 ( .A1(n4781), .A2(n5705), .ZN(n7128) );
  NAND2_X1 U5598 ( .A1(n4400), .A2(n4398), .ZN(n7518) );
  AND2_X1 U5599 ( .A1(n4399), .A2(n4765), .ZN(n4398) );
  AOI21_X1 U5600 ( .B1(n4768), .B2(n4770), .A(n4766), .ZN(n4765) );
  XNOR2_X1 U5601 ( .A(n5910), .B(n5908), .ZN(n8246) );
  NAND2_X1 U5602 ( .A1(n4401), .A2(n5738), .ZN(n7297) );
  NAND2_X1 U5603 ( .A1(n7125), .A2(n4405), .ZN(n4401) );
  XNOR2_X1 U5604 ( .A(n4382), .B(n5602), .ZN(n6723) );
  NAND2_X1 U5605 ( .A1(n4383), .A2(n4387), .ZN(n8264) );
  OR2_X1 U5606 ( .A1(n8149), .A2(n4389), .ZN(n4383) );
  OR2_X1 U5607 ( .A1(n6043), .A2(n6042), .ZN(n8273) );
  INV_X1 U5608 ( .A(n8259), .ZN(n8282) );
  NAND2_X1 U5609 ( .A1(n7985), .A2(n7982), .ZN(n4370) );
  NAND2_X1 U5610 ( .A1(n4316), .A2(n4569), .ZN(n4369) );
  INV_X1 U5611 ( .A(n8133), .ZN(n7991) );
  OR2_X1 U5612 ( .A1(n6044), .A2(n5985), .ZN(n5992) );
  OR2_X1 U5613 ( .A1(n6429), .A2(n10022), .ZN(n8303) );
  OAI211_X1 U5614 ( .C1(n5989), .C2(n6440), .A(n5624), .B(n4558), .ZN(n8321)
         );
  AND2_X1 U5615 ( .A1(n5623), .A2(n5622), .ZN(n4558) );
  INV_X1 U5616 ( .A(n7832), .ZN(n8322) );
  XNOR2_X1 U5617 ( .A(n5578), .B(P2_IR_REG_1__SCAN_IN), .ZN(n9656) );
  INV_X1 U5618 ( .A(n4527), .ZN(n6490) );
  NAND2_X1 U5619 ( .A1(n6452), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4526) );
  NAND2_X1 U5620 ( .A1(n4365), .A2(n4282), .ZN(n6457) );
  AND2_X1 U5621 ( .A1(n4535), .A2(n4534), .ZN(n6473) );
  INV_X1 U5622 ( .A(n6460), .ZN(n4534) );
  INV_X1 U5623 ( .A(n4535), .ZN(n6461) );
  NOR2_X1 U5624 ( .A1(n6473), .A2(n4533), .ZN(n6505) );
  AND2_X1 U5625 ( .A1(n6480), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4533) );
  NOR2_X1 U5626 ( .A1(n6505), .A2(n6504), .ZN(n6503) );
  INV_X1 U5627 ( .A(n4523), .ZN(n6537) );
  INV_X1 U5628 ( .A(n4521), .ZN(n6734) );
  NAND2_X1 U5629 ( .A1(n4594), .A2(n8455), .ZN(n8442) );
  NAND2_X1 U5630 ( .A1(n4559), .A2(n4563), .ZN(n8577) );
  OAI22_X1 U5631 ( .A1(n7576), .A2(n4513), .B1(n4514), .B2(n6073), .ZN(n7763)
         );
  NAND2_X1 U5632 ( .A1(n4584), .A2(n6106), .ZN(n7581) );
  AND2_X1 U5633 ( .A1(n7408), .A2(n6070), .ZN(n7555) );
  AND2_X1 U5634 ( .A1(n7283), .A2(n6068), .ZN(n7409) );
  NAND2_X1 U5635 ( .A1(n7167), .A2(n7845), .ZN(n9948) );
  INV_X2 U5636 ( .A(n10009), .ZN(n10011) );
  AND2_X1 U5637 ( .A1(n10009), .A2(n6091), .ZN(n10006) );
  INV_X1 U5638 ( .A(n10120), .ZN(n10117) );
  AOI21_X1 U5639 ( .B1(n8758), .B2(n5706), .A(n7799), .ZN(n8689) );
  OAI21_X1 U5640 ( .B1(n4493), .B2(n7974), .A(n4485), .ZN(n4484) );
  NAND2_X1 U5641 ( .A1(n8454), .A2(n4300), .ZN(n4487) );
  NAND2_X1 U5642 ( .A1(n4492), .A2(n4499), .ZN(n8425) );
  NAND2_X1 U5643 ( .A1(n5864), .A2(n5863), .ZN(n8737) );
  NAND2_X1 U5644 ( .A1(n5850), .A2(n5849), .ZN(n8742) );
  NAND2_X1 U5645 ( .A1(n5834), .A2(n5833), .ZN(n8747) );
  NOR2_X1 U5646 ( .A1(n5812), .A2(n4835), .ZN(n6001) );
  XNOR2_X1 U5647 ( .A(n5997), .B(P2_IR_REG_24__SCAN_IN), .ZN(n7400) );
  XNOR2_X1 U5648 ( .A(n5995), .B(n5994), .ZN(n8133) );
  INV_X1 U5649 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6226) );
  INV_X1 U5650 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6231) );
  INV_X1 U5651 ( .A(n8150), .ZN(n4658) );
  INV_X1 U5652 ( .A(n4652), .ZN(n4651) );
  NAND2_X1 U5653 ( .A1(n4620), .A2(n4627), .ZN(n8777) );
  NAND2_X1 U5654 ( .A1(n4626), .A2(n4624), .ZN(n8780) );
  INV_X1 U5655 ( .A(n4631), .ZN(n8788) );
  AOI21_X1 U5656 ( .B1(n8065), .B2(n4642), .A(n4635), .ZN(n4631) );
  INV_X1 U5657 ( .A(n7087), .ZN(n6824) );
  NAND2_X1 U5658 ( .A1(n5427), .A2(n5426), .ZN(n9530) );
  NAND2_X1 U5659 ( .A1(n5254), .A2(n5253), .ZN(n9594) );
  NAND2_X1 U5660 ( .A1(n7030), .A2(n7258), .ZN(n7032) );
  INV_X1 U5661 ( .A(n4637), .ZN(n4634) );
  NOR2_X1 U5662 ( .A1(n5057), .A2(n5056), .ZN(n7156) );
  NOR2_X1 U5663 ( .A1(n5332), .A2(n5055), .ZN(n5056) );
  AND2_X1 U5664 ( .A1(n6567), .A2(n9736), .ZN(n8936) );
  NOR2_X1 U5665 ( .A1(n8065), .A2(n8066), .ZN(n8895) );
  NAND2_X1 U5666 ( .A1(n5285), .A2(n5284), .ZN(n9582) );
  OAI21_X1 U5667 ( .B1(n7689), .B2(n4623), .A(n4621), .ZN(n7996) );
  INV_X1 U5668 ( .A(n8945), .ZN(n8928) );
  NAND2_X1 U5669 ( .A1(n5460), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5462) );
  NAND2_X1 U5670 ( .A1(n5439), .A2(n5438), .ZN(n9245) );
  NAND2_X1 U5671 ( .A1(n5422), .A2(n5421), .ZN(n9356) );
  NAND2_X1 U5672 ( .A1(n5387), .A2(n5386), .ZN(n9355) );
  OR2_X1 U5673 ( .A1(n9364), .A2(n5049), .ZN(n5387) );
  NAND4_X1 U5674 ( .A1(n5029), .A2(n5028), .A3(n5027), .A4(n5026), .ZN(n9260)
         );
  AND2_X1 U5675 ( .A1(n6170), .A2(n6169), .ZN(n6628) );
  AND2_X1 U5676 ( .A1(n6680), .A2(n6679), .ZN(n6682) );
  INV_X1 U5677 ( .A(n4461), .ZN(n9815) );
  INV_X1 U5678 ( .A(n9267), .ZN(n4460) );
  OAI21_X1 U5679 ( .B1(n9280), .B2(n9279), .A(n9832), .ZN(n9848) );
  AND2_X1 U5680 ( .A1(n6189), .A2(n6188), .ZN(n9847) );
  NAND2_X1 U5681 ( .A1(n8113), .A2(n8112), .ZN(n9525) );
  XNOR2_X1 U5682 ( .A(n9296), .B(n4549), .ZN(n9527) );
  INV_X1 U5683 ( .A(n9525), .ZN(n4549) );
  NAND2_X1 U5684 ( .A1(n4693), .A2(n4690), .ZN(n9314) );
  NAND2_X1 U5685 ( .A1(n9392), .A2(n9217), .ZN(n9369) );
  INV_X1 U5686 ( .A(n9550), .ZN(n9387) );
  NAND2_X1 U5687 ( .A1(n5340), .A2(n5339), .ZN(n9560) );
  NAND2_X1 U5688 ( .A1(n4661), .A2(n4664), .ZN(n9407) );
  NAND2_X1 U5689 ( .A1(n9438), .A2(n4667), .ZN(n4661) );
  NAND2_X1 U5690 ( .A1(n5326), .A2(n5325), .ZN(n9429) );
  NAND2_X1 U5691 ( .A1(n4669), .A2(n4667), .ZN(n9421) );
  NAND2_X1 U5692 ( .A1(n4669), .A2(n4671), .ZN(n9419) );
  NAND2_X1 U5693 ( .A1(n4672), .A2(n4675), .ZN(n9452) );
  NAND2_X1 U5694 ( .A1(n9487), .A2(n4677), .ZN(n4672) );
  NAND2_X1 U5695 ( .A1(n4679), .A2(n4677), .ZN(n9581) );
  NAND2_X1 U5696 ( .A1(n4679), .A2(n5276), .ZN(n9482) );
  NAND2_X1 U5697 ( .A1(n4824), .A2(n9140), .ZN(n9507) );
  NAND2_X1 U5698 ( .A1(n5236), .A2(n5235), .ZN(n9599) );
  NAND2_X1 U5699 ( .A1(n5219), .A2(n5218), .ZN(n8977) );
  INV_X1 U5700 ( .A(n9308), .ZN(n9504) );
  NAND2_X1 U5701 ( .A1(n5169), .A2(n4704), .ZN(n4845) );
  NAND2_X1 U5702 ( .A1(n5169), .A2(n5168), .ZN(n7219) );
  NAND2_X1 U5703 ( .A1(n7041), .A2(n5137), .ZN(n7104) );
  NAND2_X1 U5704 ( .A1(n4830), .A2(n5473), .ZN(n6992) );
  AND3_X1 U5705 ( .A1(n4711), .A2(n4712), .A3(n5080), .ZN(n7146) );
  AND2_X1 U5706 ( .A1(n4711), .A2(n4712), .ZN(n6847) );
  INV_X1 U5707 ( .A(n9912), .ZN(n6947) );
  AND2_X1 U5708 ( .A1(n9885), .A2(n6937), .ZN(n9693) );
  NOR2_X1 U5709 ( .A1(n9311), .A2(n5499), .ZN(n5500) );
  INV_X2 U5710 ( .A(n9927), .ZN(n9929) );
  INV_X1 U5711 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9631) );
  NOR2_X1 U5712 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n4799) );
  XNOR2_X1 U5713 ( .A(n5441), .B(n5440), .ZN(n7743) );
  NAND2_X1 U5714 ( .A1(n4724), .A2(n5425), .ZN(n5441) );
  NAND2_X1 U5715 ( .A1(n5423), .A2(n5424), .ZN(n4724) );
  XNOR2_X1 U5716 ( .A(n4976), .B(n4991), .ZN(n7745) );
  XNOR2_X1 U5717 ( .A(n5423), .B(n5424), .ZN(n7728) );
  OR2_X1 U5718 ( .A1(n5457), .A2(n5456), .ZN(n5458) );
  OAI21_X1 U5719 ( .B1(n4893), .B2(n4284), .A(n4744), .ZN(n5199) );
  INV_X1 U5720 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6229) );
  XNOR2_X1 U5721 ( .A(n5092), .B(n5067), .ZN(n6220) );
  XNOR2_X1 U5722 ( .A(n5035), .B(n5034), .ZN(n6604) );
  OAI21_X1 U5723 ( .B1(n5021), .B2(n5020), .A(n5033), .ZN(n6636) );
  XNOR2_X1 U5724 ( .A(n5006), .B(n4464), .ZN(n6223) );
  NAND2_X1 U5725 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4464) );
  NAND2_X1 U5726 ( .A1(n8699), .A2(n8290), .ZN(n6150) );
  INV_X1 U5727 ( .A(n4531), .ZN(n8380) );
  MUX2_X1 U5728 ( .A(n8407), .B(n8406), .S(n8405), .Z(n8409) );
  OAI211_X1 U5729 ( .C1(n4660), .C2(n4650), .A(n4649), .B(n4645), .ZN(P1_U3212) );
  NAND2_X1 U5730 ( .A1(n4286), .A2(n4651), .ZN(n4650) );
  INV_X1 U5731 ( .A(n4646), .ZN(n4645) );
  OR2_X1 U5732 ( .A1(n8933), .A2(n4273), .ZN(n4649) );
  NAND2_X1 U5733 ( .A1(n4368), .A2(n4366), .ZN(n9294) );
  INV_X1 U5734 ( .A(n7936), .ZN(n7976) );
  NAND2_X1 U5735 ( .A1(n7939), .A2(n7930), .ZN(n7936) );
  OR3_X1 U5736 ( .A1(n9695), .A2(n8830), .A3(n4540), .ZN(n4270) );
  OR3_X1 U5737 ( .A1(n7412), .A2(n4474), .A3(n8291), .ZN(n4271) );
  NAND2_X1 U5738 ( .A1(n5592), .A2(n7794), .ZN(n5610) );
  AND2_X1 U5739 ( .A1(n10057), .A2(n10062), .ZN(n4272) );
  NAND2_X1 U5740 ( .A1(n4326), .A2(n4651), .ZN(n4273) );
  AND2_X1 U5741 ( .A1(n7893), .A2(n7807), .ZN(n4274) );
  AND2_X1 U5742 ( .A1(n9582), .A2(n9500), .ZN(n4275) );
  OR3_X1 U5743 ( .A1(n8550), .A2(n4469), .A3(n8647), .ZN(n4276) );
  INV_X1 U5744 ( .A(n7887), .ZN(n4561) );
  INV_X1 U5745 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6000) );
  NAND2_X1 U5746 ( .A1(n5314), .A2(n5313), .ZN(n9570) );
  AND2_X1 U5747 ( .A1(n4538), .A2(n4537), .ZN(n4277) );
  INV_X1 U5748 ( .A(n6870), .ZN(n4395) );
  INV_X1 U5749 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5549) );
  AND2_X1 U5750 ( .A1(n4634), .A2(n4635), .ZN(n4278) );
  AND2_X1 U5751 ( .A1(n4272), .A2(n4467), .ZN(n4280) );
  NAND2_X1 U5752 ( .A1(n5577), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4281) );
  NAND2_X1 U5753 ( .A1(n5979), .A2(n5978), .ZN(n8616) );
  INV_X1 U5754 ( .A(n8616), .ZN(n4481) );
  INV_X1 U5755 ( .A(n6082), .ZN(n8298) );
  AND2_X1 U5756 ( .A1(n5960), .A2(n5959), .ZN(n6082) );
  INV_X1 U5757 ( .A(n7947), .ZN(n7979) );
  XNOR2_X1 U5758 ( .A(n5570), .B(n5569), .ZN(n7947) );
  NAND2_X1 U5759 ( .A1(n5913), .A2(n5912), .ZN(n8715) );
  AND2_X1 U5760 ( .A1(n5932), .A2(n5931), .ZN(n8226) );
  AND2_X1 U5761 ( .A1(n6424), .A2(n6696), .ZN(n8935) );
  INV_X1 U5762 ( .A(n8935), .ZN(n4653) );
  XOR2_X1 U5763 ( .A(n6465), .B(n6447), .Z(n4282) );
  NOR2_X1 U5764 ( .A1(n5196), .A2(n9101), .ZN(n4283) );
  OR2_X1 U5765 ( .A1(n5183), .A2(n4746), .ZN(n4284) );
  AND2_X1 U5766 ( .A1(n9424), .A2(n9085), .ZN(n4285) );
  OR2_X1 U5767 ( .A1(n8892), .A2(n8066), .ZN(n4642) );
  AND2_X1 U5768 ( .A1(n4658), .A2(n4655), .ZN(n4286) );
  NOR2_X1 U5769 ( .A1(n7690), .A2(n8772), .ZN(n4287) );
  AND2_X1 U5770 ( .A1(n4521), .A2(n4520), .ZN(n4288) );
  OR2_X1 U5771 ( .A1(n7181), .A2(n7959), .ZN(n4289) );
  AND2_X1 U5772 ( .A1(n4656), .A2(n4286), .ZN(n4290) );
  NAND2_X1 U5773 ( .A1(n9570), .A2(n9463), .ZN(n4291) );
  AND2_X1 U5774 ( .A1(n7957), .A2(n7842), .ZN(n4292) );
  AND3_X1 U5775 ( .A1(n4607), .A2(n4608), .A3(n4609), .ZN(n5089) );
  NAND2_X1 U5776 ( .A1(n7663), .A2(n7662), .ZN(n4293) );
  NAND2_X1 U5777 ( .A1(n9530), .A2(n9245), .ZN(n4294) );
  INV_X1 U5778 ( .A(n7946), .ZN(n4516) );
  XNOR2_X1 U5779 ( .A(n8699), .B(n8162), .ZN(n8439) );
  INV_X1 U5780 ( .A(n9033), .ZN(n4805) );
  AND2_X1 U5781 ( .A1(n8039), .A2(n4614), .ZN(n4295) );
  AND2_X1 U5782 ( .A1(n4768), .A2(n4402), .ZN(n4296) );
  NAND2_X1 U5783 ( .A1(n5694), .A2(n5693), .ZN(n7176) );
  NAND2_X1 U5784 ( .A1(n5552), .A2(n5550), .ZN(n5555) );
  OR3_X1 U5785 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .A3(
        P2_IR_REG_1__SCAN_IN), .ZN(n4297) );
  OR2_X1 U5786 ( .A1(n8893), .A2(n8892), .ZN(n4298) );
  AND3_X1 U5787 ( .A1(n7902), .A2(n8499), .A3(n7904), .ZN(n4299) );
  AND2_X1 U5788 ( .A1(n4493), .A2(n4488), .ZN(n4300) );
  NOR3_X1 U5789 ( .A1(n8550), .A2(n4469), .A3(n4468), .ZN(n4470) );
  AND3_X1 U5790 ( .A1(n5606), .A2(n5605), .A3(n5604), .ZN(n4301) );
  OR3_X1 U5791 ( .A1(n10027), .A2(n7979), .A3(n8480), .ZN(n5643) );
  NAND2_X1 U5792 ( .A1(n4790), .A2(n5019), .ZN(n5068) );
  AND2_X1 U5793 ( .A1(n9667), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4302) );
  NAND2_X1 U5794 ( .A1(n5268), .A2(n5267), .ZN(n9587) );
  NAND2_X1 U5795 ( .A1(n5804), .A2(n5803), .ZN(n8291) );
  XNOR2_X1 U5796 ( .A(n4865), .B(SI_6_), .ZN(n5095) );
  INV_X1 U5797 ( .A(n9555), .ZN(n9404) );
  NAND2_X1 U5798 ( .A1(n5355), .A2(n5354), .ZN(n9555) );
  INV_X1 U5799 ( .A(n4551), .ZN(n9322) );
  NOR2_X1 U5800 ( .A1(n9338), .A2(n9530), .ZN(n4551) );
  INV_X1 U5801 ( .A(n5607), .ZN(n5989) );
  NAND2_X1 U5802 ( .A1(n6084), .A2(n6083), .ZN(n8130) );
  INV_X1 U5803 ( .A(n7038), .ZN(n9874) );
  NAND2_X1 U5804 ( .A1(n4720), .A2(n4719), .ZN(n7038) );
  AND2_X1 U5805 ( .A1(n8038), .A2(n8866), .ZN(n4303) );
  AND2_X1 U5806 ( .A1(n5480), .A2(n9033), .ZN(n4304) );
  INV_X1 U5807 ( .A(n5277), .ZN(n4680) );
  OR2_X1 U5808 ( .A1(n5592), .A2(n6465), .ZN(n4305) );
  AND2_X1 U5809 ( .A1(n5723), .A2(n5705), .ZN(n4306) );
  NAND2_X1 U5810 ( .A1(n5377), .A2(n5376), .ZN(n9543) );
  NOR2_X1 U5811 ( .A1(n7956), .A2(n6064), .ZN(n4307) );
  AND2_X1 U5812 ( .A1(n4590), .A2(n7899), .ZN(n4308) );
  AND2_X1 U5813 ( .A1(n7852), .A2(n7847), .ZN(n9954) );
  NAND2_X1 U5814 ( .A1(n6108), .A2(n6107), .ZN(n4309) );
  NAND2_X1 U5815 ( .A1(n4370), .A2(n4369), .ZN(n4310) );
  AND2_X1 U5816 ( .A1(n7908), .A2(n4425), .ZN(n4311) );
  AND2_X1 U5817 ( .A1(n8446), .A2(n8162), .ZN(n4312) );
  NOR2_X1 U5818 ( .A1(n9575), .A2(n9472), .ZN(n4313) );
  NOR2_X1 U5819 ( .A1(n9565), .A2(n9411), .ZN(n4314) );
  INV_X1 U5820 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5294) );
  AND2_X1 U5821 ( .A1(n6616), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4315) );
  AND3_X1 U5822 ( .A1(n4568), .A2(n4570), .A3(n7987), .ZN(n4316) );
  OR2_X1 U5823 ( .A1(n8236), .A2(n8189), .ZN(n4317) );
  OR2_X1 U5824 ( .A1(n4641), .A2(n4639), .ZN(n4318) );
  NOR2_X1 U5825 ( .A1(n9605), .A2(n9249), .ZN(n4319) );
  NOR2_X1 U5826 ( .A1(n9560), .A2(n9426), .ZN(n4320) );
  AND2_X1 U5827 ( .A1(n7846), .A2(n7847), .ZN(n4321) );
  AND2_X1 U5828 ( .A1(n5217), .A2(n4603), .ZN(n5454) );
  OR2_X1 U5829 ( .A1(n4427), .A2(n4426), .ZN(n4322) );
  INV_X1 U5830 ( .A(n4545), .ZN(n4544) );
  NAND2_X1 U5831 ( .A1(n4547), .A2(n4546), .ZN(n4545) );
  INV_X1 U5832 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4473) );
  INV_X1 U5833 ( .A(n4968), .ZN(n4969) );
  NOR2_X1 U5834 ( .A1(n4967), .A2(n4966), .ZN(n4968) );
  INV_X1 U5835 ( .A(n4828), .ZN(n4827) );
  NAND2_X1 U5836 ( .A1(n4829), .A2(n5473), .ZN(n4828) );
  OR3_X1 U5837 ( .A1(n5812), .A2(P2_IR_REG_16__SCAN_IN), .A3(n4407), .ZN(n4323) );
  AND2_X1 U5838 ( .A1(n4633), .A2(n4632), .ZN(n4324) );
  AND2_X1 U5839 ( .A1(n6844), .A2(n6843), .ZN(n5079) );
  INV_X1 U5840 ( .A(n5592), .ZN(n4454) );
  AND2_X1 U5841 ( .A1(n4654), .A2(n4657), .ZN(n4325) );
  AND2_X1 U5842 ( .A1(n4659), .A2(n8150), .ZN(n4326) );
  INV_X1 U5843 ( .A(n4565), .ZN(n4564) );
  NAND2_X1 U5844 ( .A1(n6110), .A2(n7803), .ZN(n4565) );
  AND2_X1 U5845 ( .A1(n4394), .A2(n4393), .ZN(n4327) );
  AND2_X1 U5846 ( .A1(n7997), .A2(n7995), .ZN(n4328) );
  INV_X1 U5847 ( .A(n7941), .ZN(n4578) );
  NAND2_X1 U5848 ( .A1(n5058), .A2(n4864), .ZN(n4329) );
  OR2_X1 U5849 ( .A1(n7936), .A2(n8420), .ZN(n4330) );
  OR2_X1 U5850 ( .A1(n9344), .A2(n8945), .ZN(n4331) );
  OR2_X1 U5851 ( .A1(n8914), .A2(n9251), .ZN(n4332) );
  AND2_X1 U5852 ( .A1(n6119), .A2(n6115), .ZN(n4333) );
  AND2_X1 U5853 ( .A1(n4424), .A2(n4421), .ZN(n4334) );
  AND2_X1 U5854 ( .A1(n4424), .A2(n4299), .ZN(n4335) );
  NAND2_X1 U5855 ( .A1(n5786), .A2(n5785), .ZN(n7722) );
  AND2_X1 U5856 ( .A1(n4693), .A2(n4691), .ZN(n4336) );
  AND2_X1 U5857 ( .A1(n9316), .A2(n9059), .ZN(n9333) );
  INV_X1 U5858 ( .A(n9333), .ZN(n9329) );
  INV_X1 U5859 ( .A(n8776), .ZN(n4625) );
  AND2_X1 U5860 ( .A1(n5280), .A2(n5294), .ZN(n4337) );
  AND2_X1 U5861 ( .A1(n4392), .A2(n4395), .ZN(n4338) );
  NAND3_X1 U5862 ( .A1(n8647), .A2(n8196), .A3(n7904), .ZN(n4339) );
  INV_X1 U5863 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4964) );
  INV_X1 U5864 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n4414) );
  INV_X1 U5865 ( .A(n4595), .ZN(n4594) );
  NAND2_X1 U5866 ( .A1(n8437), .A2(n7916), .ZN(n4595) );
  OR2_X2 U5867 ( .A1(n7991), .A2(n7802), .ZN(n7807) );
  INV_X1 U5868 ( .A(n6245), .ZN(n5332) );
  INV_X1 U5869 ( .A(n5332), .ZN(n5491) );
  NAND2_X1 U5870 ( .A1(n7788), .A2(n7787), .ZN(n8420) );
  INV_X1 U5871 ( .A(n8420), .ZN(n4579) );
  NAND2_X1 U5872 ( .A1(n5904), .A2(n5903), .ZN(n8647) );
  AND2_X1 U5873 ( .A1(n8598), .A2(n6061), .ZN(n7161) );
  OR2_X1 U5874 ( .A1(n8550), .A2(n8728), .ZN(n4340) );
  AND2_X1 U5875 ( .A1(n4779), .A2(n8204), .ZN(n4341) );
  XNOR2_X1 U5876 ( .A(n8616), .B(n8296), .ZN(n8427) );
  NAND2_X1 U5877 ( .A1(n5891), .A2(n5890), .ZN(n8728) );
  NAND2_X1 U5878 ( .A1(n7633), .A2(n7632), .ZN(n7689) );
  AND2_X1 U5879 ( .A1(n6601), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4342) );
  NAND2_X1 U5880 ( .A1(n7577), .A2(n6072), .ZN(n7707) );
  INV_X1 U5881 ( .A(n9120), .ZN(n4819) );
  NAND2_X1 U5882 ( .A1(n5952), .A2(n5951), .ZN(n8626) );
  INV_X1 U5883 ( .A(n8626), .ZN(n4504) );
  OR2_X1 U5884 ( .A1(n9555), .A2(n9246), .ZN(n4343) );
  NAND2_X1 U5885 ( .A1(n5446), .A2(n5445), .ZN(n9306) );
  INV_X1 U5886 ( .A(n9306), .ZN(n4550) );
  INV_X1 U5887 ( .A(n4677), .ZN(n4676) );
  NOR2_X1 U5888 ( .A1(n9481), .A2(n4678), .ZN(n4677) );
  INV_X1 U5889 ( .A(n4667), .ZN(n4666) );
  NOR2_X1 U5890 ( .A1(n9424), .A2(n4668), .ZN(n4667) );
  NAND2_X1 U5891 ( .A1(n5185), .A2(n4964), .ZN(n5215) );
  NAND2_X1 U5892 ( .A1(n5217), .A2(n5216), .ZN(n5251) );
  NAND2_X1 U5893 ( .A1(n5941), .A2(n5940), .ZN(n8708) );
  NAND2_X1 U5894 ( .A1(n9516), .A2(n4544), .ZN(n4548) );
  NAND2_X1 U5895 ( .A1(n9413), .A2(n4556), .ZN(n4557) );
  NOR2_X1 U5896 ( .A1(n9538), .A2(n9372), .ZN(n9082) );
  AND3_X1 U5897 ( .A1(n5921), .A2(n5920), .A3(n5919), .ZN(n8250) );
  AND2_X1 U5898 ( .A1(n4461), .A2(n4460), .ZN(n4344) );
  AND2_X1 U5899 ( .A1(n4824), .A2(n4822), .ZN(n4345) );
  AND2_X1 U5900 ( .A1(n4780), .A2(n5798), .ZN(n4346) );
  OR2_X1 U5901 ( .A1(n9404), .A2(n9412), .ZN(n4347) );
  OR2_X1 U5902 ( .A1(n9750), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4348) );
  INV_X1 U5903 ( .A(n8151), .ZN(n4655) );
  NAND2_X1 U5904 ( .A1(n9952), .A2(n9951), .ZN(n4349) );
  AND2_X1 U5905 ( .A1(n5217), .A2(n4605), .ZN(n4350) );
  NAND2_X1 U5906 ( .A1(n5398), .A2(n5397), .ZN(n9538) );
  INV_X1 U5907 ( .A(n9538), .ZN(n4553) );
  NAND2_X1 U5908 ( .A1(n7220), .A2(n9002), .ZN(n4351) );
  AND2_X1 U5909 ( .A1(n4626), .A2(n7683), .ZN(n4352) );
  NAND2_X1 U5910 ( .A1(n5300), .A2(n5299), .ZN(n9575) );
  INV_X1 U5911 ( .A(n9575), .ZN(n4546) );
  NAND2_X1 U5912 ( .A1(n5923), .A2(n5922), .ZN(n8636) );
  INV_X1 U5913 ( .A(n8636), .ZN(n4506) );
  AND2_X1 U5914 ( .A1(n9979), .A2(n4280), .ZN(n4353) );
  AND2_X1 U5915 ( .A1(n9786), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4354) );
  INV_X1 U5916 ( .A(n8914), .ZN(n4542) );
  AND2_X1 U5917 ( .A1(n9801), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4355) );
  AND2_X1 U5918 ( .A1(n7009), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4356) );
  NAND2_X1 U5919 ( .A1(n7340), .A2(n7339), .ZN(n7486) );
  AND2_X1 U5920 ( .A1(n4397), .A2(n4396), .ZN(n4357) );
  NAND2_X1 U5921 ( .A1(n7283), .A2(n4519), .ZN(n7408) );
  OR2_X1 U5922 ( .A1(n7412), .A2(n7416), .ZN(n4358) );
  AND3_X1 U5923 ( .A1(n7030), .A2(n7258), .A3(n7031), .ZN(n4359) );
  AND2_X1 U5924 ( .A1(n6066), .A2(n9952), .ZN(n7179) );
  NAND2_X1 U5925 ( .A1(n4599), .A2(n4596), .ZN(n5998) );
  XNOR2_X1 U5926 ( .A(n5462), .B(P1_IR_REG_22__SCAN_IN), .ZN(n5488) );
  NAND2_X1 U5927 ( .A1(n7269), .A2(n7270), .ZN(n7340) );
  NOR2_X1 U5928 ( .A1(n8414), .A2(n5579), .ZN(n4360) );
  INV_X1 U5929 ( .A(n4539), .ZN(n7547) );
  NOR3_X1 U5930 ( .A1(n9695), .A2(n8830), .A3(n4541), .ZN(n4539) );
  AND2_X1 U5931 ( .A1(n4830), .A2(n4827), .ZN(n4361) );
  NAND2_X1 U5932 ( .A1(n5847), .A2(n6279), .ZN(n4362) );
  AND2_X1 U5933 ( .A1(n8971), .A2(n9123), .ZN(n9098) );
  AND2_X1 U5934 ( .A1(n5443), .A2(n5442), .ZN(n4363) );
  AND2_X1 U5935 ( .A1(n9969), .A2(n7842), .ZN(n4364) );
  XNOR2_X1 U5936 ( .A(n5572), .B(n5571), .ZN(n8405) );
  INV_X1 U5937 ( .A(n7350), .ZN(n4537) );
  XNOR2_X1 U5938 ( .A(n5574), .B(n5573), .ZN(n6034) );
  AND2_X1 U5939 ( .A1(n5593), .A2(n5586), .ZN(n6746) );
  INV_X1 U5940 ( .A(n9878), .ZN(n9434) );
  INV_X2 U5941 ( .A(n7794), .ZN(n6203) );
  NAND2_X1 U5942 ( .A1(n5579), .A2(n8133), .ZN(n10027) );
  NAND2_X1 U5943 ( .A1(n4527), .A2(n4526), .ZN(n4365) );
  NOR2_X1 U5944 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n7447) );
  INV_X1 U5945 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4606) );
  INV_X1 U5946 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n4457) );
  INV_X1 U5947 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n4417) );
  AOI21_X1 U5948 ( .B1(n6128), .B2(n9968), .A(n6127), .ZN(n8123) );
  NAND3_X1 U5949 ( .A1(n9287), .A2(n4367), .A3(n9434), .ZN(n4366) );
  NOR2_X1 U5950 ( .A1(n6182), .A2(n6515), .ZN(n9780) );
  NOR2_X1 U5951 ( .A1(n6620), .A2(n6619), .ZN(n6624) );
  AOI21_X1 U5952 ( .B1(n6212), .B2(n5081), .A(n6590), .ZN(n6517) );
  AOI21_X1 U5953 ( .B1(n6219), .B2(n6180), .A(n9751), .ZN(n9767) );
  AOI21_X1 U5954 ( .B1(n9275), .B2(n9721), .A(n9274), .ZN(n9277) );
  AOI21_X1 U5955 ( .B1(n7357), .B2(n7356), .A(n9808), .ZN(n7359) );
  AOI21_X1 U5956 ( .B1(n7353), .B2(n7383), .A(n7352), .ZN(n9795) );
  AOI21_X1 U5957 ( .B1(n7355), .B2(n9728), .A(n9793), .ZN(n9809) );
  NAND2_X1 U5958 ( .A1(n5758), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5772) );
  NAND2_X1 U5959 ( .A1(n5729), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5744) );
  NOR2_X1 U5960 ( .A1(n9663), .A2(n4302), .ZN(n6492) );
  NOR2_X1 U5961 ( .A1(n7323), .A2(n4525), .ZN(n7327) );
  NOR2_X1 U5962 ( .A1(n8359), .A2(n4532), .ZN(n8362) );
  NOR2_X1 U5963 ( .A1(n6913), .A2(n4528), .ZN(n6916) );
  AOI21_X1 U5964 ( .B1(n4621), .B2(n4623), .A(n4328), .ZN(n4618) );
  NOR2_X1 U5965 ( .A1(n8858), .A2(n8077), .ZN(n8834) );
  NOR2_X1 U5966 ( .A1(n8859), .A2(n8860), .ZN(n8858) );
  NAND2_X1 U5967 ( .A1(n4660), .A2(n4659), .ZN(n4656) );
  NAND2_X1 U5968 ( .A1(n4747), .A2(n4896), .ZN(n5184) );
  NAND2_X1 U5969 ( .A1(n5139), .A2(n4876), .ZN(n4886) );
  MUX2_X1 U5970 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n7794), .Z(n4860) );
  NAND2_X1 U5971 ( .A1(n4619), .A2(n4618), .ZN(n8001) );
  NAND2_X1 U5972 ( .A1(n6746), .A2(n6748), .ZN(n6747) );
  NAND2_X1 U5973 ( .A1(n6747), .A2(n5593), .ZN(n6724) );
  NAND2_X1 U5974 ( .A1(n6730), .A2(n6729), .ZN(n5620) );
  NAND2_X1 U5975 ( .A1(n8149), .A2(n4387), .ZN(n4386) );
  NAND2_X1 U5976 ( .A1(n6794), .A2(n4338), .ZN(n4391) );
  NAND2_X1 U5977 ( .A1(n7125), .A2(n4296), .ZN(n4400) );
  INV_X1 U5978 ( .A(n10027), .ZN(n4415) );
  XNOR2_X1 U5979 ( .A(n4849), .B(SI_1_), .ZN(n5005) );
  NAND2_X1 U5980 ( .A1(n7891), .A2(n4334), .ZN(n4419) );
  NAND2_X1 U5981 ( .A1(n7903), .A2(n4335), .ZN(n4418) );
  NAND3_X1 U5982 ( .A1(n4419), .A2(n4418), .A3(n4420), .ZN(n7909) );
  OAI21_X1 U5983 ( .B1(n7894), .B2(n4274), .A(n4423), .ZN(n4422) );
  INV_X1 U5984 ( .A(n7890), .ZN(n4427) );
  NAND2_X1 U5985 ( .A1(n4432), .A2(n4431), .ZN(n4430) );
  INV_X1 U5986 ( .A(n7839), .ZN(n4432) );
  NAND2_X1 U5987 ( .A1(n4859), .A2(n4437), .ZN(n4438) );
  INV_X1 U5988 ( .A(n5031), .ZN(n4437) );
  NAND3_X1 U5989 ( .A1(n4439), .A2(n4438), .A3(n5067), .ZN(n5059) );
  NAND3_X1 U5990 ( .A1(n4859), .A2(n4856), .A3(n4855), .ZN(n4439) );
  NAND2_X1 U5991 ( .A1(n5032), .A2(n5031), .ZN(n4440) );
  XNOR2_X1 U5992 ( .A(n9266), .B(n9276), .ZN(n9816) );
  INV_X1 U5993 ( .A(n4470), .ZN(n8493) );
  AND3_X1 U5994 ( .A1(n4599), .A2(n4596), .A3(n4473), .ZN(n5575) );
  NAND3_X1 U5995 ( .A1(n4599), .A2(n4596), .A3(n4472), .ZN(n4471) );
  AND2_X1 U5996 ( .A1(n8463), .A2(n4478), .ZN(n8431) );
  NAND2_X1 U5997 ( .A1(n8463), .A2(n4479), .ZN(n8419) );
  NAND2_X1 U5998 ( .A1(n8463), .A2(n8446), .ZN(n8445) );
  OAI21_X1 U5999 ( .B1(n6222), .B2(n6203), .A(n4281), .ZN(n4482) );
  NAND2_X2 U6000 ( .A1(n5592), .A2(n5577), .ZN(n7798) );
  OR2_X1 U6001 ( .A1(n8454), .A2(n4490), .ZN(n4489) );
  NAND2_X1 U6002 ( .A1(n8454), .A2(n4497), .ZN(n4492) );
  NAND3_X1 U6003 ( .A1(n4489), .A2(n4487), .A3(n4484), .ZN(n8127) );
  MUX2_X1 U6004 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n7794), .Z(n5004) );
  OAI22_X2 U6005 ( .A1(n7576), .A2(n4511), .B1(n4514), .B2(n4510), .ZN(n7765)
         );
  INV_X1 U6006 ( .A(n6073), .ZN(n4517) );
  NAND2_X1 U6007 ( .A1(n6060), .A2(n6059), .ZN(n8598) );
  INV_X1 U6008 ( .A(n9984), .ZN(n6881) );
  OAI211_X2 U6009 ( .C1(n6220), .C2(n5610), .A(n5629), .B(n4305), .ZN(n9984)
         );
  NAND2_X1 U6010 ( .A1(n7408), .A2(n4518), .ZN(n7553) );
  NOR2_X2 U6011 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5249) );
  NAND2_X1 U6012 ( .A1(n9516), .A2(n4543), .ZN(n9439) );
  INV_X1 U6013 ( .A(n4548), .ZN(n9453) );
  INV_X1 U6014 ( .A(n4557), .ZN(n9383) );
  OAI21_X1 U6015 ( .B1(n7708), .B2(n4562), .A(n4560), .ZN(n8560) );
  AND2_X1 U6016 ( .A1(n5575), .A2(n4567), .ZN(n5552) );
  NAND2_X1 U6017 ( .A1(n7789), .A2(n4572), .ZN(n4568) );
  OR2_X1 U6018 ( .A1(n7789), .A2(n4573), .ZN(n4569) );
  INV_X1 U6019 ( .A(n4581), .ZN(n4580) );
  OAI21_X1 U6020 ( .B1(n4292), .B2(n4582), .A(n9954), .ZN(n4581) );
  NAND2_X1 U6021 ( .A1(n4584), .A2(n4583), .ZN(n7579) );
  AOI21_X1 U6022 ( .B1(n6116), .B2(n4333), .A(n4585), .ZN(n8490) );
  OAI21_X1 U6023 ( .B1(n8469), .B2(n4595), .A(n4591), .ZN(n8428) );
  XNOR2_X1 U6024 ( .A(n5061), .B(n5060), .ZN(n5646) );
  OAI21_X1 U6025 ( .B1(n6423), .B2(n4600), .A(n6555), .ZN(n6653) );
  NAND2_X1 U6026 ( .A1(n6423), .A2(n4600), .ZN(n6555) );
  NAND2_X1 U6027 ( .A1(n6421), .A2(n6422), .ZN(n4600) );
  NAND3_X1 U6028 ( .A1(n4601), .A2(n6563), .A3(n6668), .ZN(n6669) );
  NAND2_X1 U6029 ( .A1(n6562), .A2(n6561), .ZN(n6668) );
  NAND2_X1 U6030 ( .A1(n4601), .A2(n6668), .ZN(n6565) );
  NAND2_X1 U6031 ( .A1(n6560), .A2(n6559), .ZN(n4601) );
  NAND2_X1 U6032 ( .A1(n7030), .A2(n7031), .ZN(n4602) );
  NAND2_X1 U6033 ( .A1(n5455), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5459) );
  NAND3_X1 U6034 ( .A1(n4610), .A2(n5034), .A3(n5019), .ZN(n5063) );
  INV_X1 U6035 ( .A(n4611), .ZN(n8050) );
  AOI21_X1 U6036 ( .B1(n8850), .B2(n4295), .A(n4612), .ZN(n4611) );
  NAND2_X1 U6037 ( .A1(n7689), .A2(n4621), .ZN(n4619) );
  NOR2_X1 U6038 ( .A1(n7684), .A2(n4625), .ZN(n4624) );
  NAND2_X1 U6039 ( .A1(n7689), .A2(n7688), .ZN(n8818) );
  INV_X1 U6040 ( .A(n8071), .ZN(n4640) );
  INV_X1 U6041 ( .A(n8933), .ZN(n4660) );
  NOR2_X1 U6042 ( .A1(n8931), .A2(n8932), .ZN(n4659) );
  OAI21_X1 U6043 ( .B1(n9438), .B2(n4663), .A(n4662), .ZN(n5348) );
  OAI21_X1 U6044 ( .B1(n9487), .B2(n4674), .A(n4673), .ZN(n5310) );
  INV_X1 U6045 ( .A(n9347), .ZN(n4685) );
  OR2_X1 U6046 ( .A1(n9347), .A2(n9082), .ZN(n4694) );
  NAND2_X1 U6047 ( .A1(n4694), .A2(n9080), .ZN(n9330) );
  NAND2_X1 U6048 ( .A1(n4694), .A2(n4689), .ZN(n4693) );
  NAND2_X1 U6049 ( .A1(n5116), .A2(n4708), .ZN(n4705) );
  NAND2_X1 U6050 ( .A1(n4705), .A2(n4706), .ZN(n9675) );
  INV_X1 U6051 ( .A(n5116), .ZN(n7042) );
  NAND3_X1 U6052 ( .A1(n4711), .A2(n4712), .A3(n4710), .ZN(n7145) );
  NAND2_X1 U6053 ( .A1(n4713), .A2(n6842), .ZN(n4711) );
  NAND2_X1 U6054 ( .A1(n5079), .A2(n4714), .ZN(n4712) );
  NAND2_X1 U6055 ( .A1(n5214), .A2(n4732), .ZN(n4728) );
  NAND2_X1 U6056 ( .A1(n4728), .A2(n4729), .ZN(n5265) );
  NAND2_X1 U6057 ( .A1(n4893), .A2(n4744), .ZN(n4743) );
  NAND2_X1 U6058 ( .A1(n4758), .A2(n4757), .ZN(n5392) );
  NAND3_X1 U6059 ( .A1(n5091), .A2(n5095), .A3(n5092), .ZN(n4762) );
  NAND3_X1 U6060 ( .A1(n5939), .A2(n4772), .A3(n5938), .ZN(n4771) );
  NAND2_X1 U6061 ( .A1(n7620), .A2(n5798), .ZN(n5810) );
  NAND2_X1 U6062 ( .A1(n8280), .A2(n8281), .ZN(n5811) );
  INV_X1 U6063 ( .A(n5809), .ZN(n4780) );
  NAND2_X1 U6064 ( .A1(n4786), .A2(n6050), .ZN(P2_U3222) );
  OAI211_X1 U6065 ( .C1(n6023), .C2(n6017), .A(n4787), .B(n6033), .ZN(n4786)
         );
  NAND2_X1 U6066 ( .A1(n6023), .A2(n6022), .ZN(n4787) );
  OAI21_X1 U6067 ( .B1(n5469), .B2(n7054), .A(n9189), .ZN(n8954) );
  AOI21_X1 U6068 ( .B1(n9189), .B2(n7054), .A(n4792), .ZN(n4791) );
  NAND2_X1 U6069 ( .A1(n5469), .A2(n9189), .ZN(n4793) );
  NAND2_X1 U6070 ( .A1(n4794), .A2(n9193), .ZN(n6932) );
  NAND2_X1 U6071 ( .A1(n9446), .A2(n4285), .ZN(n4797) );
  NAND2_X1 U6072 ( .A1(n4992), .A2(n4991), .ZN(n4994) );
  NAND2_X1 U6073 ( .A1(n4992), .A2(n4799), .ZN(n9632) );
  XNOR2_X2 U6074 ( .A(n6556), .B(n6557), .ZN(n9093) );
  AND3_X2 U6075 ( .A1(n4808), .A2(n4807), .A3(n4806), .ZN(n6557) );
  NAND2_X1 U6076 ( .A1(n7105), .A2(n4813), .ZN(n4812) );
  NAND2_X1 U6077 ( .A1(n4812), .A2(n4815), .ZN(n5475) );
  OAI21_X1 U6078 ( .B1(n7594), .B2(n4821), .A(n4818), .ZN(n9496) );
  INV_X1 U6079 ( .A(n9088), .ZN(n4829) );
  NAND2_X1 U6080 ( .A1(n5089), .A2(n4833), .ZN(n4832) );
  NAND3_X1 U6081 ( .A1(n4968), .A2(n4831), .A3(n5089), .ZN(n4990) );
  AND2_X2 U6082 ( .A1(n4963), .A2(n4964), .ZN(n4833) );
  NOR2_X2 U6083 ( .A1(n4832), .A2(n4969), .ZN(n5512) );
  NAND2_X1 U6084 ( .A1(n7786), .A2(n7785), .ZN(n7792) );
  MUX2_X1 U6085 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n6156), .S(n9935), .Z(
        P1_U3552) );
  INV_X1 U6086 ( .A(n6849), .ZN(n9258) );
  NAND2_X2 U6087 ( .A1(n9189), .A2(n9191), .ZN(n7054) );
  XNOR2_X1 U6088 ( .A(n5388), .B(n5389), .ZN(n7568) );
  NAND2_X1 U6089 ( .A1(n4263), .A2(n7794), .ZN(n5062) );
  XNOR2_X1 U6090 ( .A(n8425), .B(n8424), .ZN(n8696) );
  OR2_X1 U6091 ( .A1(n6152), .A2(n6151), .ZN(P2_U3216) );
  NAND2_X1 U6092 ( .A1(n7828), .A2(n7068), .ZN(n7829) );
  NAND2_X1 U6093 ( .A1(n8324), .A2(n6052), .ZN(n6093) );
  NOR2_X1 U6094 ( .A1(n6051), .A2(n4266), .ZN(n5585) );
  OR2_X1 U6095 ( .A1(n5989), .A2(n5634), .ZN(n5642) );
  OR2_X1 U6096 ( .A1(n5989), .A2(n5608), .ZN(n5609) );
  NAND2_X1 U6097 ( .A1(n7068), .A2(n7806), .ZN(n6097) );
  NAND2_X1 U6098 ( .A1(n5310), .A2(n5309), .ZN(n9438) );
  NAND2_X1 U6099 ( .A1(n5477), .A2(n8953), .ZN(n9469) );
  INV_X1 U6100 ( .A(n9496), .ZN(n5477) );
  NOR2_X2 U6101 ( .A1(n8834), .A2(n8833), .ZN(n8933) );
  INV_X1 U6102 ( .A(n7048), .ZN(n5474) );
  INV_X1 U6103 ( .A(n7980), .ZN(n5579) );
  AND2_X2 U6105 ( .A1(n5558), .A2(n5557), .ZN(n5649) );
  NAND2_X1 U6106 ( .A1(n5557), .A2(n8767), .ZN(n5648) );
  INV_X1 U6107 ( .A(n5557), .ZN(n8764) );
  INV_X1 U6108 ( .A(n5097), .ZN(n5122) );
  INV_X1 U6109 ( .A(n4997), .ZN(n9637) );
  CLKBUF_X1 U6110 ( .A(n5489), .Z(n6649) );
  OAI21_X1 U6111 ( .B1(n7546), .B2(n5228), .A(n5227), .ZN(n7592) );
  AND2_X1 U6112 ( .A1(n6420), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n4834) );
  OR2_X1 U6113 ( .A1(n5547), .A2(n5546), .ZN(n4835) );
  AND4_X1 U6114 ( .A1(n5689), .A2(n5538), .A3(n6389), .A4(n5537), .ZN(n4836)
         );
  OR2_X1 U6115 ( .A1(n5592), .A2(n6197), .ZN(n4837) );
  AND4_X1 U6116 ( .A1(n4975), .A2(n4974), .A3(n4970), .A4(n4973), .ZN(n4838)
         );
  OR2_X1 U6117 ( .A1(n8224), .A2(n8228), .ZN(n4839) );
  OR2_X1 U6118 ( .A1(n8902), .A2(n8813), .ZN(n4840) );
  OR2_X1 U6119 ( .A1(n9929), .A2(n6157), .ZN(n4841) );
  AND2_X1 U6120 ( .A1(n5948), .A2(n5947), .ZN(n8158) );
  INV_X1 U6121 ( .A(n8158), .ZN(n8299) );
  AND2_X1 U6122 ( .A1(n5893), .A2(n5881), .ZN(n4843) );
  INV_X1 U6123 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5461) );
  NOR2_X1 U6124 ( .A1(n6951), .A2(n5664), .ZN(n4844) );
  AND2_X1 U6125 ( .A1(n6136), .A2(n6135), .ZN(n4846) );
  NOR2_X1 U6126 ( .A1(n8877), .A2(n7681), .ZN(n4848) );
  INV_X1 U6127 ( .A(n7829), .ZN(n7830) );
  INV_X1 U6128 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5537) );
  INV_X1 U6129 ( .A(n5759), .ZN(n5758) );
  INV_X1 U6130 ( .A(n7259), .ZN(n6658) );
  OAI22_X1 U6131 ( .A1(n6658), .A2(n6673), .B1(n6898), .B2(n7263), .ZN(n6659)
         );
  INV_X1 U6132 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5216) );
  INV_X1 U6133 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n4960) );
  INV_X1 U6134 ( .A(n5820), .ZN(n5817) );
  OR2_X1 U6135 ( .A1(n5772), .A2(n7328), .ZN(n5787) );
  INV_X1 U6136 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5689) );
  INV_X1 U6137 ( .A(n6566), .ZN(n6563) );
  XNOR2_X1 U6138 ( .A(n8063), .B(n6659), .ZN(n6662) );
  INV_X1 U6139 ( .A(n5380), .ZN(n5378) );
  INV_X1 U6140 ( .A(n5357), .ZN(n4987) );
  INV_X1 U6141 ( .A(n5109), .ZN(n4980) );
  INV_X1 U6142 ( .A(n6844), .ZN(n6848) );
  INV_X1 U6143 ( .A(n6894), .ZN(n5014) );
  INV_X1 U6144 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5453) );
  INV_X1 U6145 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5280) );
  AND2_X1 U6146 ( .A1(n5138), .A2(n5142), .ZN(n4876) );
  INV_X1 U6147 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5104) );
  INV_X1 U6148 ( .A(n6090), .ZN(n5580) );
  OR2_X1 U6149 ( .A1(n5936), .A2(n8300), .ZN(n5933) );
  INV_X1 U6150 ( .A(n7127), .ZN(n5723) );
  AND2_X1 U6151 ( .A1(n8191), .A2(n5901), .ZN(n5902) );
  INV_X1 U6152 ( .A(n5918), .ZN(n5929) );
  INV_X1 U6153 ( .A(n8130), .ZN(n6132) );
  INV_X1 U6154 ( .A(n7964), .ZN(n6069) );
  INV_X1 U6155 ( .A(n5730), .ZN(n5729) );
  NAND2_X1 U6156 ( .A1(n7832), .A2(n7831), .ZN(n7809) );
  OR2_X1 U6157 ( .A1(n6861), .A2(n9984), .ZN(n7075) );
  INV_X1 U6158 ( .A(n8843), .ZN(n8012) );
  AND2_X1 U6159 ( .A1(n9232), .A2(n9878), .ZN(n6415) );
  OR2_X1 U6160 ( .A1(n5399), .A2(n8940), .ZN(n5430) );
  NAND2_X1 U6161 ( .A1(n5378), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5399) );
  OR2_X1 U6162 ( .A1(n5315), .A2(n8872), .ZN(n5328) );
  NAND2_X1 U6163 ( .A1(n5286), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5315) );
  AOI21_X1 U6164 ( .B1(n7259), .B2(n6900), .A(n4834), .ZN(n6421) );
  NOR2_X1 U6165 ( .A1(n9788), .A2(n9789), .ZN(n9787) );
  OR2_X1 U6166 ( .A1(n5238), .A2(n5237), .ZN(n5256) );
  OR2_X1 U6167 ( .A1(n5162), .A2(n6625), .ZN(n5177) );
  NAND2_X1 U6168 ( .A1(n4980), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5130) );
  NAND2_X1 U6169 ( .A1(n5408), .A2(n5407), .ZN(n5410) );
  NAND2_X1 U6170 ( .A1(n4900), .A2(n4899), .ZN(n4903) );
  AND2_X1 U6171 ( .A1(n5067), .A2(n4861), .ZN(n5091) );
  AND2_X1 U6172 ( .A1(n5977), .A2(n5976), .ZN(n6140) );
  OR2_X1 U6173 ( .A1(n5744), .A2(n5743), .ZN(n5759) );
  OR2_X1 U6174 ( .A1(n6832), .A2(n6086), .ZN(n6045) );
  NAND2_X1 U6175 ( .A1(n7179), .A2(n7959), .ZN(n7180) );
  OR2_X1 U6176 ( .A1(n6428), .A2(n6454), .ZN(n8249) );
  OR2_X1 U6177 ( .A1(n8747), .A2(n8308), .ZN(n6077) );
  OR2_X1 U6178 ( .A1(n5328), .A2(n5327), .ZN(n5341) );
  NAND2_X1 U6179 ( .A1(n8013), .A2(n8012), .ZN(n8841) );
  INV_X1 U6180 ( .A(n9252), .ZN(n7512) );
  NOR2_X1 U6181 ( .A1(n8083), .A2(n8082), .ZN(n8932) );
  AND2_X1 U6182 ( .A1(n5430), .A2(n5400), .ZN(n9349) );
  OR2_X1 U6183 ( .A1(n5074), .A2(n6180), .ZN(n5077) );
  OR2_X1 U6184 ( .A1(n6624), .A2(n6623), .ZN(n6680) );
  OR2_X1 U6185 ( .A1(n6187), .A2(n7704), .ZN(n9288) );
  NAND2_X1 U6186 ( .A1(n9168), .A2(n9223), .ZN(n9114) );
  INV_X1 U6187 ( .A(n9245), .ZN(n9337) );
  AND2_X1 U6188 ( .A1(n9149), .A2(n9031), .ZN(n9424) );
  AND2_X1 U6189 ( .A1(n9140), .A2(n9138), .ZN(n9105) );
  AND2_X1 U6190 ( .A1(n8992), .A2(n9000), .ZN(n9087) );
  INV_X1 U6191 ( .A(n9911), .ZN(n9606) );
  OR2_X1 U6192 ( .A1(n9068), .A2(n9183), .ZN(n9609) );
  NAND2_X1 U6193 ( .A1(n5410), .A2(n5409), .ZN(n5423) );
  INV_X1 U6194 ( .A(n8275), .ZN(n8287) );
  AND2_X1 U6195 ( .A1(n6725), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8275) );
  INV_X1 U6196 ( .A(n8278), .ZN(n8290) );
  AND4_X1 U6197 ( .A1(n5885), .A2(n5884), .A3(n5883), .A4(n5882), .ZN(n8197)
         );
  AND4_X1 U6198 ( .A1(n5808), .A2(n5807), .A3(n5806), .A4(n5805), .ZN(n7768)
         );
  INV_X1 U6199 ( .A(n9937), .ZN(n9662) );
  AND2_X1 U6200 ( .A1(n9938), .A2(n6454), .ZN(n9937) );
  INV_X1 U6201 ( .A(n8588), .ZN(n9993) );
  AND2_X1 U6202 ( .A1(n10120), .A2(n10069), .ZN(n8670) );
  AND2_X1 U6203 ( .A1(n10101), .A2(n10069), .ZN(n8748) );
  AND2_X1 U6204 ( .A1(n6429), .A2(n6029), .ZN(n10013) );
  AND2_X1 U6205 ( .A1(n8090), .A2(n8089), .ZN(n8151) );
  OR2_X1 U6206 ( .A1(n6943), .A2(n6415), .ZN(n9911) );
  OR2_X1 U6207 ( .A1(n8102), .A2(n5049), .ZN(n5439) );
  OR3_X1 U6208 ( .A1(n9609), .A2(n9186), .A3(n9629), .ZN(n9876) );
  INV_X1 U6209 ( .A(n9682), .ZN(n9497) );
  OR2_X1 U6210 ( .A1(n6943), .A2(n9183), .ZN(n9921) );
  INV_X1 U6211 ( .A(n9926), .ZN(n9597) );
  INV_X1 U6212 ( .A(n5488), .ZN(n6414) );
  AND2_X1 U6213 ( .A1(n5127), .A2(n5126), .ZN(n9772) );
  XNOR2_X1 U6214 ( .A(n4862), .B(SI_4_), .ZN(n5067) );
  INV_X1 U6215 ( .A(n9650), .ZN(n9943) );
  OR3_X1 U6216 ( .A1(n6043), .A2(n6257), .A3(n10069), .ZN(n8259) );
  NAND2_X1 U6217 ( .A1(n5992), .A2(n5991), .ZN(n8296) );
  INV_X1 U6218 ( .A(n9668), .ZN(n9939) );
  INV_X1 U6219 ( .A(n9990), .ZN(n10004) );
  INV_X1 U6220 ( .A(n10006), .ZN(n8592) );
  INV_X1 U6221 ( .A(n8639), .ZN(n8672) );
  INV_X1 U6222 ( .A(n8716), .ZN(n8750) );
  INV_X1 U6223 ( .A(n10101), .ZN(n10099) );
  INV_X1 U6224 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6237) );
  AND2_X1 U6225 ( .A1(n6703), .A2(n6702), .ZN(n8926) );
  OR2_X1 U6226 ( .A1(n7252), .A2(n9911), .ZN(n8945) );
  AND2_X1 U6227 ( .A1(n5451), .A2(n5450), .ZN(n9321) );
  INV_X1 U6228 ( .A(n9773), .ZN(n9870) );
  INV_X1 U6229 ( .A(n9693), .ZN(n9519) );
  OR2_X1 U6230 ( .A1(n6155), .A2(n6409), .ZN(n9933) );
  OR3_X1 U6231 ( .A1(n9604), .A2(n9603), .A3(n9602), .ZN(n9627) );
  OR2_X1 U6232 ( .A1(n6155), .A2(n6907), .ZN(n9927) );
  INV_X1 U6233 ( .A(n9891), .ZN(n9892) );
  INV_X1 U6234 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6205) );
  NAND2_X1 U6235 ( .A1(n5005), .A2(n5004), .ZN(n4852) );
  INV_X1 U6236 ( .A(n4849), .ZN(n4850) );
  NAND2_X1 U6237 ( .A1(n4850), .A2(SI_1_), .ZN(n4851) );
  NAND2_X1 U6238 ( .A1(n4852), .A2(n4851), .ZN(n5018) );
  INV_X1 U6239 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6218) );
  INV_X1 U6240 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6199) );
  MUX2_X1 U6241 ( .A(n6218), .B(n6199), .S(n7794), .Z(n4853) );
  XNOR2_X1 U6242 ( .A(n4853), .B(SI_2_), .ZN(n5017) );
  NAND2_X1 U6243 ( .A1(n5018), .A2(n5017), .ZN(n4856) );
  INV_X1 U6244 ( .A(n4853), .ZN(n4854) );
  NAND2_X1 U6245 ( .A1(n4854), .A2(SI_2_), .ZN(n4855) );
  INV_X1 U6246 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6198) );
  INV_X1 U6247 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6216) );
  MUX2_X1 U6248 ( .A(n6198), .B(n6216), .S(n5577), .Z(n4857) );
  XNOR2_X1 U6249 ( .A(n4857), .B(SI_3_), .ZN(n5031) );
  INV_X1 U6250 ( .A(n4857), .ZN(n4858) );
  NAND2_X1 U6251 ( .A1(n4858), .A2(SI_3_), .ZN(n4859) );
  INV_X1 U6252 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6200) );
  INV_X1 U6253 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6221) );
  MUX2_X1 U6254 ( .A(n6200), .B(n6221), .S(n5577), .Z(n4862) );
  NAND2_X1 U6255 ( .A1(n4860), .A2(SI_5_), .ZN(n4864) );
  INV_X1 U6256 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6201) );
  INV_X1 U6257 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6214) );
  MUX2_X1 U6258 ( .A(n6201), .B(n6214), .S(n5577), .Z(n4865) );
  INV_X1 U6259 ( .A(n4862), .ZN(n4863) );
  NAND2_X1 U6260 ( .A1(n4863), .A2(SI_4_), .ZN(n5058) );
  INV_X1 U6261 ( .A(n4865), .ZN(n4866) );
  NAND2_X1 U6262 ( .A1(n4866), .A2(SI_6_), .ZN(n5101) );
  MUX2_X1 U6263 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n7794), .Z(n4878) );
  NAND2_X1 U6264 ( .A1(n4878), .A2(SI_7_), .ZN(n4877) );
  AND2_X1 U6265 ( .A1(n5101), .A2(n4877), .ZN(n5117) );
  MUX2_X1 U6266 ( .A(n6231), .B(n6229), .S(n6203), .Z(n4868) );
  INV_X1 U6267 ( .A(SI_8_), .ZN(n4867) );
  INV_X1 U6268 ( .A(n4868), .ZN(n4869) );
  NAND2_X1 U6269 ( .A1(n4869), .A2(SI_8_), .ZN(n4870) );
  INV_X1 U6270 ( .A(n5120), .ZN(n4871) );
  MUX2_X1 U6271 ( .A(n6226), .B(n6205), .S(n6203), .Z(n4873) );
  INV_X1 U6272 ( .A(SI_9_), .ZN(n4872) );
  INV_X1 U6273 ( .A(n4873), .ZN(n4874) );
  NAND2_X1 U6274 ( .A1(n4874), .A2(SI_9_), .ZN(n4875) );
  INV_X1 U6275 ( .A(n5142), .ZN(n4883) );
  INV_X1 U6276 ( .A(n4877), .ZN(n4880) );
  INV_X1 U6277 ( .A(n5102), .ZN(n4879) );
  NAND3_X1 U6278 ( .A1(n4886), .A2(n4885), .A3(n4884), .ZN(n5156) );
  INV_X1 U6279 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n4887) );
  MUX2_X1 U6280 ( .A(n6237), .B(n4887), .S(n5577), .Z(n4889) );
  INV_X1 U6281 ( .A(SI_10_), .ZN(n4888) );
  NAND2_X1 U6282 ( .A1(n4889), .A2(n4888), .ZN(n4892) );
  INV_X1 U6283 ( .A(n4889), .ZN(n4890) );
  NAND2_X1 U6284 ( .A1(n4890), .A2(SI_10_), .ZN(n4891) );
  INV_X1 U6285 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6241) );
  INV_X1 U6286 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6239) );
  MUX2_X1 U6287 ( .A(n6241), .B(n6239), .S(n6203), .Z(n4894) );
  INV_X1 U6288 ( .A(n4894), .ZN(n4895) );
  INV_X1 U6289 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6253) );
  INV_X1 U6290 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n4898) );
  MUX2_X1 U6291 ( .A(n6253), .B(n4898), .S(n5577), .Z(n4900) );
  INV_X1 U6292 ( .A(SI_12_), .ZN(n4899) );
  INV_X1 U6293 ( .A(n4900), .ZN(n4901) );
  NAND2_X1 U6294 ( .A1(n4901), .A2(SI_12_), .ZN(n4902) );
  INV_X1 U6295 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6256) );
  INV_X1 U6296 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n4904) );
  MUX2_X1 U6297 ( .A(n6256), .B(n4904), .S(n5577), .Z(n4906) );
  INV_X1 U6298 ( .A(SI_13_), .ZN(n4905) );
  NAND2_X1 U6299 ( .A1(n4906), .A2(n4905), .ZN(n4909) );
  INV_X1 U6300 ( .A(n4906), .ZN(n4907) );
  NAND2_X1 U6301 ( .A1(n4907), .A2(SI_13_), .ZN(n4908) );
  INV_X1 U6302 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6274) );
  INV_X1 U6303 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6265) );
  MUX2_X1 U6304 ( .A(n6274), .B(n6265), .S(n5577), .Z(n4910) );
  XNOR2_X1 U6305 ( .A(n4910), .B(SI_14_), .ZN(n5213) );
  INV_X1 U6306 ( .A(n4910), .ZN(n4911) );
  NAND2_X1 U6307 ( .A1(n4911), .A2(SI_14_), .ZN(n4912) );
  INV_X1 U6308 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6408) );
  INV_X1 U6309 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6406) );
  MUX2_X1 U6310 ( .A(n6408), .B(n6406), .S(n6203), .Z(n4914) );
  INV_X1 U6311 ( .A(SI_15_), .ZN(n4913) );
  NAND2_X1 U6312 ( .A1(n4914), .A2(n4913), .ZN(n4917) );
  INV_X1 U6313 ( .A(n4914), .ZN(n4915) );
  NAND2_X1 U6314 ( .A1(n4915), .A2(SI_15_), .ZN(n4916) );
  NAND2_X1 U6315 ( .A1(n4917), .A2(n4916), .ZN(n5229) );
  INV_X1 U6316 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n4919) );
  INV_X1 U6317 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n4918) );
  MUX2_X1 U6318 ( .A(n4919), .B(n4918), .S(n5577), .Z(n4921) );
  INV_X1 U6319 ( .A(SI_16_), .ZN(n4920) );
  NAND2_X1 U6320 ( .A1(n4921), .A2(n4920), .ZN(n4924) );
  INV_X1 U6321 ( .A(n4921), .ZN(n4922) );
  NAND2_X1 U6322 ( .A1(n4922), .A2(SI_16_), .ZN(n4923) );
  INV_X1 U6323 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6695) );
  INV_X1 U6324 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n4925) );
  MUX2_X1 U6325 ( .A(n6695), .B(n4925), .S(n6203), .Z(n4926) );
  XNOR2_X1 U6326 ( .A(n4926), .B(SI_17_), .ZN(n5264) );
  INV_X1 U6327 ( .A(n5264), .ZN(n4929) );
  INV_X1 U6328 ( .A(n4926), .ZN(n4927) );
  NAND2_X1 U6329 ( .A1(n4927), .A2(SI_17_), .ZN(n4928) );
  MUX2_X1 U6330 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5577), .Z(n4931) );
  XNOR2_X1 U6331 ( .A(n4931), .B(SI_18_), .ZN(n5278) );
  INV_X1 U6332 ( .A(n5278), .ZN(n4930) );
  NAND2_X1 U6333 ( .A1(n4931), .A2(SI_18_), .ZN(n4932) );
  INV_X1 U6334 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n8137) );
  INV_X1 U6335 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6891) );
  MUX2_X1 U6336 ( .A(n8137), .B(n6891), .S(n5577), .Z(n4935) );
  INV_X1 U6337 ( .A(SI_19_), .ZN(n4934) );
  NAND2_X1 U6338 ( .A1(n4935), .A2(n4934), .ZN(n4938) );
  INV_X1 U6339 ( .A(n4935), .ZN(n4936) );
  NAND2_X1 U6340 ( .A1(n4936), .A2(SI_19_), .ZN(n4937) );
  NAND2_X1 U6341 ( .A1(n4938), .A2(n4937), .ZN(n5292) );
  INV_X1 U6342 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6980) );
  INV_X1 U6343 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6966) );
  MUX2_X1 U6344 ( .A(n6980), .B(n6966), .S(n6203), .Z(n4940) );
  INV_X1 U6345 ( .A(SI_20_), .ZN(n4939) );
  NAND2_X1 U6346 ( .A1(n4940), .A2(n4939), .ZN(n4943) );
  INV_X1 U6347 ( .A(n4940), .ZN(n4941) );
  NAND2_X1 U6348 ( .A1(n4941), .A2(SI_20_), .ZN(n4942) );
  AND2_X1 U6349 ( .A1(n4943), .A2(n4942), .ZN(n5311) );
  INV_X1 U6350 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7019) );
  INV_X1 U6351 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7066) );
  MUX2_X1 U6352 ( .A(n7019), .B(n7066), .S(n6203), .Z(n4945) );
  XNOR2_X1 U6353 ( .A(n4945), .B(SI_21_), .ZN(n5323) );
  INV_X1 U6354 ( .A(n5323), .ZN(n4948) );
  INV_X1 U6355 ( .A(n4945), .ZN(n4946) );
  NAND2_X1 U6356 ( .A1(n4946), .A2(SI_21_), .ZN(n4947) );
  INV_X1 U6357 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8135) );
  INV_X1 U6358 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7778) );
  MUX2_X1 U6359 ( .A(n8135), .B(n7778), .S(n6203), .Z(n4949) );
  INV_X1 U6360 ( .A(SI_22_), .ZN(n6324) );
  NAND2_X1 U6361 ( .A1(n4949), .A2(n6324), .ZN(n4952) );
  INV_X1 U6362 ( .A(n4949), .ZN(n4950) );
  NAND2_X1 U6363 ( .A1(n4950), .A2(SI_22_), .ZN(n4951) );
  NAND2_X1 U6364 ( .A1(n4952), .A2(n4951), .ZN(n5337) );
  INV_X1 U6365 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7278) );
  INV_X1 U6366 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7282) );
  MUX2_X1 U6367 ( .A(n7278), .B(n7282), .S(n5577), .Z(n4954) );
  INV_X1 U6368 ( .A(SI_23_), .ZN(n4953) );
  NAND2_X1 U6369 ( .A1(n4954), .A2(n4953), .ZN(n4958) );
  INV_X1 U6370 ( .A(n4954), .ZN(n4955) );
  NAND2_X1 U6371 ( .A1(n4955), .A2(SI_23_), .ZN(n4956) );
  NAND2_X1 U6372 ( .A1(n4958), .A2(n4956), .ZN(n5350) );
  INV_X1 U6373 ( .A(n5350), .ZN(n4957) );
  INV_X1 U6374 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7401) );
  INV_X1 U6375 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7386) );
  MUX2_X1 U6376 ( .A(n7401), .B(n7386), .S(n6203), .Z(n5367) );
  XNOR2_X1 U6377 ( .A(n5367), .B(SI_24_), .ZN(n5366) );
  XNOR2_X1 U6378 ( .A(n5371), .B(n5366), .ZN(n7385) );
  NOR2_X1 U6379 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n4962) );
  NOR2_X1 U6380 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4961) );
  NOR2_X1 U6381 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n4965) );
  NAND4_X1 U6382 ( .A1(n5249), .A2(n4965), .A3(n5453), .A4(n5280), .ZN(n4967)
         );
  INV_X1 U6383 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5266) );
  NAND4_X1 U6384 ( .A1(n5266), .A2(n5216), .A3(n5294), .A4(n5461), .ZN(n4966)
         );
  INV_X1 U6385 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4970) );
  INV_X1 U6386 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4974) );
  NAND2_X1 U6387 ( .A1(n5505), .A2(n4974), .ZN(n5508) );
  INV_X1 U6388 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n6392) );
  INV_X1 U6389 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5502) );
  NAND2_X1 U6390 ( .A1(n6392), .A2(n5502), .ZN(n4972) );
  INV_X1 U6391 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4973) );
  INV_X1 U6392 ( .A(n4972), .ZN(n4975) );
  NAND2_X1 U6393 ( .A1(n4990), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4976) );
  INV_X1 U6394 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4991) );
  NAND2_X2 U6395 ( .A1(n4263), .A2(n6203), .ZN(n5097) );
  NAND2_X1 U6396 ( .A1(n7385), .A2(n8114), .ZN(n4978) );
  OR2_X1 U6397 ( .A1(n8115), .A2(n7386), .ZN(n4977) );
  NAND3_X1 U6398 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5082) );
  INV_X1 U6399 ( .A(n5082), .ZN(n4979) );
  INV_X1 U6400 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5147) );
  INV_X1 U6401 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6625) );
  INV_X1 U6402 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5205) );
  INV_X1 U6403 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5237) );
  INV_X1 U6404 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5269) );
  INV_X1 U6405 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5287) );
  INV_X1 U6406 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8872) );
  INV_X1 U6407 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5327) );
  INV_X1 U6408 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n4988) );
  NAND2_X1 U6409 ( .A1(n5359), .A2(n4988), .ZN(n4989) );
  AND2_X1 U6410 ( .A1(n5380), .A2(n4989), .ZN(n9384) );
  INV_X1 U6411 ( .A(n4990), .ZN(n4992) );
  XNOR2_X2 U6412 ( .A(n4993), .B(P1_IR_REG_30__SCAN_IN), .ZN(n4997) );
  NAND2_X1 U6413 ( .A1(n4994), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4995) );
  XNOR2_X2 U6414 ( .A(n4995), .B(P1_IR_REG_29__SCAN_IN), .ZN(n4996) );
  NAND2_X1 U6415 ( .A1(n9384), .A2(n5416), .ZN(n5003) );
  INV_X1 U6416 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n5000) );
  AND2_X2 U6417 ( .A1(n9637), .A2(n9643), .ZN(n5051) );
  NAND2_X1 U6418 ( .A1(n5492), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n4999) );
  NAND2_X1 U6419 ( .A1(n5491), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n4998) );
  OAI211_X1 U6420 ( .C1(n5074), .C2(n5000), .A(n4999), .B(n4998), .ZN(n5001)
         );
  INV_X1 U6421 ( .A(n5001), .ZN(n5002) );
  INV_X1 U6422 ( .A(n9394), .ZN(n5481) );
  INV_X1 U6423 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6224) );
  XNOR2_X1 U6424 ( .A(n5005), .B(n5004), .ZN(n6222) );
  INV_X1 U6425 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5006) );
  OR2_X1 U6426 ( .A1(n5088), .A2(n6223), .ZN(n5007) );
  INV_X1 U6427 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6903) );
  INV_X1 U6428 ( .A(n9093), .ZN(n5015) );
  INV_X1 U6429 ( .A(SI_0_), .ZN(n6383) );
  NOR2_X1 U6430 ( .A1(n7794), .A2(n6383), .ZN(n5009) );
  INV_X1 U6431 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5008) );
  XNOR2_X1 U6432 ( .A(n5009), .B(n5008), .ZN(n9647) );
  MUX2_X1 U6433 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9647), .S(n5088), .Z(n6900) );
  NAND2_X1 U6434 ( .A1(n5416), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5013) );
  NAND2_X1 U6435 ( .A1(n5051), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5012) );
  NAND2_X1 U6436 ( .A1(n6245), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5011) );
  NAND2_X1 U6437 ( .A1(n5050), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5010) );
  NAND2_X1 U6438 ( .A1(n6900), .A2(n6568), .ZN(n6894) );
  INV_X1 U6439 ( .A(n6556), .ZN(n6901) );
  INV_X1 U6440 ( .A(n6557), .ZN(n9262) );
  NAND2_X1 U6441 ( .A1(n6901), .A2(n9262), .ZN(n5016) );
  XNOR2_X1 U6442 ( .A(n5018), .B(n5017), .ZN(n6217) );
  OR2_X1 U6443 ( .A1(n5097), .A2(n6217), .ZN(n5024) );
  OR2_X1 U6444 ( .A1(n5062), .A2(n6218), .ZN(n5023) );
  INV_X1 U6445 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5020) );
  NAND2_X1 U6446 ( .A1(n5021), .A2(n5020), .ZN(n5033) );
  OR2_X1 U6447 ( .A1(n5088), .A2(n6636), .ZN(n5022) );
  NAND2_X1 U6448 ( .A1(n5492), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5029) );
  INV_X1 U6449 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6176) );
  OR2_X1 U6450 ( .A1(n5074), .A2(n6176), .ZN(n5028) );
  INV_X1 U6451 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5025) );
  INV_X1 U6452 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7062) );
  AND4_X2 U6453 ( .A1(n5029), .A2(n5028), .A3(n5027), .A4(n5026), .ZN(n6898)
         );
  NAND2_X2 U6454 ( .A1(n7059), .A2(n6898), .ZN(n9189) );
  NAND2_X1 U6455 ( .A1(n9260), .A2(n6673), .ZN(n9191) );
  NAND2_X1 U6456 ( .A1(n7055), .A2(n7054), .ZN(n7053) );
  NAND2_X1 U6457 ( .A1(n6673), .A2(n6898), .ZN(n5030) );
  NAND2_X1 U6458 ( .A1(n7053), .A2(n5030), .ZN(n6818) );
  OR2_X1 U6459 ( .A1(n8115), .A2(n6216), .ZN(n5039) );
  XNOR2_X1 U6460 ( .A(n5032), .B(n5031), .ZN(n6215) );
  OR2_X1 U6461 ( .A1(n5097), .A2(n6215), .ZN(n5037) );
  NAND2_X1 U6462 ( .A1(n5033), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5035) );
  INV_X1 U6463 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5034) );
  OR2_X1 U6464 ( .A1(n5088), .A2(n6604), .ZN(n5036) );
  NAND2_X1 U6465 ( .A1(n5051), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5045) );
  INV_X1 U6466 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6179) );
  OR2_X1 U6467 ( .A1(n5074), .A2(n6179), .ZN(n5044) );
  INV_X1 U6468 ( .A(n6245), .ZN(n5041) );
  INV_X1 U6469 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n5040) );
  OR2_X1 U6470 ( .A1(n5041), .A2(n5040), .ZN(n5043) );
  OR2_X1 U6471 ( .A1(n5049), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5042) );
  NAND2_X1 U6472 ( .A1(n9193), .A2(n9192), .ZN(n9089) );
  NAND2_X1 U6473 ( .A1(n7087), .A2(n6933), .ZN(n6841) );
  INV_X1 U6474 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5047) );
  NAND2_X1 U6475 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5046) );
  NAND2_X1 U6476 ( .A1(n5047), .A2(n5046), .ZN(n5048) );
  NAND2_X1 U6477 ( .A1(n5082), .A2(n5048), .ZN(n9875) );
  OR2_X1 U6478 ( .A1(n5049), .A2(n9875), .ZN(n5054) );
  NAND2_X1 U6479 ( .A1(n5050), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5053) );
  NAND2_X1 U6480 ( .A1(n5051), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5052) );
  NAND3_X1 U6481 ( .A1(n5054), .A2(n5053), .A3(n5052), .ZN(n5057) );
  INV_X1 U6482 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5055) );
  NAND2_X1 U6483 ( .A1(n5059), .A2(n5058), .ZN(n5061) );
  INV_X1 U6484 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6233) );
  OR2_X1 U6485 ( .A1(n5062), .A2(n6233), .ZN(n5066) );
  NAND2_X1 U6486 ( .A1(n5063), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5064) );
  XNOR2_X1 U6487 ( .A(n5064), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9760) );
  INV_X1 U6488 ( .A(n9760), .ZN(n6232) );
  OR2_X1 U6489 ( .A1(n5088), .A2(n6232), .ZN(n5065) );
  NAND2_X1 U6490 ( .A1(n9257), .A2(n9874), .ZN(n8955) );
  NAND2_X1 U6491 ( .A1(n7038), .A2(n7156), .ZN(n7153) );
  NAND2_X1 U6492 ( .A1(n8955), .A2(n7153), .ZN(n6844) );
  OR2_X1 U6493 ( .A1(n5097), .A2(n6220), .ZN(n5073) );
  OR2_X1 U6494 ( .A1(n8115), .A2(n6221), .ZN(n5072) );
  NAND2_X1 U6495 ( .A1(n5068), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5069) );
  MUX2_X1 U6496 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5069), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5070) );
  NAND2_X1 U6497 ( .A1(n5070), .A2(n5063), .ZN(n6219) );
  OR2_X1 U6498 ( .A1(n5088), .A2(n6219), .ZN(n5071) );
  NAND2_X1 U6499 ( .A1(n5492), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5078) );
  INV_X1 U6500 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6180) );
  XNOR2_X1 U6501 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6938) );
  OR2_X1 U6502 ( .A1(n5049), .A2(n6938), .ZN(n5076) );
  INV_X1 U6503 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6939) );
  OR2_X1 U6504 ( .A1(n5332), .A2(n6939), .ZN(n5075) );
  NAND2_X1 U6505 ( .A1(n9912), .A2(n6849), .ZN(n6843) );
  NAND2_X1 U6506 ( .A1(n7038), .A2(n9257), .ZN(n5080) );
  NAND2_X1 U6507 ( .A1(n5492), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5087) );
  INV_X1 U6508 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n5081) );
  OR2_X1 U6509 ( .A1(n5074), .A2(n5081), .ZN(n5086) );
  INV_X1 U6510 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6593) );
  NAND2_X1 U6511 ( .A1(n5082), .A2(n6593), .ZN(n5083) );
  NAND2_X1 U6512 ( .A1(n5109), .A2(n5083), .ZN(n7257) );
  OR2_X1 U6513 ( .A1(n5049), .A2(n7257), .ZN(n5085) );
  INV_X1 U6514 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6165) );
  OR2_X1 U6515 ( .A1(n5332), .A2(n6165), .ZN(n5084) );
  OR2_X1 U6516 ( .A1(n5089), .A2(n9631), .ZN(n5090) );
  XNOR2_X1 U6517 ( .A(n5090), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6601) );
  AOI22_X1 U6518 ( .A1(n5298), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6161), .B2(
        n6601), .ZN(n5099) );
  NAND2_X1 U6519 ( .A1(n5092), .A2(n5091), .ZN(n5094) );
  NAND2_X1 U6520 ( .A1(n5094), .A2(n5093), .ZN(n5096) );
  XNOR2_X1 U6521 ( .A(n5096), .B(n5095), .ZN(n6213) );
  OR2_X1 U6522 ( .A1(n6213), .A2(n5097), .ZN(n5098) );
  NAND2_X1 U6523 ( .A1(n5099), .A2(n5098), .ZN(n7264) );
  OR2_X1 U6524 ( .A1(n7262), .A2(n7264), .ZN(n8958) );
  NAND2_X1 U6525 ( .A1(n7264), .A2(n7262), .ZN(n8965) );
  NAND2_X1 U6526 ( .A1(n8958), .A2(n8965), .ZN(n9095) );
  INV_X1 U6527 ( .A(n7264), .ZN(n7253) );
  NAND2_X1 U6528 ( .A1(n7253), .A2(n7262), .ZN(n5100) );
  NAND2_X1 U6529 ( .A1(n5139), .A2(n5101), .ZN(n5103) );
  XNOR2_X1 U6530 ( .A(n5103), .B(n5102), .ZN(n6207) );
  NAND2_X1 U6531 ( .A1(n6207), .A2(n5122), .ZN(n5107) );
  NAND2_X1 U6532 ( .A1(n5089), .A2(n5104), .ZN(n5123) );
  NAND2_X1 U6533 ( .A1(n5123), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5105) );
  XNOR2_X1 U6534 ( .A(n5105), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6522) );
  AOI22_X1 U6535 ( .A1(n5298), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6161), .B2(
        n6522), .ZN(n5106) );
  NAND2_X2 U6536 ( .A1(n5107), .A2(n5106), .ZN(n7350) );
  INV_X1 U6537 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5108) );
  NAND2_X1 U6538 ( .A1(n5109), .A2(n5108), .ZN(n5110) );
  NAND2_X1 U6539 ( .A1(n5130), .A2(n5110), .ZN(n7338) );
  OR2_X1 U6540 ( .A1(n5049), .A2(n7338), .ZN(n5114) );
  NAND2_X1 U6541 ( .A1(n5492), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5113) );
  NAND2_X1 U6542 ( .A1(n6245), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5112) );
  NAND2_X1 U6543 ( .A1(n6244), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5111) );
  NAND4_X1 U6544 ( .A1(n5114), .A2(n5113), .A3(n5112), .A4(n5111), .ZN(n9255)
         );
  OR2_X1 U6545 ( .A1(n7350), .A2(n7157), .ZN(n8967) );
  NAND2_X1 U6546 ( .A1(n7350), .A2(n7157), .ZN(n9122) );
  NAND2_X1 U6547 ( .A1(n8967), .A2(n9122), .ZN(n9088) );
  NAND2_X1 U6548 ( .A1(n6990), .A2(n9088), .ZN(n6989) );
  OR2_X1 U6549 ( .A1(n7350), .A2(n9255), .ZN(n5115) );
  NAND2_X1 U6550 ( .A1(n6989), .A2(n5115), .ZN(n5116) );
  NAND2_X1 U6551 ( .A1(n5139), .A2(n5117), .ZN(n5119) );
  AND2_X1 U6552 ( .A1(n5119), .A2(n5118), .ZN(n5121) );
  XNOR2_X1 U6553 ( .A(n5121), .B(n5120), .ZN(n6227) );
  NAND2_X1 U6554 ( .A1(n6227), .A2(n5122), .ZN(n5129) );
  NOR2_X1 U6555 ( .A1(n5124), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5158) );
  INV_X1 U6556 ( .A(n5158), .ZN(n5127) );
  NAND2_X1 U6557 ( .A1(n5124), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5125) );
  MUX2_X1 U6558 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5125), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n5126) );
  AOI22_X1 U6559 ( .A1(n5298), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6161), .B2(
        n9772), .ZN(n5128) );
  INV_X1 U6560 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7528) );
  NAND2_X1 U6561 ( .A1(n5130), .A2(n7528), .ZN(n5131) );
  NAND2_X1 U6562 ( .A1(n5148), .A2(n5131), .ZN(n7531) );
  OR2_X1 U6563 ( .A1(n5049), .A2(n7531), .ZN(n5135) );
  NAND2_X1 U6564 ( .A1(n6244), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5134) );
  NAND2_X1 U6565 ( .A1(n5492), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5133) );
  NAND2_X1 U6566 ( .A1(n6245), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5132) );
  NAND4_X1 U6567 ( .A1(n5135), .A2(n5134), .A3(n5133), .A4(n5132), .ZN(n9254)
         );
  INV_X1 U6568 ( .A(n9254), .ZN(n6994) );
  OR2_X1 U6569 ( .A1(n7540), .A2(n6994), .ZN(n8971) );
  NAND2_X1 U6570 ( .A1(n7540), .A2(n6994), .ZN(n9123) );
  INV_X1 U6571 ( .A(n9098), .ZN(n5136) );
  NAND2_X1 U6572 ( .A1(n7540), .A2(n9254), .ZN(n5137) );
  NAND2_X1 U6573 ( .A1(n5139), .A2(n5138), .ZN(n5141) );
  NAND2_X1 U6574 ( .A1(n5141), .A2(n5140), .ZN(n5143) );
  XNOR2_X1 U6575 ( .A(n5143), .B(n5142), .ZN(n6204) );
  NAND2_X1 U6576 ( .A1(n6204), .A2(n8114), .ZN(n5146) );
  OR2_X1 U6577 ( .A1(n5158), .A2(n9631), .ZN(n5144) );
  XNOR2_X1 U6578 ( .A(n5144), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6629) );
  AOI22_X1 U6579 ( .A1(n5298), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6161), .B2(
        n6629), .ZN(n5145) );
  NAND2_X1 U6580 ( .A1(n5146), .A2(n5145), .ZN(n7494) );
  NAND2_X1 U6581 ( .A1(n5148), .A2(n5147), .ZN(n5149) );
  NAND2_X1 U6582 ( .A1(n5162), .A2(n5149), .ZN(n7113) );
  OR2_X1 U6583 ( .A1(n5049), .A2(n7113), .ZN(n5153) );
  NAND2_X1 U6584 ( .A1(n5492), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5152) );
  NAND2_X1 U6585 ( .A1(n6245), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5151) );
  NAND2_X1 U6586 ( .A1(n6244), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5150) );
  NAND4_X1 U6587 ( .A1(n5153), .A2(n5152), .A3(n5151), .A4(n5150), .ZN(n9253)
         );
  AND2_X1 U6588 ( .A1(n7494), .A2(n9253), .ZN(n5154) );
  XNOR2_X1 U6589 ( .A(n5156), .B(n5155), .ZN(n6234) );
  NAND2_X1 U6590 ( .A1(n6234), .A2(n8114), .ZN(n5161) );
  INV_X1 U6591 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5157) );
  NAND2_X1 U6592 ( .A1(n5158), .A2(n5157), .ZN(n5172) );
  NAND2_X1 U6593 ( .A1(n5172), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5159) );
  XNOR2_X1 U6594 ( .A(n5159), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6684) );
  AOI22_X1 U6595 ( .A1(n5298), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6161), .B2(
        n6684), .ZN(n5160) );
  NAND2_X1 U6596 ( .A1(n5161), .A2(n5160), .ZN(n9694) );
  NAND2_X1 U6597 ( .A1(n5162), .A2(n6625), .ZN(n5163) );
  NAND2_X1 U6598 ( .A1(n5177), .A2(n5163), .ZN(n9689) );
  OR2_X1 U6599 ( .A1(n5049), .A2(n9689), .ZN(n5167) );
  NAND2_X1 U6600 ( .A1(n6244), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5166) );
  NAND2_X1 U6601 ( .A1(n5492), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5165) );
  NAND2_X1 U6602 ( .A1(n5491), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5164) );
  NAND4_X1 U6603 ( .A1(n5167), .A2(n5166), .A3(n5165), .A4(n5164), .ZN(n9252)
         );
  NAND2_X1 U6604 ( .A1(n9694), .A2(n7512), .ZN(n8978) );
  NAND2_X1 U6605 ( .A1(n9130), .A2(n8978), .ZN(n9676) );
  NAND2_X1 U6606 ( .A1(n9675), .A2(n9676), .ZN(n5169) );
  OR2_X1 U6607 ( .A1(n9694), .A2(n9252), .ZN(n5168) );
  NAND2_X1 U6608 ( .A1(n6238), .A2(n8114), .ZN(n5175) );
  OAI21_X1 U6609 ( .B1(n5172), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5173) );
  XNOR2_X1 U6610 ( .A(n5173), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7362) );
  AOI22_X1 U6611 ( .A1(n5298), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6161), .B2(
        n7362), .ZN(n5174) );
  INV_X1 U6612 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5176) );
  NAND2_X1 U6613 ( .A1(n5177), .A2(n5176), .ZN(n5178) );
  NAND2_X1 U6614 ( .A1(n5189), .A2(n5178), .ZN(n8907) );
  OR2_X1 U6615 ( .A1(n5049), .A2(n8907), .ZN(n5182) );
  NAND2_X1 U6616 ( .A1(n6244), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5181) );
  NAND2_X1 U6617 ( .A1(n5492), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5180) );
  NAND2_X1 U6618 ( .A1(n6245), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5179) );
  NAND4_X1 U6619 ( .A1(n5182), .A2(n5181), .A3(n5180), .A4(n5179), .ZN(n9251)
         );
  NAND2_X1 U6620 ( .A1(n8914), .A2(n9251), .ZN(n7304) );
  XNOR2_X1 U6621 ( .A(n5184), .B(n5183), .ZN(n6242) );
  NAND2_X1 U6622 ( .A1(n6242), .A2(n8114), .ZN(n5188) );
  OR2_X1 U6623 ( .A1(n5185), .A2(n9631), .ZN(n5186) );
  XNOR2_X1 U6624 ( .A(n5186), .B(P1_IR_REG_12__SCAN_IN), .ZN(n9786) );
  AOI22_X1 U6625 ( .A1(n5298), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6161), .B2(
        n9786), .ZN(n5187) );
  INV_X1 U6626 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n8824) );
  NAND2_X1 U6627 ( .A1(n5189), .A2(n8824), .ZN(n5190) );
  NAND2_X1 U6628 ( .A1(n5206), .A2(n5190), .ZN(n8828) );
  OR2_X1 U6629 ( .A1(n5049), .A2(n8828), .ZN(n5194) );
  NAND2_X1 U6630 ( .A1(n5051), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5193) );
  NAND2_X1 U6631 ( .A1(n5491), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5192) );
  NAND2_X1 U6632 ( .A1(n6244), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5191) );
  NAND4_X1 U6633 ( .A1(n5194), .A2(n5193), .A3(n5192), .A4(n5191), .ZN(n9250)
         );
  NAND2_X1 U6634 ( .A1(n8830), .A2(n9250), .ZN(n5195) );
  AND2_X1 U6635 ( .A1(n7304), .A2(n5195), .ZN(n5197) );
  INV_X1 U6636 ( .A(n5195), .ZN(n5196) );
  OR2_X1 U6637 ( .A1(n8830), .A2(n8885), .ZN(n8990) );
  NAND2_X1 U6638 ( .A1(n8830), .A2(n8885), .ZN(n9125) );
  NAND2_X1 U6639 ( .A1(n8990), .A2(n9125), .ZN(n9101) );
  OR2_X1 U6640 ( .A1(n5199), .A2(n5198), .ZN(n5200) );
  NAND2_X1 U6641 ( .A1(n5201), .A2(n5200), .ZN(n6275) );
  NAND2_X1 U6642 ( .A1(n6275), .A2(n8114), .ZN(n5204) );
  NAND2_X1 U6643 ( .A1(n5215), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5202) );
  XNOR2_X1 U6644 ( .A(n5202), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9801) );
  AOI22_X1 U6645 ( .A1(n5298), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6161), .B2(
        n9801), .ZN(n5203) );
  NAND2_X1 U6646 ( .A1(n5206), .A2(n5205), .ZN(n5207) );
  NAND2_X1 U6647 ( .A1(n5221), .A2(n5207), .ZN(n8888) );
  OR2_X1 U6648 ( .A1(n5049), .A2(n8888), .ZN(n5211) );
  NAND2_X1 U6649 ( .A1(n6244), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5210) );
  NAND2_X1 U6650 ( .A1(n5492), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5209) );
  NAND2_X1 U6651 ( .A1(n6245), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5208) );
  NAND4_X1 U6652 ( .A1(n5211), .A2(n5210), .A3(n5209), .A4(n5208), .ZN(n9249)
         );
  AND2_X1 U6653 ( .A1(n9605), .A2(n9249), .ZN(n5212) );
  XNOR2_X1 U6654 ( .A(n5214), .B(n5213), .ZN(n6264) );
  NAND2_X1 U6655 ( .A1(n6264), .A2(n8114), .ZN(n5219) );
  INV_X1 U6656 ( .A(n5215), .ZN(n5217) );
  NAND2_X1 U6657 ( .A1(n5251), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5232) );
  XNOR2_X1 U6658 ( .A(n5232), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7371) );
  AOI22_X1 U6659 ( .A1(n5298), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6161), .B2(
        n7371), .ZN(n5218) );
  INV_X1 U6660 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5220) );
  NAND2_X1 U6661 ( .A1(n5221), .A2(n5220), .ZN(n5222) );
  NAND2_X1 U6662 ( .A1(n5238), .A2(n5222), .ZN(n8782) );
  OR2_X1 U6663 ( .A1(n5049), .A2(n8782), .ZN(n5226) );
  NAND2_X1 U6664 ( .A1(n5492), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5225) );
  NAND2_X1 U6665 ( .A1(n6245), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5224) );
  NAND2_X1 U6666 ( .A1(n6244), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5223) );
  NAND4_X1 U6667 ( .A1(n5226), .A2(n5225), .A3(n5224), .A4(n5223), .ZN(n9248)
         );
  NOR2_X1 U6668 ( .A1(n8977), .A2(n9248), .ZN(n5228) );
  NAND2_X1 U6669 ( .A1(n8977), .A2(n9248), .ZN(n5227) );
  XNOR2_X1 U6670 ( .A(n5230), .B(n5229), .ZN(n6405) );
  NAND2_X1 U6671 ( .A1(n6405), .A2(n8114), .ZN(n5236) );
  INV_X1 U6672 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5231) );
  NAND2_X1 U6673 ( .A1(n5232), .A2(n5231), .ZN(n5233) );
  NAND2_X1 U6674 ( .A1(n5233), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5234) );
  XNOR2_X1 U6675 ( .A(n5234), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9819) );
  AOI22_X1 U6676 ( .A1(n5298), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6161), .B2(
        n9819), .ZN(n5235) );
  NAND2_X1 U6677 ( .A1(n5238), .A2(n5237), .ZN(n5239) );
  NAND2_X1 U6678 ( .A1(n5256), .A2(n5239), .ZN(n7699) );
  OR2_X1 U6679 ( .A1(n5049), .A2(n7699), .ZN(n5243) );
  NAND2_X1 U6680 ( .A1(n6244), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5242) );
  NAND2_X1 U6681 ( .A1(n5051), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5241) );
  NAND2_X1 U6682 ( .A1(n5491), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5240) );
  NAND4_X1 U6683 ( .A1(n5243), .A2(n5242), .A3(n5241), .A4(n5240), .ZN(n9247)
         );
  OR2_X1 U6684 ( .A1(n9599), .A2(n9247), .ZN(n5244) );
  NAND2_X1 U6685 ( .A1(n7592), .A2(n5244), .ZN(n5246) );
  NAND2_X1 U6686 ( .A1(n9599), .A2(n9247), .ZN(n5245) );
  NAND2_X1 U6687 ( .A1(n5246), .A2(n5245), .ZN(n9506) );
  XNOR2_X1 U6688 ( .A(n5248), .B(n5247), .ZN(n6574) );
  NAND2_X1 U6689 ( .A1(n6574), .A2(n8114), .ZN(n5254) );
  INV_X1 U6690 ( .A(n5249), .ZN(n5250) );
  OR2_X1 U6691 ( .A1(n4350), .A2(n9631), .ZN(n5252) );
  XNOR2_X1 U6692 ( .A(n5252), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9831) );
  AOI22_X1 U6693 ( .A1(n5298), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6161), .B2(
        n9831), .ZN(n5253) );
  INV_X1 U6694 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5255) );
  NAND2_X1 U6695 ( .A1(n5256), .A2(n5255), .ZN(n5257) );
  NAND2_X1 U6696 ( .A1(n5270), .A2(n5257), .ZN(n9513) );
  OR2_X1 U6697 ( .A1(n9513), .A2(n5049), .ZN(n5261) );
  NAND2_X1 U6698 ( .A1(n5492), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5260) );
  NAND2_X1 U6699 ( .A1(n5491), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5259) );
  NAND2_X1 U6700 ( .A1(n6244), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5258) );
  NAND4_X1 U6701 ( .A1(n5261), .A2(n5260), .A3(n5259), .A4(n5258), .ZN(n9498)
         );
  INV_X1 U6702 ( .A(n9498), .ZN(n8005) );
  OR2_X1 U6703 ( .A1(n9594), .A2(n8005), .ZN(n9141) );
  NAND2_X1 U6704 ( .A1(n9594), .A2(n8005), .ZN(n9120) );
  NAND2_X1 U6705 ( .A1(n9506), .A2(n9508), .ZN(n5263) );
  NAND2_X1 U6706 ( .A1(n9594), .A2(n9498), .ZN(n5262) );
  NAND2_X1 U6707 ( .A1(n5263), .A2(n5262), .ZN(n9487) );
  XNOR2_X1 U6708 ( .A(n5265), .B(n5264), .ZN(n6656) );
  NAND2_X1 U6709 ( .A1(n6656), .A2(n8114), .ZN(n5268) );
  NAND2_X1 U6710 ( .A1(n5295), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5281) );
  XNOR2_X1 U6711 ( .A(n5281), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9842) );
  AOI22_X1 U6712 ( .A1(n5298), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6161), .B2(
        n9842), .ZN(n5267) );
  NAND2_X1 U6713 ( .A1(n5270), .A2(n5269), .ZN(n5271) );
  NAND2_X1 U6714 ( .A1(n5288), .A2(n5271), .ZN(n9491) );
  NAND2_X1 U6715 ( .A1(n5492), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5273) );
  NAND2_X1 U6716 ( .A1(n6244), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5272) );
  AND2_X1 U6717 ( .A1(n5273), .A2(n5272), .ZN(n5275) );
  NAND2_X1 U6718 ( .A1(n6245), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5274) );
  OAI211_X1 U6719 ( .C1(n9491), .C2(n5049), .A(n5275), .B(n5274), .ZN(n9471)
         );
  AND2_X1 U6720 ( .A1(n9587), .A2(n9471), .ZN(n5277) );
  OR2_X1 U6721 ( .A1(n9587), .A2(n9471), .ZN(n5276) );
  XNOR2_X1 U6722 ( .A(n5279), .B(n5278), .ZN(n6814) );
  NAND2_X1 U6723 ( .A1(n6814), .A2(n8114), .ZN(n5285) );
  NAND2_X1 U6724 ( .A1(n5281), .A2(n5280), .ZN(n5282) );
  NAND2_X1 U6725 ( .A1(n5282), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5283) );
  XNOR2_X1 U6726 ( .A(n5283), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9858) );
  AOI22_X1 U6727 ( .A1(n5298), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6161), .B2(
        n9858), .ZN(n5284) );
  INV_X1 U6728 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9478) );
  INV_X1 U6729 ( .A(n5286), .ZN(n5302) );
  NAND2_X1 U6730 ( .A1(n5288), .A2(n5287), .ZN(n5289) );
  NAND2_X1 U6731 ( .A1(n5302), .A2(n5289), .ZN(n9477) );
  OR2_X1 U6732 ( .A1(n9477), .A2(n5049), .ZN(n5291) );
  AOI22_X1 U6733 ( .A1(n6244), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n5492), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n5290) );
  OAI211_X1 U6734 ( .C1(n5041), .C2(n9478), .A(n5291), .B(n5290), .ZN(n9500)
         );
  INV_X1 U6735 ( .A(n9500), .ZN(n8853) );
  OR2_X1 U6736 ( .A1(n9582), .A2(n8853), .ZN(n8951) );
  NAND2_X1 U6737 ( .A1(n9582), .A2(n8853), .ZN(n9458) );
  XNOR2_X1 U6738 ( .A(n5293), .B(n5292), .ZN(n6890) );
  NAND2_X1 U6739 ( .A1(n6890), .A2(n8114), .ZN(n5300) );
  INV_X1 U6740 ( .A(n5454), .ZN(n5296) );
  NAND2_X1 U6741 ( .A1(n5296), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5297) );
  AOI22_X1 U6742 ( .A1(n5298), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9434), .B2(
        n6161), .ZN(n5299) );
  INV_X1 U6743 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5301) );
  NAND2_X1 U6744 ( .A1(n5302), .A2(n5301), .ZN(n5303) );
  NAND2_X1 U6745 ( .A1(n5315), .A2(n5303), .ZN(n9454) );
  OR2_X1 U6746 ( .A1(n9454), .A2(n5049), .ZN(n5308) );
  INV_X1 U6747 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9285) );
  NAND2_X1 U6748 ( .A1(n5051), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5305) );
  NAND2_X1 U6749 ( .A1(n5491), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5304) );
  OAI211_X1 U6750 ( .C1(n9285), .C2(n5074), .A(n5305), .B(n5304), .ZN(n5306)
         );
  INV_X1 U6751 ( .A(n5306), .ZN(n5307) );
  NAND2_X1 U6752 ( .A1(n5308), .A2(n5307), .ZN(n9472) );
  NAND2_X1 U6753 ( .A1(n9575), .A2(n9472), .ZN(n5309) );
  XNOR2_X1 U6754 ( .A(n5312), .B(n5311), .ZN(n6965) );
  NAND2_X1 U6755 ( .A1(n6965), .A2(n8114), .ZN(n5314) );
  OR2_X1 U6756 ( .A1(n8115), .A2(n6966), .ZN(n5313) );
  NAND2_X1 U6757 ( .A1(n5315), .A2(n8872), .ZN(n5316) );
  NAND2_X1 U6758 ( .A1(n5328), .A2(n5316), .ZN(n9441) );
  OR2_X1 U6759 ( .A1(n9441), .A2(n5049), .ZN(n5322) );
  INV_X1 U6760 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n5319) );
  NAND2_X1 U6761 ( .A1(n5492), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5318) );
  NAND2_X1 U6762 ( .A1(n5491), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5317) );
  OAI211_X1 U6763 ( .C1(n5319), .C2(n5074), .A(n5318), .B(n5317), .ZN(n5320)
         );
  INV_X1 U6764 ( .A(n5320), .ZN(n5321) );
  NAND2_X1 U6765 ( .A1(n5322), .A2(n5321), .ZN(n9463) );
  XNOR2_X1 U6766 ( .A(n5324), .B(n5323), .ZN(n7018) );
  NAND2_X1 U6767 ( .A1(n7018), .A2(n8114), .ZN(n5326) );
  OR2_X1 U6768 ( .A1(n8115), .A2(n7066), .ZN(n5325) );
  NAND2_X1 U6769 ( .A1(n5328), .A2(n5327), .ZN(n5329) );
  AND2_X1 U6770 ( .A1(n5341), .A2(n5329), .ZN(n9432) );
  NAND2_X1 U6771 ( .A1(n9432), .A2(n5416), .ZN(n5336) );
  INV_X1 U6772 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n5333) );
  NAND2_X1 U6773 ( .A1(n6244), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5331) );
  NAND2_X1 U6774 ( .A1(n5051), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5330) );
  OAI211_X1 U6775 ( .C1(n5333), .C2(n5332), .A(n5331), .B(n5330), .ZN(n5334)
         );
  INV_X1 U6776 ( .A(n5334), .ZN(n5335) );
  NAND2_X1 U6777 ( .A1(n5336), .A2(n5335), .ZN(n9447) );
  NAND2_X1 U6778 ( .A1(n9429), .A2(n9411), .ZN(n9031) );
  INV_X1 U6779 ( .A(n9429), .ZN(n9565) );
  XNOR2_X1 U6780 ( .A(n5338), .B(n5337), .ZN(n7777) );
  NAND2_X1 U6781 ( .A1(n7777), .A2(n8114), .ZN(n5340) );
  OR2_X1 U6782 ( .A1(n8115), .A2(n7778), .ZN(n5339) );
  INV_X1 U6783 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8896) );
  NAND2_X1 U6784 ( .A1(n5341), .A2(n8896), .ZN(n5342) );
  NAND2_X1 U6785 ( .A1(n5357), .A2(n5342), .ZN(n9414) );
  OR2_X1 U6786 ( .A1(n9414), .A2(n5049), .ZN(n5347) );
  INV_X1 U6787 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n6355) );
  NAND2_X1 U6788 ( .A1(n5491), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5344) );
  NAND2_X1 U6789 ( .A1(n5492), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5343) );
  OAI211_X1 U6790 ( .C1(n5074), .C2(n6355), .A(n5344), .B(n5343), .ZN(n5345)
         );
  INV_X1 U6791 ( .A(n5345), .ZN(n5346) );
  NAND2_X1 U6792 ( .A1(n5347), .A2(n5346), .ZN(n9426) );
  INV_X1 U6793 ( .A(n9560), .ZN(n8902) );
  INV_X1 U6794 ( .A(n9426), .ZN(n8813) );
  NAND2_X1 U6795 ( .A1(n5348), .A2(n4840), .ZN(n9390) );
  INV_X1 U6796 ( .A(n5349), .ZN(n5351) );
  NAND2_X1 U6797 ( .A1(n5351), .A2(n5350), .ZN(n5353) );
  NAND2_X1 U6798 ( .A1(n5353), .A2(n5352), .ZN(n7279) );
  NAND2_X1 U6799 ( .A1(n7279), .A2(n8114), .ZN(n5355) );
  OR2_X1 U6800 ( .A1(n8115), .A2(n7282), .ZN(n5354) );
  INV_X1 U6801 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5356) );
  NAND2_X1 U6802 ( .A1(n5357), .A2(n5356), .ZN(n5358) );
  NAND2_X1 U6803 ( .A1(n5359), .A2(n5358), .ZN(n9400) );
  OR2_X1 U6804 ( .A1(n9400), .A2(n5049), .ZN(n5365) );
  INV_X1 U6805 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n5362) );
  NAND2_X1 U6806 ( .A1(n5051), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U6807 ( .A1(n5491), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5360) );
  OAI211_X1 U6808 ( .C1(n5074), .C2(n5362), .A(n5361), .B(n5360), .ZN(n5363)
         );
  INV_X1 U6809 ( .A(n5363), .ZN(n5364) );
  NAND2_X1 U6810 ( .A1(n5365), .A2(n5364), .ZN(n9246) );
  INV_X1 U6811 ( .A(n5366), .ZN(n5370) );
  INV_X1 U6812 ( .A(n5367), .ZN(n5368) );
  NAND2_X1 U6813 ( .A1(n5368), .A2(SI_24_), .ZN(n5369) );
  INV_X1 U6814 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7575) );
  INV_X1 U6815 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7571) );
  MUX2_X1 U6816 ( .A(n7575), .B(n7571), .S(n5577), .Z(n5373) );
  INV_X1 U6817 ( .A(SI_25_), .ZN(n5372) );
  NAND2_X1 U6818 ( .A1(n5373), .A2(n5372), .ZN(n5391) );
  INV_X1 U6819 ( .A(n5373), .ZN(n5374) );
  NAND2_X1 U6820 ( .A1(n5374), .A2(SI_25_), .ZN(n5375) );
  NAND2_X1 U6821 ( .A1(n5391), .A2(n5375), .ZN(n5389) );
  NAND2_X1 U6822 ( .A1(n7568), .A2(n8114), .ZN(n5377) );
  OR2_X1 U6823 ( .A1(n8115), .A2(n7571), .ZN(n5376) );
  INV_X1 U6824 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5379) );
  NAND2_X1 U6825 ( .A1(n5380), .A2(n5379), .ZN(n5381) );
  NAND2_X1 U6826 ( .A1(n5399), .A2(n5381), .ZN(n9364) );
  INV_X1 U6827 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n5384) );
  NAND2_X1 U6828 ( .A1(n5051), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5383) );
  NAND2_X1 U6829 ( .A1(n5491), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5382) );
  OAI211_X1 U6830 ( .C1(n5384), .C2(n5074), .A(n5383), .B(n5382), .ZN(n5385)
         );
  INV_X1 U6831 ( .A(n5385), .ZN(n5386) );
  NAND2_X1 U6832 ( .A1(n9543), .A2(n9382), .ZN(n9043) );
  OAI22_X1 U6833 ( .A1(n9361), .A2(n9370), .B1(n9355), .B2(n9543), .ZN(n9347)
         );
  INV_X1 U6834 ( .A(n5389), .ZN(n5390) );
  INV_X1 U6835 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7649) );
  INV_X1 U6836 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7609) );
  MUX2_X1 U6837 ( .A(n7649), .B(n7609), .S(n6203), .Z(n5394) );
  INV_X1 U6838 ( .A(SI_26_), .ZN(n5393) );
  NAND2_X1 U6839 ( .A1(n5394), .A2(n5393), .ZN(n5409) );
  INV_X1 U6840 ( .A(n5394), .ZN(n5395) );
  NAND2_X1 U6841 ( .A1(n5395), .A2(SI_26_), .ZN(n5396) );
  AND2_X1 U6842 ( .A1(n5409), .A2(n5396), .ZN(n5407) );
  OR2_X1 U6843 ( .A1(n8115), .A2(n7609), .ZN(n5397) );
  INV_X1 U6844 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8940) );
  NAND2_X1 U6845 ( .A1(n5399), .A2(n8940), .ZN(n5400) );
  NAND2_X1 U6846 ( .A1(n9349), .A2(n5416), .ZN(n5406) );
  INV_X1 U6847 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n5403) );
  NAND2_X1 U6848 ( .A1(n5492), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5402) );
  NAND2_X1 U6849 ( .A1(n6244), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5401) );
  OAI211_X1 U6850 ( .C1(n5332), .C2(n5403), .A(n5402), .B(n5401), .ZN(n5404)
         );
  INV_X1 U6851 ( .A(n5404), .ZN(n5405) );
  NAND2_X1 U6852 ( .A1(n9538), .A2(n9372), .ZN(n9080) );
  INV_X1 U6853 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7730) );
  INV_X1 U6854 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7706) );
  MUX2_X1 U6855 ( .A(n7730), .B(n7706), .S(n5577), .Z(n5411) );
  INV_X1 U6856 ( .A(SI_27_), .ZN(n6278) );
  NAND2_X1 U6857 ( .A1(n5411), .A2(n6278), .ZN(n5425) );
  INV_X1 U6858 ( .A(n5411), .ZN(n5412) );
  NAND2_X1 U6859 ( .A1(n5412), .A2(SI_27_), .ZN(n5413) );
  AND2_X1 U6860 ( .A1(n5425), .A2(n5413), .ZN(n5424) );
  NAND2_X1 U6861 ( .A1(n7728), .A2(n8114), .ZN(n5415) );
  OR2_X1 U6862 ( .A1(n8115), .A2(n7706), .ZN(n5414) );
  XNOR2_X1 U6863 ( .A(n5430), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9341) );
  NAND2_X1 U6864 ( .A1(n9341), .A2(n5416), .ZN(n5422) );
  INV_X1 U6865 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n5419) );
  NAND2_X1 U6866 ( .A1(n5051), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5418) );
  NAND2_X1 U6867 ( .A1(n5491), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5417) );
  OAI211_X1 U6868 ( .C1(n5419), .C2(n5074), .A(n5418), .B(n5417), .ZN(n5420)
         );
  INV_X1 U6869 ( .A(n5420), .ZN(n5421) );
  NAND2_X1 U6870 ( .A1(n9535), .A2(n9320), .ZN(n9059) );
  INV_X1 U6871 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7742) );
  INV_X1 U6872 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7744) );
  MUX2_X1 U6873 ( .A(n7742), .B(n7744), .S(n6203), .Z(n5443) );
  XNOR2_X1 U6874 ( .A(n5443), .B(SI_28_), .ZN(n5440) );
  NAND2_X1 U6875 ( .A1(n7743), .A2(n8114), .ZN(n5427) );
  OR2_X1 U6876 ( .A1(n8115), .A2(n7744), .ZN(n5426) );
  INV_X1 U6877 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5429) );
  INV_X1 U6878 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5428) );
  OAI21_X1 U6879 ( .B1(n5430), .B2(n5429), .A(n5428), .ZN(n5433) );
  INV_X1 U6880 ( .A(n5430), .ZN(n5432) );
  AND2_X1 U6881 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5431) );
  NAND2_X1 U6882 ( .A1(n5432), .A2(n5431), .ZN(n9304) );
  NAND2_X1 U6883 ( .A1(n5433), .A2(n9304), .ZN(n8102) );
  INV_X1 U6884 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U6885 ( .A1(n5491), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5435) );
  NAND2_X1 U6886 ( .A1(n5492), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5434) );
  OAI211_X1 U6887 ( .C1(n5074), .C2(n5436), .A(n5435), .B(n5434), .ZN(n5437)
         );
  INV_X1 U6888 ( .A(n5437), .ZN(n5438) );
  NAND2_X1 U6889 ( .A1(n9530), .A2(n9337), .ZN(n9060) );
  INV_X1 U6890 ( .A(SI_28_), .ZN(n5442) );
  MUX2_X1 U6891 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n5577), .Z(n7783) );
  INV_X1 U6892 ( .A(SI_29_), .ZN(n7781) );
  XNOR2_X1 U6893 ( .A(n7783), .B(n7781), .ZN(n5444) );
  NAND2_X1 U6894 ( .A1(n8766), .A2(n8114), .ZN(n5446) );
  INV_X1 U6895 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9642) );
  OR2_X1 U6896 ( .A1(n8115), .A2(n9642), .ZN(n5445) );
  OR2_X1 U6897 ( .A1(n9304), .A2(n5049), .ZN(n5451) );
  NAND2_X1 U6898 ( .A1(n6244), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5449) );
  NAND2_X1 U6899 ( .A1(n5051), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5448) );
  NAND2_X1 U6900 ( .A1(n6245), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5447) );
  AND3_X1 U6901 ( .A1(n5449), .A2(n5448), .A3(n5447), .ZN(n5450) );
  NAND2_X1 U6902 ( .A1(n9306), .A2(n9321), .ZN(n9223) );
  XNOR2_X1 U6903 ( .A(n5452), .B(n9114), .ZN(n9302) );
  NAND2_X1 U6904 ( .A1(n5454), .A2(n5453), .ZN(n5455) );
  INV_X1 U6905 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5456) );
  NAND2_X1 U6906 ( .A1(n5457), .A2(n5456), .ZN(n5460) );
  NAND2_X1 U6907 ( .A1(n5460), .A2(n5458), .ZN(n5464) );
  XNOR2_X1 U6908 ( .A(n5459), .B(P1_IR_REG_20__SCAN_IN), .ZN(n9183) );
  INV_X1 U6909 ( .A(n6417), .ZN(n5463) );
  OR2_X1 U6910 ( .A1(n5463), .A2(n6554), .ZN(n5466) );
  INV_X1 U6911 ( .A(n9183), .ZN(n9232) );
  NAND3_X1 U6912 ( .A1(n6414), .A2(n9186), .A3(n6415), .ZN(n5465) );
  AND2_X1 U6913 ( .A1(n5466), .A2(n5465), .ZN(n6819) );
  NAND2_X1 U6914 ( .A1(n6819), .A2(n9609), .ZN(n9926) );
  NAND2_X1 U6915 ( .A1(n9302), .A2(n9926), .ZN(n5501) );
  AND2_X1 U6916 ( .A1(n6897), .A2(n6900), .ZN(n6895) );
  NAND2_X1 U6917 ( .A1(n9093), .A2(n6895), .ZN(n5468) );
  NAND2_X1 U6918 ( .A1(n6901), .A2(n6557), .ZN(n5467) );
  INV_X1 U6919 ( .A(n9198), .ZN(n5469) );
  INV_X1 U6920 ( .A(n9199), .ZN(n5470) );
  AND2_X1 U6922 ( .A1(n7153), .A2(n8965), .ZN(n9200) );
  INV_X1 U6923 ( .A(n8955), .ZN(n5472) );
  NAND2_X1 U6924 ( .A1(n5472), .A2(n8965), .ZN(n9202) );
  AND2_X1 U6925 ( .A1(n9202), .A2(n8958), .ZN(n5473) );
  INV_X1 U6926 ( .A(n9123), .ZN(n8981) );
  INV_X1 U6927 ( .A(n9253), .ZN(n9683) );
  OR2_X1 U6928 ( .A1(n7494), .A2(n9683), .ZN(n8974) );
  AND2_X1 U6929 ( .A1(n8974), .A2(n8971), .ZN(n9129) );
  NAND2_X1 U6930 ( .A1(n7494), .A2(n9683), .ZN(n8972) );
  INV_X1 U6931 ( .A(n9676), .ZN(n9679) );
  NAND2_X1 U6932 ( .A1(n8978), .A2(n8972), .ZN(n8983) );
  NAND2_X1 U6933 ( .A1(n8983), .A2(n9130), .ZN(n7220) );
  INV_X1 U6934 ( .A(n9251), .ZN(n9680) );
  NAND2_X1 U6935 ( .A1(n8914), .A2(n9680), .ZN(n9002) );
  OR2_X1 U6936 ( .A1(n8914), .A2(n9680), .ZN(n8989) );
  NAND2_X1 U6937 ( .A1(n5475), .A2(n8989), .ZN(n7307) );
  INV_X1 U6938 ( .A(n8990), .ZN(n5476) );
  OAI21_X2 U6939 ( .B1(n7307), .B2(n5476), .A(n9125), .ZN(n7454) );
  INV_X1 U6940 ( .A(n9249), .ZN(n8825) );
  OR2_X1 U6941 ( .A1(n9605), .A2(n8825), .ZN(n8992) );
  NAND2_X1 U6942 ( .A1(n9605), .A2(n8825), .ZN(n9000) );
  NAND2_X1 U6943 ( .A1(n7454), .A2(n9087), .ZN(n7453) );
  NAND2_X1 U6944 ( .A1(n7453), .A2(n9000), .ZN(n7543) );
  INV_X1 U6945 ( .A(n9248), .ZN(n8976) );
  XNOR2_X1 U6946 ( .A(n8977), .B(n8976), .ZN(n9107) );
  INV_X1 U6947 ( .A(n9247), .ZN(n9511) );
  NAND2_X1 U6948 ( .A1(n9599), .A2(n9511), .ZN(n9138) );
  OR2_X1 U6949 ( .A1(n9599), .A2(n9511), .ZN(n9140) );
  INV_X1 U6950 ( .A(n9471), .ZN(n9512) );
  AND2_X1 U6951 ( .A1(n9587), .A2(n9512), .ZN(n9121) );
  OR2_X1 U6952 ( .A1(n9587), .A2(n9512), .ZN(n9468) );
  AND2_X1 U6953 ( .A1(n8951), .A2(n9468), .ZN(n9151) );
  NAND2_X1 U6954 ( .A1(n9469), .A2(n9151), .ZN(n9460) );
  NAND2_X1 U6955 ( .A1(n9460), .A2(n9458), .ZN(n5478) );
  INV_X1 U6956 ( .A(n9472), .ZN(n8922) );
  OR2_X1 U6957 ( .A1(n9575), .A2(n8922), .ZN(n9023) );
  NAND2_X1 U6958 ( .A1(n9575), .A2(n8922), .ZN(n9022) );
  NAND2_X1 U6959 ( .A1(n5478), .A2(n9457), .ZN(n9462) );
  NAND2_X1 U6960 ( .A1(n9462), .A2(n9022), .ZN(n9446) );
  INV_X1 U6961 ( .A(n9463), .ZN(n5479) );
  AND2_X1 U6962 ( .A1(n9570), .A2(n5479), .ZN(n9084) );
  OR2_X1 U6963 ( .A1(n9560), .A2(n8813), .ZN(n9155) );
  NAND2_X1 U6964 ( .A1(n9560), .A2(n8813), .ZN(n9033) );
  NAND2_X1 U6965 ( .A1(n9409), .A2(n9083), .ZN(n5480) );
  NAND2_X1 U6966 ( .A1(n9555), .A2(n9412), .ZN(n9214) );
  NAND2_X1 U6967 ( .A1(n9378), .A2(n9214), .ZN(n9391) );
  OR2_X1 U6968 ( .A1(n9550), .A2(n5481), .ZN(n8946) );
  NAND2_X1 U6969 ( .A1(n9550), .A2(n5481), .ZN(n9368) );
  INV_X1 U6970 ( .A(n9372), .ZN(n5482) );
  OR2_X1 U6971 ( .A1(n9538), .A2(n5482), .ZN(n9041) );
  NAND2_X1 U6972 ( .A1(n9352), .A2(n9169), .ZN(n5483) );
  NAND2_X1 U6973 ( .A1(n9538), .A2(n5482), .ZN(n9162) );
  NAND2_X1 U6974 ( .A1(n5483), .A2(n9162), .ZN(n9331) );
  AND2_X1 U6975 ( .A1(n9167), .A2(n9316), .ZN(n9056) );
  INV_X1 U6976 ( .A(n9060), .ZN(n9055) );
  AOI21_X1 U6977 ( .B1(n9332), .B2(n9056), .A(n9055), .ZN(n5484) );
  XNOR2_X1 U6978 ( .A(n5484), .B(n9114), .ZN(n5487) );
  OR2_X1 U6979 ( .A1(n6414), .A2(n9878), .ZN(n5486) );
  OR2_X1 U6980 ( .A1(n5464), .A2(n9232), .ZN(n5485) );
  NAND2_X1 U6981 ( .A1(n5486), .A2(n5485), .ZN(n9685) );
  NAND2_X1 U6982 ( .A1(n5487), .A2(n9685), .ZN(n5497) );
  NAND2_X1 U6983 ( .A1(n5488), .A2(n9186), .ZN(n9079) );
  OR2_X1 U6984 ( .A1(n9079), .A2(n7745), .ZN(n9682) );
  INV_X1 U6985 ( .A(n7745), .ZN(n9736) );
  INV_X1 U6986 ( .A(P1_B_REG_SCAN_IN), .ZN(n5516) );
  NOR2_X1 U6987 ( .A1(n6649), .A2(n5516), .ZN(n5490) );
  NOR2_X1 U6988 ( .A1(n9681), .A2(n5490), .ZN(n8119) );
  NAND2_X1 U6989 ( .A1(n6244), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5495) );
  NAND2_X1 U6990 ( .A1(n5491), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5494) );
  NAND2_X1 U6991 ( .A1(n5492), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5493) );
  NAND3_X1 U6992 ( .A1(n5495), .A2(n5494), .A3(n5493), .ZN(n9244) );
  AOI22_X1 U6993 ( .A1(n9245), .A2(n9497), .B1(n8119), .B2(n9244), .ZN(n5496)
         );
  NAND2_X1 U6994 ( .A1(n5497), .A2(n5496), .ZN(n9311) );
  INV_X1 U6995 ( .A(n9535), .ZN(n9344) );
  INV_X1 U6996 ( .A(n9543), .ZN(n9367) );
  INV_X1 U6997 ( .A(n6900), .ZN(n6984) );
  NAND2_X1 U6998 ( .A1(n6984), .A2(n6556), .ZN(n7056) );
  INV_X1 U6999 ( .A(n7494), .ZN(n7517) );
  NAND2_X1 U7000 ( .A1(n7110), .A2(n7517), .ZN(n7111) );
  INV_X1 U7001 ( .A(n8830), .ZN(n9723) );
  INV_X1 U7002 ( .A(n9605), .ZN(n7461) );
  INV_X1 U7003 ( .A(n9594), .ZN(n9520) );
  INV_X1 U7004 ( .A(n9587), .ZN(n9494) );
  INV_X1 U7005 ( .A(n9570), .ZN(n9444) );
  NAND2_X1 U7006 ( .A1(n9344), .A2(n9348), .ZN(n9338) );
  NAND2_X1 U7007 ( .A1(n9306), .A2(n9322), .ZN(n5498) );
  NAND2_X1 U7008 ( .A1(n9297), .A2(n5498), .ZN(n9309) );
  NAND2_X1 U7009 ( .A1(n6414), .A2(n5464), .ZN(n6943) );
  OAI22_X1 U7010 ( .A1(n9309), .A2(n9921), .B1(n4550), .B2(n9911), .ZN(n5499)
         );
  NAND2_X1 U7011 ( .A1(n5501), .A2(n5500), .ZN(n6156) );
  OR2_X1 U7012 ( .A1(n9079), .A2(n6415), .ZN(n6908) );
  NAND2_X1 U7013 ( .A1(n5508), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5510) );
  NAND2_X1 U7014 ( .A1(n5510), .A2(n5502), .ZN(n5503) );
  NAND2_X1 U7015 ( .A1(n5503), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5504) );
  XNOR2_X1 U7016 ( .A(n5504), .B(P1_IR_REG_26__SCAN_IN), .ZN(n7608) );
  INV_X1 U7017 ( .A(n5505), .ZN(n5506) );
  NAND2_X1 U7018 ( .A1(n5506), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5507) );
  MUX2_X1 U7019 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5507), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n5509) );
  NAND2_X1 U7020 ( .A1(n5509), .A2(n5508), .ZN(n7387) );
  INV_X1 U7021 ( .A(n7387), .ZN(n5521) );
  XNOR2_X1 U7022 ( .A(n5510), .B(P1_IR_REG_25__SCAN_IN), .ZN(n7569) );
  AND2_X1 U7023 ( .A1(n5521), .A2(n7569), .ZN(n5511) );
  INV_X1 U7024 ( .A(n5512), .ZN(n5513) );
  NAND2_X1 U7025 ( .A1(n5513), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5514) );
  XNOR2_X1 U7026 ( .A(n5514), .B(n4970), .ZN(n7280) );
  AND2_X1 U7027 ( .A1(n7280), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5515) );
  AND2_X1 U7028 ( .A1(n6697), .A2(n5515), .ZN(n9895) );
  AND2_X1 U7029 ( .A1(n6908), .A2(n9895), .ZN(n6412) );
  NAND2_X1 U7030 ( .A1(n7387), .A2(P1_B_REG_SCAN_IN), .ZN(n5518) );
  NAND2_X1 U7031 ( .A1(n5521), .A2(n5516), .ZN(n5517) );
  OAI211_X1 U7032 ( .C1(n7569), .C2(n5518), .A(n7608), .B(n5517), .ZN(n9888)
         );
  OR2_X1 U7033 ( .A1(n9888), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5520) );
  OR2_X1 U7034 ( .A1(n7608), .A2(n7569), .ZN(n5519) );
  NAND2_X1 U7035 ( .A1(n5520), .A2(n5519), .ZN(n6905) );
  OAI211_X1 U7036 ( .C1(n9186), .C2(n9609), .A(n6412), .B(n6905), .ZN(n6155)
         );
  OR2_X1 U7037 ( .A1(n9888), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5523) );
  OR2_X1 U7038 ( .A1(n5521), .A2(n7608), .ZN(n5522) );
  AND2_X1 U7039 ( .A1(n5523), .A2(n5522), .ZN(n9630) );
  NOR4_X1 U7040 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n5527) );
  NOR4_X1 U7041 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n5526) );
  NOR4_X1 U7042 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5525) );
  NOR4_X1 U7043 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5524) );
  NAND4_X1 U7044 ( .A1(n5527), .A2(n5526), .A3(n5525), .A4(n5524), .ZN(n5533)
         );
  NOR2_X1 U7045 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .ZN(
        n5531) );
  NOR4_X1 U7046 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n5530) );
  NOR4_X1 U7047 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n5529) );
  NOR4_X1 U7048 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n5528) );
  NAND4_X1 U7049 ( .A1(n5531), .A2(n5530), .A3(n5529), .A4(n5528), .ZN(n5532)
         );
  NOR2_X1 U7050 ( .A1(n5533), .A2(n5532), .ZN(n5534) );
  OR2_X1 U7051 ( .A1(n9888), .A2(n5534), .ZN(n6153) );
  NAND2_X1 U7052 ( .A1(n9630), .A2(n6153), .ZN(n6409) );
  INV_X2 U7053 ( .A(n9933), .ZN(n9935) );
  NAND3_X1 U7054 ( .A1(n5598), .A2(n5536), .A3(n5535), .ZN(n5658) );
  INV_X1 U7055 ( .A(n5658), .ZN(n5539) );
  NOR3_X1 U7056 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .A3(
        P2_IR_REG_14__SCAN_IN), .ZN(n5542) );
  INV_X1 U7057 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5563) );
  NAND4_X1 U7058 ( .A1(n5565), .A2(n5563), .A3(n6279), .A4(n6025), .ZN(n5547)
         );
  INV_X1 U7059 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5545) );
  INV_X1 U7060 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5994) );
  INV_X1 U7061 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5544) );
  INV_X1 U7062 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5543) );
  NAND4_X1 U7063 ( .A1(n5545), .A2(n5994), .A3(n5544), .A4(n5543), .ZN(n5546)
         );
  INV_X1 U7064 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5548) );
  INV_X1 U7065 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5573) );
  INV_X1 U7066 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5550) );
  XNOR2_X2 U7067 ( .A(n5551), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5557) );
  OAI21_X1 U7068 ( .B1(n5552), .B2(n6000), .A(P2_IR_REG_29__SCAN_IN), .ZN(
        n5554) );
  NAND2_X1 U7069 ( .A1(n5918), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5562) );
  NAND2_X1 U7070 ( .A1(n5607), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U7071 ( .A1(n5603), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5560) );
  NAND2_X1 U7072 ( .A1(n5649), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5559) );
  NAND4_X1 U7073 ( .A1(n5562), .A2(n5561), .A3(n5560), .A4(n5559), .ZN(n8324)
         );
  INV_X1 U7074 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n6279) );
  NAND2_X1 U7075 ( .A1(n4323), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5566) );
  NAND2_X1 U7076 ( .A1(n5572), .A2(n5571), .ZN(n5568) );
  NAND2_X1 U7077 ( .A1(n5568), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5570) );
  INV_X1 U7078 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5569) );
  INV_X1 U7079 ( .A(n5585), .ZN(n5583) );
  INV_X1 U7080 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6390) );
  NAND2_X1 U7081 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5578) );
  INV_X1 U7082 ( .A(n9656), .ZN(n6197) );
  INV_X1 U7083 ( .A(n6052), .ZN(n7101) );
  NAND3_X1 U7084 ( .A1(n7983), .A2(n10027), .A3(n5579), .ZN(n5581) );
  XNOR2_X1 U7085 ( .A(n7101), .B(n5968), .ZN(n5584) );
  INV_X1 U7086 ( .A(n5584), .ZN(n5582) );
  NAND2_X1 U7087 ( .A1(n5585), .A2(n5584), .ZN(n5586) );
  NAND2_X1 U7088 ( .A1(n5603), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5590) );
  NAND2_X1 U7089 ( .A1(n5918), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5589) );
  NAND2_X1 U7090 ( .A1(n5607), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U7091 ( .A1(n5649), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5587) );
  NAND4_X1 U7092 ( .A1(n5590), .A2(n5589), .A3(n5588), .A4(n5587), .ZN(n6756)
         );
  NAND2_X1 U7093 ( .A1(n6756), .A2(n5643), .ZN(n6754) );
  NAND2_X1 U7094 ( .A1(n7794), .A2(SI_0_), .ZN(n5591) );
  XNOR2_X1 U7095 ( .A(n5591), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8770) );
  MUX2_X1 U7096 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8770), .S(n5592), .Z(n7096) );
  MUX2_X1 U7097 ( .A(n5968), .B(n6754), .S(n7096), .Z(n6748) );
  NAND2_X1 U7098 ( .A1(n5918), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5597) );
  NAND2_X1 U7099 ( .A1(n5607), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5596) );
  NAND2_X1 U7100 ( .A1(n5649), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U7101 ( .A1(n5603), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5594) );
  NAND4_X1 U7102 ( .A1(n5597), .A2(n5596), .A3(n5595), .A4(n5594), .ZN(n8323)
         );
  INV_X1 U7103 ( .A(n8323), .ZN(n6750) );
  OR2_X1 U7104 ( .A1(n6750), .A2(n4266), .ZN(n5602) );
  OR2_X1 U7105 ( .A1(n5598), .A2(n6000), .ZN(n5599) );
  XNOR2_X1 U7106 ( .A(n5599), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9667) );
  INV_X1 U7107 ( .A(n9667), .ZN(n6438) );
  OR2_X1 U7108 ( .A1(n5610), .A2(n6217), .ZN(n5601) );
  INV_X1 U7109 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6493) );
  NAND2_X1 U7110 ( .A1(n5649), .A2(n6493), .ZN(n5606) );
  NAND2_X1 U7111 ( .A1(n5918), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5605) );
  NAND2_X1 U7112 ( .A1(n4265), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5604) );
  INV_X1 U7113 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5608) );
  NAND2_X1 U7114 ( .A1(n8322), .A2(n5643), .ZN(n5616) );
  OR2_X1 U7115 ( .A1(n5610), .A2(n6215), .ZN(n5614) );
  OR2_X1 U7116 ( .A1(n7798), .A2(n6198), .ZN(n5613) );
  NAND2_X1 U7117 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4297), .ZN(n5611) );
  XNOR2_X1 U7118 ( .A(n5611), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6452) );
  INV_X1 U7119 ( .A(n6452), .ZN(n6500) );
  OR2_X1 U7120 ( .A1(n5592), .A2(n6500), .ZN(n5612) );
  XNOR2_X1 U7121 ( .A(n7247), .B(n5615), .ZN(n5617) );
  XNOR2_X1 U7122 ( .A(n5616), .B(n5617), .ZN(n6729) );
  INV_X1 U7123 ( .A(n5616), .ZN(n5618) );
  NAND2_X1 U7124 ( .A1(n5618), .A2(n5617), .ZN(n5619) );
  NAND2_X1 U7125 ( .A1(n5603), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5624) );
  NAND2_X1 U7126 ( .A1(n5918), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5623) );
  INV_X1 U7127 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6434) );
  NAND2_X1 U7128 ( .A1(n6493), .A2(n6434), .ZN(n5621) );
  NAND2_X1 U7129 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5637) );
  AND2_X1 U7130 ( .A1(n5621), .A2(n5637), .ZN(n9983) );
  NAND2_X1 U7131 ( .A1(n5649), .A2(n9983), .ZN(n5622) );
  OR2_X1 U7132 ( .A1(n6807), .A2(n4266), .ZN(n5631) );
  NOR2_X1 U7133 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5625) );
  NAND2_X1 U7134 ( .A1(n5598), .A2(n5625), .ZN(n5627) );
  NAND2_X1 U7135 ( .A1(n5627), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5626) );
  MUX2_X1 U7136 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5626), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5628) );
  OR2_X1 U7137 ( .A1(n5627), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5644) );
  NAND2_X1 U7138 ( .A1(n5628), .A2(n5644), .ZN(n6465) );
  OR2_X1 U7139 ( .A1(n7798), .A2(n6200), .ZN(n5629) );
  XNOR2_X1 U7140 ( .A(n5615), .B(n9984), .ZN(n5630) );
  NAND2_X1 U7141 ( .A1(n5631), .A2(n5630), .ZN(n5633) );
  OAI21_X1 U7142 ( .B1(n5631), .B2(n5630), .A(n5633), .ZN(n6796) );
  INV_X1 U7143 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5634) );
  NAND2_X1 U7144 ( .A1(n5603), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5641) );
  INV_X1 U7145 ( .A(n5637), .ZN(n5635) );
  NAND2_X1 U7146 ( .A1(n5635), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5652) );
  INV_X1 U7147 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5636) );
  NAND2_X1 U7148 ( .A1(n5637), .A2(n5636), .ZN(n5638) );
  AND2_X1 U7149 ( .A1(n5652), .A2(n5638), .ZN(n6806) );
  NAND2_X1 U7150 ( .A1(n5649), .A2(n6806), .ZN(n5640) );
  NAND2_X1 U7151 ( .A1(n5918), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5639) );
  OR2_X1 U7152 ( .A1(n6798), .A2(n4266), .ZN(n5668) );
  NAND2_X1 U7153 ( .A1(n5644), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5645) );
  XNOR2_X1 U7154 ( .A(n5645), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6480) );
  INV_X1 U7155 ( .A(n6480), .ZN(n6470) );
  INV_X1 U7156 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6202) );
  OR2_X1 U7157 ( .A1(n7798), .A2(n6202), .ZN(n5647) );
  XNOR2_X1 U7158 ( .A(n5615), .B(n7079), .ZN(n5669) );
  XNOR2_X1 U7159 ( .A(n5668), .B(n5669), .ZN(n6951) );
  NAND2_X1 U7160 ( .A1(n4265), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5657) );
  NAND2_X1 U7161 ( .A1(n6266), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5656) );
  INV_X1 U7162 ( .A(n5652), .ZN(n5650) );
  NAND2_X1 U7163 ( .A1(n5650), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5676) );
  INV_X1 U7164 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5651) );
  NAND2_X1 U7165 ( .A1(n5652), .A2(n5651), .ZN(n5653) );
  AND2_X1 U7166 ( .A1(n5676), .A2(n5653), .ZN(n8597) );
  NAND2_X1 U7167 ( .A1(n6038), .A2(n8597), .ZN(n5655) );
  NAND2_X1 U7168 ( .A1(n5918), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5654) );
  NOR2_X1 U7169 ( .A1(n6871), .A2(n4266), .ZN(n5666) );
  INV_X1 U7170 ( .A(n5666), .ZN(n5663) );
  NAND2_X1 U7171 ( .A1(n5658), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5659) );
  XNOR2_X1 U7172 ( .A(n5659), .B(n6389), .ZN(n6512) );
  OR2_X1 U7173 ( .A1(n5610), .A2(n6213), .ZN(n5661) );
  OR2_X1 U7174 ( .A1(n7798), .A2(n6201), .ZN(n5660) );
  XNOR2_X1 U7175 ( .A(n10048), .B(n5968), .ZN(n5665) );
  INV_X1 U7176 ( .A(n5665), .ZN(n5662) );
  NAND2_X1 U7177 ( .A1(n5663), .A2(n5662), .ZN(n5673) );
  INV_X1 U7178 ( .A(n5673), .ZN(n5664) );
  NAND2_X1 U7179 ( .A1(n5666), .A2(n5665), .ZN(n5667) );
  AND2_X1 U7180 ( .A1(n5667), .A2(n5673), .ZN(n6958) );
  INV_X1 U7181 ( .A(n6958), .ZN(n5672) );
  INV_X1 U7182 ( .A(n5668), .ZN(n5671) );
  INV_X1 U7183 ( .A(n5669), .ZN(n5670) );
  AND2_X1 U7184 ( .A1(n5671), .A2(n5670), .ZN(n6953) );
  OR2_X1 U7185 ( .A1(n5672), .A2(n6953), .ZN(n6954) );
  AND2_X1 U7186 ( .A1(n5673), .A2(n6954), .ZN(n5674) );
  NAND2_X1 U7187 ( .A1(n6266), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5681) );
  NAND2_X1 U7188 ( .A1(n4265), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5680) );
  NAND2_X1 U7189 ( .A1(n5676), .A2(n5675), .ZN(n5677) );
  AND2_X1 U7190 ( .A1(n5696), .A2(n5677), .ZN(n9974) );
  NAND2_X1 U7191 ( .A1(n6038), .A2(n9974), .ZN(n5679) );
  NAND2_X1 U7192 ( .A1(n6267), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5678) );
  OR2_X1 U7193 ( .A1(n6970), .A2(n4266), .ZN(n5685) );
  OR2_X1 U7194 ( .A1(n5658), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5687) );
  NAND2_X1 U7195 ( .A1(n5687), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5682) );
  XNOR2_X1 U7196 ( .A(n5682), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6538) );
  INV_X1 U7197 ( .A(n6538), .ZN(n6487) );
  INV_X2 U7198 ( .A(n5610), .ZN(n5706) );
  NAND2_X1 U7199 ( .A1(n6207), .A2(n5706), .ZN(n5684) );
  INV_X1 U7200 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6211) );
  OR2_X1 U7201 ( .A1(n7798), .A2(n6211), .ZN(n5683) );
  OAI211_X1 U7202 ( .C1(n5592), .C2(n6487), .A(n5684), .B(n5683), .ZN(n9975)
         );
  XNOR2_X1 U7203 ( .A(n9975), .B(n5615), .ZN(n5686) );
  XNOR2_X1 U7204 ( .A(n5685), .B(n5686), .ZN(n6870) );
  NAND2_X1 U7205 ( .A1(n6227), .A2(n5706), .ZN(n5694) );
  NOR2_X1 U7206 ( .A1(n5687), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5690) );
  NOR2_X1 U7207 ( .A1(n5690), .A2(n6000), .ZN(n5688) );
  MUX2_X1 U7208 ( .A(n6000), .B(n5688), .S(P2_IR_REG_8__SCAN_IN), .Z(n5692) );
  NAND2_X1 U7209 ( .A1(n5690), .A2(n5689), .ZN(n5707) );
  INV_X1 U7210 ( .A(n5707), .ZN(n5691) );
  NOR2_X1 U7211 ( .A1(n5692), .A2(n5691), .ZN(n6738) );
  AOI22_X1 U7212 ( .A1(n5862), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n4454), .B2(
        n6738), .ZN(n5693) );
  XNOR2_X1 U7213 ( .A(n7176), .B(n5968), .ZN(n5703) );
  INV_X1 U7214 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5695) );
  NAND2_X1 U7215 ( .A1(n5696), .A2(n5695), .ZN(n5697) );
  NAND2_X1 U7216 ( .A1(n5712), .A2(n5697), .ZN(n7171) );
  INV_X1 U7217 ( .A(n7171), .ZN(n6973) );
  NAND2_X1 U7218 ( .A1(n6038), .A2(n6973), .ZN(n5701) );
  NAND2_X1 U7219 ( .A1(n4265), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5700) );
  NAND2_X1 U7220 ( .A1(n5918), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5699) );
  INV_X2 U7221 ( .A(n5989), .ZN(n6266) );
  NAND2_X1 U7222 ( .A1(n6266), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5698) );
  OR2_X1 U7223 ( .A1(n7129), .A2(n4266), .ZN(n5702) );
  XNOR2_X1 U7224 ( .A(n5703), .B(n5702), .ZN(n6967) );
  INV_X1 U7225 ( .A(n5702), .ZN(n5704) );
  NAND2_X1 U7226 ( .A1(n5704), .A2(n5703), .ZN(n5705) );
  NAND2_X1 U7227 ( .A1(n6204), .A2(n5706), .ZN(n5710) );
  NAND2_X1 U7228 ( .A1(n5707), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5708) );
  XNOR2_X1 U7229 ( .A(n5708), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6914) );
  AOI22_X1 U7230 ( .A1(n5862), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n4454), .B2(
        n6914), .ZN(n5709) );
  XNOR2_X1 U7231 ( .A(n10070), .B(n5615), .ZN(n5718) );
  NAND2_X1 U7232 ( .A1(n4265), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5717) );
  NAND2_X1 U7233 ( .A1(n6267), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5716) );
  INV_X1 U7234 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5711) );
  NAND2_X1 U7235 ( .A1(n5712), .A2(n5711), .ZN(n5713) );
  AND2_X1 U7236 ( .A1(n5730), .A2(n5713), .ZN(n9959) );
  NAND2_X1 U7237 ( .A1(n6038), .A2(n9959), .ZN(n5715) );
  NAND2_X1 U7238 ( .A1(n6266), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5714) );
  OR2_X1 U7239 ( .A1(n6969), .A2(n4266), .ZN(n5719) );
  NAND2_X1 U7240 ( .A1(n5718), .A2(n5719), .ZN(n5724) );
  INV_X1 U7241 ( .A(n5718), .ZN(n5721) );
  INV_X1 U7242 ( .A(n5719), .ZN(n5720) );
  NAND2_X1 U7243 ( .A1(n5721), .A2(n5720), .ZN(n5722) );
  NAND2_X1 U7244 ( .A1(n5724), .A2(n5722), .ZN(n7127) );
  NAND2_X1 U7245 ( .A1(n6234), .A2(n5706), .ZN(n5728) );
  NAND2_X1 U7246 ( .A1(n5725), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5726) );
  XNOR2_X1 U7247 ( .A(n5726), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7009) );
  AOI22_X1 U7248 ( .A1(n5862), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n4454), .B2(
        n7009), .ZN(n5727) );
  NAND2_X1 U7249 ( .A1(n5728), .A2(n5727), .ZN(n7189) );
  XNOR2_X1 U7250 ( .A(n7189), .B(n5968), .ZN(n5737) );
  NAND2_X1 U7251 ( .A1(n4265), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5735) );
  NAND2_X1 U7252 ( .A1(n6266), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5734) );
  INV_X1 U7253 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7120) );
  NAND2_X1 U7254 ( .A1(n5730), .A2(n7120), .ZN(n5731) );
  AND2_X1 U7255 ( .A1(n5744), .A2(n5731), .ZN(n7186) );
  NAND2_X1 U7256 ( .A1(n6038), .A2(n7186), .ZN(n5733) );
  NAND2_X1 U7257 ( .A1(n6267), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5732) );
  NOR2_X1 U7258 ( .A1(n7286), .A2(n4266), .ZN(n5736) );
  XNOR2_X1 U7259 ( .A(n5737), .B(n5736), .ZN(n7118) );
  NAND2_X1 U7260 ( .A1(n5737), .A2(n5736), .ZN(n5738) );
  NAND2_X1 U7261 ( .A1(n6238), .A2(n5706), .ZN(n5742) );
  OR2_X1 U7262 ( .A1(n5739), .A2(n6000), .ZN(n5740) );
  XNOR2_X1 U7263 ( .A(n5740), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7212) );
  AOI22_X1 U7264 ( .A1(n5862), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n4454), .B2(
        n7212), .ZN(n5741) );
  NAND2_X1 U7265 ( .A1(n5742), .A2(n5741), .ZN(n7291) );
  XNOR2_X1 U7266 ( .A(n7291), .B(n5615), .ZN(n5750) );
  NAND2_X1 U7267 ( .A1(n6266), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5749) );
  NAND2_X1 U7268 ( .A1(n4265), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5748) );
  INV_X1 U7269 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5743) );
  NAND2_X1 U7270 ( .A1(n5744), .A2(n5743), .ZN(n5745) );
  AND2_X1 U7271 ( .A1(n5759), .A2(n5745), .ZN(n7301) );
  NAND2_X1 U7272 ( .A1(n6038), .A2(n7301), .ZN(n5747) );
  NAND2_X1 U7273 ( .A1(n6267), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5746) );
  NOR2_X1 U7274 ( .A1(n7393), .A2(n4266), .ZN(n5751) );
  XNOR2_X1 U7275 ( .A(n5750), .B(n5751), .ZN(n7296) );
  INV_X1 U7276 ( .A(n5750), .ZN(n5752) );
  NAND2_X1 U7277 ( .A1(n5752), .A2(n5751), .ZN(n5753) );
  NAND2_X1 U7278 ( .A1(n6242), .A2(n5706), .ZN(n5757) );
  OR2_X1 U7279 ( .A1(n5754), .A2(n6000), .ZN(n5755) );
  XNOR2_X1 U7280 ( .A(n5755), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7324) );
  AOI22_X1 U7281 ( .A1(n5862), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n4454), .B2(
        n7324), .ZN(n5756) );
  NAND2_X1 U7282 ( .A1(n5757), .A2(n5756), .ZN(n7416) );
  XNOR2_X1 U7283 ( .A(n7416), .B(n5615), .ZN(n5765) );
  NAND2_X1 U7284 ( .A1(n6266), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5764) );
  NAND2_X1 U7285 ( .A1(n4265), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5763) );
  INV_X1 U7286 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7208) );
  NAND2_X1 U7287 ( .A1(n5759), .A2(n7208), .ZN(n5760) );
  AND2_X1 U7288 ( .A1(n5772), .A2(n5760), .ZN(n7392) );
  NAND2_X1 U7289 ( .A1(n6038), .A2(n7392), .ZN(n5762) );
  NAND2_X1 U7290 ( .A1(n5918), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5761) );
  OR2_X1 U7291 ( .A1(n7520), .A2(n4266), .ZN(n5766) );
  NAND2_X1 U7292 ( .A1(n5765), .A2(n5766), .ZN(n7388) );
  INV_X1 U7293 ( .A(n5765), .ZN(n5768) );
  INV_X1 U7294 ( .A(n5766), .ZN(n5767) );
  NAND2_X1 U7295 ( .A1(n5768), .A2(n5767), .ZN(n7389) );
  NAND2_X1 U7296 ( .A1(n6275), .A2(n5706), .ZN(n5771) );
  OR2_X1 U7297 ( .A1(n5769), .A2(n6000), .ZN(n5783) );
  XNOR2_X1 U7298 ( .A(n5783), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7474) );
  AOI22_X1 U7299 ( .A1(n5862), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n4454), .B2(
        n7474), .ZN(n5770) );
  XNOR2_X1 U7300 ( .A(n8680), .B(n5968), .ZN(n5778) );
  NAND2_X1 U7301 ( .A1(n6266), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5777) );
  NAND2_X1 U7302 ( .A1(n4265), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5776) );
  INV_X1 U7303 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7328) );
  NAND2_X1 U7304 ( .A1(n5772), .A2(n7328), .ZN(n5773) );
  AND2_X1 U7305 ( .A1(n5787), .A2(n5773), .ZN(n7562) );
  NAND2_X1 U7306 ( .A1(n6038), .A2(n7562), .ZN(n5775) );
  NAND2_X1 U7307 ( .A1(n5918), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5774) );
  NOR2_X1 U7308 ( .A1(n7868), .A2(n4266), .ZN(n5779) );
  NAND2_X1 U7309 ( .A1(n5778), .A2(n5779), .ZN(n5793) );
  INV_X1 U7310 ( .A(n5778), .ZN(n7612) );
  INV_X1 U7311 ( .A(n5779), .ZN(n5780) );
  NAND2_X1 U7312 ( .A1(n7612), .A2(n5780), .ZN(n5781) );
  AND2_X1 U7313 ( .A1(n5793), .A2(n5781), .ZN(n7519) );
  NAND2_X1 U7314 ( .A1(n6264), .A2(n5706), .ZN(n5786) );
  INV_X1 U7315 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5782) );
  NAND2_X1 U7316 ( .A1(n5783), .A2(n5782), .ZN(n5784) );
  NAND2_X1 U7317 ( .A1(n5784), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5800) );
  XNOR2_X1 U7318 ( .A(n5800), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8330) );
  AOI22_X1 U7319 ( .A1(n5862), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n4454), .B2(
        n8330), .ZN(n5785) );
  XNOR2_X1 U7320 ( .A(n7722), .B(n5615), .ZN(n5797) );
  NAND2_X1 U7321 ( .A1(n6266), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5792) );
  NAND2_X1 U7322 ( .A1(n4265), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5791) );
  INV_X1 U7323 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7477) );
  NAND2_X1 U7324 ( .A1(n5787), .A2(n7477), .ZN(n5788) );
  AND2_X1 U7325 ( .A1(n5820), .A2(n5788), .ZN(n7615) );
  NAND2_X1 U7326 ( .A1(n6038), .A2(n7615), .ZN(n5790) );
  NAND2_X1 U7327 ( .A1(n6267), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5789) );
  NOR2_X1 U7328 ( .A1(n7709), .A2(n4266), .ZN(n5795) );
  XNOR2_X1 U7329 ( .A(n5797), .B(n5795), .ZN(n7624) );
  AND2_X1 U7330 ( .A1(n7624), .A2(n5793), .ZN(n5794) );
  INV_X1 U7331 ( .A(n5795), .ZN(n5796) );
  NAND2_X1 U7332 ( .A1(n5797), .A2(n5796), .ZN(n5798) );
  NAND2_X1 U7333 ( .A1(n6405), .A2(n5706), .ZN(n5804) );
  INV_X1 U7334 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5799) );
  NAND2_X1 U7335 ( .A1(n5800), .A2(n5799), .ZN(n5801) );
  NAND2_X1 U7336 ( .A1(n5801), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5802) );
  XNOR2_X1 U7337 ( .A(n5802), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8340) );
  AOI22_X1 U7338 ( .A1(n5862), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n4454), .B2(
        n8340), .ZN(n5803) );
  XNOR2_X1 U7339 ( .A(n8291), .B(n5615), .ZN(n5809) );
  NAND2_X1 U7340 ( .A1(n6266), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5808) );
  NAND2_X1 U7341 ( .A1(n4265), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5807) );
  XNOR2_X1 U7342 ( .A(n5820), .B(P2_REG3_REG_15__SCAN_IN), .ZN(n8283) );
  NAND2_X1 U7343 ( .A1(n6038), .A2(n8283), .ZN(n5806) );
  NAND2_X1 U7344 ( .A1(n6267), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5805) );
  OR2_X1 U7345 ( .A1(n7768), .A2(n4266), .ZN(n8281) );
  NAND2_X1 U7346 ( .A1(n5810), .A2(n5809), .ZN(n8279) );
  NAND2_X1 U7347 ( .A1(n5811), .A2(n8279), .ZN(n5826) );
  NAND2_X1 U7348 ( .A1(n6574), .A2(n5706), .ZN(n5815) );
  NAND2_X1 U7349 ( .A1(n5812), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5813) );
  XNOR2_X1 U7350 ( .A(n5813), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8365) );
  AOI22_X1 U7351 ( .A1(n5862), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n4454), .B2(
        n8365), .ZN(n5814) );
  XNOR2_X1 U7352 ( .A(n8143), .B(n5968), .ZN(n5827) );
  NAND2_X1 U7353 ( .A1(n6266), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5825) );
  NAND2_X1 U7354 ( .A1(n4265), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5824) );
  AND2_X1 U7355 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_REG3_REG_15__SCAN_IN), 
        .ZN(n5816) );
  INV_X1 U7356 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5819) );
  INV_X1 U7357 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5818) );
  OAI21_X1 U7358 ( .B1(n5820), .B2(n5819), .A(n5818), .ZN(n5821) );
  AND2_X1 U7359 ( .A1(n5835), .A2(n5821), .ZN(n8138) );
  NAND2_X1 U7360 ( .A1(n6038), .A2(n8138), .ZN(n5823) );
  NAND2_X1 U7361 ( .A1(n6267), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5822) );
  NAND4_X1 U7362 ( .A1(n5825), .A2(n5824), .A3(n5823), .A4(n5822), .ZN(n8309)
         );
  NAND2_X1 U7363 ( .A1(n8309), .A2(n5643), .ZN(n5828) );
  XNOR2_X1 U7364 ( .A(n5827), .B(n5828), .ZN(n8144) );
  INV_X1 U7365 ( .A(n5827), .ZN(n5829) );
  NAND2_X1 U7366 ( .A1(n5829), .A2(n5828), .ZN(n5830) );
  NAND2_X1 U7367 ( .A1(n6656), .A2(n5706), .ZN(n5834) );
  INV_X1 U7368 ( .A(n5847), .ZN(n5831) );
  NAND2_X1 U7369 ( .A1(n5831), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5832) );
  XNOR2_X1 U7370 ( .A(n5832), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8381) );
  AOI22_X1 U7371 ( .A1(n5862), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n4454), .B2(
        n8381), .ZN(n5833) );
  XNOR2_X1 U7372 ( .A(n8747), .B(n5968), .ZN(n5841) );
  NAND2_X1 U7373 ( .A1(n6266), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5840) );
  NAND2_X1 U7374 ( .A1(n4265), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5839) );
  INV_X1 U7375 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8363) );
  NAND2_X1 U7376 ( .A1(n5835), .A2(n8363), .ZN(n5836) );
  AND2_X1 U7377 ( .A1(n5852), .A2(n5836), .ZN(n8218) );
  NAND2_X1 U7378 ( .A1(n6038), .A2(n8218), .ZN(n5838) );
  NAND2_X1 U7379 ( .A1(n6267), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5837) );
  NOR2_X1 U7380 ( .A1(n8268), .A2(n4266), .ZN(n5842) );
  NAND2_X1 U7381 ( .A1(n5841), .A2(n5842), .ZN(n5846) );
  INV_X1 U7382 ( .A(n5841), .ZN(n8263) );
  INV_X1 U7383 ( .A(n5842), .ZN(n5843) );
  NAND2_X1 U7384 ( .A1(n8263), .A2(n5843), .ZN(n5844) );
  NAND2_X1 U7385 ( .A1(n5846), .A2(n5844), .ZN(n8212) );
  NAND2_X1 U7386 ( .A1(n6814), .A2(n5706), .ZN(n5850) );
  NAND2_X1 U7387 ( .A1(n4362), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5848) );
  XNOR2_X1 U7388 ( .A(n5848), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8387) );
  AOI22_X1 U7389 ( .A1(n5862), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n4454), .B2(
        n8387), .ZN(n5849) );
  XNOR2_X1 U7390 ( .A(n8742), .B(n5968), .ZN(n5858) );
  NAND2_X1 U7391 ( .A1(n6266), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5857) );
  NAND2_X1 U7392 ( .A1(n4265), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5856) );
  INV_X1 U7393 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5851) );
  NAND2_X1 U7394 ( .A1(n5852), .A2(n5851), .ZN(n5853) );
  AND2_X1 U7395 ( .A1(n5866), .A2(n5853), .ZN(n8585) );
  NAND2_X1 U7396 ( .A1(n6038), .A2(n8585), .ZN(n5855) );
  NAND2_X1 U7397 ( .A1(n6267), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5854) );
  NAND4_X1 U7398 ( .A1(n5857), .A2(n5856), .A3(n5855), .A4(n5854), .ZN(n8307)
         );
  AND2_X1 U7399 ( .A1(n8307), .A2(n5643), .ZN(n5859) );
  NAND2_X1 U7400 ( .A1(n5858), .A2(n5859), .ZN(n5872) );
  INV_X1 U7401 ( .A(n5858), .ZN(n8176) );
  INV_X1 U7402 ( .A(n5859), .ZN(n5860) );
  NAND2_X1 U7403 ( .A1(n8176), .A2(n5860), .ZN(n5861) );
  NAND2_X1 U7404 ( .A1(n6890), .A2(n5706), .ZN(n5864) );
  AOI22_X1 U7405 ( .A1(n5862), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8480), .B2(
        n4454), .ZN(n5863) );
  XNOR2_X1 U7406 ( .A(n8737), .B(n5968), .ZN(n5874) );
  NAND2_X1 U7407 ( .A1(n6266), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5871) );
  NAND2_X1 U7408 ( .A1(n4265), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5870) );
  INV_X1 U7409 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5865) );
  NAND2_X1 U7410 ( .A1(n5866), .A2(n5865), .ZN(n5867) );
  AND2_X1 U7411 ( .A1(n5880), .A2(n5867), .ZN(n8568) );
  NAND2_X1 U7412 ( .A1(n6038), .A2(n8568), .ZN(n5869) );
  NAND2_X1 U7413 ( .A1(n6267), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5868) );
  NAND4_X1 U7414 ( .A1(n5871), .A2(n5870), .A3(n5869), .A4(n5868), .ZN(n8306)
         );
  NAND2_X1 U7415 ( .A1(n8306), .A2(n5643), .ZN(n5875) );
  XNOR2_X1 U7416 ( .A(n5874), .B(n5875), .ZN(n8187) );
  AND2_X1 U7417 ( .A1(n8187), .A2(n5872), .ZN(n5873) );
  INV_X1 U7418 ( .A(n5874), .ZN(n5876) );
  NAND2_X1 U7419 ( .A1(n5876), .A2(n5875), .ZN(n5877) );
  NAND2_X1 U7420 ( .A1(n6965), .A2(n5706), .ZN(n5879) );
  OR2_X1 U7421 ( .A1(n7798), .A2(n6980), .ZN(n5878) );
  XNOR2_X1 U7422 ( .A(n8549), .B(n5968), .ZN(n5886) );
  INV_X1 U7423 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8240) );
  NAND2_X1 U7424 ( .A1(n5880), .A2(n8240), .ZN(n5881) );
  NAND2_X1 U7425 ( .A1(n4843), .A2(n6038), .ZN(n5885) );
  NAND2_X1 U7426 ( .A1(n6266), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5884) );
  NAND2_X1 U7427 ( .A1(n4265), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5883) );
  NAND2_X1 U7428 ( .A1(n6267), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5882) );
  NOR2_X1 U7429 ( .A1(n8197), .A2(n4266), .ZN(n5887) );
  NAND2_X1 U7430 ( .A1(n5886), .A2(n5887), .ZN(n5897) );
  INV_X1 U7431 ( .A(n5886), .ZN(n8190) );
  INV_X1 U7432 ( .A(n5887), .ZN(n5888) );
  NAND2_X1 U7433 ( .A1(n8190), .A2(n5888), .ZN(n5889) );
  NAND2_X1 U7434 ( .A1(n5897), .A2(n5889), .ZN(n8236) );
  NAND2_X1 U7435 ( .A1(n7018), .A2(n5706), .ZN(n5891) );
  OR2_X1 U7436 ( .A1(n7798), .A2(n7019), .ZN(n5890) );
  XNOR2_X1 U7437 ( .A(n8728), .B(n5968), .ZN(n5900) );
  INV_X1 U7438 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5892) );
  NAND2_X1 U7439 ( .A1(n5893), .A2(n5892), .ZN(n5894) );
  NAND2_X1 U7440 ( .A1(n5916), .A2(n5894), .ZN(n8534) );
  INV_X1 U7441 ( .A(n6038), .ZN(n5985) );
  AOI22_X1 U7442 ( .A1(n6266), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n4265), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n5896) );
  NAND2_X1 U7443 ( .A1(n5918), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5895) );
  OAI211_X1 U7444 ( .C1(n8534), .C2(n5985), .A(n5896), .B(n5895), .ZN(n8304)
         );
  NAND2_X1 U7445 ( .A1(n8304), .A2(n5643), .ZN(n5898) );
  XOR2_X1 U7446 ( .A(n5900), .B(n5898), .Z(n8189) );
  INV_X1 U7447 ( .A(n5898), .ZN(n5899) );
  NAND2_X1 U7448 ( .A1(n5900), .A2(n5899), .ZN(n5901) );
  NAND2_X1 U7449 ( .A1(n7777), .A2(n5706), .ZN(n5904) );
  OR2_X1 U7450 ( .A1(n7798), .A2(n8135), .ZN(n5903) );
  XNOR2_X1 U7451 ( .A(n8647), .B(n5615), .ZN(n5908) );
  XNOR2_X1 U7452 ( .A(n5916), .B(P2_REG3_REG_22__SCAN_IN), .ZN(n8521) );
  INV_X1 U7453 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8648) );
  NAND2_X1 U7454 ( .A1(n6267), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5906) );
  NAND2_X1 U7455 ( .A1(n4265), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5905) );
  OAI211_X1 U7456 ( .C1(n5989), .C2(n8648), .A(n5906), .B(n5905), .ZN(n5907)
         );
  AOI21_X1 U7457 ( .B1(n8521), .B2(n6038), .A(n5907), .ZN(n8196) );
  OR2_X1 U7458 ( .A1(n8196), .A2(n4266), .ZN(n8245) );
  INV_X1 U7459 ( .A(n5908), .ZN(n5909) );
  NOR2_X1 U7460 ( .A1(n5910), .A2(n5909), .ZN(n5911) );
  NAND2_X1 U7461 ( .A1(n7279), .A2(n5706), .ZN(n5913) );
  OR2_X1 U7462 ( .A1(n7798), .A2(n7278), .ZN(n5912) );
  XNOR2_X1 U7463 ( .A(n8715), .B(n5968), .ZN(n5934) );
  INV_X1 U7464 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8254) );
  INV_X1 U7465 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n5915) );
  OAI21_X1 U7466 ( .B1(n5916), .B2(n8254), .A(n5915), .ZN(n5917) );
  AND2_X1 U7467 ( .A1(n5917), .A2(n5925), .ZN(n8507) );
  NAND2_X1 U7468 ( .A1(n8507), .A2(n6038), .ZN(n5921) );
  AOI22_X1 U7469 ( .A1(n6266), .A2(P2_REG1_REG_23__SCAN_IN), .B1(n4265), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n5920) );
  NAND2_X1 U7470 ( .A1(n5918), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5919) );
  NOR2_X1 U7471 ( .A1(n8250), .A2(n4266), .ZN(n8168) );
  NAND2_X1 U7472 ( .A1(n7385), .A2(n5706), .ZN(n5923) );
  OR2_X1 U7473 ( .A1(n7798), .A2(n7401), .ZN(n5922) );
  XNOR2_X1 U7474 ( .A(n8636), .B(n5968), .ZN(n5936) );
  INV_X1 U7475 ( .A(n5925), .ZN(n5924) );
  NAND2_X1 U7476 ( .A1(n5924), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5942) );
  INV_X1 U7477 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8232) );
  NAND2_X1 U7478 ( .A1(n5925), .A2(n8232), .ZN(n5926) );
  NAND2_X1 U7479 ( .A1(n5942), .A2(n5926), .ZN(n8230) );
  OR2_X1 U7480 ( .A1(n8230), .A2(n5985), .ZN(n5932) );
  INV_X1 U7481 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8712) );
  NAND2_X1 U7482 ( .A1(n6266), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U7483 ( .A1(n4265), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5927) );
  OAI211_X1 U7484 ( .C1(n8712), .C2(n5929), .A(n5928), .B(n5927), .ZN(n5930)
         );
  INV_X1 U7485 ( .A(n5930), .ZN(n5931) );
  INV_X1 U7486 ( .A(n8226), .ZN(n8300) );
  NAND3_X1 U7487 ( .A1(n8169), .A2(n8168), .A3(n5933), .ZN(n5939) );
  INV_X1 U7488 ( .A(n5936), .ZN(n8224) );
  NOR2_X1 U7489 ( .A1(n8226), .A2(n4266), .ZN(n5937) );
  INV_X1 U7490 ( .A(n5937), .ZN(n8228) );
  NAND2_X1 U7491 ( .A1(n7568), .A2(n5706), .ZN(n5941) );
  OR2_X1 U7492 ( .A1(n7798), .A2(n7575), .ZN(n5940) );
  XNOR2_X1 U7493 ( .A(n8708), .B(n5615), .ZN(n8159) );
  INV_X1 U7494 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8207) );
  NAND2_X1 U7495 ( .A1(n5942), .A2(n8207), .ZN(n5943) );
  AND2_X1 U7496 ( .A1(n5954), .A2(n5943), .ZN(n8477) );
  NAND2_X1 U7497 ( .A1(n8477), .A2(n6038), .ZN(n5948) );
  INV_X1 U7498 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n6346) );
  NAND2_X1 U7499 ( .A1(n6267), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U7500 ( .A1(n4265), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5944) );
  OAI211_X1 U7501 ( .C1(n5989), .C2(n6346), .A(n5945), .B(n5944), .ZN(n5946)
         );
  INV_X1 U7502 ( .A(n5946), .ZN(n5947) );
  NAND2_X1 U7503 ( .A1(n8299), .A2(n5643), .ZN(n5949) );
  NOR2_X1 U7504 ( .A1(n8159), .A2(n5949), .ZN(n5950) );
  AOI21_X1 U7505 ( .B1(n8159), .B2(n5949), .A(n5950), .ZN(n8204) );
  NAND2_X1 U7506 ( .A1(n7607), .A2(n5706), .ZN(n5952) );
  OR2_X1 U7507 ( .A1(n7798), .A2(n7649), .ZN(n5951) );
  XNOR2_X1 U7508 ( .A(n8626), .B(n5968), .ZN(n6138) );
  INV_X1 U7509 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n5953) );
  NAND2_X1 U7510 ( .A1(n5954), .A2(n5953), .ZN(n5955) );
  NAND2_X1 U7511 ( .A1(n5983), .A2(n5955), .ZN(n8464) );
  OR2_X1 U7512 ( .A1(n8464), .A2(n5985), .ZN(n5960) );
  INV_X1 U7513 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8703) );
  NAND2_X1 U7514 ( .A1(n6266), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5957) );
  NAND2_X1 U7515 ( .A1(n4265), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5956) );
  OAI211_X1 U7516 ( .C1(n8703), .C2(n5929), .A(n5957), .B(n5956), .ZN(n5958)
         );
  INV_X1 U7517 ( .A(n5958), .ZN(n5959) );
  NOR2_X1 U7518 ( .A1(n6082), .A2(n4266), .ZN(n5961) );
  NAND2_X1 U7519 ( .A1(n6138), .A2(n5961), .ZN(n5965) );
  INV_X1 U7520 ( .A(n6138), .ZN(n5963) );
  INV_X1 U7521 ( .A(n5961), .ZN(n5962) );
  NAND2_X1 U7522 ( .A1(n5963), .A2(n5962), .ZN(n5964) );
  NAND2_X1 U7523 ( .A1(n5965), .A2(n5964), .ZN(n8157) );
  OR2_X1 U7524 ( .A1(n7798), .A2(n7730), .ZN(n5966) );
  XNOR2_X1 U7525 ( .A(n8699), .B(n5968), .ZN(n5972) );
  XNOR2_X1 U7526 ( .A(n5983), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8447) );
  INV_X1 U7527 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n6348) );
  NAND2_X1 U7528 ( .A1(n6266), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5970) );
  NAND2_X1 U7529 ( .A1(n4265), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5969) );
  OAI211_X1 U7530 ( .C1(n6348), .C2(n5929), .A(n5970), .B(n5969), .ZN(n5971)
         );
  NOR2_X1 U7531 ( .A1(n8162), .A2(n4266), .ZN(n5973) );
  NAND2_X1 U7532 ( .A1(n5972), .A2(n5973), .ZN(n5977) );
  INV_X1 U7533 ( .A(n5972), .ZN(n5975) );
  INV_X1 U7534 ( .A(n5973), .ZN(n5974) );
  NAND2_X1 U7535 ( .A1(n5975), .A2(n5974), .ZN(n5976) );
  NAND2_X1 U7536 ( .A1(n6141), .A2(n5977), .ZN(n6023) );
  OR2_X1 U7537 ( .A1(n7798), .A2(n7742), .ZN(n5978) );
  INV_X1 U7538 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5981) );
  INV_X1 U7539 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5980) );
  OAI21_X1 U7540 ( .B1(n5983), .B2(n5981), .A(n5980), .ZN(n5984) );
  NAND2_X1 U7541 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n5982) );
  NAND2_X1 U7542 ( .A1(n5984), .A2(n6131), .ZN(n6044) );
  INV_X1 U7543 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8617) );
  NAND2_X1 U7544 ( .A1(n6267), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5988) );
  NAND2_X1 U7545 ( .A1(n4265), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5987) );
  OAI211_X1 U7546 ( .C1(n5989), .C2(n8617), .A(n5988), .B(n5987), .ZN(n5990)
         );
  INV_X1 U7547 ( .A(n5990), .ZN(n5991) );
  NAND2_X1 U7548 ( .A1(n8296), .A2(n5643), .ZN(n5993) );
  XNOR2_X1 U7549 ( .A(n5993), .B(n5615), .ZN(n6018) );
  INV_X1 U7550 ( .A(n6018), .ZN(n6019) );
  NAND2_X1 U7551 ( .A1(n5995), .A2(n5994), .ZN(n5996) );
  NAND2_X1 U7552 ( .A1(n5996), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6026) );
  NAND2_X1 U7553 ( .A1(n6026), .A2(n6025), .ZN(n6028) );
  NAND2_X1 U7554 ( .A1(n6028), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5997) );
  NAND2_X1 U7555 ( .A1(n5998), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5999) );
  XNOR2_X1 U7556 ( .A(n5999), .B(P2_IR_REG_26__SCAN_IN), .ZN(n7648) );
  OR2_X1 U7557 ( .A1(n7400), .A2(n7648), .ZN(n10019) );
  OR2_X1 U7558 ( .A1(n6001), .A2(n6000), .ZN(n6002) );
  XNOR2_X1 U7559 ( .A(n6002), .B(P2_IR_REG_25__SCAN_IN), .ZN(n7572) );
  XNOR2_X1 U7560 ( .A(n7400), .B(P2_B_REG_SCAN_IN), .ZN(n6003) );
  INV_X1 U7561 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6005) );
  NAND2_X1 U7562 ( .A1(n10012), .A2(n6005), .ZN(n6006) );
  NAND2_X1 U7563 ( .A1(n10019), .A2(n6006), .ZN(n6832) );
  INV_X1 U7564 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10024) );
  NOR2_X1 U7565 ( .A1(n7572), .A2(n7648), .ZN(n10026) );
  AOI21_X1 U7566 ( .B1(n10012), .B2(n10024), .A(n10026), .ZN(n6770) );
  NOR4_X1 U7567 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n6010) );
  NOR4_X1 U7568 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n6009) );
  NOR4_X1 U7569 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n6008) );
  NOR4_X1 U7570 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6007) );
  NAND4_X1 U7571 ( .A1(n6010), .A2(n6009), .A3(n6008), .A4(n6007), .ZN(n6015)
         );
  NOR2_X1 U7572 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .ZN(
        n6387) );
  NOR4_X1 U7573 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6013) );
  NOR4_X1 U7574 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n6012) );
  NOR4_X1 U7575 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n6011) );
  NAND4_X1 U7576 ( .A1(n6387), .A2(n6013), .A3(n6012), .A4(n6011), .ZN(n6014)
         );
  OAI21_X1 U7577 ( .B1(n6015), .B2(n6014), .A(n10012), .ZN(n6836) );
  NAND2_X1 U7578 ( .A1(n6770), .A2(n6836), .ZN(n6086) );
  OR2_X1 U7579 ( .A1(n10027), .A2(n7947), .ZN(n6129) );
  NOR2_X1 U7580 ( .A1(n10086), .A2(n8405), .ZN(n6767) );
  INV_X1 U7581 ( .A(n6767), .ZN(n6831) );
  OAI21_X1 U7582 ( .B1(n6045), .B2(n6129), .A(n6831), .ZN(n6030) );
  NOR3_X1 U7583 ( .A1(n4481), .A2(n6030), .A3(n6019), .ZN(n6016) );
  AOI21_X1 U7584 ( .B1(n4481), .B2(n6019), .A(n6016), .ZN(n6017) );
  NOR3_X1 U7585 ( .A1(n4481), .A2(n6018), .A3(n6030), .ZN(n6021) );
  NOR2_X1 U7586 ( .A1(n8616), .A2(n6019), .ZN(n6020) );
  AND2_X1 U7587 ( .A1(n7648), .A2(n7572), .ZN(n6024) );
  NAND2_X1 U7588 ( .A1(n7400), .A2(n6024), .ZN(n6429) );
  OR2_X1 U7589 ( .A1(n6026), .A2(n6025), .ZN(n6027) );
  NAND2_X1 U7590 ( .A1(n6028), .A2(n6027), .ZN(n6259) );
  AND2_X1 U7591 ( .A1(n6259), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6029) );
  NAND2_X1 U7592 ( .A1(n6030), .A2(n10013), .ZN(n8278) );
  INV_X1 U7593 ( .A(n6045), .ZN(n6031) );
  NAND2_X1 U7594 ( .A1(n6031), .A2(n10013), .ZN(n6043) );
  NAND2_X1 U7595 ( .A1(n7991), .A2(n7980), .ZN(n6428) );
  INV_X1 U7596 ( .A(n6428), .ZN(n6257) );
  OR2_X1 U7597 ( .A1(n10027), .A2(n8405), .ZN(n6032) );
  NAND2_X1 U7598 ( .A1(n6129), .A2(n6032), .ZN(n10069) );
  OAI21_X1 U7599 ( .B1(n4481), .B2(n8278), .A(n8259), .ZN(n6033) );
  OR2_X1 U7600 ( .A1(n6428), .A2(n6034), .ZN(n8267) );
  OR2_X1 U7601 ( .A1(n8162), .A2(n8267), .ZN(n6041) );
  INV_X1 U7602 ( .A(n6131), .ZN(n6039) );
  INV_X1 U7603 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n6130) );
  NAND2_X1 U7604 ( .A1(n6267), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6036) );
  NAND2_X1 U7605 ( .A1(n6266), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6035) );
  OAI211_X1 U7606 ( .C1(n5648), .C2(n6130), .A(n6036), .B(n6035), .ZN(n6037)
         );
  AOI21_X1 U7607 ( .B1(n6039), .B2(n6038), .A(n6037), .ZN(n6782) );
  INV_X1 U7608 ( .A(n6034), .ZN(n6454) );
  OR2_X1 U7609 ( .A1(n6782), .A2(n8249), .ZN(n6040) );
  AND2_X1 U7610 ( .A1(n6041), .A2(n6040), .ZN(n8429) );
  AND2_X1 U7611 ( .A1(n7947), .A2(n8405), .ZN(n7988) );
  INV_X1 U7612 ( .A(n7988), .ZN(n6042) );
  INV_X1 U7613 ( .A(n6044), .ZN(n8432) );
  NAND2_X1 U7614 ( .A1(n6045), .A2(n6831), .ZN(n6047) );
  OR2_X1 U7615 ( .A1(n6428), .A2(n7988), .ZN(n6085) );
  AND3_X1 U7616 ( .A1(n6429), .A2(n6259), .A3(n6085), .ZN(n6046) );
  NAND2_X1 U7617 ( .A1(n6047), .A2(n6046), .ZN(n6725) );
  AOI22_X1 U7618 ( .A1(n8432), .A2(n8275), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        n4262), .ZN(n6048) );
  OAI21_X1 U7619 ( .B1(n8429), .B2(n8273), .A(n6048), .ZN(n6049) );
  INV_X1 U7620 ( .A(n6049), .ZN(n6050) );
  INV_X1 U7621 ( .A(n8250), .ZN(n8301) );
  INV_X1 U7622 ( .A(n8737), .ZN(n8567) );
  INV_X1 U7623 ( .A(n8306), .ZN(n6111) );
  NAND2_X1 U7624 ( .A1(n6756), .A2(n7096), .ZN(n7100) );
  NAND2_X1 U7625 ( .A1(n7092), .A2(n7100), .ZN(n7099) );
  NAND2_X1 U7626 ( .A1(n6051), .A2(n6052), .ZN(n6053) );
  NAND2_X1 U7627 ( .A1(n7099), .A2(n6053), .ZN(n6762) );
  NAND2_X1 U7628 ( .A1(n6750), .A2(n9991), .ZN(n7821) );
  INV_X1 U7629 ( .A(n9991), .ZN(n6886) );
  NAND2_X1 U7630 ( .A1(n6886), .A2(n8323), .ZN(n7819) );
  NAND2_X1 U7631 ( .A1(n6762), .A2(n7948), .ZN(n6761) );
  NAND2_X1 U7632 ( .A1(n6750), .A2(n6886), .ZN(n6054) );
  NAND2_X1 U7633 ( .A1(n6761), .A2(n6054), .ZN(n6774) );
  XNOR2_X2 U7634 ( .A(n7832), .B(n7831), .ZN(n7954) );
  NAND2_X1 U7635 ( .A1(n7832), .A2(n7247), .ZN(n6055) );
  NAND2_X1 U7636 ( .A1(n6773), .A2(n6055), .ZN(n6859) );
  NAND2_X1 U7637 ( .A1(n8321), .A2(n6881), .ZN(n7068) );
  NAND2_X1 U7638 ( .A1(n6807), .A2(n9984), .ZN(n7806) );
  NAND2_X1 U7639 ( .A1(n6859), .A2(n6097), .ZN(n6858) );
  NAND2_X1 U7640 ( .A1(n6807), .A2(n6881), .ZN(n6056) );
  NAND2_X1 U7641 ( .A1(n6858), .A2(n6056), .ZN(n7080) );
  NAND2_X1 U7642 ( .A1(n6798), .A2(n7079), .ZN(n7811) );
  INV_X1 U7643 ( .A(n6798), .ZN(n8320) );
  NAND2_X1 U7644 ( .A1(n7811), .A2(n7828), .ZN(n7953) );
  NAND2_X1 U7645 ( .A1(n7080), .A2(n7953), .ZN(n6058) );
  NAND2_X1 U7646 ( .A1(n6798), .A2(n10043), .ZN(n6057) );
  NAND2_X1 U7647 ( .A1(n6058), .A2(n6057), .ZN(n8599) );
  INV_X1 U7648 ( .A(n8599), .ZN(n6060) );
  NAND2_X1 U7649 ( .A1(n6871), .A2(n10048), .ZN(n9965) );
  INV_X1 U7650 ( .A(n6871), .ZN(n8319) );
  INV_X1 U7651 ( .A(n10048), .ZN(n6964) );
  NAND2_X1 U7652 ( .A1(n8319), .A2(n6964), .ZN(n7837) );
  INV_X1 U7653 ( .A(n8600), .ZN(n6059) );
  NAND2_X1 U7654 ( .A1(n8319), .A2(n10048), .ZN(n6061) );
  NAND2_X1 U7655 ( .A1(n6970), .A2(n9975), .ZN(n7841) );
  INV_X1 U7656 ( .A(n6970), .ZN(n8318) );
  INV_X1 U7657 ( .A(n9975), .ZN(n10057) );
  NAND2_X1 U7658 ( .A1(n8318), .A2(n10057), .ZN(n7842) );
  OR2_X1 U7659 ( .A1(n6969), .A2(n10070), .ZN(n7852) );
  NAND2_X1 U7660 ( .A1(n10070), .A2(n6969), .ZN(n7847) );
  INV_X1 U7661 ( .A(n9954), .ZN(n6062) );
  INV_X1 U7662 ( .A(n7129), .ZN(n8317) );
  NAND2_X1 U7663 ( .A1(n8317), .A2(n7176), .ZN(n9949) );
  NAND2_X1 U7664 ( .A1(n6062), .A2(n9949), .ZN(n6064) );
  INV_X1 U7665 ( .A(n6969), .ZN(n8316) );
  OR2_X1 U7666 ( .A1(n8316), .A2(n10070), .ZN(n6065) );
  NAND2_X1 U7667 ( .A1(n7129), .A2(n7176), .ZN(n7845) );
  INV_X1 U7668 ( .A(n7176), .ZN(n10062) );
  NAND2_X1 U7669 ( .A1(n10062), .A2(n8317), .ZN(n7844) );
  INV_X1 U7670 ( .A(n7957), .ZN(n6103) );
  NAND2_X1 U7671 ( .A1(n6970), .A2(n10057), .ZN(n7163) );
  AND2_X1 U7672 ( .A1(n6103), .A2(n7163), .ZN(n6063) );
  AND2_X1 U7673 ( .A1(n6065), .A2(n9951), .ZN(n6066) );
  NAND2_X1 U7674 ( .A1(n7189), .A2(n7286), .ZN(n7849) );
  NAND2_X1 U7675 ( .A1(n7850), .A2(n7849), .ZN(n7959) );
  INV_X1 U7676 ( .A(n7286), .ZN(n8315) );
  NAND2_X1 U7677 ( .A1(n7189), .A2(n8315), .ZN(n6067) );
  NAND2_X1 U7678 ( .A1(n7180), .A2(n6067), .ZN(n7284) );
  OR2_X1 U7679 ( .A1(n7291), .A2(n7393), .ZN(n7851) );
  NAND2_X1 U7680 ( .A1(n7291), .A2(n7393), .ZN(n7859) );
  NAND2_X1 U7681 ( .A1(n7851), .A2(n7859), .ZN(n7960) );
  NAND2_X1 U7682 ( .A1(n7284), .A2(n7960), .ZN(n7283) );
  INV_X1 U7683 ( .A(n7393), .ZN(n8314) );
  NAND2_X1 U7684 ( .A1(n7291), .A2(n8314), .ZN(n6068) );
  OR2_X1 U7685 ( .A1(n7416), .A2(n7520), .ZN(n7862) );
  NAND2_X1 U7686 ( .A1(n7416), .A2(n7520), .ZN(n7863) );
  INV_X1 U7687 ( .A(n7520), .ZN(n8313) );
  OR2_X1 U7688 ( .A1(n7416), .A2(n8313), .ZN(n6070) );
  XNOR2_X1 U7689 ( .A(n8680), .B(n7868), .ZN(n7554) );
  INV_X1 U7690 ( .A(n7868), .ZN(n8312) );
  NAND2_X1 U7691 ( .A1(n8680), .A2(n8312), .ZN(n6071) );
  OR2_X1 U7692 ( .A1(n7722), .A2(n7709), .ZN(n7873) );
  NAND2_X1 U7693 ( .A1(n7722), .A2(n7709), .ZN(n7872) );
  NAND2_X1 U7694 ( .A1(n7873), .A2(n7872), .ZN(n7946) );
  INV_X1 U7695 ( .A(n7709), .ZN(n8311) );
  OR2_X1 U7696 ( .A1(n7722), .A2(n8311), .ZN(n6072) );
  OR2_X1 U7697 ( .A1(n8291), .A2(n7768), .ZN(n6107) );
  NAND2_X1 U7698 ( .A1(n8291), .A2(n7768), .ZN(n7803) );
  NAND2_X1 U7699 ( .A1(n6107), .A2(n7803), .ZN(n7966) );
  INV_X1 U7700 ( .A(n7768), .ZN(n8310) );
  NOR2_X1 U7701 ( .A1(n8291), .A2(n8310), .ZN(n6073) );
  NAND2_X1 U7702 ( .A1(n8143), .A2(n8309), .ZN(n6075) );
  OR2_X1 U7703 ( .A1(n8143), .A2(n8309), .ZN(n6074) );
  INV_X1 U7704 ( .A(n6075), .ZN(n6076) );
  NOR2_X2 U7705 ( .A1(n7765), .A2(n6076), .ZN(n7748) );
  OR2_X1 U7706 ( .A1(n8747), .A2(n8268), .ZN(n6109) );
  NAND2_X1 U7707 ( .A1(n8747), .A2(n8268), .ZN(n7881) );
  NAND2_X1 U7708 ( .A1(n6109), .A2(n7881), .ZN(n7968) );
  NAND2_X1 U7709 ( .A1(n7748), .A2(n7968), .ZN(n7747) );
  INV_X1 U7710 ( .A(n8268), .ZN(n8308) );
  NAND2_X1 U7711 ( .A1(n8742), .A2(n8307), .ZN(n6078) );
  INV_X1 U7712 ( .A(n8307), .ZN(n8175) );
  INV_X1 U7713 ( .A(n8742), .ZN(n8584) );
  AOI22_X1 U7714 ( .A1(n8574), .A2(n6078), .B1(n8175), .B2(n8584), .ZN(n8557)
         );
  OAI21_X1 U7715 ( .B1(n8737), .B2(n8306), .A(n8557), .ZN(n6079) );
  NAND2_X1 U7716 ( .A1(n8549), .A2(n8197), .ZN(n7900) );
  NAND2_X1 U7717 ( .A1(n7897), .A2(n7900), .ZN(n7945) );
  INV_X1 U7718 ( .A(n8197), .ZN(n8305) );
  AOI22_X2 U7719 ( .A1(n8541), .A2(n7945), .B1(n8549), .B2(n8305), .ZN(n8527)
         );
  NAND2_X1 U7720 ( .A1(n8728), .A2(n8304), .ZN(n6080) );
  INV_X1 U7721 ( .A(n8304), .ZN(n6117) );
  INV_X1 U7722 ( .A(n8728), .ZN(n8533) );
  NAND2_X1 U7723 ( .A1(n8647), .A2(n8196), .ZN(n7890) );
  INV_X1 U7724 ( .A(n8196), .ZN(n8302) );
  OR2_X1 U7725 ( .A1(n8715), .A2(n8250), .ZN(n7906) );
  NAND2_X1 U7726 ( .A1(n8715), .A2(n8250), .ZN(n6118) );
  NAND2_X1 U7727 ( .A1(n8636), .A2(n8226), .ZN(n7905) );
  NAND2_X1 U7728 ( .A1(n7908), .A2(n7905), .ZN(n8485) );
  NAND2_X1 U7729 ( .A1(n8708), .A2(n8158), .ZN(n7912) );
  NAND2_X1 U7730 ( .A1(n8457), .A2(n7912), .ZN(n7910) );
  INV_X1 U7731 ( .A(n8708), .ZN(n8211) );
  AOI21_X2 U7732 ( .B1(n8468), .B2(n7910), .A(n6081), .ZN(n8454) );
  NAND2_X1 U7733 ( .A1(n8626), .A2(n6082), .ZN(n7916) );
  NAND2_X1 U7734 ( .A1(n8766), .A2(n5706), .ZN(n6084) );
  INV_X1 U7735 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8769) );
  OR2_X1 U7736 ( .A1(n7798), .A2(n8769), .ZN(n6083) );
  NAND2_X1 U7737 ( .A1(n8130), .A2(n6782), .ZN(n7925) );
  NAND2_X1 U7738 ( .A1(n10013), .A2(n6085), .ZN(n6834) );
  INV_X1 U7739 ( .A(n6086), .ZN(n6087) );
  NAND2_X1 U7740 ( .A1(n6832), .A2(n6087), .ZN(n6088) );
  NAND2_X1 U7741 ( .A1(n10013), .A2(n6767), .ZN(n8479) );
  OR2_X1 U7742 ( .A1(n7991), .A2(n6090), .ZN(n6089) );
  NAND3_X1 U7743 ( .A1(n6089), .A2(n6428), .A3(n8405), .ZN(n9955) );
  NAND2_X1 U7744 ( .A1(n6090), .A2(n8480), .ZN(n7166) );
  NAND2_X1 U7745 ( .A1(n9955), .A2(n7166), .ZN(n6091) );
  NAND2_X1 U7746 ( .A1(n8127), .A2(n10006), .ZN(n6137) );
  INV_X1 U7747 ( .A(n6756), .ZN(n6751) );
  NAND2_X1 U7748 ( .A1(n6751), .A2(n7096), .ZN(n7950) );
  NAND2_X1 U7749 ( .A1(n6092), .A2(n7950), .ZN(n7814) );
  NAND2_X1 U7750 ( .A1(n7814), .A2(n6093), .ZN(n6763) );
  INV_X1 U7751 ( .A(n6763), .ZN(n6095) );
  INV_X1 U7752 ( .A(n7948), .ZN(n6094) );
  NAND2_X1 U7753 ( .A1(n6095), .A2(n6094), .ZN(n6096) );
  NAND2_X1 U7754 ( .A1(n6096), .A2(n7821), .ZN(n6863) );
  INV_X1 U7755 ( .A(n6097), .ZN(n6098) );
  INV_X1 U7756 ( .A(n7247), .ZN(n7831) );
  NOR2_X1 U7757 ( .A1(n7829), .A2(n4842), .ZN(n6099) );
  AOI21_X1 U7758 ( .B1(n6863), .B2(n6100), .A(n6099), .ZN(n6101) );
  NAND2_X1 U7759 ( .A1(n6101), .A2(n7811), .ZN(n8593) );
  NAND2_X1 U7760 ( .A1(n8593), .A2(n8600), .ZN(n9966) );
  INV_X1 U7761 ( .A(n7956), .ZN(n9977) );
  INV_X1 U7762 ( .A(n9965), .ZN(n7812) );
  NOR2_X1 U7763 ( .A1(n9977), .A2(n7812), .ZN(n6102) );
  NAND2_X1 U7764 ( .A1(n9966), .A2(n6102), .ZN(n9969) );
  NAND2_X1 U7765 ( .A1(n6104), .A2(n7847), .ZN(n7181) );
  NAND2_X1 U7766 ( .A1(n4289), .A2(n7850), .ZN(n7285) );
  NAND2_X1 U7767 ( .A1(n7285), .A2(n7859), .ZN(n7404) );
  AND2_X1 U7768 ( .A1(n7862), .A2(n7851), .ZN(n7858) );
  NAND2_X1 U7769 ( .A1(n7404), .A2(n7858), .ZN(n6105) );
  NAND2_X1 U7770 ( .A1(n6105), .A2(n7863), .ZN(n7556) );
  INV_X1 U7771 ( .A(n7554), .ZN(n7962) );
  NAND2_X1 U7772 ( .A1(n8680), .A2(n7868), .ZN(n6106) );
  NAND2_X1 U7773 ( .A1(n7579), .A2(n7873), .ZN(n7708) );
  INV_X1 U7774 ( .A(n6107), .ZN(n7805) );
  INV_X1 U7775 ( .A(n7967), .ZN(n7766) );
  AND2_X1 U7776 ( .A1(n7766), .A2(n6109), .ZN(n6108) );
  INV_X1 U7777 ( .A(n6109), .ZN(n7883) );
  INV_X1 U7778 ( .A(n8309), .ZN(n7880) );
  NAND2_X1 U7779 ( .A1(n8143), .A2(n7880), .ZN(n7882) );
  INV_X1 U7780 ( .A(n7968), .ZN(n7886) );
  AND2_X1 U7781 ( .A1(n7882), .A2(n7886), .ZN(n7751) );
  OR2_X1 U7782 ( .A1(n7883), .A2(n7751), .ZN(n6110) );
  NAND2_X1 U7783 ( .A1(n8742), .A2(n8175), .ZN(n7887) );
  OR2_X1 U7784 ( .A1(n8737), .A2(n6111), .ZN(n7896) );
  NAND2_X1 U7785 ( .A1(n8737), .A2(n6111), .ZN(n8545) );
  NAND2_X1 U7786 ( .A1(n7896), .A2(n8545), .ZN(n8561) );
  AND2_X1 U7787 ( .A1(n8584), .A2(n8307), .ZN(n8558) );
  NOR2_X1 U7788 ( .A1(n8561), .A2(n8558), .ZN(n6112) );
  NAND2_X1 U7789 ( .A1(n8560), .A2(n6112), .ZN(n8543) );
  INV_X1 U7790 ( .A(n8545), .ZN(n6113) );
  NOR2_X1 U7791 ( .A1(n7945), .A2(n6113), .ZN(n6114) );
  NAND2_X1 U7792 ( .A1(n8543), .A2(n6114), .ZN(n8542) );
  NAND2_X1 U7793 ( .A1(n8542), .A2(n7897), .ZN(n8529) );
  INV_X1 U7794 ( .A(n8529), .ZN(n6116) );
  XNOR2_X1 U7795 ( .A(n8728), .B(n6117), .ZN(n8528) );
  INV_X1 U7796 ( .A(n8528), .ZN(n6115) );
  NAND2_X1 U7797 ( .A1(n8728), .A2(n6117), .ZN(n7899) );
  INV_X1 U7798 ( .A(n8506), .ZN(n8500) );
  INV_X1 U7799 ( .A(n8499), .ZN(n7892) );
  NOR2_X1 U7800 ( .A1(n8500), .A2(n7892), .ZN(n6119) );
  INV_X1 U7801 ( .A(n6118), .ZN(n7893) );
  INV_X1 U7802 ( .A(n8485), .ZN(n8489) );
  NAND2_X1 U7803 ( .A1(n8490), .A2(n8489), .ZN(n8488) );
  NAND2_X1 U7804 ( .A1(n8488), .A2(n7908), .ZN(n8470) );
  INV_X1 U7805 ( .A(n7910), .ZN(n8471) );
  INV_X1 U7806 ( .A(n8456), .ZN(n8453) );
  INV_X1 U7807 ( .A(n8457), .ZN(n6120) );
  NOR2_X1 U7808 ( .A1(n8453), .A2(n6120), .ZN(n6121) );
  OR2_X1 U7809 ( .A1(n8699), .A2(n8162), .ZN(n7921) );
  NAND2_X1 U7810 ( .A1(n8428), .A2(n8427), .ZN(n8426) );
  INV_X1 U7811 ( .A(n8296), .ZN(n7927) );
  OR2_X1 U7812 ( .A1(n8616), .A2(n7927), .ZN(n7922) );
  NAND2_X1 U7813 ( .A1(n8426), .A2(n7922), .ZN(n7779) );
  XNOR2_X1 U7814 ( .A(n7779), .B(n7974), .ZN(n6128) );
  NAND2_X1 U7815 ( .A1(n7979), .A2(n7980), .ZN(n7801) );
  NAND2_X1 U7816 ( .A1(n7983), .A2(n7801), .ZN(n9968) );
  NAND2_X1 U7817 ( .A1(n6266), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6124) );
  NAND2_X1 U7818 ( .A1(n4265), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6123) );
  NAND2_X1 U7819 ( .A1(n6267), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6122) );
  AND3_X1 U7820 ( .A1(n6124), .A2(n6123), .A3(n6122), .ZN(n7800) );
  INV_X1 U7821 ( .A(n8249), .ZN(n8269) );
  INV_X1 U7822 ( .A(n6125), .ZN(n7989) );
  NAND2_X1 U7823 ( .A1(n7989), .A2(P2_B_REG_SCAN_IN), .ZN(n6126) );
  NAND2_X1 U7824 ( .A1(n8269), .A2(n6126), .ZN(n8412) );
  OAI22_X1 U7825 ( .A1(n7927), .A2(n8267), .B1(n7800), .B2(n8412), .ZN(n6127)
         );
  OR2_X1 U7826 ( .A1(n8123), .A2(n10011), .ZN(n6136) );
  NOR2_X2 U7827 ( .A1(n10011), .A2(n6129), .ZN(n9990) );
  OAI22_X1 U7828 ( .A1(n6131), .A2(n8479), .B1(n10009), .B2(n6130), .ZN(n6134)
         );
  NAND2_X1 U7829 ( .A1(n6775), .A2(n7247), .ZN(n6861) );
  NOR2_X2 U7830 ( .A1(n8601), .A2(n10048), .ZN(n9979) );
  INV_X1 U7831 ( .A(n7189), .ZN(n10078) );
  INV_X1 U7832 ( .A(n7291), .ZN(n10085) );
  INV_X1 U7833 ( .A(n7722), .ZN(n7589) );
  INV_X1 U7834 ( .A(n8291), .ZN(n7713) );
  NAND2_X1 U7835 ( .A1(n8581), .A2(n8567), .ZN(n8566) );
  INV_X1 U7836 ( .A(n8647), .ZN(n8524) );
  INV_X1 U7837 ( .A(n8715), .ZN(n8509) );
  INV_X1 U7838 ( .A(n10086), .ZN(n10049) );
  OAI211_X1 U7839 ( .C1(n8431), .C2(n6132), .A(n10049), .B(n8419), .ZN(n8122)
         );
  OR2_X1 U7840 ( .A1(n7095), .A2(n8480), .ZN(n8588) );
  NOR2_X1 U7841 ( .A1(n8122), .A2(n8588), .ZN(n6133) );
  AOI211_X1 U7842 ( .C1(n9990), .C2(n8130), .A(n6134), .B(n6133), .ZN(n6135)
         );
  NAND2_X1 U7843 ( .A1(n6137), .A2(n4846), .ZN(P2_U3267) );
  NOR2_X1 U7844 ( .A1(n8259), .A2(n4266), .ZN(n8244) );
  NAND3_X1 U7845 ( .A1(n6138), .A2(n8244), .A3(n8298), .ZN(n6144) );
  OAI21_X1 U7846 ( .B1(n6139), .B2(n6140), .A(n8282), .ZN(n6143) );
  INV_X1 U7847 ( .A(n6141), .ZN(n6142) );
  AOI21_X1 U7848 ( .B1(n6144), .B2(n6143), .A(n6142), .ZN(n6152) );
  NAND2_X1 U7849 ( .A1(n8296), .A2(n8269), .ZN(n6146) );
  INV_X1 U7850 ( .A(n8267), .ZN(n8251) );
  NAND2_X1 U7851 ( .A1(n8298), .A2(n8251), .ZN(n6145) );
  AND2_X1 U7852 ( .A1(n6146), .A2(n6145), .ZN(n8443) );
  AOI22_X1 U7853 ( .A1(n8447), .A2(n8275), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n6147) );
  OAI21_X1 U7854 ( .B1(n8443), .B2(n8273), .A(n6147), .ZN(n6148) );
  INV_X1 U7855 ( .A(n6148), .ZN(n6149) );
  NAND2_X1 U7856 ( .A1(n6150), .A2(n6149), .ZN(n6151) );
  INV_X1 U7857 ( .A(n9630), .ZN(n6154) );
  NAND2_X1 U7858 ( .A1(n6154), .A2(n6153), .ZN(n6907) );
  NAND2_X1 U7859 ( .A1(n6156), .A2(n9929), .ZN(n6158) );
  INV_X1 U7860 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6157) );
  NAND2_X1 U7861 ( .A1(n6158), .A2(n4841), .ZN(P1_U3520) );
  NAND2_X1 U7862 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6259), .ZN(n10022) );
  INV_X1 U7863 ( .A(n7280), .ZN(n6159) );
  OR2_X1 U7864 ( .A1(n9079), .A2(n6159), .ZN(n6160) );
  NAND2_X1 U7865 ( .A1(n6420), .A2(n7280), .ZN(n6191) );
  NAND2_X1 U7866 ( .A1(n6160), .A2(n6191), .ZN(n6187) );
  OR2_X1 U7867 ( .A1(n6187), .A2(n6161), .ZN(n6162) );
  NAND2_X1 U7868 ( .A1(n6162), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  OR2_X2 U7869 ( .A1(n6191), .A2(P1_U3084), .ZN(n9261) );
  INV_X1 U7870 ( .A(n9261), .ZN(P1_U4006) );
  AND2_X1 U7871 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7510) );
  NOR2_X1 U7872 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6522), .ZN(n6163) );
  AOI21_X1 U7873 ( .B1(n6522), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6163), .ZN(
        n6520) );
  NOR2_X1 U7874 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n9760), .ZN(n6164) );
  AOI21_X1 U7875 ( .B1(n9760), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6164), .ZN(
        n9762) );
  INV_X1 U7876 ( .A(n6219), .ZN(n9750) );
  INV_X1 U7877 ( .A(n6604), .ZN(n6616) );
  INV_X1 U7878 ( .A(n6636), .ZN(n6648) );
  INV_X1 U7879 ( .A(n6223), .ZN(n6582) );
  NAND2_X1 U7880 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9739) );
  NOR2_X1 U7881 ( .A1(n6580), .A2(n9739), .ZN(n6579) );
  AOI21_X1 U7882 ( .B1(P1_REG2_REG_1__SCAN_IN), .B2(n6582), .A(n6579), .ZN(
        n6645) );
  XOR2_X1 U7883 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6636), .Z(n6644) );
  NOR2_X1 U7884 ( .A1(n6645), .A2(n6644), .ZN(n6643) );
  AOI21_X1 U7885 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(n6648), .A(n6643), .ZN(
        n6613) );
  XOR2_X1 U7886 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6604), .Z(n6612) );
  NOR2_X1 U7887 ( .A1(n6613), .A2(n6612), .ZN(n6611) );
  XNOR2_X1 U7888 ( .A(n6219), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n9748) );
  OAI21_X1 U7889 ( .B1(n9760), .B2(P1_REG2_REG_5__SCAN_IN), .A(n9761), .ZN(
        n6598) );
  MUX2_X1 U7890 ( .A(n6165), .B(P1_REG2_REG_6__SCAN_IN), .S(n6601), .Z(n6597)
         );
  NOR2_X1 U7891 ( .A1(n6598), .A2(n6597), .ZN(n6596) );
  INV_X1 U7892 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7045) );
  XNOR2_X1 U7893 ( .A(n9772), .B(n7045), .ZN(n9775) );
  NOR2_X1 U7894 ( .A1(n9772), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6166) );
  OR2_X1 U7895 ( .A1(n6629), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6168) );
  NAND2_X1 U7896 ( .A1(n6629), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6167) );
  AND2_X1 U7897 ( .A1(n6168), .A2(n6167), .ZN(n6169) );
  OR2_X1 U7898 ( .A1(n6649), .A2(P1_U3084), .ZN(n7704) );
  NOR2_X1 U7899 ( .A1(n9288), .A2(n7745), .ZN(n9857) );
  OAI21_X1 U7900 ( .B1(n6170), .B2(n6169), .A(n9857), .ZN(n6171) );
  NOR2_X1 U7901 ( .A1(n6171), .A2(n6628), .ZN(n6196) );
  NAND2_X1 U7902 ( .A1(n9772), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6184) );
  NOR2_X1 U7903 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6522), .ZN(n6182) );
  INV_X1 U7904 ( .A(n6601), .ZN(n6212) );
  NAND2_X1 U7905 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n9760), .ZN(n6181) );
  INV_X1 U7906 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6172) );
  MUX2_X1 U7907 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6172), .S(n9760), .Z(n9766)
         );
  MUX2_X1 U7908 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6180), .S(n6219), .Z(n9752)
         );
  INV_X1 U7909 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6173) );
  MUX2_X1 U7910 ( .A(n6173), .B(P1_REG1_REG_1__SCAN_IN), .S(n6223), .Z(n6583)
         );
  AND2_X1 U7911 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6584) );
  NAND2_X1 U7912 ( .A1(n6583), .A2(n6584), .ZN(n6638) );
  OR2_X1 U7913 ( .A1(n6223), .A2(n6173), .ZN(n6637) );
  NAND2_X1 U7914 ( .A1(n6638), .A2(n6637), .ZN(n6175) );
  MUX2_X1 U7915 ( .A(n6176), .B(P1_REG1_REG_2__SCAN_IN), .S(n6636), .Z(n6174)
         );
  OR2_X1 U7916 ( .A1(n6636), .A2(n6176), .ZN(n6605) );
  MUX2_X1 U7917 ( .A(n6179), .B(P1_REG1_REG_3__SCAN_IN), .S(n6604), .Z(n6177)
         );
  NAND2_X1 U7918 ( .A1(n6178), .A2(n6177), .ZN(n6608) );
  OAI21_X1 U7919 ( .B1(n6179), .B2(n6604), .A(n6608), .ZN(n9753) );
  NOR2_X1 U7920 ( .A1(n9752), .A2(n9753), .ZN(n9751) );
  NAND2_X1 U7921 ( .A1(n9766), .A2(n9767), .ZN(n9765) );
  NAND2_X1 U7922 ( .A1(n6181), .A2(n9765), .ZN(n6592) );
  AOI22_X1 U7923 ( .A1(n6601), .A2(n5081), .B1(P1_REG1_REG_6__SCAN_IN), .B2(
        n6212), .ZN(n6591) );
  NOR2_X1 U7924 ( .A1(n6592), .A2(n6591), .ZN(n6590) );
  INV_X1 U7925 ( .A(n6522), .ZN(n6208) );
  INV_X1 U7926 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7144) );
  AOI22_X1 U7927 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6208), .B1(n6522), .B2(
        n7144), .ZN(n6516) );
  NOR2_X1 U7928 ( .A1(n6517), .A2(n6516), .ZN(n6515) );
  INV_X1 U7929 ( .A(n9772), .ZN(n6228) );
  INV_X1 U7930 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7238) );
  NAND2_X1 U7931 ( .A1(n6228), .A2(n7238), .ZN(n6183) );
  AND2_X1 U7932 ( .A1(n6183), .A2(n6184), .ZN(n9779) );
  NAND2_X1 U7933 ( .A1(n9780), .A2(n9779), .ZN(n9778) );
  NAND2_X1 U7934 ( .A1(n6184), .A2(n9778), .ZN(n6186) );
  INV_X1 U7935 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7200) );
  INV_X1 U7936 ( .A(n6629), .ZN(n6206) );
  AOI22_X1 U7937 ( .A1(n6629), .A2(n7200), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n6206), .ZN(n6185) );
  NOR2_X1 U7938 ( .A1(n6186), .A2(n6185), .ZN(n6619) );
  AOI21_X1 U7939 ( .B1(n6186), .B2(n6185), .A(n6619), .ZN(n6190) );
  INV_X1 U7940 ( .A(n6187), .ZN(n6189) );
  NAND2_X1 U7941 ( .A1(n6649), .A2(n9736), .ZN(n6652) );
  NOR2_X1 U7942 ( .A1(n6652), .A2(P1_U3084), .ZN(n6188) );
  INV_X1 U7943 ( .A(n9847), .ZN(n9867) );
  NOR2_X1 U7944 ( .A1(n6190), .A2(n9867), .ZN(n6195) );
  INV_X1 U7945 ( .A(n6191), .ZN(n6192) );
  NOR2_X1 U7946 ( .A1(P1_U3083), .A2(n6192), .ZN(n9773) );
  INV_X1 U7947 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10163) );
  NOR2_X2 U7948 ( .A1(n9288), .A2(n9736), .ZN(n9859) );
  INV_X1 U7949 ( .A(n9859), .ZN(n6193) );
  OAI22_X1 U7950 ( .A1(n9870), .A2(n10163), .B1(n6206), .B2(n6193), .ZN(n6194)
         );
  OR4_X1 U7951 ( .A1(n7510), .A2(n6196), .A3(n6195), .A4(n6194), .ZN(P1_U3250)
         );
  XNOR2_X1 U7952 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AND2_X1 U7953 ( .A1(n6203), .A2(n4262), .ZN(n6576) );
  AND2_X1 U7954 ( .A1(n7794), .A2(n4262), .ZN(n7739) );
  INV_X2 U7955 ( .A(n7739), .ZN(n8768) );
  OAI222_X1 U7956 ( .A1(n4268), .A2(n6390), .B1(n8768), .B2(n6222), .C1(n6197), 
        .C2(P2_U3152), .ZN(P2_U3357) );
  OAI222_X1 U7957 ( .A1(n4268), .A2(n6198), .B1(n8768), .B2(n6215), .C1(n4262), 
        .C2(n6500), .ZN(P2_U3355) );
  OAI222_X1 U7958 ( .A1(n4268), .A2(n6199), .B1(n8768), .B2(n6217), .C1(
        P2_U3152), .C2(n6438), .ZN(P2_U3356) );
  OAI222_X1 U7959 ( .A1(n4268), .A2(n6200), .B1(n8768), .B2(n6220), .C1(n4262), 
        .C2(n6465), .ZN(P2_U3354) );
  OAI222_X1 U7960 ( .A1(n4268), .A2(n6201), .B1(n8768), .B2(n6213), .C1(
        P2_U3152), .C2(n6512), .ZN(P2_U3352) );
  OAI222_X1 U7961 ( .A1(n4268), .A2(n6202), .B1(n8768), .B2(n5646), .C1(n4262), 
        .C2(n6470), .ZN(P2_U3353) );
  NAND2_X1 U7962 ( .A1(n6203), .A2(P1_U3084), .ZN(n9645) );
  INV_X1 U7963 ( .A(n6204), .ZN(n6225) );
  AND2_X1 U7964 ( .A1(n7794), .A2(P1_U3084), .ZN(n9634) );
  INV_X1 U7965 ( .A(n9634), .ZN(n9641) );
  OAI222_X1 U7966 ( .A1(n9645), .A2(n6225), .B1(n6206), .B2(P1_U3084), .C1(
        n6205), .C2(n9641), .ZN(P1_U3344) );
  INV_X1 U7967 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6209) );
  INV_X1 U7968 ( .A(n6207), .ZN(n6210) );
  OAI222_X1 U7969 ( .A1(n9641), .A2(n6209), .B1(n9645), .B2(n6210), .C1(
        P1_U3084), .C2(n6208), .ZN(P1_U3346) );
  OAI222_X1 U7970 ( .A1(n4268), .A2(n6211), .B1(n8768), .B2(n6210), .C1(
        P2_U3152), .C2(n6487), .ZN(P2_U3351) );
  INV_X1 U7971 ( .A(n9645), .ZN(n7703) );
  INV_X1 U7972 ( .A(n7703), .ZN(n9639) );
  OAI222_X1 U7973 ( .A1(n9641), .A2(n6214), .B1(n9639), .B2(n6213), .C1(
        P1_U3084), .C2(n6212), .ZN(P1_U3347) );
  OAI222_X1 U7974 ( .A1(n9641), .A2(n6216), .B1(n9639), .B2(n6215), .C1(
        P1_U3084), .C2(n6604), .ZN(P1_U3350) );
  OAI222_X1 U7975 ( .A1(n9641), .A2(n6218), .B1(n9639), .B2(n6217), .C1(
        P1_U3084), .C2(n6636), .ZN(P1_U3351) );
  OAI222_X1 U7976 ( .A1(n9641), .A2(n6221), .B1(n9639), .B2(n6220), .C1(
        P1_U3084), .C2(n6219), .ZN(P1_U3349) );
  OAI222_X1 U7977 ( .A1(n9641), .A2(n6224), .B1(n6223), .B2(P1_U3084), .C1(
        n9639), .C2(n6222), .ZN(P1_U3352) );
  INV_X1 U7978 ( .A(n6914), .ZN(n6918) );
  OAI222_X1 U7979 ( .A1(n4268), .A2(n6226), .B1(n8768), .B2(n6225), .C1(n6918), 
        .C2(n4262), .ZN(P2_U3349) );
  INV_X1 U7980 ( .A(n6227), .ZN(n6230) );
  OAI222_X1 U7981 ( .A1(n9641), .A2(n6229), .B1(n9645), .B2(n6230), .C1(
        P1_U3084), .C2(n6228), .ZN(P1_U3345) );
  INV_X1 U7982 ( .A(n6738), .ZN(n6544) );
  OAI222_X1 U7983 ( .A1(n4268), .A2(n6231), .B1(n8768), .B2(n6230), .C1(
        P2_U3152), .C2(n6544), .ZN(P2_U3350) );
  OAI222_X1 U7984 ( .A1(n9641), .A2(n6233), .B1(n9639), .B2(n5646), .C1(
        P1_U3084), .C2(n6232), .ZN(P1_U3348) );
  INV_X1 U7985 ( .A(n6234), .ZN(n6236) );
  AOI22_X1 U7986 ( .A1(n6684), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9634), .ZN(n6235) );
  OAI21_X1 U7987 ( .B1(n6236), .B2(n9639), .A(n6235), .ZN(P1_U3343) );
  INV_X1 U7988 ( .A(n7009), .ZN(n6929) );
  OAI222_X1 U7989 ( .A1(n4268), .A2(n6237), .B1(n8768), .B2(n6236), .C1(n6929), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U7990 ( .A(n6238), .ZN(n6240) );
  INV_X1 U7991 ( .A(n7362), .ZN(n7353) );
  OAI222_X1 U7992 ( .A1(n9645), .A2(n6240), .B1(n7353), .B2(P1_U3084), .C1(
        n6239), .C2(n9641), .ZN(P1_U3342) );
  INV_X1 U7993 ( .A(n7212), .ZN(n7005) );
  OAI222_X1 U7994 ( .A1(n4268), .A2(n6241), .B1(n8768), .B2(n6240), .C1(n7005), 
        .C2(n4262), .ZN(P2_U3347) );
  INV_X1 U7995 ( .A(n6242), .ZN(n6252) );
  AOI22_X1 U7996 ( .A1(n9786), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n9634), .ZN(n6243) );
  OAI21_X1 U7997 ( .B1(n6252), .B2(n9639), .A(n6243), .ZN(P1_U3341) );
  INV_X1 U7998 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6250) );
  NAND2_X1 U7999 ( .A1(n6244), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6248) );
  NAND2_X1 U8000 ( .A1(n5051), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6247) );
  NAND2_X1 U8001 ( .A1(n6245), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6246) );
  AND3_X1 U8002 ( .A1(n6248), .A2(n6247), .A3(n6246), .ZN(n9075) );
  INV_X1 U8003 ( .A(n9075), .ZN(n8118) );
  NAND2_X1 U8004 ( .A1(P1_U4006), .A2(n8118), .ZN(n6249) );
  OAI21_X1 U8005 ( .B1(P1_U4006), .B2(n6250), .A(n6249), .ZN(P1_U3586) );
  NAND2_X1 U8006 ( .A1(P1_U4006), .A2(n6568), .ZN(n6251) );
  OAI21_X1 U8007 ( .B1(P1_U4006), .B2(n4417), .A(n6251), .ZN(P1_U3555) );
  INV_X1 U8008 ( .A(n7324), .ZN(n7320) );
  OAI222_X1 U8009 ( .A1(n4268), .A2(n6253), .B1(n8768), .B2(n6252), .C1(n4262), 
        .C2(n7320), .ZN(P2_U3346) );
  NAND2_X1 U8010 ( .A1(n8303), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n6254) );
  OAI21_X1 U8011 ( .B1(n8303), .B2(n7800), .A(n6254), .ZN(P2_U3582) );
  INV_X1 U8012 ( .A(n6275), .ZN(n6255) );
  INV_X1 U8013 ( .A(n7474), .ZN(n7469) );
  OAI222_X1 U8014 ( .A1(n4268), .A2(n6256), .B1(n8768), .B2(n6255), .C1(
        P2_U3152), .C2(n7469), .ZN(P2_U3345) );
  NAND2_X1 U8015 ( .A1(n10013), .A2(n6257), .ZN(n6258) );
  NAND2_X1 U8016 ( .A1(n6258), .A2(n5592), .ZN(n6263) );
  INV_X1 U8017 ( .A(n6259), .ZN(n6260) );
  NAND2_X1 U8018 ( .A1(n6260), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7993) );
  INV_X1 U8019 ( .A(n7993), .ZN(n6261) );
  OR2_X1 U8020 ( .A1(n10013), .A2(n6261), .ZN(n6262) );
  NAND2_X1 U8021 ( .A1(n6263), .A2(n6262), .ZN(n9650) );
  NOR2_X1 U8022 ( .A1(n9943), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8023 ( .A(n6264), .ZN(n6273) );
  INV_X1 U8024 ( .A(n7371), .ZN(n9275) );
  OAI222_X1 U8025 ( .A1(n9645), .A2(n6273), .B1(n9275), .B2(P1_U3084), .C1(
        n6265), .C2(n9641), .ZN(P1_U3339) );
  INV_X1 U8026 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6369) );
  NAND2_X1 U8027 ( .A1(n6266), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6270) );
  NAND2_X1 U8028 ( .A1(n4265), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6269) );
  NAND2_X1 U8029 ( .A1(n6267), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6268) );
  NAND3_X1 U8030 ( .A1(n6270), .A2(n6269), .A3(n6268), .ZN(n8414) );
  NAND2_X1 U8031 ( .A1(P2_U3966), .A2(n8414), .ZN(n6271) );
  OAI21_X1 U8032 ( .B1(P2_U3966), .B2(n6369), .A(n6271), .ZN(P2_U3583) );
  NAND2_X1 U8033 ( .A1(P2_U3966), .A2(n6756), .ZN(n6272) );
  OAI21_X1 U8034 ( .B1(P2_U3966), .B2(n5008), .A(n6272), .ZN(P2_U3552) );
  INV_X1 U8035 ( .A(n8330), .ZN(n8327) );
  OAI222_X1 U8036 ( .A1(n4268), .A2(n6274), .B1(n8768), .B2(n6273), .C1(n8327), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  AOI222_X1 U8037 ( .A1(n6275), .A2(n7703), .B1(P2_DATAO_REG_13__SCAN_IN), 
        .B2(n9634), .C1(P1_STATE_REG_SCAN_IN), .C2(n9801), .ZN(n6404) );
  INV_X1 U8038 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10112) );
  AOI22_X1 U8039 ( .A1(n10112), .A2(keyinput15), .B1(keyinput32), .B2(n8648), 
        .ZN(n6276) );
  OAI221_X1 U8040 ( .B1(n10112), .B2(keyinput15), .C1(n8648), .C2(keyinput32), 
        .A(n6276), .ZN(n6286) );
  AOI22_X1 U8041 ( .A1(n5538), .A2(keyinput51), .B1(n6278), .B2(keyinput18), 
        .ZN(n6277) );
  OAI221_X1 U8042 ( .B1(n5538), .B2(keyinput51), .C1(n6278), .C2(keyinput18), 
        .A(n6277), .ZN(n6285) );
  XOR2_X1 U8043 ( .A(n6279), .B(keyinput33), .Z(n6283) );
  XNOR2_X1 U8044 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(keyinput60), .ZN(n6282) );
  XNOR2_X1 U8045 ( .A(P2_IR_REG_6__SCAN_IN), .B(keyinput5), .ZN(n6281) );
  XNOR2_X1 U8046 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(keyinput42), .ZN(n6280) );
  NAND4_X1 U8047 ( .A1(n6283), .A2(n6282), .A3(n6281), .A4(n6280), .ZN(n6284)
         );
  NOR3_X1 U8048 ( .A1(n6286), .A2(n6285), .A3(n6284), .ZN(n6322) );
  INV_X1 U8049 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n6289) );
  INV_X1 U8050 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n6288) );
  AOI22_X1 U8051 ( .A1(n6289), .A2(keyinput19), .B1(keyinput43), .B2(n6288), 
        .ZN(n6287) );
  OAI221_X1 U8052 ( .B1(n6289), .B2(keyinput19), .C1(n6288), .C2(keyinput43), 
        .A(n6287), .ZN(n6297) );
  AOI22_X1 U8053 ( .A1(n5994), .A2(keyinput63), .B1(n6980), .B2(keyinput36), 
        .ZN(n6290) );
  OAI221_X1 U8054 ( .B1(n5994), .B2(keyinput63), .C1(n6980), .C2(keyinput36), 
        .A(n6290), .ZN(n6296) );
  INV_X1 U8055 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n9890) );
  AOI22_X1 U8056 ( .A1(n8232), .A2(keyinput58), .B1(n9890), .B2(keyinput12), 
        .ZN(n6291) );
  OAI221_X1 U8057 ( .B1(n8232), .B2(keyinput58), .C1(n9890), .C2(keyinput12), 
        .A(n6291), .ZN(n6295) );
  INV_X1 U8058 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10108) );
  INV_X1 U8059 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6293) );
  AOI22_X1 U8060 ( .A1(n10108), .A2(keyinput39), .B1(keyinput20), .B2(n6293), 
        .ZN(n6292) );
  OAI221_X1 U8061 ( .B1(n10108), .B2(keyinput39), .C1(n6293), .C2(keyinput20), 
        .A(n6292), .ZN(n6294) );
  NOR4_X1 U8062 ( .A1(n6297), .A2(n6296), .A3(n6295), .A4(n6294), .ZN(n6321)
         );
  INV_X1 U8063 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6385) );
  AOI22_X1 U8064 ( .A1(n6385), .A2(keyinput8), .B1(n6383), .B2(keyinput44), 
        .ZN(n6298) );
  OAI221_X1 U8065 ( .B1(n6385), .B2(keyinput8), .C1(n6383), .C2(keyinput44), 
        .A(n6298), .ZN(n6307) );
  INV_X1 U8066 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n10018) );
  INV_X1 U8067 ( .A(SI_4_), .ZN(n6384) );
  AOI22_X1 U8068 ( .A1(n10018), .A2(keyinput14), .B1(n6384), .B2(keyinput29), 
        .ZN(n6299) );
  OAI221_X1 U8069 ( .B1(n10018), .B2(keyinput14), .C1(n6384), .C2(keyinput29), 
        .A(n6299), .ZN(n6306) );
  INV_X1 U8070 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6301) );
  INV_X1 U8071 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9281) );
  AOI22_X1 U8072 ( .A1(n6301), .A2(keyinput10), .B1(n9281), .B2(keyinput34), 
        .ZN(n6300) );
  OAI221_X1 U8073 ( .B1(n6301), .B2(keyinput10), .C1(n9281), .C2(keyinput34), 
        .A(n6300), .ZN(n6305) );
  XNOR2_X1 U8074 ( .A(P2_REG1_REG_26__SCAN_IN), .B(keyinput62), .ZN(n6303) );
  XNOR2_X1 U8075 ( .A(SI_1_), .B(keyinput37), .ZN(n6302) );
  NAND2_X1 U8076 ( .A1(n6303), .A2(n6302), .ZN(n6304) );
  NOR4_X1 U8077 ( .A1(n6307), .A2(n6306), .A3(n6305), .A4(n6304), .ZN(n6320)
         );
  INV_X1 U8078 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6309) );
  AOI22_X1 U8079 ( .A1(n7571), .A2(keyinput35), .B1(keyinput27), .B2(n6309), 
        .ZN(n6308) );
  OAI221_X1 U8080 ( .B1(n7571), .B2(keyinput35), .C1(n6309), .C2(keyinput27), 
        .A(n6308), .ZN(n6318) );
  INV_X1 U8081 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n10016) );
  INV_X1 U8082 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6311) );
  AOI22_X1 U8083 ( .A1(n10016), .A2(keyinput40), .B1(keyinput16), .B2(n6311), 
        .ZN(n6310) );
  OAI221_X1 U8084 ( .B1(n10016), .B2(keyinput40), .C1(n6311), .C2(keyinput16), 
        .A(n6310), .ZN(n6317) );
  AOI22_X1 U8085 ( .A1(n7781), .A2(keyinput52), .B1(n5403), .B2(keyinput41), 
        .ZN(n6312) );
  OAI221_X1 U8086 ( .B1(n7781), .B2(keyinput52), .C1(n5403), .C2(keyinput41), 
        .A(n6312), .ZN(n6316) );
  INV_X1 U8087 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6685) );
  XOR2_X1 U8088 ( .A(n6685), .B(keyinput30), .Z(n6314) );
  XNOR2_X1 U8089 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput59), .ZN(n6313) );
  NAND2_X1 U8090 ( .A1(n6314), .A2(n6313), .ZN(n6315) );
  NOR4_X1 U8091 ( .A1(n6318), .A2(n6317), .A3(n6316), .A4(n6315), .ZN(n6319)
         );
  NAND4_X1 U8092 ( .A1(n6322), .A2(n6321), .A3(n6320), .A4(n6319), .ZN(n6368)
         );
  INV_X1 U8093 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8691) );
  AOI22_X1 U8094 ( .A1(n8691), .A2(keyinput38), .B1(n6324), .B2(keyinput31), 
        .ZN(n6323) );
  OAI221_X1 U8095 ( .B1(n8691), .B2(keyinput38), .C1(n6324), .C2(keyinput31), 
        .A(n6323), .ZN(n6332) );
  AOI22_X1 U8096 ( .A1(n6406), .A2(keyinput9), .B1(keyinput49), .B2(n6493), 
        .ZN(n6325) );
  OAI221_X1 U8097 ( .B1(n6406), .B2(keyinput9), .C1(n6493), .C2(keyinput49), 
        .A(n6325), .ZN(n6331) );
  INV_X1 U8098 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8765) );
  AOI22_X1 U8099 ( .A1(n5711), .A2(keyinput57), .B1(keyinput55), .B2(n8765), 
        .ZN(n6326) );
  OAI221_X1 U8100 ( .B1(n5711), .B2(keyinput57), .C1(n8765), .C2(keyinput55), 
        .A(n6326), .ZN(n6330) );
  INV_X1 U8101 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n10015) );
  INV_X1 U8102 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n6328) );
  AOI22_X1 U8103 ( .A1(n10015), .A2(keyinput7), .B1(keyinput4), .B2(n6328), 
        .ZN(n6327) );
  OAI221_X1 U8104 ( .B1(n10015), .B2(keyinput7), .C1(n6328), .C2(keyinput4), 
        .A(n6327), .ZN(n6329) );
  NOR4_X1 U8105 ( .A1(n6332), .A2(n6331), .A3(n6330), .A4(n6329), .ZN(n6366)
         );
  AOI22_X1 U8106 ( .A1(n6165), .A2(keyinput0), .B1(n6334), .B2(keyinput25), 
        .ZN(n6333) );
  OAI221_X1 U8107 ( .B1(n6165), .B2(keyinput0), .C1(n6334), .C2(keyinput25), 
        .A(n6333), .ZN(n6337) );
  INV_X1 U8108 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9824) );
  XNOR2_X1 U8109 ( .A(n9824), .B(keyinput2), .ZN(n6336) );
  XNOR2_X1 U8110 ( .A(n6391), .B(keyinput26), .ZN(n6335) );
  OR3_X1 U8111 ( .A1(n6337), .A2(n6336), .A3(n6335), .ZN(n6342) );
  INV_X1 U8112 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6689) );
  INV_X1 U8113 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n10017) );
  AOI22_X1 U8114 ( .A1(n6689), .A2(keyinput45), .B1(n10017), .B2(keyinput21), 
        .ZN(n6338) );
  OAI221_X1 U8115 ( .B1(n6689), .B2(keyinput45), .C1(n10017), .C2(keyinput21), 
        .A(n6338), .ZN(n6341) );
  AOI22_X1 U8116 ( .A1(n6130), .A2(keyinput53), .B1(n5571), .B2(keyinput1), 
        .ZN(n6339) );
  OAI221_X1 U8117 ( .B1(n6130), .B2(keyinput53), .C1(n5571), .C2(keyinput1), 
        .A(n6339), .ZN(n6340) );
  NOR3_X1 U8118 ( .A1(n6342), .A2(n6341), .A3(n6340), .ZN(n6365) );
  INV_X1 U8119 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8608) );
  INV_X1 U8120 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n6388) );
  AOI22_X1 U8121 ( .A1(n8608), .A2(keyinput3), .B1(keyinput24), .B2(n6388), 
        .ZN(n6343) );
  OAI221_X1 U8122 ( .B1(n8608), .B2(keyinput3), .C1(n6388), .C2(keyinput24), 
        .A(n6343), .ZN(n6352) );
  INV_X1 U8123 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n9889) );
  AOI22_X1 U8124 ( .A1(n9889), .A2(keyinput28), .B1(keyinput17), .B2(n5333), 
        .ZN(n6344) );
  OAI221_X1 U8125 ( .B1(n9889), .B2(keyinput28), .C1(n5333), .C2(keyinput17), 
        .A(n6344), .ZN(n6351) );
  AOI22_X1 U8126 ( .A1(n5081), .A2(keyinput46), .B1(keyinput50), .B2(n6346), 
        .ZN(n6345) );
  OAI221_X1 U8127 ( .B1(n5081), .B2(keyinput46), .C1(n6346), .C2(keyinput50), 
        .A(n6345), .ZN(n6350) );
  AOI22_X1 U8128 ( .A1(n6348), .A2(keyinput54), .B1(n8896), .B2(keyinput11), 
        .ZN(n6347) );
  OAI221_X1 U8129 ( .B1(n6348), .B2(keyinput54), .C1(n8896), .C2(keyinput11), 
        .A(n6347), .ZN(n6349) );
  NOR4_X1 U8130 ( .A1(n6352), .A2(n6351), .A3(n6350), .A4(n6349), .ZN(n6364)
         );
  INV_X1 U8131 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9946) );
  AOI22_X1 U8132 ( .A1(n8712), .A2(keyinput48), .B1(n9946), .B2(keyinput56), 
        .ZN(n6353) );
  OAI221_X1 U8133 ( .B1(n8712), .B2(keyinput48), .C1(n9946), .C2(keyinput56), 
        .A(n6353), .ZN(n6362) );
  AOI22_X1 U8134 ( .A1(n6369), .A2(keyinput61), .B1(n6355), .B2(keyinput13), 
        .ZN(n6354) );
  OAI221_X1 U8135 ( .B1(n6369), .B2(keyinput61), .C1(n6355), .C2(keyinput13), 
        .A(n6354), .ZN(n6361) );
  INV_X1 U8136 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n6371) );
  AOI22_X1 U8137 ( .A1(n8703), .A2(keyinput6), .B1(n6371), .B2(keyinput47), 
        .ZN(n6356) );
  OAI221_X1 U8138 ( .B1(n8703), .B2(keyinput6), .C1(n6371), .C2(keyinput47), 
        .A(n6356), .ZN(n6360) );
  XNOR2_X1 U8139 ( .A(P1_REG1_REG_15__SCAN_IN), .B(keyinput22), .ZN(n6358) );
  XNOR2_X1 U8140 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput23), .ZN(n6357) );
  NAND2_X1 U8141 ( .A1(n6358), .A2(n6357), .ZN(n6359) );
  NOR4_X1 U8142 ( .A1(n6362), .A2(n6361), .A3(n6360), .A4(n6359), .ZN(n6363)
         );
  NAND4_X1 U8143 ( .A1(n6366), .A2(n6365), .A3(n6364), .A4(n6363), .ZN(n6367)
         );
  NOR2_X1 U8144 ( .A1(n6368), .A2(n6367), .ZN(n6402) );
  NOR4_X1 U8145 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(P1_REG2_REG_26__SCAN_IN), 
        .A3(P1_REG2_REG_11__SCAN_IN), .A4(P2_REG2_REG_24__SCAN_IN), .ZN(n6400)
         );
  INV_X1 U8146 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n6370) );
  NAND3_X1 U8147 ( .A1(n6371), .A2(n6370), .A3(n6369), .ZN(n6374) );
  NAND4_X1 U8148 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), 
        .A3(P2_IR_REG_17__SCAN_IN), .A4(P1_DATAO_REG_29__SCAN_IN), .ZN(n6373)
         );
  NAND4_X1 U8149 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_REG0_REG_27__SCAN_IN), 
        .A3(P2_REG0_REG_26__SCAN_IN), .A4(P2_REG1_REG_22__SCAN_IN), .ZN(n6372)
         );
  NOR4_X1 U8150 ( .A1(SI_29_), .A2(n6374), .A3(n6373), .A4(n6372), .ZN(n6399)
         );
  NAND4_X1 U8151 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_REG3_REG_9__SCAN_IN), 
        .A3(P2_REG1_REG_9__SCAN_IN), .A4(P2_REG2_REG_3__SCAN_IN), .ZN(n6378)
         );
  NAND4_X1 U8152 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_REG2_REG_6__SCAN_IN), 
        .A3(P1_REG1_REG_6__SCAN_IN), .A4(P2_REG1_REG_7__SCAN_IN), .ZN(n6377)
         );
  NAND4_X1 U8153 ( .A1(P1_REG2_REG_21__SCAN_IN), .A2(P1_REG1_REG_17__SCAN_IN), 
        .A3(P2_REG2_REG_26__SCAN_IN), .A4(P1_DATAO_REG_30__SCAN_IN), .ZN(n6376) );
  NAND4_X1 U8154 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG3_REG_24__SCAN_IN), 
        .A3(P2_REG2_REG_20__SCAN_IN), .A4(P2_REG2_REG_29__SCAN_IN), .ZN(n6375)
         );
  NOR4_X1 U8155 ( .A1(n6378), .A2(n6377), .A3(n6376), .A4(n6375), .ZN(n6398)
         );
  NOR4_X1 U8156 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(SI_22_), .A3(
        P2_DATAO_REG_15__SCAN_IN), .A4(P2_IR_REG_7__SCAN_IN), .ZN(n6382) );
  NOR4_X1 U8157 ( .A1(P2_REG1_REG_26__SCAN_IN), .A2(P2_REG1_REG_25__SCAN_IN), 
        .A3(P2_REG1_REG_31__SCAN_IN), .A4(P2_REG0_REG_30__SCAN_IN), .ZN(n6381)
         );
  NOR4_X1 U8158 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), .A3(
        P2_REG0_REG_3__SCAN_IN), .A4(P2_REG0_REG_24__SCAN_IN), .ZN(n6380) );
  NOR4_X1 U8159 ( .A1(P1_D_REG_12__SCAN_IN), .A2(SI_27_), .A3(
        P1_REG1_REG_22__SCAN_IN), .A4(P1_REG1_REG_31__SCAN_IN), .ZN(n6379) );
  NAND4_X1 U8160 ( .A1(n6382), .A2(n6381), .A3(n6380), .A4(n6379), .ZN(n6396)
         );
  NOR4_X1 U8161 ( .A1(SI_5_), .A2(SI_1_), .A3(n6384), .A4(n6383), .ZN(n6386)
         );
  NAND4_X1 U8162 ( .A1(n6387), .A2(n6386), .A3(n6385), .A4(n9824), .ZN(n6395)
         );
  NAND4_X1 U8163 ( .A1(n6391), .A2(n6390), .A3(n6389), .A4(n6388), .ZN(n6394)
         );
  NAND4_X1 U8164 ( .A1(n6392), .A2(P1_IR_REG_6__SCAN_IN), .A3(
        P2_ADDR_REG_13__SCAN_IN), .A4(P1_ADDR_REG_11__SCAN_IN), .ZN(n6393) );
  NOR4_X1 U8165 ( .A1(n6396), .A2(n6395), .A3(n6394), .A4(n6393), .ZN(n6397)
         );
  NAND4_X1 U8166 ( .A1(n6400), .A2(n6399), .A3(n6398), .A4(n6397), .ZN(n6401)
         );
  XNOR2_X1 U8167 ( .A(n6402), .B(n6401), .ZN(n6403) );
  XNOR2_X1 U8168 ( .A(n6404), .B(n6403), .ZN(P1_U3340) );
  INV_X1 U8169 ( .A(n6405), .ZN(n6407) );
  INV_X1 U8170 ( .A(n9819), .ZN(n9276) );
  OAI222_X1 U8171 ( .A1(n9641), .A2(n6406), .B1(n9645), .B2(n6407), .C1(
        P1_U3084), .C2(n9276), .ZN(P1_U3338) );
  INV_X1 U8172 ( .A(n8340), .ZN(n8349) );
  OAI222_X1 U8173 ( .A1(n4268), .A2(n6408), .B1(n8768), .B2(n6407), .C1(n4262), 
        .C2(n8349), .ZN(P2_U3343) );
  OR2_X1 U8174 ( .A1(n6943), .A2(n9232), .ZN(n9873) );
  OR2_X1 U8175 ( .A1(n6554), .A2(n6417), .ZN(n9238) );
  NAND2_X1 U8176 ( .A1(n9873), .A2(n9238), .ZN(n6411) );
  NOR2_X1 U8177 ( .A1(n6409), .A2(n6905), .ZN(n6699) );
  INV_X1 U8178 ( .A(n6699), .ZN(n6410) );
  NAND3_X1 U8179 ( .A1(n6411), .A2(n9895), .A3(n6410), .ZN(n6702) );
  NAND2_X1 U8180 ( .A1(n6702), .A2(n6412), .ZN(n7252) );
  NOR2_X1 U8181 ( .A1(n9606), .A2(n6699), .ZN(n6413) );
  NOR2_X1 U8182 ( .A1(n7252), .A2(n6413), .ZN(n6676) );
  INV_X1 U8183 ( .A(n6676), .ZN(n6571) );
  AOI22_X1 U8184 ( .A1(n6571), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n6900), .B2(
        n8928), .ZN(n6427) );
  AND2_X1 U8185 ( .A1(n6699), .A2(n9895), .ZN(n6424) );
  AND2_X1 U8186 ( .A1(n9911), .A2(n9079), .ZN(n6696) );
  NAND2_X1 U8187 ( .A1(n6415), .A2(n6414), .ZN(n6416) );
  NAND2_X1 U8188 ( .A1(n6553), .A2(n6568), .ZN(n6419) );
  AOI22_X1 U8189 ( .A1(n6661), .A2(n6900), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n6420), .ZN(n6418) );
  AND2_X1 U8190 ( .A1(n6419), .A2(n6418), .ZN(n6423) );
  NAND2_X1 U8191 ( .A1(n6661), .A2(n6568), .ZN(n6422) );
  INV_X1 U8192 ( .A(n6424), .ZN(n6425) );
  NOR2_X1 U8193 ( .A1(n6425), .A2(n9238), .ZN(n6567) );
  AND2_X1 U8194 ( .A1(n6567), .A2(n7745), .ZN(n8942) );
  AOI22_X1 U8195 ( .A1(n8935), .A2(n6653), .B1(n8942), .B2(n9262), .ZN(n6426)
         );
  NAND2_X1 U8196 ( .A1(n6427), .A2(n6426), .ZN(P1_U3230) );
  NAND2_X1 U8197 ( .A1(n10013), .A2(n6428), .ZN(n6432) );
  OR2_X1 U8198 ( .A1(n6034), .A2(P2_U3152), .ZN(n7740) );
  OAI21_X1 U8199 ( .B1(n6429), .B2(n7740), .A(n7993), .ZN(n6430) );
  INV_X1 U8200 ( .A(n6430), .ZN(n6431) );
  NAND2_X1 U8201 ( .A1(n6432), .A2(n6431), .ZN(n6433) );
  NAND2_X1 U8202 ( .A1(n6433), .A2(n5592), .ZN(n6441) );
  NAND2_X1 U8203 ( .A1(n8303), .A2(n6441), .ZN(n6453) );
  AND2_X1 U8204 ( .A1(n6034), .A2(n6453), .ZN(n9668) );
  NOR2_X1 U8205 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6434), .ZN(n6446) );
  NAND2_X1 U8206 ( .A1(n6452), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6439) );
  MUX2_X1 U8207 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n5608), .S(n6452), .Z(n6497)
         );
  INV_X1 U8208 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6437) );
  XNOR2_X1 U8209 ( .A(n6438), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n9670) );
  NAND2_X1 U8210 ( .A1(n9656), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6436) );
  INV_X1 U8211 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6435) );
  MUX2_X1 U8212 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6435), .S(n9656), .Z(n9658)
         );
  NAND3_X1 U8213 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .A3(n9658), .ZN(n9657) );
  NAND2_X1 U8214 ( .A1(n6436), .A2(n9657), .ZN(n9671) );
  NAND2_X1 U8215 ( .A1(n9670), .A2(n9671), .ZN(n9669) );
  OAI21_X1 U8216 ( .B1(n6438), .B2(n6437), .A(n9669), .ZN(n6496) );
  NAND2_X1 U8217 ( .A1(n6497), .A2(n6496), .ZN(n6495) );
  AND2_X1 U8218 ( .A1(n6439), .A2(n6495), .ZN(n6444) );
  INV_X1 U8219 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6440) );
  MUX2_X1 U8220 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6440), .S(n6465), .Z(n6443)
         );
  NOR2_X1 U8221 ( .A1(n6444), .A2(n6443), .ZN(n6463) );
  INV_X1 U8222 ( .A(n6441), .ZN(n6442) );
  AND2_X1 U8223 ( .A1(n6125), .A2(n6442), .ZN(n9936) );
  INV_X1 U8224 ( .A(n9936), .ZN(n9941) );
  AOI211_X1 U8225 ( .C1(n6444), .C2(n6443), .A(n6463), .B(n9941), .ZN(n6445)
         );
  AOI211_X1 U8226 ( .C1(n9943), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n6446), .B(
        n6445), .ZN(n6456) );
  INV_X1 U8227 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6447) );
  INV_X1 U8228 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10008) );
  NAND2_X1 U8229 ( .A1(n9656), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6448) );
  OAI21_X1 U8230 ( .B1(n9656), .B2(P2_REG2_REG_1__SCAN_IN), .A(n6448), .ZN(
        n9652) );
  AND2_X1 U8231 ( .A1(n9656), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6449) );
  NOR2_X1 U8232 ( .A1(n9651), .A2(n6449), .ZN(n9665) );
  NAND2_X1 U8233 ( .A1(n9667), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6450) );
  OAI21_X1 U8234 ( .B1(n9667), .B2(P2_REG2_REG_2__SCAN_IN), .A(n6450), .ZN(
        n9664) );
  NAND2_X1 U8235 ( .A1(n6452), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6451) );
  OAI21_X1 U8236 ( .B1(n6452), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6451), .ZN(
        n6491) );
  AND2_X1 U8237 ( .A1(n6453), .A2(n7989), .ZN(n9938) );
  OAI211_X1 U8238 ( .C1(n4282), .C2(n4365), .A(n9937), .B(n6457), .ZN(n6455)
         );
  OAI211_X1 U8239 ( .C1(n9939), .C2(n6465), .A(n6456), .B(n6455), .ZN(P2_U3249) );
  INV_X1 U8240 ( .A(n6465), .ZN(n6458) );
  NAND2_X1 U8241 ( .A1(n6480), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6459) );
  OAI21_X1 U8242 ( .B1(n6480), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6459), .ZN(
        n6460) );
  AOI211_X1 U8243 ( .C1(n6461), .C2(n6460), .A(n6473), .B(n9662), .ZN(n6472)
         );
  AND2_X1 U8244 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6462) );
  AOI21_X1 U8245 ( .B1(n9943), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6462), .ZN(
        n6469) );
  MUX2_X1 U8246 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n5634), .S(n6480), .Z(n6467)
         );
  INV_X1 U8247 ( .A(n6463), .ZN(n6464) );
  OAI21_X1 U8248 ( .B1(n6440), .B2(n6465), .A(n6464), .ZN(n6466) );
  NAND2_X1 U8249 ( .A1(n6467), .A2(n6466), .ZN(n6481) );
  OAI211_X1 U8250 ( .C1(n6467), .C2(n6466), .A(n9936), .B(n6481), .ZN(n6468)
         );
  OAI211_X1 U8251 ( .C1(n9939), .C2(n6470), .A(n6469), .B(n6468), .ZN(n6471)
         );
  OR2_X1 U8252 ( .A1(n6472), .A2(n6471), .ZN(P2_U3250) );
  INV_X1 U8253 ( .A(n6512), .ZN(n6476) );
  INV_X1 U8254 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6474) );
  MUX2_X1 U8255 ( .A(n6474), .B(P2_REG2_REG_6__SCAN_IN), .S(n6512), .Z(n6475)
         );
  INV_X1 U8256 ( .A(n6475), .ZN(n6504) );
  AOI21_X1 U8257 ( .B1(n6476), .B2(P2_REG2_REG_6__SCAN_IN), .A(n6503), .ZN(
        n6479) );
  NAND2_X1 U8258 ( .A1(n6538), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6477) );
  OAI21_X1 U8259 ( .B1(n6538), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6477), .ZN(
        n6478) );
  AOI211_X1 U8260 ( .C1(n6479), .C2(n6478), .A(n6537), .B(n9662), .ZN(n6489)
         );
  AND2_X1 U8261 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6874) );
  AOI21_X1 U8262 ( .B1(n9943), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n6874), .ZN(
        n6486) );
  MUX2_X1 U8263 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10108), .S(n6538), .Z(n6484)
         );
  INV_X1 U8264 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10106) );
  MUX2_X1 U8265 ( .A(n10106), .B(P2_REG1_REG_6__SCAN_IN), .S(n6512), .Z(n6508)
         );
  NAND2_X1 U8266 ( .A1(n6480), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6482) );
  NAND2_X1 U8267 ( .A1(n6482), .A2(n6481), .ZN(n6509) );
  NAND2_X1 U8268 ( .A1(n6508), .A2(n6509), .ZN(n6507) );
  OAI21_X1 U8269 ( .B1(n6512), .B2(n10106), .A(n6507), .ZN(n6483) );
  NAND2_X1 U8270 ( .A1(n6484), .A2(n6483), .ZN(n6528) );
  OAI211_X1 U8271 ( .C1(n6484), .C2(n6483), .A(n9936), .B(n6528), .ZN(n6485)
         );
  OAI211_X1 U8272 ( .C1(n9939), .C2(n6487), .A(n6486), .B(n6485), .ZN(n6488)
         );
  OR2_X1 U8273 ( .A1(n6489), .A2(n6488), .ZN(P2_U3252) );
  AOI211_X1 U8274 ( .C1(n6492), .C2(n6491), .A(n6490), .B(n9662), .ZN(n6502)
         );
  NOR2_X1 U8275 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6493), .ZN(n6494) );
  AOI21_X1 U8276 ( .B1(n9943), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n6494), .ZN(
        n6499) );
  OAI211_X1 U8277 ( .C1(n6497), .C2(n6496), .A(n9936), .B(n6495), .ZN(n6498)
         );
  OAI211_X1 U8278 ( .C1(n9939), .C2(n6500), .A(n6499), .B(n6498), .ZN(n6501)
         );
  OR2_X1 U8279 ( .A1(n6502), .A2(n6501), .ZN(P2_U3248) );
  AOI211_X1 U8280 ( .C1(n6505), .C2(n6504), .A(n6503), .B(n9662), .ZN(n6514)
         );
  NAND2_X1 U8281 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(n4262), .ZN(n6960) );
  INV_X1 U8282 ( .A(n6960), .ZN(n6506) );
  AOI21_X1 U8283 ( .B1(n9943), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n6506), .ZN(
        n6511) );
  OAI211_X1 U8284 ( .C1(n6509), .C2(n6508), .A(n9936), .B(n6507), .ZN(n6510)
         );
  OAI211_X1 U8285 ( .C1(n9939), .C2(n6512), .A(n6511), .B(n6510), .ZN(n6513)
         );
  OR2_X1 U8286 ( .A1(n6514), .A2(n6513), .ZN(P2_U3251) );
  INV_X1 U8287 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6527) );
  AOI21_X1 U8288 ( .B1(n6517), .B2(n6516), .A(n6515), .ZN(n6524) );
  OAI21_X1 U8289 ( .B1(n6520), .B2(n6519), .A(n6518), .ZN(n6521) );
  AOI22_X1 U8290 ( .A1(n6522), .A2(n9859), .B1(n9857), .B2(n6521), .ZN(n6523)
         );
  NAND2_X1 U8291 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7334) );
  OAI211_X1 U8292 ( .C1(n6524), .C2(n9867), .A(n6523), .B(n7334), .ZN(n6525)
         );
  INV_X1 U8293 ( .A(n6525), .ZN(n6526) );
  OAI21_X1 U8294 ( .B1(n6527), .B2(n9870), .A(n6526), .ZN(P1_U3248) );
  NAND2_X1 U8295 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(n4262), .ZN(n6974) );
  INV_X1 U8296 ( .A(n6974), .ZN(n6536) );
  NAND2_X1 U8297 ( .A1(n6538), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6529) );
  NAND2_X1 U8298 ( .A1(n6529), .A2(n6528), .ZN(n6531) );
  INV_X1 U8299 ( .A(n6531), .ZN(n6534) );
  INV_X1 U8300 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10110) );
  MUX2_X1 U8301 ( .A(n10110), .B(P2_REG1_REG_8__SCAN_IN), .S(n6738), .Z(n6533)
         );
  MUX2_X1 U8302 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n10110), .S(n6738), .Z(n6530)
         );
  NAND2_X1 U8303 ( .A1(n6531), .A2(n6530), .ZN(n6741) );
  INV_X1 U8304 ( .A(n6741), .ZN(n6532) );
  AOI211_X1 U8305 ( .C1(n6534), .C2(n6533), .A(n6532), .B(n9941), .ZN(n6535)
         );
  AOI211_X1 U8306 ( .C1(n9943), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n6536), .B(
        n6535), .ZN(n6543) );
  XNOR2_X1 U8307 ( .A(n6738), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n6539) );
  AOI211_X1 U8308 ( .C1(n6540), .C2(n6539), .A(n6734), .B(n9662), .ZN(n6541)
         );
  INV_X1 U8309 ( .A(n6541), .ZN(n6542) );
  OAI211_X1 U8310 ( .C1(n9939), .C2(n6544), .A(n6543), .B(n6542), .ZN(P2_U3253) );
  INV_X1 U8311 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9737) );
  NAND2_X1 U8312 ( .A1(n9238), .A2(n6943), .ZN(n6545) );
  AND2_X1 U8313 ( .A1(n6984), .A2(n6568), .ZN(n9185) );
  NOR2_X1 U8314 ( .A1(n9185), .A2(n6895), .ZN(n9090) );
  OR2_X1 U8315 ( .A1(n6545), .A2(n9090), .ZN(n6547) );
  OR2_X1 U8316 ( .A1(n9681), .A2(n6557), .ZN(n6546) );
  NAND2_X1 U8317 ( .A1(n6547), .A2(n6546), .ZN(n6987) );
  INV_X1 U8318 ( .A(n6987), .ZN(n6548) );
  OAI21_X1 U8319 ( .B1(n6984), .B2(n6943), .A(n6548), .ZN(n6550) );
  NAND2_X1 U8320 ( .A1(n6550), .A2(n9935), .ZN(n6549) );
  OAI21_X1 U8321 ( .B1(n9935), .B2(n9737), .A(n6549), .ZN(P1_U3523) );
  INV_X1 U8322 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6552) );
  NAND2_X1 U8323 ( .A1(n6550), .A2(n9929), .ZN(n6551) );
  OAI21_X1 U8324 ( .B1(n9929), .B2(n6552), .A(n6551), .ZN(P1_U3454) );
  OAI22_X1 U8325 ( .A1(n6660), .A2(n6557), .B1(n7263), .B2(n6556), .ZN(n6566)
         );
  NAND2_X1 U8326 ( .A1(n6555), .A2(n4847), .ZN(n6562) );
  INV_X1 U8327 ( .A(n6562), .ZN(n6560) );
  XNOR2_X1 U8328 ( .A(n6558), .B(n8063), .ZN(n6561) );
  INV_X1 U8329 ( .A(n6561), .ZN(n6559) );
  INV_X1 U8330 ( .A(n6669), .ZN(n6564) );
  AOI21_X1 U8331 ( .B1(n6566), .B2(n6565), .A(n6564), .ZN(n6573) );
  OR2_X1 U8332 ( .A1(n9911), .A2(n6556), .ZN(n9897) );
  AOI22_X1 U8333 ( .A1(n8936), .A2(n6568), .B1(n8942), .B2(n9260), .ZN(n6569)
         );
  OAI21_X1 U8334 ( .B1(n6571), .B2(n9897), .A(n6569), .ZN(n6570) );
  AOI21_X1 U8335 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n6571), .A(n6570), .ZN(
        n6572) );
  OAI21_X1 U8336 ( .B1(n6573), .B2(n4653), .A(n6572), .ZN(P1_U3220) );
  INV_X1 U8337 ( .A(n6574), .ZN(n6578) );
  AOI22_X1 U8338 ( .A1(n9831), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n9634), .ZN(n6575) );
  OAI21_X1 U8339 ( .B1(n6578), .B2(n9639), .A(n6575), .ZN(P1_U3337) );
  AOI22_X1 U8340 ( .A1(n8365), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n6576), .ZN(n6577) );
  OAI21_X1 U8341 ( .B1(n6578), .B2(n8768), .A(n6577), .ZN(P2_U3342) );
  INV_X1 U8342 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6589) );
  INV_X1 U8343 ( .A(n9857), .ZN(n9826) );
  AOI211_X1 U8344 ( .C1(n9739), .C2(n6580), .A(n6579), .B(n9826), .ZN(n6581)
         );
  AOI21_X1 U8345 ( .B1(n9859), .B2(n6582), .A(n6581), .ZN(n6588) );
  OAI211_X1 U8346 ( .C1(n6584), .C2(n6583), .A(n9847), .B(n6638), .ZN(n6585)
         );
  OAI21_X1 U8347 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6903), .A(n6585), .ZN(n6586) );
  INV_X1 U8348 ( .A(n6586), .ZN(n6587) );
  OAI211_X1 U8349 ( .C1(n9870), .C2(n6589), .A(n6588), .B(n6587), .ZN(P1_U3242) );
  INV_X1 U8350 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6603) );
  AOI21_X1 U8351 ( .B1(n6592), .B2(n6591), .A(n6590), .ZN(n6595) );
  NOR2_X1 U8352 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6593), .ZN(n7254) );
  INV_X1 U8353 ( .A(n7254), .ZN(n6594) );
  OAI21_X1 U8354 ( .B1(n9867), .B2(n6595), .A(n6594), .ZN(n6600) );
  AOI211_X1 U8355 ( .C1(n6598), .C2(n6597), .A(n6596), .B(n9826), .ZN(n6599)
         );
  AOI211_X1 U8356 ( .C1(n9859), .C2(n6601), .A(n6600), .B(n6599), .ZN(n6602)
         );
  OAI21_X1 U8357 ( .B1(n9870), .B2(n6603), .A(n6602), .ZN(P1_U3247) );
  INV_X1 U8358 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6618) );
  MUX2_X1 U8359 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6179), .S(n6604), .Z(n6606)
         );
  NAND3_X1 U8360 ( .A1(n6606), .A2(n6641), .A3(n6605), .ZN(n6607) );
  NAND3_X1 U8361 ( .A1(n9847), .A2(n6608), .A3(n6607), .ZN(n6610) );
  INV_X1 U8362 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7084) );
  NOR2_X1 U8363 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7084), .ZN(n6718) );
  INV_X1 U8364 ( .A(n6718), .ZN(n6609) );
  NAND2_X1 U8365 ( .A1(n6610), .A2(n6609), .ZN(n6615) );
  AOI211_X1 U8366 ( .C1(n6613), .C2(n6612), .A(n6611), .B(n9826), .ZN(n6614)
         );
  AOI211_X1 U8367 ( .C1(n9859), .C2(n6616), .A(n6615), .B(n6614), .ZN(n6617)
         );
  OAI21_X1 U8368 ( .B1(n9870), .B2(n6618), .A(n6617), .ZN(P1_U3244) );
  NOR2_X1 U8369 ( .A1(n6629), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6620) );
  INV_X1 U8370 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6621) );
  MUX2_X1 U8371 ( .A(n6621), .B(P1_REG1_REG_10__SCAN_IN), .S(n6684), .Z(n6623)
         );
  INV_X1 U8372 ( .A(n6680), .ZN(n6622) );
  AOI21_X1 U8373 ( .B1(n6624), .B2(n6623), .A(n6622), .ZN(n6635) );
  NAND2_X1 U8374 ( .A1(n9859), .A2(n6684), .ZN(n6627) );
  NOR2_X1 U8375 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6625), .ZN(n7626) );
  INV_X1 U8376 ( .A(n7626), .ZN(n6626) );
  NAND2_X1 U8377 ( .A1(n6627), .A2(n6626), .ZN(n6633) );
  XNOR2_X1 U8378 ( .A(n6684), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n6630) );
  AOI211_X1 U8379 ( .C1(n6631), .C2(n6630), .A(n9826), .B(n6683), .ZN(n6632)
         );
  AOI211_X1 U8380 ( .C1(n9773), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n6633), .B(
        n6632), .ZN(n6634) );
  OAI21_X1 U8381 ( .B1(n6635), .B2(n9867), .A(n6634), .ZN(P1_U3251) );
  INV_X1 U8382 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6655) );
  MUX2_X1 U8383 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6176), .S(n6636), .Z(n6639)
         );
  NAND3_X1 U8384 ( .A1(n6639), .A2(n6638), .A3(n6637), .ZN(n6640) );
  NAND3_X1 U8385 ( .A1(n9847), .A2(n6641), .A3(n6640), .ZN(n6642) );
  OAI21_X1 U8386 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n7062), .A(n6642), .ZN(n6647) );
  AOI211_X1 U8387 ( .C1(n6645), .C2(n6644), .A(n6643), .B(n9826), .ZN(n6646)
         );
  AOI211_X1 U8388 ( .C1(n9859), .C2(n6648), .A(n6647), .B(n6646), .ZN(n6654)
         );
  INV_X1 U8389 ( .A(n6649), .ZN(n9740) );
  NAND2_X1 U8390 ( .A1(n9740), .A2(n9736), .ZN(n9237) );
  INV_X1 U8391 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6983) );
  OAI211_X1 U8392 ( .C1(n6983), .C2(n7745), .A(n6652), .B(n4606), .ZN(n9735)
         );
  OAI211_X1 U8393 ( .C1(n9739), .C2(n9237), .A(P1_U4006), .B(n9735), .ZN(n6650) );
  INV_X1 U8394 ( .A(n6650), .ZN(n6651) );
  OAI21_X1 U8395 ( .B1(n6653), .B2(n6652), .A(n6651), .ZN(n9757) );
  OAI211_X1 U8396 ( .C1(n6655), .C2(n9870), .A(n6654), .B(n9757), .ZN(P1_U3243) );
  INV_X1 U8397 ( .A(n6656), .ZN(n6694) );
  AOI22_X1 U8398 ( .A1(n9842), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9634), .ZN(n6657) );
  OAI21_X1 U8399 ( .B1(n6694), .B2(n9639), .A(n6657), .ZN(P1_U3336) );
  INV_X1 U8400 ( .A(n6668), .ZN(n6667) );
  AOI22_X1 U8401 ( .A1(n6553), .A2(n9260), .B1(n6661), .B2(n7059), .ZN(n6663)
         );
  NAND2_X1 U8402 ( .A1(n6662), .A2(n6663), .ZN(n6712) );
  INV_X1 U8403 ( .A(n6662), .ZN(n6665) );
  INV_X1 U8404 ( .A(n6663), .ZN(n6664) );
  NAND2_X1 U8405 ( .A1(n6665), .A2(n6664), .ZN(n6666) );
  AND2_X1 U8406 ( .A1(n6712), .A2(n6666), .ZN(n6670) );
  NOR2_X1 U8407 ( .A1(n6667), .A2(n6670), .ZN(n6672) );
  NAND2_X1 U8408 ( .A1(n6669), .A2(n6668), .ZN(n6671) );
  NAND2_X1 U8409 ( .A1(n6671), .A2(n6670), .ZN(n6713) );
  INV_X1 U8410 ( .A(n6713), .ZN(n6711) );
  AOI21_X1 U8411 ( .B1(n6672), .B2(n6669), .A(n6711), .ZN(n6678) );
  NOR2_X1 U8412 ( .A1(n9911), .A2(n6673), .ZN(n9903) );
  AOI22_X1 U8413 ( .A1(n8942), .A2(n9259), .B1(n8936), .B2(n9262), .ZN(n6674)
         );
  OAI21_X1 U8414 ( .B1(n6676), .B2(n7062), .A(n6674), .ZN(n6675) );
  AOI21_X1 U8415 ( .B1(n6676), .B2(n9903), .A(n6675), .ZN(n6677) );
  OAI21_X1 U8416 ( .B1(n6678), .B2(n4653), .A(n6677), .ZN(P1_U3235) );
  OR2_X1 U8417 ( .A1(n6684), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6679) );
  INV_X1 U8418 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7383) );
  AOI22_X1 U8419 ( .A1(n7362), .A2(n7383), .B1(P1_REG1_REG_11__SCAN_IN), .B2(
        n7353), .ZN(n6681) );
  NOR2_X1 U8420 ( .A1(n6682), .A2(n6681), .ZN(n7352) );
  AOI21_X1 U8421 ( .B1(n6682), .B2(n6681), .A(n7352), .ZN(n6693) );
  AOI22_X1 U8422 ( .A1(n7362), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n6685), .B2(
        n7353), .ZN(n6686) );
  OAI21_X1 U8423 ( .B1(n6687), .B2(n6686), .A(n7363), .ZN(n6691) );
  NAND2_X1 U8424 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8903) );
  NAND2_X1 U8425 ( .A1(n9859), .A2(n7362), .ZN(n6688) );
  OAI211_X1 U8426 ( .C1(n9870), .C2(n6689), .A(n8903), .B(n6688), .ZN(n6690)
         );
  AOI21_X1 U8427 ( .B1(n6691), .B2(n9857), .A(n6690), .ZN(n6692) );
  OAI21_X1 U8428 ( .B1(n6693), .B2(n9867), .A(n6692), .ZN(P1_U3252) );
  INV_X1 U8429 ( .A(n8381), .ZN(n8376) );
  OAI222_X1 U8430 ( .A1(n4268), .A2(n6695), .B1(n8768), .B2(n6694), .C1(n8376), 
        .C2(n4262), .ZN(P2_U3341) );
  INV_X1 U8431 ( .A(n6696), .ZN(n6700) );
  AND3_X1 U8432 ( .A1(n6908), .A2(n6697), .A3(n7280), .ZN(n6698) );
  OAI21_X1 U8433 ( .B1(n6700), .B2(n6699), .A(n6698), .ZN(n6701) );
  NAND2_X1 U8434 ( .A1(n6701), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6703) );
  INV_X1 U8435 ( .A(n6712), .ZN(n6710) );
  OAI22_X1 U8436 ( .A1(n7263), .A2(n6933), .B1(n7087), .B2(n6658), .ZN(n6704)
         );
  XNOR2_X1 U8437 ( .A(n6704), .B(n8063), .ZN(n6705) );
  AOI22_X1 U8438 ( .A1(n8073), .A2(n9259), .B1(n6661), .B2(n6824), .ZN(n6706)
         );
  NAND2_X1 U8439 ( .A1(n6705), .A2(n6706), .ZN(n6784) );
  INV_X1 U8440 ( .A(n6705), .ZN(n6708) );
  INV_X1 U8441 ( .A(n6706), .ZN(n6707) );
  NAND2_X1 U8442 ( .A1(n6708), .A2(n6707), .ZN(n6709) );
  AND2_X1 U8443 ( .A1(n6784), .A2(n6709), .ZN(n6714) );
  NOR3_X1 U8444 ( .A1(n6711), .A2(n6710), .A3(n6714), .ZN(n6717) );
  NAND2_X1 U8445 ( .A1(n6713), .A2(n6712), .ZN(n6715) );
  NAND2_X1 U8446 ( .A1(n6715), .A2(n6714), .ZN(n6785) );
  INV_X1 U8447 ( .A(n6785), .ZN(n6716) );
  OAI21_X1 U8448 ( .B1(n6717), .B2(n6716), .A(n8935), .ZN(n6722) );
  INV_X1 U8449 ( .A(n8942), .ZN(n8923) );
  AOI21_X1 U8450 ( .B1(n8936), .B2(n9260), .A(n6718), .ZN(n6719) );
  OAI21_X1 U8451 ( .B1(n8923), .B2(n6849), .A(n6719), .ZN(n6720) );
  AOI21_X1 U8452 ( .B1(n8928), .B2(n6824), .A(n6720), .ZN(n6721) );
  OAI211_X1 U8453 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n8926), .A(n6722), .B(
        n6721), .ZN(P1_U3216) );
  XNOR2_X1 U8454 ( .A(n6724), .B(n6723), .ZN(n6728) );
  OAI22_X1 U8455 ( .A1(n7832), .A2(n8249), .B1(n6051), .B2(n8267), .ZN(n6764)
         );
  OR2_X1 U8456 ( .A1(n6725), .A2(n4262), .ZN(n6755) );
  AOI22_X1 U8457 ( .A1(n8285), .A2(n6764), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n6755), .ZN(n6727) );
  NAND2_X1 U8458 ( .A1(n8290), .A2(n9991), .ZN(n6726) );
  OAI211_X1 U8459 ( .C1(n6728), .C2(n8259), .A(n6727), .B(n6726), .ZN(P2_U3239) );
  XNOR2_X1 U8460 ( .A(n6730), .B(n6729), .ZN(n6733) );
  OAI22_X1 U8461 ( .A1(n6750), .A2(n8267), .B1(n6807), .B2(n8249), .ZN(n6777)
         );
  AOI22_X1 U8462 ( .A1(n8290), .A2(n7831), .B1(n8285), .B2(n6777), .ZN(n6732)
         );
  MUX2_X1 U8463 ( .A(n8287), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n6731) );
  OAI211_X1 U8464 ( .C1(n6733), .C2(n8259), .A(n6732), .B(n6731), .ZN(P2_U3220) );
  NAND2_X1 U8465 ( .A1(n6914), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6735) );
  OAI21_X1 U8466 ( .B1(n6914), .B2(P2_REG2_REG_9__SCAN_IN), .A(n6735), .ZN(
        n6736) );
  NOR2_X1 U8467 ( .A1(n4288), .A2(n6736), .ZN(n6913) );
  AOI211_X1 U8468 ( .C1(n4288), .C2(n6736), .A(n6913), .B(n9662), .ZN(n6737)
         );
  INV_X1 U8469 ( .A(n6737), .ZN(n6745) );
  NOR2_X1 U8470 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5711), .ZN(n7130) );
  NAND2_X1 U8471 ( .A1(n6738), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6740) );
  MUX2_X1 U8472 ( .A(n10112), .B(P2_REG1_REG_9__SCAN_IN), .S(n6914), .Z(n6739)
         );
  AOI21_X1 U8473 ( .B1(n6741), .B2(n6740), .A(n6739), .ZN(n6922) );
  AND3_X1 U8474 ( .A1(n6741), .A2(n6740), .A3(n6739), .ZN(n6742) );
  NOR3_X1 U8475 ( .A1(n9941), .A2(n6922), .A3(n6742), .ZN(n6743) );
  AOI211_X1 U8476 ( .C1(n9943), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n7130), .B(
        n6743), .ZN(n6744) );
  OAI211_X1 U8477 ( .C1(n9939), .C2(n6918), .A(n6745), .B(n6744), .ZN(P2_U3254) );
  OAI21_X1 U8478 ( .B1(n6746), .B2(n6748), .A(n6747), .ZN(n6749) );
  NAND2_X1 U8479 ( .A1(n6749), .A2(n8282), .ZN(n6753) );
  OAI22_X1 U8480 ( .A1(n6751), .A2(n8267), .B1(n6750), .B2(n8249), .ZN(n7093)
         );
  AOI22_X1 U8481 ( .A1(n8285), .A2(n7093), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n6755), .ZN(n6752) );
  OAI211_X1 U8482 ( .C1(n6052), .C2(n8278), .A(n6753), .B(n6752), .ZN(P2_U3224) );
  AOI21_X1 U8483 ( .B1(n8282), .B2(n6754), .A(n8290), .ZN(n6759) );
  INV_X1 U8484 ( .A(n7096), .ZN(n10028) );
  NOR2_X1 U8485 ( .A1(n6051), .A2(n8249), .ZN(n9998) );
  AOI22_X1 U8486 ( .A1(n8285), .A2(n9998), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n6755), .ZN(n6758) );
  NAND2_X1 U8487 ( .A1(n6756), .A2(n10028), .ZN(n7949) );
  INV_X1 U8488 ( .A(n7949), .ZN(n7822) );
  NAND2_X1 U8489 ( .A1(n8244), .A2(n7822), .ZN(n6757) );
  OAI211_X1 U8490 ( .C1(n6759), .C2(n10028), .A(n6758), .B(n6757), .ZN(
        P2_U3234) );
  NAND2_X1 U8491 ( .A1(n7947), .A2(n8480), .ZN(n6760) );
  OR2_X1 U8492 ( .A1(n7991), .A2(n6760), .ZN(n10073) );
  NAND2_X1 U8493 ( .A1(n9955), .A2(n10073), .ZN(n10097) );
  OAI21_X1 U8494 ( .B1(n6762), .B2(n7948), .A(n6761), .ZN(n9994) );
  AOI211_X1 U8495 ( .C1(n9991), .C2(n10034), .A(n10086), .B(n6775), .ZN(n9992)
         );
  XNOR2_X1 U8496 ( .A(n6763), .B(n7948), .ZN(n6765) );
  AOI21_X1 U8497 ( .B1(n6765), .B2(n9968), .A(n6764), .ZN(n9997) );
  INV_X1 U8498 ( .A(n9997), .ZN(n6766) );
  AOI211_X1 U8499 ( .C1(n10097), .C2(n9994), .A(n9992), .B(n6766), .ZN(n6889)
         );
  OR2_X1 U8500 ( .A1(n6832), .A2(n6767), .ZN(n6768) );
  NOR2_X1 U8501 ( .A1(n6834), .A2(n6768), .ZN(n6769) );
  AND2_X1 U8502 ( .A1(n6836), .A2(n6769), .ZN(n6771) );
  INV_X1 U8503 ( .A(n6770), .ZN(n6837) );
  AND2_X2 U8504 ( .A1(n6771), .A2(n6837), .ZN(n10120) );
  AOI22_X1 U8505 ( .A1(n8670), .A2(n9991), .B1(n10117), .B2(
        P2_REG1_REG_2__SCAN_IN), .ZN(n6772) );
  OAI21_X1 U8506 ( .B1(n6889), .B2(n10117), .A(n6772), .ZN(P2_U3522) );
  OAI21_X1 U8507 ( .B1(n6774), .B2(n7954), .A(n6773), .ZN(n7249) );
  OR2_X1 U8508 ( .A1(n6775), .A2(n7247), .ZN(n6776) );
  AND3_X1 U8509 ( .A1(n6861), .A2(n10049), .A3(n6776), .ZN(n7244) );
  XNOR2_X1 U8510 ( .A(n6863), .B(n7954), .ZN(n6779) );
  INV_X1 U8511 ( .A(n9968), .ZN(n10000) );
  INV_X1 U8512 ( .A(n6777), .ZN(n6778) );
  OAI21_X1 U8513 ( .B1(n6779), .B2(n10000), .A(n6778), .ZN(n7242) );
  AOI211_X1 U8514 ( .C1(n10097), .C2(n7249), .A(n7244), .B(n7242), .ZN(n6840)
         );
  AOI22_X1 U8515 ( .A1(n8670), .A2(n7831), .B1(n10117), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n6780) );
  OAI21_X1 U8516 ( .B1(n6840), .B2(n10117), .A(n6780), .ZN(P2_U3523) );
  NAND2_X1 U8517 ( .A1(n8303), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6781) );
  OAI21_X1 U8518 ( .B1(n6782), .B2(n8303), .A(n6781), .ZN(P2_U3581) );
  OAI22_X1 U8519 ( .A1(n7263), .A2(n6849), .B1(n9912), .B2(n6658), .ZN(n6783)
         );
  XNOR2_X1 U8520 ( .A(n6783), .B(n8096), .ZN(n7020) );
  AOI22_X1 U8521 ( .A1(n8073), .A2(n9258), .B1(n4269), .B2(n6947), .ZN(n7021)
         );
  XNOR2_X1 U8522 ( .A(n7020), .B(n7021), .ZN(n6787) );
  NAND2_X1 U8523 ( .A1(n6785), .A2(n6784), .ZN(n6786) );
  NAND2_X1 U8524 ( .A1(n6786), .A2(n6787), .ZN(n7024) );
  OAI21_X1 U8525 ( .B1(n6787), .B2(n6786), .A(n7024), .ZN(n6788) );
  NAND2_X1 U8526 ( .A1(n6788), .A2(n8935), .ZN(n6792) );
  AND2_X1 U8527 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9756) );
  AOI21_X1 U8528 ( .B1(n8936), .B2(n9259), .A(n9756), .ZN(n6789) );
  OAI21_X1 U8529 ( .B1(n8923), .B2(n7156), .A(n6789), .ZN(n6790) );
  AOI21_X1 U8530 ( .B1(n8928), .B2(n6947), .A(n6790), .ZN(n6791) );
  OAI211_X1 U8531 ( .C1(n8926), .C2(n6938), .A(n6792), .B(n6791), .ZN(P1_U3228) );
  NAND2_X1 U8532 ( .A1(n9261), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6793) );
  OAI21_X1 U8533 ( .B1(n9321), .B2(n9261), .A(n6793), .ZN(P1_U3584) );
  INV_X1 U8534 ( .A(n6794), .ZN(n6795) );
  AOI21_X1 U8535 ( .B1(n6797), .B2(n6796), .A(n6795), .ZN(n6805) );
  INV_X1 U8536 ( .A(n9983), .ZN(n6802) );
  OR2_X1 U8537 ( .A1(n6798), .A2(n8249), .ZN(n6800) );
  NAND2_X1 U8538 ( .A1(n8322), .A2(n8251), .ZN(n6799) );
  NAND2_X1 U8539 ( .A1(n6800), .A2(n6799), .ZN(n6866) );
  AOI22_X1 U8540 ( .A1(n8285), .A2(n6866), .B1(P2_REG3_REG_4__SCAN_IN), .B2(
        P2_U3152), .ZN(n6801) );
  OAI21_X1 U8541 ( .B1(n6802), .B2(n8287), .A(n6801), .ZN(n6803) );
  AOI21_X1 U8542 ( .B1(n8290), .B2(n9984), .A(n6803), .ZN(n6804) );
  OAI21_X1 U8543 ( .B1(n6805), .B2(n8259), .A(n6804), .ZN(P2_U3232) );
  XNOR2_X1 U8544 ( .A(n6952), .B(n6951), .ZN(n6813) );
  INV_X1 U8545 ( .A(n6806), .ZN(n7073) );
  OR2_X1 U8546 ( .A1(n6807), .A2(n8267), .ZN(n6809) );
  OR2_X1 U8547 ( .A1(n6871), .A2(n8249), .ZN(n6808) );
  NAND2_X1 U8548 ( .A1(n6809), .A2(n6808), .ZN(n7071) );
  AOI22_X1 U8549 ( .A1(n8285), .A2(n7071), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        n4262), .ZN(n6810) );
  OAI21_X1 U8550 ( .B1(n7073), .B2(n8287), .A(n6810), .ZN(n6811) );
  AOI21_X1 U8551 ( .B1(n8290), .B2(n7079), .A(n6811), .ZN(n6812) );
  OAI21_X1 U8552 ( .B1(n6813), .B2(n8259), .A(n6812), .ZN(P2_U3229) );
  INV_X1 U8553 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6815) );
  INV_X1 U8554 ( .A(n6814), .ZN(n6816) );
  INV_X1 U8555 ( .A(n8387), .ZN(n8396) );
  OAI222_X1 U8556 ( .A1(n4268), .A2(n6815), .B1(n8768), .B2(n6816), .C1(
        P2_U3152), .C2(n8396), .ZN(P2_U3340) );
  INV_X1 U8557 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6817) );
  INV_X1 U8558 ( .A(n9858), .ZN(n9283) );
  OAI222_X1 U8559 ( .A1(n9641), .A2(n6817), .B1(n9645), .B2(n6816), .C1(
        P1_U3084), .C2(n9283), .ZN(P1_U3335) );
  OAI21_X1 U8560 ( .B1(n6818), .B2(n9089), .A(n6842), .ZN(n7089) );
  INV_X1 U8561 ( .A(n7089), .ZN(n6826) );
  INV_X1 U8562 ( .A(n6819), .ZN(n9688) );
  OAI22_X1 U8563 ( .A1(n6898), .A2(n9682), .B1(n9681), .B2(n6849), .ZN(n6822)
         );
  XNOR2_X1 U8564 ( .A(n8954), .B(n9089), .ZN(n6820) );
  NOR2_X1 U8565 ( .A1(n6820), .A2(n9510), .ZN(n6821) );
  AOI211_X1 U8566 ( .C1(n9688), .C2(n7089), .A(n6822), .B(n6821), .ZN(n7091)
         );
  INV_X1 U8567 ( .A(n6823), .ZN(n6942) );
  AOI21_X1 U8568 ( .B1(n6824), .B2(n7058), .A(n6942), .ZN(n7083) );
  AOI22_X1 U8569 ( .A1(n7083), .A2(n9713), .B1(n9606), .B2(n6824), .ZN(n6825)
         );
  OAI211_X1 U8570 ( .C1(n6826), .C2(n9609), .A(n7091), .B(n6825), .ZN(n6828)
         );
  NAND2_X1 U8571 ( .A1(n6828), .A2(n9935), .ZN(n6827) );
  OAI21_X1 U8572 ( .B1(n9935), .B2(n6179), .A(n6827), .ZN(P1_U3526) );
  INV_X1 U8573 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6830) );
  NAND2_X1 U8574 ( .A1(n6828), .A2(n9929), .ZN(n6829) );
  OAI21_X1 U8575 ( .B1(n9929), .B2(n6830), .A(n6829), .ZN(P1_U3463) );
  NAND2_X1 U8576 ( .A1(n6832), .A2(n6831), .ZN(n6833) );
  NOR2_X1 U8577 ( .A1(n6834), .A2(n6833), .ZN(n6835) );
  AND2_X1 U8578 ( .A1(n6836), .A2(n6835), .ZN(n6838) );
  AND2_X2 U8579 ( .A1(n6838), .A2(n6837), .ZN(n10101) );
  AOI22_X1 U8580 ( .A1(n8748), .A2(n7831), .B1(n10099), .B2(
        P2_REG0_REG_3__SCAN_IN), .ZN(n6839) );
  OAI21_X1 U8581 ( .B1(n6840), .B2(n10099), .A(n6839), .ZN(P2_U3460) );
  INV_X1 U8582 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6855) );
  NAND2_X1 U8583 ( .A1(n6842), .A2(n6841), .ZN(n6931) );
  NAND2_X1 U8584 ( .A1(n6931), .A2(n9094), .ZN(n6930) );
  NAND2_X1 U8585 ( .A1(n6930), .A2(n6843), .ZN(n6845) );
  NAND2_X1 U8586 ( .A1(n6845), .A2(n6848), .ZN(n6846) );
  NAND2_X1 U8587 ( .A1(n6847), .A2(n6846), .ZN(n9883) );
  XNOR2_X1 U8588 ( .A(n7152), .B(n6844), .ZN(n6851) );
  OAI22_X1 U8589 ( .A1(n6849), .A2(n9682), .B1(n9681), .B2(n7262), .ZN(n6850)
         );
  AOI21_X1 U8590 ( .B1(n6851), .B2(n9685), .A(n6850), .ZN(n9881) );
  OR2_X1 U8591 ( .A1(n6940), .A2(n9874), .ZN(n6852) );
  AND3_X1 U8592 ( .A1(n7147), .A2(n9713), .A3(n6852), .ZN(n9879) );
  AOI21_X1 U8593 ( .B1(n9606), .B2(n7038), .A(n9879), .ZN(n6853) );
  OAI211_X1 U8594 ( .C1(n9883), .C2(n9597), .A(n9881), .B(n6853), .ZN(n6856)
         );
  NAND2_X1 U8595 ( .A1(n6856), .A2(n9929), .ZN(n6854) );
  OAI21_X1 U8596 ( .B1(n9929), .B2(n6855), .A(n6854), .ZN(P1_U3469) );
  NAND2_X1 U8597 ( .A1(n6856), .A2(n9935), .ZN(n6857) );
  OAI21_X1 U8598 ( .B1(n9935), .B2(n6172), .A(n6857), .ZN(P1_U3528) );
  OAI21_X1 U8599 ( .B1(n6859), .B2(n6097), .A(n6858), .ZN(n9986) );
  INV_X1 U8600 ( .A(n7075), .ZN(n6860) );
  AOI211_X1 U8601 ( .C1(n9984), .C2(n6861), .A(n10086), .B(n6860), .ZN(n9985)
         );
  INV_X1 U8602 ( .A(n7954), .ZN(n6862) );
  NAND2_X1 U8603 ( .A1(n6863), .A2(n6862), .ZN(n6864) );
  NAND2_X1 U8604 ( .A1(n6864), .A2(n7809), .ZN(n6865) );
  AOI21_X1 U8605 ( .B1(n6865), .B2(n6097), .A(n10000), .ZN(n6867) );
  OR2_X1 U8606 ( .A1(n6865), .A2(n6097), .ZN(n7069) );
  AOI21_X1 U8607 ( .B1(n6867), .B2(n7069), .A(n6866), .ZN(n9989) );
  INV_X1 U8608 ( .A(n9989), .ZN(n6868) );
  AOI211_X1 U8609 ( .C1(n10097), .C2(n9986), .A(n9985), .B(n6868), .ZN(n6884)
         );
  AOI22_X1 U8610 ( .A1(n8670), .A2(n9984), .B1(n10117), .B2(
        P2_REG1_REG_4__SCAN_IN), .ZN(n6869) );
  OAI21_X1 U8611 ( .B1(n6884), .B2(n10117), .A(n6869), .ZN(P2_U3524) );
  XNOR2_X1 U8612 ( .A(n4357), .B(n6870), .ZN(n6879) );
  INV_X1 U8613 ( .A(n9974), .ZN(n6876) );
  OR2_X1 U8614 ( .A1(n7129), .A2(n8249), .ZN(n6873) );
  OR2_X1 U8615 ( .A1(n6871), .A2(n8267), .ZN(n6872) );
  NAND2_X1 U8616 ( .A1(n6873), .A2(n6872), .ZN(n9971) );
  AOI21_X1 U8617 ( .B1(n8285), .B2(n9971), .A(n6874), .ZN(n6875) );
  OAI21_X1 U8618 ( .B1(n6876), .B2(n8287), .A(n6875), .ZN(n6877) );
  AOI21_X1 U8619 ( .B1(n8290), .B2(n9975), .A(n6877), .ZN(n6878) );
  OAI21_X1 U8620 ( .B1(n6879), .B2(n8259), .A(n6878), .ZN(P2_U3215) );
  INV_X1 U8621 ( .A(n8748), .ZN(n8755) );
  INV_X1 U8622 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n6880) );
  OAI22_X1 U8623 ( .A1(n8755), .A2(n6881), .B1(n10101), .B2(n6880), .ZN(n6882)
         );
  INV_X1 U8624 ( .A(n6882), .ZN(n6883) );
  OAI21_X1 U8625 ( .B1(n6884), .B2(n10099), .A(n6883), .ZN(P2_U3463) );
  INV_X1 U8626 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6885) );
  OAI22_X1 U8627 ( .A1(n8755), .A2(n6886), .B1(n10101), .B2(n6885), .ZN(n6887)
         );
  INV_X1 U8628 ( .A(n6887), .ZN(n6888) );
  OAI21_X1 U8629 ( .B1(n6889), .B2(n10099), .A(n6888), .ZN(P2_U3457) );
  INV_X1 U8630 ( .A(n6890), .ZN(n8136) );
  OAI222_X1 U8631 ( .A1(n9641), .A2(n6891), .B1(n9639), .B2(n8136), .C1(n9878), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  INV_X1 U8632 ( .A(n6892), .ZN(n6893) );
  AOI21_X1 U8633 ( .B1(n9093), .B2(n6894), .A(n6893), .ZN(n9901) );
  XOR2_X1 U8634 ( .A(n9093), .B(n6895), .Z(n6896) );
  OAI222_X1 U8635 ( .A1(n9681), .A2(n6898), .B1(n9682), .B2(n6897), .C1(n6896), 
        .C2(n9510), .ZN(n9899) );
  INV_X1 U8636 ( .A(n9895), .ZN(n9629) );
  INV_X1 U8637 ( .A(n7056), .ZN(n6899) );
  AOI211_X1 U8638 ( .C1(n6900), .C2(n6901), .A(n9921), .B(n6899), .ZN(n9896)
         );
  INV_X1 U8639 ( .A(n9873), .ZN(n6937) );
  AOI22_X1 U8640 ( .A1(n9896), .A2(n9878), .B1(n6937), .B2(n6901), .ZN(n6902)
         );
  OAI21_X1 U8641 ( .B1(n6903), .B2(n9876), .A(n6902), .ZN(n6904) );
  AOI211_X1 U8642 ( .C1(n9901), .C2(n9688), .A(n9899), .B(n6904), .ZN(n6912)
         );
  INV_X1 U8643 ( .A(n6905), .ZN(n6906) );
  NAND2_X1 U8644 ( .A1(n6906), .A2(n9895), .ZN(n9893) );
  NOR2_X1 U8645 ( .A1(n6907), .A2(n9893), .ZN(n6909) );
  NAND2_X1 U8646 ( .A1(n6909), .A2(n6908), .ZN(n6996) );
  NAND2_X2 U8647 ( .A1(n6996), .A2(n9876), .ZN(n9885) );
  NOR2_X1 U8648 ( .A1(n6417), .A2(n9878), .ZN(n6910) );
  NAND2_X1 U8649 ( .A1(n9885), .A2(n6910), .ZN(n7605) );
  INV_X1 U8650 ( .A(n7605), .ZN(n9699) );
  AOI22_X1 U8651 ( .A1(n9901), .A2(n9699), .B1(P1_REG2_REG_1__SCAN_IN), .B2(
        n9887), .ZN(n6911) );
  OAI21_X1 U8652 ( .B1(n6912), .B2(n9692), .A(n6911), .ZN(P1_U3290) );
  XNOR2_X1 U8653 ( .A(n7009), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n6915) );
  AOI211_X1 U8654 ( .C1(n6916), .C2(n6915), .A(n7008), .B(n9662), .ZN(n6917)
         );
  INV_X1 U8655 ( .A(n6917), .ZN(n6928) );
  NOR2_X1 U8656 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7120), .ZN(n6926) );
  NOR2_X1 U8657 ( .A1(n6918), .A2(n10112), .ZN(n6921) );
  INV_X1 U8658 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6919) );
  MUX2_X1 U8659 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n6919), .S(n7009), .Z(n6920)
         );
  OAI21_X1 U8660 ( .B1(n6922), .B2(n6921), .A(n6920), .ZN(n7003) );
  INV_X1 U8661 ( .A(n7003), .ZN(n6924) );
  NOR3_X1 U8662 ( .A1(n6922), .A2(n6921), .A3(n6920), .ZN(n6923) );
  NOR3_X1 U8663 ( .A1(n9941), .A2(n6924), .A3(n6923), .ZN(n6925) );
  AOI211_X1 U8664 ( .C1(n9943), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n6926), .B(
        n6925), .ZN(n6927) );
  OAI211_X1 U8665 ( .C1(n9939), .C2(n6929), .A(n6928), .B(n6927), .ZN(P2_U3255) );
  OAI21_X1 U8666 ( .B1(n6931), .B2(n9094), .A(n6930), .ZN(n9916) );
  INV_X1 U8667 ( .A(n9916), .ZN(n6950) );
  XNOR2_X1 U8668 ( .A(n6932), .B(n9094), .ZN(n6936) );
  OAI22_X1 U8669 ( .A1(n6933), .A2(n9682), .B1(n9681), .B2(n7156), .ZN(n6934)
         );
  AOI21_X1 U8670 ( .B1(n9916), .B2(n9688), .A(n6934), .ZN(n6935) );
  OAI21_X1 U8671 ( .B1(n9510), .B2(n6936), .A(n6935), .ZN(n9914) );
  NAND2_X1 U8672 ( .A1(n9914), .A2(n9885), .ZN(n6949) );
  OAI22_X1 U8673 ( .A1(n9885), .A2(n6939), .B1(n6938), .B2(n9876), .ZN(n6946)
         );
  INV_X1 U8674 ( .A(n6940), .ZN(n6941) );
  OAI21_X1 U8675 ( .B1(n9912), .B2(n6942), .A(n6941), .ZN(n9913) );
  INV_X1 U8676 ( .A(n6415), .ZN(n9235) );
  NOR2_X1 U8677 ( .A1(n6943), .A2(n9235), .ZN(n6944) );
  NAND2_X1 U8678 ( .A1(n9885), .A2(n6944), .ZN(n9308) );
  NOR2_X1 U8679 ( .A1(n9913), .A2(n9308), .ZN(n6945) );
  AOI211_X1 U8680 ( .C1(n9693), .C2(n6947), .A(n6946), .B(n6945), .ZN(n6948)
         );
  OAI211_X1 U8681 ( .C1(n6950), .C2(n7605), .A(n6949), .B(n6948), .ZN(P1_U3287) );
  NOR2_X1 U8682 ( .A1(n6952), .A2(n6951), .ZN(n6955) );
  NOR2_X1 U8683 ( .A1(n6955), .A2(n6953), .ZN(n6957) );
  OR2_X1 U8684 ( .A1(n6955), .A2(n6954), .ZN(n6956) );
  OAI21_X1 U8685 ( .B1(n6958), .B2(n6957), .A(n6956), .ZN(n6959) );
  NAND2_X1 U8686 ( .A1(n6959), .A2(n8282), .ZN(n6963) );
  AOI22_X1 U8687 ( .A1(n8251), .A2(n8320), .B1(n8318), .B2(n8269), .ZN(n8594)
         );
  OAI21_X1 U8688 ( .B1(n8594), .B2(n8273), .A(n6960), .ZN(n6961) );
  AOI21_X1 U8689 ( .B1(n8597), .B2(n8275), .A(n6961), .ZN(n6962) );
  OAI211_X1 U8690 ( .C1(n6964), .C2(n8278), .A(n6963), .B(n6962), .ZN(P2_U3241) );
  INV_X1 U8691 ( .A(n6965), .ZN(n6981) );
  OAI222_X1 U8692 ( .A1(n9645), .A2(n6981), .B1(P1_U3084), .B2(n9232), .C1(
        n6966), .C2(n9641), .ZN(P1_U3333) );
  XNOR2_X1 U8693 ( .A(n6968), .B(n6967), .ZN(n6979) );
  OR2_X1 U8694 ( .A1(n6969), .A2(n8249), .ZN(n6972) );
  OR2_X1 U8695 ( .A1(n6970), .A2(n8267), .ZN(n6971) );
  NAND2_X1 U8696 ( .A1(n6972), .A2(n6971), .ZN(n7168) );
  INV_X1 U8697 ( .A(n7168), .ZN(n6976) );
  NAND2_X1 U8698 ( .A1(n8275), .A2(n6973), .ZN(n6975) );
  OAI211_X1 U8699 ( .C1(n8273), .C2(n6976), .A(n6975), .B(n6974), .ZN(n6977)
         );
  AOI21_X1 U8700 ( .B1(n8290), .B2(n7176), .A(n6977), .ZN(n6978) );
  OAI21_X1 U8701 ( .B1(n6979), .B2(n8259), .A(n6978), .ZN(P2_U3223) );
  OAI222_X1 U8702 ( .A1(n4262), .A2(n7947), .B1(n8768), .B2(n6981), .C1(n6980), 
        .C2(n4268), .ZN(P2_U3338) );
  INV_X1 U8703 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6982) );
  OAI22_X1 U8704 ( .A1(n9885), .A2(n6983), .B1(n6982), .B2(n9876), .ZN(n6986)
         );
  AOI21_X1 U8705 ( .B1(n9519), .B2(n9308), .A(n6984), .ZN(n6985) );
  AOI211_X1 U8706 ( .C1(n9885), .C2(n6987), .A(n6986), .B(n6985), .ZN(n6988)
         );
  INV_X1 U8707 ( .A(n6988), .ZN(P1_U3291) );
  OAI21_X1 U8708 ( .B1(n6990), .B2(n9088), .A(n6989), .ZN(n6991) );
  INV_X1 U8709 ( .A(n6991), .ZN(n7139) );
  AND2_X1 U8710 ( .A1(n8096), .A2(n9238), .ZN(n9872) );
  NAND2_X1 U8711 ( .A1(n9872), .A2(n9885), .ZN(n9524) );
  AOI21_X1 U8712 ( .B1(n9088), .B2(n6992), .A(n4361), .ZN(n6993) );
  OAI222_X1 U8713 ( .A1(n9681), .A2(n6994), .B1(n9682), .B2(n7262), .C1(n9510), 
        .C2(n6993), .ZN(n7136) );
  NAND2_X1 U8714 ( .A1(n7136), .A2(n9885), .ZN(n7000) );
  INV_X1 U8715 ( .A(n7043), .ZN(n6995) );
  AOI211_X1 U8716 ( .C1(n7350), .C2(n7149), .A(n9921), .B(n6995), .ZN(n7137)
         );
  NOR2_X1 U8717 ( .A1(n6996), .A2(n9434), .ZN(n9698) );
  NOR2_X1 U8718 ( .A1(n9519), .A2(n4537), .ZN(n6998) );
  OAI22_X1 U8719 ( .A1(n9885), .A2(n4457), .B1(n7338), .B2(n9876), .ZN(n6997)
         );
  AOI211_X1 U8720 ( .C1(n7137), .C2(n9698), .A(n6998), .B(n6997), .ZN(n6999)
         );
  OAI211_X1 U8721 ( .C1(n7139), .C2(n9524), .A(n7000), .B(n6999), .ZN(P1_U3284) );
  NAND2_X1 U8722 ( .A1(n7009), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7002) );
  INV_X1 U8723 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10115) );
  MUX2_X1 U8724 ( .A(n10115), .B(P2_REG1_REG_11__SCAN_IN), .S(n7212), .Z(n7001) );
  AOI21_X1 U8725 ( .B1(n7003), .B2(n7002), .A(n7001), .ZN(n7204) );
  NAND3_X1 U8726 ( .A1(n7003), .A2(n7002), .A3(n7001), .ZN(n7004) );
  NAND2_X1 U8727 ( .A1(n9936), .A2(n7004), .ZN(n7017) );
  NOR2_X1 U8728 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5743), .ZN(n7007) );
  NOR2_X1 U8729 ( .A1(n9939), .A2(n7005), .ZN(n7006) );
  AOI211_X1 U8730 ( .C1(n9943), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n7007), .B(
        n7006), .ZN(n7016) );
  INV_X1 U8731 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7010) );
  MUX2_X1 U8732 ( .A(n7010), .B(P2_REG2_REG_11__SCAN_IN), .S(n7212), .Z(n7011)
         );
  INV_X1 U8733 ( .A(n7011), .ZN(n7012) );
  OAI21_X1 U8734 ( .B1(n7013), .B2(n7012), .A(n7211), .ZN(n7014) );
  NAND2_X1 U8735 ( .A1(n9937), .A2(n7014), .ZN(n7015) );
  OAI211_X1 U8736 ( .C1(n7204), .C2(n7017), .A(n7016), .B(n7015), .ZN(P2_U3256) );
  INV_X1 U8737 ( .A(n7018), .ZN(n7067) );
  OAI222_X1 U8738 ( .A1(n4268), .A2(n7019), .B1(n8768), .B2(n7067), .C1(n5579), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  OAI22_X1 U8739 ( .A1(n6660), .A2(n7156), .B1(n7263), .B2(n9874), .ZN(n7033)
         );
  INV_X1 U8740 ( .A(n7020), .ZN(n7022) );
  NAND2_X1 U8741 ( .A1(n7022), .A2(n7021), .ZN(n7023) );
  NAND2_X1 U8742 ( .A1(n7024), .A2(n7023), .ZN(n7029) );
  INV_X1 U8743 ( .A(n7029), .ZN(n7027) );
  OAI22_X1 U8744 ( .A1(n7263), .A2(n7156), .B1(n9874), .B2(n6658), .ZN(n7025)
         );
  XNOR2_X1 U8745 ( .A(n7025), .B(n8063), .ZN(n7028) );
  INV_X1 U8746 ( .A(n7028), .ZN(n7026) );
  NAND2_X1 U8747 ( .A1(n7027), .A2(n7026), .ZN(n7030) );
  INV_X1 U8748 ( .A(n7033), .ZN(n7031) );
  AOI21_X1 U8749 ( .B1(n7033), .B2(n7032), .A(n4359), .ZN(n7040) );
  NOR2_X1 U8750 ( .A1(n8926), .A2(n9875), .ZN(n7037) );
  NAND2_X1 U8751 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9770) );
  INV_X1 U8752 ( .A(n9770), .ZN(n7034) );
  AOI21_X1 U8753 ( .B1(n8936), .B2(n9258), .A(n7034), .ZN(n7035) );
  OAI21_X1 U8754 ( .B1(n8923), .B2(n7262), .A(n7035), .ZN(n7036) );
  AOI211_X1 U8755 ( .C1(n8928), .C2(n7038), .A(n7037), .B(n7036), .ZN(n7039)
         );
  OAI21_X1 U8756 ( .B1(n7040), .B2(n4653), .A(n7039), .ZN(P1_U3225) );
  OAI21_X1 U8757 ( .B1(n7042), .B2(n5136), .A(n7041), .ZN(n7236) );
  AOI211_X1 U8758 ( .C1(n7540), .C2(n7043), .A(n9921), .B(n7110), .ZN(n7234)
         );
  INV_X1 U8759 ( .A(n7540), .ZN(n7044) );
  NOR2_X1 U8760 ( .A1(n9519), .A2(n7044), .ZN(n7047) );
  OAI22_X1 U8761 ( .A1(n9885), .A2(n7045), .B1(n7531), .B2(n9876), .ZN(n7046)
         );
  AOI211_X1 U8762 ( .C1(n7234), .C2(n9698), .A(n7047), .B(n7046), .ZN(n7051)
         );
  XOR2_X1 U8763 ( .A(n9098), .B(n7048), .Z(n7049) );
  OAI222_X1 U8764 ( .A1(n9681), .A2(n9683), .B1(n9682), .B2(n7157), .C1(n7049), 
        .C2(n9510), .ZN(n7233) );
  NAND2_X1 U8765 ( .A1(n7233), .A2(n9885), .ZN(n7050) );
  OAI211_X1 U8766 ( .C1(n7236), .C2(n9524), .A(n7051), .B(n7050), .ZN(P1_U3283) );
  INV_X1 U8767 ( .A(n9885), .ZN(n9887) );
  INV_X1 U8768 ( .A(n7054), .ZN(n9091) );
  XNOR2_X1 U8769 ( .A(n9198), .B(n9091), .ZN(n7052) );
  AOI222_X1 U8770 ( .A1(n9685), .A2(n7052), .B1(n9262), .B2(n9497), .C1(n9259), 
        .C2(n9499), .ZN(n9906) );
  INV_X1 U8771 ( .A(n9524), .ZN(n9483) );
  OAI21_X1 U8772 ( .B1(n7055), .B2(n7054), .A(n7053), .ZN(n9909) );
  NAND2_X1 U8773 ( .A1(n7056), .A2(n7059), .ZN(n7057) );
  NAND2_X1 U8774 ( .A1(n7058), .A2(n7057), .ZN(n9905) );
  NOR2_X1 U8775 ( .A1(n9308), .A2(n9905), .ZN(n7064) );
  NAND2_X1 U8776 ( .A1(n9693), .A2(n7059), .ZN(n7061) );
  NAND2_X1 U8777 ( .A1(n9887), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7060) );
  OAI211_X1 U8778 ( .C1(n9876), .C2(n7062), .A(n7061), .B(n7060), .ZN(n7063)
         );
  AOI211_X1 U8779 ( .C1(n9483), .C2(n9909), .A(n7064), .B(n7063), .ZN(n7065)
         );
  OAI21_X1 U8780 ( .B1(n9887), .B2(n9906), .A(n7065), .ZN(P1_U3289) );
  OAI222_X1 U8781 ( .A1(n9639), .A2(n7067), .B1(P1_U3084), .B2(n5464), .C1(
        n7066), .C2(n9641), .ZN(P1_U3332) );
  NAND2_X1 U8782 ( .A1(n7069), .A2(n7068), .ZN(n7070) );
  XNOR2_X1 U8783 ( .A(n7070), .B(n7953), .ZN(n7072) );
  AOI21_X1 U8784 ( .B1(n7072), .B2(n9968), .A(n7071), .ZN(n10042) );
  INV_X1 U8785 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7074) );
  OAI22_X1 U8786 ( .A1(n10009), .A2(n7074), .B1(n7073), .B2(n8479), .ZN(n7078)
         );
  AOI21_X1 U8787 ( .B1(n7075), .B2(n7079), .A(n10086), .ZN(n7076) );
  NAND2_X1 U8788 ( .A1(n7076), .A2(n8601), .ZN(n10041) );
  NOR2_X1 U8789 ( .A1(n10041), .A2(n8588), .ZN(n7077) );
  AOI211_X1 U8790 ( .C1(n9990), .C2(n7079), .A(n7078), .B(n7077), .ZN(n7082)
         );
  XNOR2_X1 U8791 ( .A(n7080), .B(n7953), .ZN(n10045) );
  NAND2_X1 U8792 ( .A1(n10045), .A2(n10006), .ZN(n7081) );
  OAI211_X1 U8793 ( .C1(n10042), .C2(n10011), .A(n7082), .B(n7081), .ZN(
        P2_U3291) );
  NAND2_X1 U8794 ( .A1(n7083), .A2(n9504), .ZN(n7086) );
  INV_X1 U8795 ( .A(n9885), .ZN(n9692) );
  INV_X1 U8796 ( .A(n9876), .ZN(n9690) );
  AOI22_X1 U8797 ( .A1(n9692), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9690), .B2(
        n7084), .ZN(n7085) );
  OAI211_X1 U8798 ( .C1(n7087), .C2(n9519), .A(n7086), .B(n7085), .ZN(n7088)
         );
  AOI21_X1 U8799 ( .B1(n9699), .B2(n7089), .A(n7088), .ZN(n7090) );
  OAI21_X1 U8800 ( .B1(n7091), .B2(n9692), .A(n7090), .ZN(P1_U3288) );
  XNOR2_X1 U8801 ( .A(n7092), .B(n7950), .ZN(n7094) );
  AOI21_X1 U8802 ( .B1(n7094), .B2(n9968), .A(n7093), .ZN(n10036) );
  INV_X1 U8803 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9648) );
  OR2_X1 U8804 ( .A1(n7095), .A2(n5643), .ZN(n10003) );
  INV_X1 U8805 ( .A(n10003), .ZN(n8602) );
  NAND2_X1 U8806 ( .A1(n7101), .A2(n7096), .ZN(n10033) );
  NAND3_X1 U8807 ( .A1(n8602), .A2(n10034), .A3(n10033), .ZN(n7097) );
  OAI21_X1 U8808 ( .B1(n8479), .B2(n9648), .A(n7097), .ZN(n7098) );
  AOI21_X1 U8809 ( .B1(P2_REG2_REG_1__SCAN_IN), .B2(n10011), .A(n7098), .ZN(
        n7103) );
  OAI21_X1 U8810 ( .B1(n7092), .B2(n7100), .A(n7099), .ZN(n10039) );
  AOI22_X1 U8811 ( .A1(n9990), .A2(n7101), .B1(n10006), .B2(n10039), .ZN(n7102) );
  OAI211_X1 U8812 ( .C1(n10011), .C2(n10036), .A(n7103), .B(n7102), .ZN(
        P2_U3295) );
  AND2_X1 U8813 ( .A1(n8974), .A2(n8972), .ZN(n9099) );
  XNOR2_X1 U8814 ( .A(n7104), .B(n9099), .ZN(n7194) );
  NAND2_X1 U8815 ( .A1(n7105), .A2(n8971), .ZN(n7106) );
  XNOR2_X1 U8816 ( .A(n7106), .B(n9099), .ZN(n7108) );
  AOI22_X1 U8817 ( .A1(n9497), .A2(n9254), .B1(n9499), .B2(n9252), .ZN(n7107)
         );
  OAI21_X1 U8818 ( .B1(n7108), .B2(n9510), .A(n7107), .ZN(n7109) );
  AOI21_X1 U8819 ( .B1(n7194), .B2(n9688), .A(n7109), .ZN(n7197) );
  INV_X1 U8820 ( .A(n7110), .ZN(n7112) );
  INV_X1 U8821 ( .A(n7111), .ZN(n9696) );
  AOI21_X1 U8822 ( .B1(n7494), .B2(n7112), .A(n9696), .ZN(n7195) );
  NAND2_X1 U8823 ( .A1(n7195), .A2(n9504), .ZN(n7115) );
  INV_X1 U8824 ( .A(n7113), .ZN(n7514) );
  AOI22_X1 U8825 ( .A1(n9692), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7514), .B2(
        n9690), .ZN(n7114) );
  OAI211_X1 U8826 ( .C1(n7517), .C2(n9519), .A(n7115), .B(n7114), .ZN(n7116)
         );
  AOI21_X1 U8827 ( .B1(n7194), .B2(n9699), .A(n7116), .ZN(n7117) );
  OAI21_X1 U8828 ( .B1(n7197), .B2(n9887), .A(n7117), .ZN(P1_U3282) );
  XNOR2_X1 U8829 ( .A(n7119), .B(n7118), .ZN(n7124) );
  NOR2_X1 U8830 ( .A1(n8278), .A2(n10078), .ZN(n7122) );
  AOI22_X1 U8831 ( .A1(n8251), .A2(n8316), .B1(n8314), .B2(n8269), .ZN(n7185)
         );
  OAI22_X1 U8832 ( .A1(n7185), .A2(n8273), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7120), .ZN(n7121) );
  AOI211_X1 U8833 ( .C1(n8275), .C2(n7186), .A(n7122), .B(n7121), .ZN(n7123)
         );
  OAI21_X1 U8834 ( .B1(n7124), .B2(n8259), .A(n7123), .ZN(P2_U3219) );
  INV_X1 U8835 ( .A(n7125), .ZN(n7126) );
  AOI21_X1 U8836 ( .B1(n7128), .B2(n7127), .A(n7126), .ZN(n7135) );
  INV_X1 U8837 ( .A(n9959), .ZN(n7132) );
  OAI22_X1 U8838 ( .A1(n7129), .A2(n8267), .B1(n7286), .B2(n8249), .ZN(n9957)
         );
  AOI21_X1 U8839 ( .B1(n8285), .B2(n9957), .A(n7130), .ZN(n7131) );
  OAI21_X1 U8840 ( .B1(n7132), .B2(n8287), .A(n7131), .ZN(n7133) );
  AOI21_X1 U8841 ( .B1(n8290), .B2(n10070), .A(n7133), .ZN(n7134) );
  OAI21_X1 U8842 ( .B1(n7135), .B2(n8259), .A(n7134), .ZN(P2_U3233) );
  INV_X1 U8843 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7141) );
  AOI211_X1 U8844 ( .C1(n9606), .C2(n7350), .A(n7137), .B(n7136), .ZN(n7138)
         );
  OAI21_X1 U8845 ( .B1(n9597), .B2(n7139), .A(n7138), .ZN(n7142) );
  NAND2_X1 U8846 ( .A1(n7142), .A2(n9929), .ZN(n7140) );
  OAI21_X1 U8847 ( .B1(n9929), .B2(n7141), .A(n7140), .ZN(P1_U3475) );
  NAND2_X1 U8848 ( .A1(n7142), .A2(n9935), .ZN(n7143) );
  OAI21_X1 U8849 ( .B1(n9935), .B2(n7144), .A(n7143), .ZN(P1_U3530) );
  OAI21_X1 U8850 ( .B1(n7146), .B2(n9095), .A(n7145), .ZN(n9925) );
  NAND2_X1 U8851 ( .A1(n7147), .A2(n7264), .ZN(n7148) );
  NAND2_X1 U8852 ( .A1(n7149), .A2(n7148), .ZN(n9922) );
  NOR2_X1 U8853 ( .A1(n9876), .A2(n7257), .ZN(n7150) );
  AOI21_X1 U8854 ( .B1(n9693), .B2(n7264), .A(n7150), .ZN(n7151) );
  OAI21_X1 U8855 ( .B1(n9922), .B2(n9308), .A(n7151), .ZN(n7159) );
  OR2_X1 U8856 ( .A1(n7152), .A2(n6844), .ZN(n7154) );
  NAND2_X1 U8857 ( .A1(n7154), .A2(n7153), .ZN(n8964) );
  XNOR2_X1 U8858 ( .A(n8964), .B(n9095), .ZN(n7155) );
  OAI222_X1 U8859 ( .A1(n9681), .A2(n7157), .B1(n9682), .B2(n7156), .C1(n7155), 
        .C2(n9510), .ZN(n9923) );
  MUX2_X1 U8860 ( .A(n9923), .B(P1_REG2_REG_6__SCAN_IN), .S(n9887), .Z(n7158)
         );
  AOI211_X1 U8861 ( .C1(n9483), .C2(n9925), .A(n7159), .B(n7158), .ZN(n7160)
         );
  INV_X1 U8862 ( .A(n7160), .ZN(P1_U3285) );
  INV_X1 U8863 ( .A(n7161), .ZN(n7162) );
  OR2_X1 U8864 ( .A1(n7162), .A2(n7956), .ZN(n9976) );
  NAND2_X1 U8865 ( .A1(n9976), .A2(n7163), .ZN(n7164) );
  OR2_X1 U8866 ( .A1(n7164), .A2(n7957), .ZN(n9950) );
  NAND2_X1 U8867 ( .A1(n7164), .A2(n7957), .ZN(n7165) );
  NAND2_X1 U8868 ( .A1(n9950), .A2(n7165), .ZN(n10061) );
  OR2_X1 U8869 ( .A1(n10011), .A2(n7166), .ZN(n7776) );
  OAI21_X1 U8870 ( .B1(n4364), .B2(n7957), .A(n7167), .ZN(n7169) );
  AOI21_X1 U8871 ( .B1(n7169), .B2(n9968), .A(n7168), .ZN(n7170) );
  OAI21_X1 U8872 ( .B1(n10061), .B2(n9955), .A(n7170), .ZN(n10064) );
  NAND2_X1 U8873 ( .A1(n10064), .A2(n10009), .ZN(n7178) );
  INV_X1 U8874 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7172) );
  OAI22_X1 U8875 ( .A1(n10009), .A2(n7172), .B1(n7171), .B2(n8479), .ZN(n7175)
         );
  NAND2_X1 U8876 ( .A1(n9978), .A2(n7176), .ZN(n7173) );
  NAND2_X1 U8877 ( .A1(n9960), .A2(n7173), .ZN(n10063) );
  NOR2_X1 U8878 ( .A1(n10063), .A2(n10003), .ZN(n7174) );
  AOI211_X1 U8879 ( .C1(n9990), .C2(n7176), .A(n7175), .B(n7174), .ZN(n7177)
         );
  OAI211_X1 U8880 ( .C1(n10061), .C2(n7776), .A(n7178), .B(n7177), .ZN(
        P2_U3288) );
  INV_X1 U8881 ( .A(n8479), .ZN(n10001) );
  OAI21_X1 U8882 ( .B1(n7179), .B2(n7959), .A(n7180), .ZN(n7187) );
  INV_X1 U8883 ( .A(n7181), .ZN(n7183) );
  INV_X1 U8884 ( .A(n7959), .ZN(n7182) );
  OAI211_X1 U8885 ( .C1(n7183), .C2(n7182), .A(n9968), .B(n4289), .ZN(n7184)
         );
  OAI211_X1 U8886 ( .C1(n7187), .C2(n9955), .A(n7185), .B(n7184), .ZN(n10079)
         );
  AOI21_X1 U8887 ( .B1(n7186), .B2(n10001), .A(n10079), .ZN(n7193) );
  INV_X1 U8888 ( .A(n7187), .ZN(n10081) );
  INV_X1 U8889 ( .A(n7776), .ZN(n9961) );
  INV_X1 U8890 ( .A(n7290), .ZN(n7188) );
  OAI211_X1 U8891 ( .C1(n10078), .C2(n4353), .A(n7188), .B(n10049), .ZN(n10077) );
  AOI22_X1 U8892 ( .A1(n9990), .A2(n7189), .B1(n10011), .B2(
        P2_REG2_REG_10__SCAN_IN), .ZN(n7190) );
  OAI21_X1 U8893 ( .B1(n10077), .B2(n8588), .A(n7190), .ZN(n7191) );
  AOI21_X1 U8894 ( .B1(n10081), .B2(n9961), .A(n7191), .ZN(n7192) );
  OAI21_X1 U8895 ( .B1(n7193), .B2(n10011), .A(n7192), .ZN(P2_U3286) );
  INV_X1 U8896 ( .A(n7194), .ZN(n7198) );
  AOI22_X1 U8897 ( .A1(n7195), .A2(n9713), .B1(n9606), .B2(n7494), .ZN(n7196)
         );
  OAI211_X1 U8898 ( .C1(n9609), .C2(n7198), .A(n7197), .B(n7196), .ZN(n7201)
         );
  NAND2_X1 U8899 ( .A1(n7201), .A2(n9935), .ZN(n7199) );
  OAI21_X1 U8900 ( .B1(n9935), .B2(n7200), .A(n7199), .ZN(P1_U3532) );
  INV_X1 U8901 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7203) );
  NAND2_X1 U8902 ( .A1(n7201), .A2(n9929), .ZN(n7202) );
  OAI21_X1 U8903 ( .B1(n9929), .B2(n7203), .A(n7202), .ZN(P1_U3481) );
  AOI21_X1 U8904 ( .B1(n7212), .B2(P2_REG1_REG_11__SCAN_IN), .A(n7204), .ZN(
        n7207) );
  INV_X1 U8905 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10118) );
  MUX2_X1 U8906 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n10118), .S(n7324), .Z(n7206) );
  AND2_X1 U8907 ( .A1(n7207), .A2(n7206), .ZN(n7319) );
  INV_X1 U8908 ( .A(n7319), .ZN(n7205) );
  OAI21_X1 U8909 ( .B1(n7207), .B2(n7206), .A(n7205), .ZN(n7217) );
  NOR2_X1 U8910 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7208), .ZN(n7209) );
  AOI21_X1 U8911 ( .B1(n9943), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n7209), .ZN(
        n7210) );
  OAI21_X1 U8912 ( .B1(n9939), .B2(n7320), .A(n7210), .ZN(n7216) );
  OAI21_X1 U8913 ( .B1(n7212), .B2(P2_REG2_REG_11__SCAN_IN), .A(n7211), .ZN(
        n7214) );
  XNOR2_X1 U8914 ( .A(n7324), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n7213) );
  NOR2_X1 U8915 ( .A1(n7214), .A2(n7213), .ZN(n7323) );
  AOI211_X1 U8916 ( .C1(n7214), .C2(n7213), .A(n7323), .B(n9662), .ZN(n7215)
         );
  AOI211_X1 U8917 ( .C1(n9936), .C2(n7217), .A(n7216), .B(n7215), .ZN(n7218)
         );
  INV_X1 U8918 ( .A(n7218), .ZN(P2_U3257) );
  XNOR2_X1 U8919 ( .A(n8914), .B(n9251), .ZN(n9103) );
  INV_X1 U8920 ( .A(n9103), .ZN(n7221) );
  XNOR2_X1 U8921 ( .A(n7219), .B(n7221), .ZN(n7377) );
  NAND2_X1 U8922 ( .A1(n9677), .A2(n7220), .ZN(n7222) );
  XNOR2_X1 U8923 ( .A(n7222), .B(n7221), .ZN(n7225) );
  OAI22_X1 U8924 ( .A1(n7512), .A2(n9682), .B1(n9681), .B2(n8885), .ZN(n7223)
         );
  INV_X1 U8925 ( .A(n7223), .ZN(n7224) );
  OAI21_X1 U8926 ( .B1(n7225), .B2(n9510), .A(n7224), .ZN(n7226) );
  AOI21_X1 U8927 ( .B1(n7377), .B2(n9688), .A(n7226), .ZN(n7379) );
  INV_X1 U8928 ( .A(n7312), .ZN(n7228) );
  NAND2_X1 U8929 ( .A1(n9695), .A2(n8914), .ZN(n7227) );
  NAND2_X1 U8930 ( .A1(n7228), .A2(n7227), .ZN(n7375) );
  OAI22_X1 U8931 ( .A1(n9885), .A2(n6685), .B1(n8907), .B2(n9876), .ZN(n7229)
         );
  AOI21_X1 U8932 ( .B1(n8914), .B2(n9693), .A(n7229), .ZN(n7230) );
  OAI21_X1 U8933 ( .B1(n7375), .B2(n9308), .A(n7230), .ZN(n7231) );
  AOI21_X1 U8934 ( .B1(n7377), .B2(n9699), .A(n7231), .ZN(n7232) );
  OAI21_X1 U8935 ( .B1(n7379), .B2(n9692), .A(n7232), .ZN(P1_U3280) );
  AOI211_X1 U8936 ( .C1(n9606), .C2(n7540), .A(n7234), .B(n7233), .ZN(n7235)
         );
  OAI21_X1 U8937 ( .B1(n9597), .B2(n7236), .A(n7235), .ZN(n7239) );
  NAND2_X1 U8938 ( .A1(n7239), .A2(n9935), .ZN(n7237) );
  OAI21_X1 U8939 ( .B1(n9935), .B2(n7238), .A(n7237), .ZN(P1_U3531) );
  INV_X1 U8940 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7241) );
  NAND2_X1 U8941 ( .A1(n7239), .A2(n9929), .ZN(n7240) );
  OAI21_X1 U8942 ( .B1(n9929), .B2(n7241), .A(n7240), .ZN(P1_U3478) );
  INV_X1 U8943 ( .A(n7242), .ZN(n7251) );
  NOR2_X1 U8944 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(n8479), .ZN(n7243) );
  AOI21_X1 U8945 ( .B1(n9993), .B2(n7244), .A(n7243), .ZN(n7246) );
  NAND2_X1 U8946 ( .A1(n10011), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7245) );
  OAI211_X1 U8947 ( .C1(n10004), .C2(n7247), .A(n7246), .B(n7245), .ZN(n7248)
         );
  AOI21_X1 U8948 ( .B1(n10006), .B2(n7249), .A(n7248), .ZN(n7250) );
  OAI21_X1 U8949 ( .B1(n10011), .B2(n7251), .A(n7250), .ZN(P2_U3293) );
  INV_X1 U8950 ( .A(n7252), .ZN(n7275) );
  NOR2_X1 U8951 ( .A1(n9911), .A2(n7253), .ZN(n9919) );
  AOI21_X1 U8952 ( .B1(n8936), .B2(n9257), .A(n7254), .ZN(n7256) );
  NAND2_X1 U8953 ( .A1(n8942), .A2(n9255), .ZN(n7255) );
  OAI211_X1 U8954 ( .C1(n8926), .C2(n7257), .A(n7256), .B(n7255), .ZN(n7274)
         );
  NAND2_X1 U8955 ( .A1(n8098), .A2(n7264), .ZN(n7260) );
  OAI21_X1 U8956 ( .B1(n7263), .B2(n7262), .A(n7260), .ZN(n7261) );
  XNOR2_X1 U8957 ( .A(n7261), .B(n8063), .ZN(n7265) );
  INV_X1 U8958 ( .A(n7262), .ZN(n9256) );
  AOI22_X1 U8959 ( .A1(n8073), .A2(n9256), .B1(n4269), .B2(n7264), .ZN(n7266)
         );
  NAND2_X1 U8960 ( .A1(n7265), .A2(n7266), .ZN(n7270) );
  INV_X1 U8961 ( .A(n7340), .ZN(n7272) );
  INV_X1 U8962 ( .A(n7265), .ZN(n7268) );
  INV_X1 U8963 ( .A(n7266), .ZN(n7267) );
  NAND2_X1 U8964 ( .A1(n7268), .A2(n7267), .ZN(n7339) );
  AOI21_X1 U8965 ( .B1(n7339), .B2(n7270), .A(n7269), .ZN(n7271) );
  AOI211_X1 U8966 ( .C1(n7272), .C2(n7339), .A(n4653), .B(n7271), .ZN(n7273)
         );
  AOI211_X1 U8967 ( .C1(n7275), .C2(n9919), .A(n7274), .B(n7273), .ZN(n7276)
         );
  INV_X1 U8968 ( .A(n7276), .ZN(P1_U3237) );
  NAND2_X1 U8969 ( .A1(n7279), .A2(n7739), .ZN(n7277) );
  OAI211_X1 U8970 ( .C1(n7278), .C2(n4268), .A(n7277), .B(n7993), .ZN(P2_U3335) );
  NAND2_X1 U8971 ( .A1(n7279), .A2(n7703), .ZN(n7281) );
  NOR2_X1 U8972 ( .A1(n7280), .A2(P1_U3084), .ZN(n9233) );
  INV_X1 U8973 ( .A(n9233), .ZN(n9239) );
  OAI211_X1 U8974 ( .C1(n7282), .C2(n9641), .A(n7281), .B(n9239), .ZN(P1_U3330) );
  OAI21_X1 U8975 ( .B1(n7284), .B2(n7960), .A(n7283), .ZN(n10084) );
  XOR2_X1 U8976 ( .A(n7285), .B(n7960), .Z(n7289) );
  OR2_X1 U8977 ( .A1(n7520), .A2(n8249), .ZN(n7288) );
  OR2_X1 U8978 ( .A1(n7286), .A2(n8267), .ZN(n7287) );
  AND2_X1 U8979 ( .A1(n7288), .A2(n7287), .ZN(n7298) );
  OAI21_X1 U8980 ( .B1(n7289), .B2(n10000), .A(n7298), .ZN(n10089) );
  OAI21_X1 U8981 ( .B1(n7290), .B2(n10085), .A(n7412), .ZN(n10087) );
  AOI22_X1 U8982 ( .A1(n10011), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7301), .B2(
        n10001), .ZN(n7293) );
  NAND2_X1 U8983 ( .A1(n9990), .A2(n7291), .ZN(n7292) );
  OAI211_X1 U8984 ( .C1(n10087), .C2(n10003), .A(n7293), .B(n7292), .ZN(n7294)
         );
  AOI21_X1 U8985 ( .B1(n10089), .B2(n10009), .A(n7294), .ZN(n7295) );
  OAI21_X1 U8986 ( .B1(n10084), .B2(n8592), .A(n7295), .ZN(P2_U3285) );
  XNOR2_X1 U8987 ( .A(n7297), .B(n7296), .ZN(n7303) );
  OAI22_X1 U8988 ( .A1(n8273), .A2(n7298), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5743), .ZN(n7300) );
  NOR2_X1 U8989 ( .A1(n10085), .A2(n8278), .ZN(n7299) );
  AOI211_X1 U8990 ( .C1(n8275), .C2(n7301), .A(n7300), .B(n7299), .ZN(n7302)
         );
  OAI21_X1 U8991 ( .B1(n7303), .B2(n8259), .A(n7302), .ZN(P2_U3238) );
  NAND2_X1 U8992 ( .A1(n4845), .A2(n7304), .ZN(n7305) );
  INV_X1 U8993 ( .A(n9101), .ZN(n7306) );
  XNOR2_X1 U8994 ( .A(n7305), .B(n7306), .ZN(n9725) );
  XNOR2_X1 U8995 ( .A(n7307), .B(n7306), .ZN(n7310) );
  OAI22_X1 U8996 ( .A1(n8825), .A2(n9681), .B1(n9682), .B2(n9680), .ZN(n7308)
         );
  INV_X1 U8997 ( .A(n7308), .ZN(n7309) );
  OAI21_X1 U8998 ( .B1(n7310), .B2(n9510), .A(n7309), .ZN(n7311) );
  AOI21_X1 U8999 ( .B1(n9725), .B2(n9688), .A(n7311), .ZN(n9727) );
  OAI21_X1 U9000 ( .B1(n7312), .B2(n9723), .A(n9713), .ZN(n7313) );
  OR2_X1 U9001 ( .A1(n7313), .A2(n7459), .ZN(n9722) );
  INV_X1 U9002 ( .A(n9698), .ZN(n7548) );
  INV_X1 U9003 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7314) );
  OAI22_X1 U9004 ( .A1(n9885), .A2(n7314), .B1(n8828), .B2(n9876), .ZN(n7315)
         );
  AOI21_X1 U9005 ( .B1(n8830), .B2(n9693), .A(n7315), .ZN(n7316) );
  OAI21_X1 U9006 ( .B1(n9722), .B2(n7548), .A(n7316), .ZN(n7317) );
  AOI21_X1 U9007 ( .B1(n9725), .B2(n9699), .A(n7317), .ZN(n7318) );
  OAI21_X1 U9008 ( .B1(n9727), .B2(n9887), .A(n7318), .ZN(P1_U3279) );
  AOI21_X1 U9009 ( .B1(n10118), .B2(n7320), .A(n7319), .ZN(n7322) );
  INV_X1 U9010 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7468) );
  AOI22_X1 U9011 ( .A1(n7474), .A2(n7468), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n7469), .ZN(n7321) );
  NOR2_X1 U9012 ( .A1(n7322), .A2(n7321), .ZN(n7467) );
  AOI21_X1 U9013 ( .B1(n7322), .B2(n7321), .A(n7467), .ZN(n7333) );
  NOR2_X1 U9014 ( .A1(n7474), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7325) );
  AOI21_X1 U9015 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n7474), .A(n7325), .ZN(
        n7326) );
  OAI21_X1 U9016 ( .B1(n7327), .B2(n7326), .A(n7473), .ZN(n7331) );
  NOR2_X1 U9017 ( .A1(n7328), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7525) );
  AOI21_X1 U9018 ( .B1(n9943), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n7525), .ZN(
        n7329) );
  OAI21_X1 U9019 ( .B1(n9939), .B2(n7469), .A(n7329), .ZN(n7330) );
  AOI21_X1 U9020 ( .B1(n7331), .B2(n9937), .A(n7330), .ZN(n7332) );
  OAI21_X1 U9021 ( .B1(n7333), .B2(n9941), .A(n7332), .ZN(P2_U3258) );
  INV_X1 U9022 ( .A(n7334), .ZN(n7335) );
  AOI21_X1 U9023 ( .B1(n8936), .B2(n9256), .A(n7335), .ZN(n7337) );
  NAND2_X1 U9024 ( .A1(n8942), .A2(n9254), .ZN(n7336) );
  OAI211_X1 U9025 ( .C1(n8926), .C2(n7338), .A(n7337), .B(n7336), .ZN(n7349)
         );
  NAND2_X1 U9026 ( .A1(n7350), .A2(n8098), .ZN(n7342) );
  NAND2_X1 U9027 ( .A1(n4269), .A2(n9255), .ZN(n7341) );
  NAND2_X1 U9028 ( .A1(n7342), .A2(n7341), .ZN(n7343) );
  XNOR2_X1 U9029 ( .A(n7343), .B(n8063), .ZN(n7495) );
  NAND2_X1 U9030 ( .A1(n8073), .A2(n9255), .ZN(n7345) );
  NAND2_X1 U9031 ( .A1(n7350), .A2(n4269), .ZN(n7344) );
  NAND2_X1 U9032 ( .A1(n7345), .A2(n7344), .ZN(n7485) );
  XNOR2_X1 U9033 ( .A(n7495), .B(n7485), .ZN(n7346) );
  XNOR2_X1 U9034 ( .A(n7486), .B(n7346), .ZN(n7347) );
  NOR2_X1 U9035 ( .A1(n7347), .A2(n4653), .ZN(n7348) );
  AOI211_X1 U9036 ( .C1(n8928), .C2(n7350), .A(n7349), .B(n7348), .ZN(n7351)
         );
  INV_X1 U9037 ( .A(n7351), .ZN(P1_U3211) );
  INV_X1 U9038 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7357) );
  INV_X1 U9039 ( .A(n9801), .ZN(n7356) );
  INV_X1 U9040 ( .A(n9786), .ZN(n7355) );
  INV_X1 U9041 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9728) );
  NOR2_X1 U9042 ( .A1(n9786), .A2(n9728), .ZN(n7354) );
  AOI21_X1 U9043 ( .B1(n9786), .B2(n9728), .A(n7354), .ZN(n9794) );
  NOR2_X1 U9044 ( .A1(n9795), .A2(n9794), .ZN(n9793) );
  MUX2_X1 U9045 ( .A(n7357), .B(P1_REG1_REG_13__SCAN_IN), .S(n9801), .Z(n9810)
         );
  NOR2_X1 U9046 ( .A1(n9809), .A2(n9810), .ZN(n9808) );
  INV_X1 U9047 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9721) );
  AOI22_X1 U9048 ( .A1(n7371), .A2(n9721), .B1(P1_REG1_REG_14__SCAN_IN), .B2(
        n9275), .ZN(n7358) );
  NOR2_X1 U9049 ( .A1(n7359), .A2(n7358), .ZN(n9274) );
  AOI21_X1 U9050 ( .B1(n7359), .B2(n7358), .A(n9274), .ZN(n7374) );
  NAND2_X1 U9051 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8783) );
  INV_X1 U9052 ( .A(n8783), .ZN(n7370) );
  OR2_X1 U9053 ( .A1(n9786), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7361) );
  NAND2_X1 U9054 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n9786), .ZN(n7360) );
  NAND2_X1 U9055 ( .A1(n7361), .A2(n7360), .ZN(n9788) );
  OR2_X1 U9056 ( .A1(n7362), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7364) );
  NAND2_X1 U9057 ( .A1(n7364), .A2(n7363), .ZN(n9789) );
  OR2_X1 U9058 ( .A1(n9801), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7366) );
  NAND2_X1 U9059 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n9801), .ZN(n7365) );
  NAND2_X1 U9060 ( .A1(n7366), .A2(n7365), .ZN(n9804) );
  INV_X1 U9061 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7367) );
  NOR2_X1 U9062 ( .A1(n7367), .A2(n7368), .ZN(n9264) );
  AOI211_X1 U9063 ( .C1(n7368), .C2(n7367), .A(n9264), .B(n9826), .ZN(n7369)
         );
  AOI211_X1 U9064 ( .C1(n9859), .C2(n7371), .A(n7370), .B(n7369), .ZN(n7373)
         );
  NAND2_X1 U9065 ( .A1(n9773), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n7372) );
  OAI211_X1 U9066 ( .C1(n7374), .C2(n9867), .A(n7373), .B(n7372), .ZN(P1_U3255) );
  INV_X1 U9067 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7380) );
  INV_X1 U9068 ( .A(n9609), .ZN(n9917) );
  OAI22_X1 U9069 ( .A1(n7375), .A2(n9921), .B1(n4542), .B2(n9911), .ZN(n7376)
         );
  AOI21_X1 U9070 ( .B1(n7377), .B2(n9917), .A(n7376), .ZN(n7378) );
  AND2_X1 U9071 ( .A1(n7379), .A2(n7378), .ZN(n7382) );
  MUX2_X1 U9072 ( .A(n7380), .B(n7382), .S(n9929), .Z(n7381) );
  INV_X1 U9073 ( .A(n7381), .ZN(P1_U3487) );
  MUX2_X1 U9074 ( .A(n7383), .B(n7382), .S(n9935), .Z(n7384) );
  INV_X1 U9075 ( .A(n7384), .ZN(P1_U3534) );
  INV_X1 U9076 ( .A(n7385), .ZN(n7402) );
  OAI222_X1 U9077 ( .A1(n9645), .A2(n7402), .B1(P1_U3084), .B2(n7387), .C1(
        n7386), .C2(n9641), .ZN(P1_U3329) );
  NAND2_X1 U9078 ( .A1(n7389), .A2(n7388), .ZN(n7391) );
  XOR2_X1 U9079 ( .A(n7391), .B(n7390), .Z(n7399) );
  INV_X1 U9080 ( .A(n7392), .ZN(n7410) );
  OR2_X1 U9081 ( .A1(n7868), .A2(n8249), .ZN(n7395) );
  OR2_X1 U9082 ( .A1(n7393), .A2(n8267), .ZN(n7394) );
  NAND2_X1 U9083 ( .A1(n7395), .A2(n7394), .ZN(n7406) );
  AOI22_X1 U9084 ( .A1(n8285), .A2(n7406), .B1(P2_REG3_REG_12__SCAN_IN), .B2(
        P2_U3152), .ZN(n7396) );
  OAI21_X1 U9085 ( .B1(n7410), .B2(n8287), .A(n7396), .ZN(n7397) );
  AOI21_X1 U9086 ( .B1(n8290), .B2(n7416), .A(n7397), .ZN(n7398) );
  OAI21_X1 U9087 ( .B1(n7399), .B2(n8259), .A(n7398), .ZN(P2_U3226) );
  INV_X1 U9088 ( .A(n7400), .ZN(n7403) );
  OAI222_X1 U9089 ( .A1(n7403), .A2(n4262), .B1(n8768), .B2(n7402), .C1(n7401), 
        .C2(n4268), .ZN(P2_U3334) );
  NAND2_X1 U9090 ( .A1(n7404), .A2(n7851), .ZN(n7405) );
  XNOR2_X1 U9091 ( .A(n7405), .B(n6069), .ZN(n7407) );
  AOI21_X1 U9092 ( .B1(n7407), .B2(n9968), .A(n7406), .ZN(n10093) );
  OAI21_X1 U9093 ( .B1(n7409), .B2(n6069), .A(n7408), .ZN(n10098) );
  NAND2_X1 U9094 ( .A1(n10098), .A2(n10006), .ZN(n7418) );
  INV_X1 U9095 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7411) );
  OAI22_X1 U9096 ( .A1(n10009), .A2(n7411), .B1(n7410), .B2(n8479), .ZN(n7415)
         );
  INV_X1 U9097 ( .A(n7412), .ZN(n7413) );
  INV_X1 U9098 ( .A(n7416), .ZN(n10095) );
  OAI211_X1 U9099 ( .C1(n7413), .C2(n10095), .A(n10049), .B(n4358), .ZN(n10092) );
  NOR2_X1 U9100 ( .A1(n10092), .A2(n8588), .ZN(n7414) );
  AOI211_X1 U9101 ( .C1(n9990), .C2(n7416), .A(n7415), .B(n7414), .ZN(n7417)
         );
  OAI211_X1 U9102 ( .C1(n10011), .C2(n10093), .A(n7418), .B(n7417), .ZN(
        P2_U3284) );
  INV_X1 U9103 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10158) );
  NOR2_X1 U9104 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7419) );
  AOI21_X1 U9105 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7419), .ZN(n10129) );
  NOR2_X1 U9106 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7420) );
  AOI21_X1 U9107 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7420), .ZN(n10132) );
  NOR2_X1 U9108 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7421) );
  AOI21_X1 U9109 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7421), .ZN(n10135) );
  NOR2_X1 U9110 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7422) );
  AOI21_X1 U9111 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7422), .ZN(n10138) );
  NOR2_X1 U9112 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7423) );
  AOI21_X1 U9113 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7423), .ZN(n10141) );
  NOR2_X1 U9114 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7429) );
  XNOR2_X1 U9115 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10169) );
  NAND2_X1 U9116 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7427) );
  XOR2_X1 U9117 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10167) );
  NAND2_X1 U9118 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7425) );
  XOR2_X1 U9119 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10165) );
  AOI21_X1 U9120 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10121) );
  INV_X1 U9121 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9649) );
  NAND3_X1 U9122 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10123) );
  OAI21_X1 U9123 ( .B1(n10121), .B2(n9649), .A(n10123), .ZN(n10164) );
  NAND2_X1 U9124 ( .A1(n10165), .A2(n10164), .ZN(n7424) );
  NAND2_X1 U9125 ( .A1(n7425), .A2(n7424), .ZN(n10166) );
  NAND2_X1 U9126 ( .A1(n10167), .A2(n10166), .ZN(n7426) );
  NAND2_X1 U9127 ( .A1(n7427), .A2(n7426), .ZN(n10168) );
  NOR2_X1 U9128 ( .A1(n10169), .A2(n10168), .ZN(n7428) );
  NOR2_X1 U9129 ( .A1(n7429), .A2(n7428), .ZN(n7430) );
  NOR2_X1 U9130 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7430), .ZN(n10153) );
  AND2_X1 U9131 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7430), .ZN(n10152) );
  NOR2_X1 U9132 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10152), .ZN(n7431) );
  NOR2_X1 U9133 ( .A1(n10153), .A2(n7431), .ZN(n7432) );
  NAND2_X1 U9134 ( .A1(n7432), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7434) );
  XOR2_X1 U9135 ( .A(n7432), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10151) );
  NAND2_X1 U9136 ( .A1(n10151), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7433) );
  NAND2_X1 U9137 ( .A1(n7434), .A2(n7433), .ZN(n7435) );
  NAND2_X1 U9138 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7435), .ZN(n7437) );
  XOR2_X1 U9139 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7435), .Z(n10160) );
  NAND2_X1 U9140 ( .A1(n10160), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7436) );
  NAND2_X1 U9141 ( .A1(n7437), .A2(n7436), .ZN(n7438) );
  NAND2_X1 U9142 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7438), .ZN(n7440) );
  XOR2_X1 U9143 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7438), .Z(n10155) );
  NAND2_X1 U9144 ( .A1(n10155), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7439) );
  NAND2_X1 U9145 ( .A1(n7440), .A2(n7439), .ZN(n7441) );
  AND2_X1 U9146 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7441), .ZN(n7442) );
  XNOR2_X1 U9147 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7441), .ZN(n10162) );
  NOR2_X1 U9148 ( .A1(n10163), .A2(n10162), .ZN(n10161) );
  NOR2_X1 U9149 ( .A1(n7442), .A2(n10161), .ZN(n10150) );
  NAND2_X1 U9150 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7443) );
  OAI21_X1 U9151 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7443), .ZN(n10149) );
  NOR2_X1 U9152 ( .A1(n10150), .A2(n10149), .ZN(n10148) );
  AOI21_X1 U9153 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10148), .ZN(n10147) );
  NAND2_X1 U9154 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7444) );
  OAI21_X1 U9155 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7444), .ZN(n10146) );
  NOR2_X1 U9156 ( .A1(n10147), .A2(n10146), .ZN(n10145) );
  AOI21_X1 U9157 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10145), .ZN(n10144) );
  NOR2_X1 U9158 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7445) );
  AOI21_X1 U9159 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7445), .ZN(n10143) );
  NAND2_X1 U9160 ( .A1(n10144), .A2(n10143), .ZN(n10142) );
  OAI21_X1 U9161 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10142), .ZN(n10140) );
  NAND2_X1 U9162 ( .A1(n10141), .A2(n10140), .ZN(n10139) );
  OAI21_X1 U9163 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10139), .ZN(n10137) );
  NAND2_X1 U9164 ( .A1(n10138), .A2(n10137), .ZN(n10136) );
  OAI21_X1 U9165 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10136), .ZN(n10134) );
  NAND2_X1 U9166 ( .A1(n10135), .A2(n10134), .ZN(n10133) );
  OAI21_X1 U9167 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10133), .ZN(n10131) );
  NAND2_X1 U9168 ( .A1(n10132), .A2(n10131), .ZN(n10130) );
  OAI21_X1 U9169 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10130), .ZN(n10128) );
  NAND2_X1 U9170 ( .A1(n10129), .A2(n10128), .ZN(n10127) );
  OAI21_X1 U9171 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10127), .ZN(n10157) );
  NOR2_X1 U9172 ( .A1(n10158), .A2(n10157), .ZN(n7446) );
  NAND2_X1 U9173 ( .A1(n10158), .A2(n10157), .ZN(n10156) );
  OAI21_X1 U9174 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7446), .A(n10156), .ZN(
        n7450) );
  NOR2_X1 U9175 ( .A1(n7447), .A2(n7448), .ZN(n7449) );
  XNOR2_X1 U9176 ( .A(n7450), .B(n7449), .ZN(ADD_1071_U4) );
  XNOR2_X1 U9177 ( .A(n7451), .B(n9087), .ZN(n7452) );
  INV_X1 U9178 ( .A(n7452), .ZN(n9610) );
  NAND2_X1 U9179 ( .A1(n7452), .A2(n9688), .ZN(n7458) );
  OAI21_X1 U9180 ( .B1(n9087), .B2(n7454), .A(n7453), .ZN(n7456) );
  OAI22_X1 U9181 ( .A1(n8885), .A2(n9682), .B1(n9681), .B2(n8976), .ZN(n7455)
         );
  AOI21_X1 U9182 ( .B1(n7456), .B2(n9685), .A(n7455), .ZN(n7457) );
  NAND2_X1 U9183 ( .A1(n7458), .A2(n7457), .ZN(n9612) );
  NAND2_X1 U9184 ( .A1(n9612), .A2(n9885), .ZN(n7466) );
  OR2_X1 U9185 ( .A1(n7459), .A2(n7461), .ZN(n7460) );
  AND2_X1 U9186 ( .A1(n7547), .A2(n7460), .ZN(n9607) );
  NOR2_X1 U9187 ( .A1(n7461), .A2(n9519), .ZN(n7464) );
  INV_X1 U9188 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7462) );
  OAI22_X1 U9189 ( .A1(n9885), .A2(n7462), .B1(n8888), .B2(n9876), .ZN(n7463)
         );
  AOI211_X1 U9190 ( .C1(n9607), .C2(n9504), .A(n7464), .B(n7463), .ZN(n7465)
         );
  OAI211_X1 U9191 ( .C1(n9610), .C2(n7605), .A(n7466), .B(n7465), .ZN(P1_U3278) );
  AOI21_X1 U9192 ( .B1(n7469), .B2(n7468), .A(n7467), .ZN(n7471) );
  INV_X1 U9193 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8326) );
  AOI22_X1 U9194 ( .A1(n8330), .A2(n8326), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n8327), .ZN(n7470) );
  NOR2_X1 U9195 ( .A1(n7471), .A2(n7470), .ZN(n8325) );
  AOI21_X1 U9196 ( .B1(n7471), .B2(n7470), .A(n8325), .ZN(n7482) );
  NOR2_X1 U9197 ( .A1(n8330), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7472) );
  AOI21_X1 U9198 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8330), .A(n7472), .ZN(
        n7476) );
  OAI21_X1 U9199 ( .B1(n7476), .B2(n7475), .A(n8329), .ZN(n7480) );
  NOR2_X1 U9200 ( .A1(n7477), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7616) );
  AOI21_X1 U9201 ( .B1(n9943), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n7616), .ZN(
        n7478) );
  OAI21_X1 U9202 ( .B1(n9939), .B2(n8327), .A(n7478), .ZN(n7479) );
  AOI21_X1 U9203 ( .B1(n7480), .B2(n9937), .A(n7479), .ZN(n7481) );
  OAI21_X1 U9204 ( .B1(n7482), .B2(n9941), .A(n7481), .ZN(P2_U3259) );
  INV_X1 U9205 ( .A(n7486), .ZN(n7484) );
  INV_X1 U9206 ( .A(n7485), .ZN(n7483) );
  NAND2_X1 U9207 ( .A1(n7484), .A2(n7483), .ZN(n7497) );
  NAND2_X1 U9208 ( .A1(n7486), .A2(n7485), .ZN(n7500) );
  NAND2_X1 U9209 ( .A1(n7500), .A2(n7495), .ZN(n7489) );
  NAND2_X1 U9210 ( .A1(n7540), .A2(n4269), .ZN(n7488) );
  NAND2_X1 U9211 ( .A1(n8073), .A2(n9254), .ZN(n7487) );
  NAND2_X1 U9212 ( .A1(n7488), .A2(n7487), .ZN(n7498) );
  NAND2_X1 U9213 ( .A1(n7494), .A2(n8098), .ZN(n7491) );
  NAND2_X1 U9214 ( .A1(n4269), .A2(n9253), .ZN(n7490) );
  NAND2_X1 U9215 ( .A1(n7491), .A2(n7490), .ZN(n7492) );
  XNOR2_X1 U9216 ( .A(n7492), .B(n8096), .ZN(n7629) );
  NOR2_X1 U9217 ( .A1(n6660), .A2(n9683), .ZN(n7493) );
  AOI21_X1 U9218 ( .B1(n7494), .B2(n4269), .A(n7493), .ZN(n7630) );
  XNOR2_X1 U9219 ( .A(n7629), .B(n7630), .ZN(n7507) );
  INV_X1 U9220 ( .A(n7495), .ZN(n7496) );
  NAND2_X1 U9221 ( .A1(n7497), .A2(n7496), .ZN(n7502) );
  INV_X1 U9222 ( .A(n7498), .ZN(n7499) );
  AND2_X1 U9223 ( .A1(n7500), .A2(n7499), .ZN(n7501) );
  NAND2_X1 U9224 ( .A1(n7502), .A2(n7501), .ZN(n7534) );
  NAND2_X1 U9225 ( .A1(n7540), .A2(n8098), .ZN(n7504) );
  NAND2_X1 U9226 ( .A1(n4269), .A2(n9254), .ZN(n7503) );
  NAND2_X1 U9227 ( .A1(n7504), .A2(n7503), .ZN(n7505) );
  XNOR2_X1 U9228 ( .A(n7505), .B(n8096), .ZN(n7533) );
  NAND2_X1 U9229 ( .A1(n7534), .A2(n7533), .ZN(n7532) );
  NAND2_X1 U9230 ( .A1(n7506), .A2(n7532), .ZN(n7633) );
  INV_X1 U9231 ( .A(n7633), .ZN(n7509) );
  AOI21_X1 U9232 ( .B1(n7532), .B2(n7536), .A(n7507), .ZN(n7508) );
  OAI21_X1 U9233 ( .B1(n7509), .B2(n7508), .A(n8935), .ZN(n7516) );
  INV_X1 U9234 ( .A(n8926), .ZN(n8937) );
  AOI21_X1 U9235 ( .B1(n8936), .B2(n9254), .A(n7510), .ZN(n7511) );
  OAI21_X1 U9236 ( .B1(n8923), .B2(n7512), .A(n7511), .ZN(n7513) );
  AOI21_X1 U9237 ( .B1(n7514), .B2(n8937), .A(n7513), .ZN(n7515) );
  OAI211_X1 U9238 ( .C1(n7517), .C2(n8945), .A(n7516), .B(n7515), .ZN(P1_U3229) );
  INV_X1 U9239 ( .A(n8680), .ZN(n7867) );
  OAI211_X1 U9240 ( .C1(n7519), .C2(n7518), .A(n7611), .B(n8282), .ZN(n7527)
         );
  OR2_X1 U9241 ( .A1(n7709), .A2(n8249), .ZN(n7522) );
  OR2_X1 U9242 ( .A1(n7520), .A2(n8267), .ZN(n7521) );
  NAND2_X1 U9243 ( .A1(n7522), .A2(n7521), .ZN(n7557) );
  INV_X1 U9244 ( .A(n7562), .ZN(n7523) );
  NOR2_X1 U9245 ( .A1(n8287), .A2(n7523), .ZN(n7524) );
  AOI211_X1 U9246 ( .C1(n8285), .C2(n7557), .A(n7525), .B(n7524), .ZN(n7526)
         );
  OAI211_X1 U9247 ( .C1(n7867), .C2(n8278), .A(n7527), .B(n7526), .ZN(P2_U3236) );
  NOR2_X1 U9248 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7528), .ZN(n9774) );
  AOI21_X1 U9249 ( .B1(n8936), .B2(n9255), .A(n9774), .ZN(n7530) );
  NAND2_X1 U9250 ( .A1(n8942), .A2(n9253), .ZN(n7529) );
  OAI211_X1 U9251 ( .C1(n8926), .C2(n7531), .A(n7530), .B(n7529), .ZN(n7539)
         );
  INV_X1 U9252 ( .A(n7532), .ZN(n7537) );
  AOI21_X1 U9253 ( .B1(n7534), .B2(n7536), .A(n7533), .ZN(n7535) );
  AOI211_X1 U9254 ( .C1(n7537), .C2(n7536), .A(n4653), .B(n7535), .ZN(n7538)
         );
  AOI211_X1 U9255 ( .C1(n8928), .C2(n7540), .A(n7539), .B(n7538), .ZN(n7541)
         );
  INV_X1 U9256 ( .A(n7541), .ZN(P1_U3219) );
  INV_X1 U9257 ( .A(n9107), .ZN(n7542) );
  XNOR2_X1 U9258 ( .A(n7543), .B(n7542), .ZN(n7545) );
  OAI22_X1 U9259 ( .A1(n8825), .A2(n9682), .B1(n9681), .B2(n9511), .ZN(n7544)
         );
  AOI21_X1 U9260 ( .B1(n7545), .B2(n9685), .A(n7544), .ZN(n9717) );
  XNOR2_X1 U9261 ( .A(n7546), .B(n9107), .ZN(n9720) );
  NAND2_X1 U9262 ( .A1(n9720), .A2(n9483), .ZN(n7552) );
  OAI22_X1 U9263 ( .A1(n9885), .A2(n7367), .B1(n8782), .B2(n9876), .ZN(n7550)
         );
  INV_X1 U9264 ( .A(n8977), .ZN(n9718) );
  OAI211_X1 U9265 ( .C1(n4539), .C2(n9718), .A(n9713), .B(n4270), .ZN(n9716)
         );
  NOR2_X1 U9266 ( .A1(n9716), .A2(n7548), .ZN(n7549) );
  AOI211_X1 U9267 ( .C1(n9693), .C2(n8977), .A(n7550), .B(n7549), .ZN(n7551)
         );
  OAI211_X1 U9268 ( .C1(n9887), .C2(n9717), .A(n7552), .B(n7551), .ZN(P1_U3277) );
  OAI21_X1 U9269 ( .B1(n7555), .B2(n7554), .A(n7553), .ZN(n8683) );
  XNOR2_X1 U9270 ( .A(n7556), .B(n7962), .ZN(n7558) );
  AOI21_X1 U9271 ( .B1(n7558), .B2(n9968), .A(n7557), .ZN(n7559) );
  OAI21_X1 U9272 ( .B1(n8683), .B2(n9955), .A(n7559), .ZN(n8685) );
  NAND2_X1 U9273 ( .A1(n8685), .A2(n10009), .ZN(n7567) );
  NAND2_X1 U9274 ( .A1(n4358), .A2(n8680), .ZN(n7560) );
  NAND2_X1 U9275 ( .A1(n7560), .A2(n10049), .ZN(n7561) );
  OR2_X1 U9276 ( .A1(n7561), .A2(n7585), .ZN(n8681) );
  INV_X1 U9277 ( .A(n8681), .ZN(n7565) );
  AOI22_X1 U9278 ( .A1(n10011), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7562), .B2(
        n10001), .ZN(n7563) );
  OAI21_X1 U9279 ( .B1(n7867), .B2(n10004), .A(n7563), .ZN(n7564) );
  AOI21_X1 U9280 ( .B1(n7565), .B2(n9993), .A(n7564), .ZN(n7566) );
  OAI211_X1 U9281 ( .C1(n8683), .C2(n7776), .A(n7567), .B(n7566), .ZN(P2_U3283) );
  INV_X1 U9282 ( .A(n7568), .ZN(n7574) );
  INV_X1 U9283 ( .A(n7569), .ZN(n7570) );
  OAI222_X1 U9284 ( .A1(n9641), .A2(n7571), .B1(n9639), .B2(n7574), .C1(n7570), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  INV_X1 U9285 ( .A(n7572), .ZN(n7573) );
  OAI222_X1 U9286 ( .A1(n4268), .A2(n7575), .B1(n8768), .B2(n7574), .C1(n7573), 
        .C2(n4262), .ZN(P2_U3333) );
  OAI21_X1 U9287 ( .B1(n7576), .B2(n7946), .A(n7577), .ZN(n7578) );
  INV_X1 U9288 ( .A(n7578), .ZN(n7727) );
  INV_X1 U9289 ( .A(n7579), .ZN(n7580) );
  AOI211_X1 U9290 ( .C1(n7946), .C2(n7581), .A(n10000), .B(n7580), .ZN(n7584)
         );
  OR2_X1 U9291 ( .A1(n7768), .A2(n8249), .ZN(n7583) );
  OR2_X1 U9292 ( .A1(n7868), .A2(n8267), .ZN(n7582) );
  NAND2_X1 U9293 ( .A1(n7583), .A2(n7582), .ZN(n7617) );
  OR2_X1 U9294 ( .A1(n7584), .A2(n7617), .ZN(n7720) );
  INV_X1 U9295 ( .A(n7585), .ZN(n7586) );
  AOI211_X1 U9296 ( .C1(n7722), .C2(n7586), .A(n10086), .B(n7714), .ZN(n7721)
         );
  NAND2_X1 U9297 ( .A1(n7721), .A2(n9993), .ZN(n7588) );
  AOI22_X1 U9298 ( .A1(n10011), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7615), .B2(
        n10001), .ZN(n7587) );
  OAI211_X1 U9299 ( .C1(n7589), .C2(n10004), .A(n7588), .B(n7587), .ZN(n7590)
         );
  AOI21_X1 U9300 ( .B1(n7720), .B2(n10009), .A(n7590), .ZN(n7591) );
  OAI21_X1 U9301 ( .B1(n7727), .B2(n8592), .A(n7591), .ZN(P2_U3282) );
  XNOR2_X1 U9302 ( .A(n7592), .B(n9105), .ZN(n9598) );
  INV_X1 U9303 ( .A(n9598), .ZN(n7606) );
  NAND2_X1 U9304 ( .A1(n9598), .A2(n9688), .ZN(n7598) );
  INV_X1 U9305 ( .A(n9105), .ZN(n7593) );
  XNOR2_X1 U9306 ( .A(n7594), .B(n7593), .ZN(n7596) );
  OAI22_X1 U9307 ( .A1(n8976), .A2(n9682), .B1(n9681), .B2(n8005), .ZN(n7595)
         );
  AOI21_X1 U9308 ( .B1(n7596), .B2(n9685), .A(n7595), .ZN(n7597) );
  NAND2_X1 U9309 ( .A1(n7598), .A2(n7597), .ZN(n9603) );
  NAND2_X1 U9310 ( .A1(n9603), .A2(n9885), .ZN(n7604) );
  INV_X1 U9311 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7599) );
  OAI22_X1 U9312 ( .A1(n9885), .A2(n7599), .B1(n7699), .B2(n9876), .ZN(n7602)
         );
  AND2_X1 U9313 ( .A1(n4270), .A2(n9599), .ZN(n7600) );
  OR2_X1 U9314 ( .A1(n7600), .A2(n9515), .ZN(n9601) );
  NOR2_X1 U9315 ( .A1(n9601), .A2(n9308), .ZN(n7601) );
  AOI211_X1 U9316 ( .C1(n9693), .C2(n9599), .A(n7602), .B(n7601), .ZN(n7603)
         );
  OAI211_X1 U9317 ( .C1(n7606), .C2(n7605), .A(n7604), .B(n7603), .ZN(P1_U3276) );
  INV_X1 U9318 ( .A(n7607), .ZN(n7650) );
  INV_X1 U9319 ( .A(n7608), .ZN(n7610) );
  OAI222_X1 U9320 ( .A1(n9645), .A2(n7650), .B1(P1_U3084), .B2(n7610), .C1(
        n7609), .C2(n9641), .ZN(P1_U3327) );
  INV_X1 U9321 ( .A(n7611), .ZN(n7614) );
  INV_X1 U9322 ( .A(n8244), .ZN(n8262) );
  NOR3_X1 U9323 ( .A1(n7612), .A2(n7868), .A3(n8262), .ZN(n7613) );
  AOI21_X1 U9324 ( .B1(n7614), .B2(n8282), .A(n7613), .ZN(n7625) );
  INV_X1 U9325 ( .A(n7615), .ZN(n7619) );
  AOI21_X1 U9326 ( .B1(n8285), .B2(n7617), .A(n7616), .ZN(n7618) );
  OAI21_X1 U9327 ( .B1(n7619), .B2(n8287), .A(n7618), .ZN(n7622) );
  NOR2_X1 U9328 ( .A1(n7620), .A2(n8259), .ZN(n7621) );
  AOI211_X1 U9329 ( .C1(n8290), .C2(n7722), .A(n7622), .B(n7621), .ZN(n7623)
         );
  OAI21_X1 U9330 ( .B1(n7625), .B2(n7624), .A(n7623), .ZN(P2_U3217) );
  AOI21_X1 U9331 ( .B1(n8936), .B2(n9253), .A(n7626), .ZN(n7628) );
  NAND2_X1 U9332 ( .A1(n8942), .A2(n9251), .ZN(n7627) );
  OAI211_X1 U9333 ( .C1(n8926), .C2(n9689), .A(n7628), .B(n7627), .ZN(n7646)
         );
  INV_X1 U9334 ( .A(n7629), .ZN(n7631) );
  NAND2_X1 U9335 ( .A1(n7631), .A2(n7630), .ZN(n7632) );
  NAND2_X1 U9336 ( .A1(n9694), .A2(n8098), .ZN(n7635) );
  NAND2_X1 U9337 ( .A1(n4269), .A2(n9252), .ZN(n7634) );
  NAND2_X1 U9338 ( .A1(n7635), .A2(n7634), .ZN(n7636) );
  XNOR2_X1 U9339 ( .A(n7636), .B(n8096), .ZN(n7639) );
  NAND2_X1 U9340 ( .A1(n9694), .A2(n4269), .ZN(n7638) );
  NAND2_X1 U9341 ( .A1(n8073), .A2(n9252), .ZN(n7637) );
  NAND2_X1 U9342 ( .A1(n7638), .A2(n7637), .ZN(n7640) );
  NAND2_X1 U9343 ( .A1(n7639), .A2(n7640), .ZN(n7688) );
  INV_X1 U9344 ( .A(n7639), .ZN(n7642) );
  INV_X1 U9345 ( .A(n7640), .ZN(n7641) );
  NAND2_X1 U9346 ( .A1(n7642), .A2(n7641), .ZN(n8817) );
  NAND2_X1 U9347 ( .A1(n7688), .A2(n8817), .ZN(n7643) );
  XNOR2_X1 U9348 ( .A(n7689), .B(n7643), .ZN(n7644) );
  NOR2_X1 U9349 ( .A1(n7644), .A2(n4653), .ZN(n7645) );
  AOI211_X1 U9350 ( .C1(n8928), .C2(n9694), .A(n7646), .B(n7645), .ZN(n7647)
         );
  INV_X1 U9351 ( .A(n7647), .ZN(P1_U3215) );
  INV_X1 U9352 ( .A(n7648), .ZN(n7651) );
  OAI222_X1 U9353 ( .A1(n7651), .A2(P2_U3152), .B1(n8768), .B2(n7650), .C1(
        n7649), .C2(n4268), .ZN(P2_U3332) );
  NAND2_X1 U9354 ( .A1(n8977), .A2(n8098), .ZN(n7653) );
  NAND2_X1 U9355 ( .A1(n4269), .A2(n9248), .ZN(n7652) );
  NAND2_X1 U9356 ( .A1(n7653), .A2(n7652), .ZN(n7654) );
  XNOR2_X1 U9357 ( .A(n7654), .B(n8063), .ZN(n7690) );
  NAND2_X1 U9358 ( .A1(n9605), .A2(n8098), .ZN(n7656) );
  NAND2_X1 U9359 ( .A1(n4269), .A2(n9249), .ZN(n7655) );
  NAND2_X1 U9360 ( .A1(n7656), .A2(n7655), .ZN(n7657) );
  XNOR2_X1 U9361 ( .A(n7657), .B(n8096), .ZN(n7663) );
  INV_X1 U9362 ( .A(n7663), .ZN(n7661) );
  NAND2_X1 U9363 ( .A1(n9605), .A2(n4269), .ZN(n7659) );
  NAND2_X1 U9364 ( .A1(n8073), .A2(n9249), .ZN(n7658) );
  NAND2_X1 U9365 ( .A1(n7659), .A2(n7658), .ZN(n7662) );
  INV_X1 U9366 ( .A(n7662), .ZN(n7660) );
  NAND2_X1 U9367 ( .A1(n7661), .A2(n7660), .ZN(n8883) );
  INV_X1 U9368 ( .A(n8883), .ZN(n7681) );
  NAND2_X1 U9369 ( .A1(n8830), .A2(n8098), .ZN(n7665) );
  NAND2_X1 U9370 ( .A1(n4269), .A2(n9250), .ZN(n7664) );
  NAND2_X1 U9371 ( .A1(n7665), .A2(n7664), .ZN(n7666) );
  XNOR2_X1 U9372 ( .A(n7666), .B(n8063), .ZN(n8821) );
  NOR2_X1 U9373 ( .A1(n6660), .A2(n8885), .ZN(n7667) );
  AOI21_X1 U9374 ( .B1(n8830), .B2(n4269), .A(n7667), .ZN(n7674) );
  AND2_X1 U9375 ( .A1(n8821), .A2(n7674), .ZN(n7680) );
  NAND2_X1 U9376 ( .A1(n8914), .A2(n8098), .ZN(n7669) );
  NAND2_X1 U9377 ( .A1(n4269), .A2(n9251), .ZN(n7668) );
  NAND2_X1 U9378 ( .A1(n7669), .A2(n7668), .ZN(n7670) );
  XNOR2_X1 U9379 ( .A(n7670), .B(n8063), .ZN(n7679) );
  INV_X1 U9380 ( .A(n7679), .ZN(n7673) );
  NOR2_X1 U9381 ( .A1(n6660), .A2(n9680), .ZN(n7671) );
  AOI21_X1 U9382 ( .B1(n8914), .B2(n4269), .A(n7671), .ZN(n7678) );
  INV_X1 U9383 ( .A(n7678), .ZN(n7672) );
  NAND2_X1 U9384 ( .A1(n7673), .A2(n7672), .ZN(n8819) );
  INV_X1 U9385 ( .A(n8821), .ZN(n7675) );
  INV_X1 U9386 ( .A(n7674), .ZN(n8820) );
  NAND2_X1 U9387 ( .A1(n7675), .A2(n8820), .ZN(n7676) );
  AND2_X1 U9388 ( .A1(n4293), .A2(n8879), .ZN(n8878) );
  AND2_X1 U9389 ( .A1(n7688), .A2(n7677), .ZN(n7685) );
  INV_X1 U9390 ( .A(n7677), .ZN(n7682) );
  XNOR2_X1 U9391 ( .A(n7679), .B(n7678), .ZN(n8911) );
  OR2_X1 U9392 ( .A1(n8911), .A2(n7680), .ZN(n8877) );
  OR2_X1 U9393 ( .A1(n7682), .A2(n8771), .ZN(n7683) );
  INV_X1 U9394 ( .A(n7683), .ZN(n7684) );
  NAND2_X1 U9395 ( .A1(n8977), .A2(n4269), .ZN(n7687) );
  NAND2_X1 U9396 ( .A1(n8073), .A2(n9248), .ZN(n7686) );
  NAND2_X1 U9397 ( .A1(n7687), .A2(n7686), .ZN(n8776) );
  INV_X1 U9398 ( .A(n7690), .ZN(n8774) );
  AND2_X1 U9399 ( .A1(n8771), .A2(n8774), .ZN(n7691) );
  NAND2_X1 U9400 ( .A1(n9599), .A2(n8098), .ZN(n7693) );
  NAND2_X1 U9401 ( .A1(n4269), .A2(n9247), .ZN(n7692) );
  NAND2_X1 U9402 ( .A1(n7693), .A2(n7692), .ZN(n7694) );
  XNOR2_X1 U9403 ( .A(n7694), .B(n8063), .ZN(n7997) );
  NOR2_X1 U9404 ( .A1(n6660), .A2(n9511), .ZN(n7695) );
  AOI21_X1 U9405 ( .B1(n9599), .B2(n4269), .A(n7695), .ZN(n7995) );
  INV_X1 U9406 ( .A(n7995), .ZN(n7998) );
  XNOR2_X1 U9407 ( .A(n7997), .B(n7998), .ZN(n7696) );
  XNOR2_X1 U9408 ( .A(n7996), .B(n7696), .ZN(n7702) );
  AND2_X1 U9409 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9818) );
  INV_X1 U9410 ( .A(n8936), .ZN(n8897) );
  NOR2_X1 U9411 ( .A1(n8897), .A2(n8976), .ZN(n7697) );
  AOI211_X1 U9412 ( .C1(n8942), .C2(n9498), .A(n9818), .B(n7697), .ZN(n7698)
         );
  OAI21_X1 U9413 ( .B1(n8926), .B2(n7699), .A(n7698), .ZN(n7700) );
  AOI21_X1 U9414 ( .B1(n9599), .B2(n8928), .A(n7700), .ZN(n7701) );
  OAI21_X1 U9415 ( .B1(n7702), .B2(n4653), .A(n7701), .ZN(P1_U3239) );
  NAND2_X1 U9416 ( .A1(n7728), .A2(n7703), .ZN(n7705) );
  OAI211_X1 U9417 ( .C1(n9641), .C2(n7706), .A(n7705), .B(n7704), .ZN(P1_U3326) );
  XOR2_X1 U9418 ( .A(n7707), .B(n7966), .Z(n7738) );
  XNOR2_X1 U9419 ( .A(n7708), .B(n7966), .ZN(n7712) );
  OR2_X1 U9420 ( .A1(n7709), .A2(n8267), .ZN(n7711) );
  NAND2_X1 U9421 ( .A1(n8309), .A2(n8269), .ZN(n7710) );
  NAND2_X1 U9422 ( .A1(n7711), .A2(n7710), .ZN(n8284) );
  AOI21_X1 U9423 ( .B1(n7712), .B2(n9968), .A(n8284), .ZN(n7732) );
  INV_X1 U9424 ( .A(n7732), .ZN(n7718) );
  OAI211_X1 U9425 ( .C1(n7714), .C2(n7713), .A(n10049), .B(n4271), .ZN(n7731)
         );
  AOI22_X1 U9426 ( .A1(n10011), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8283), .B2(
        n10001), .ZN(n7716) );
  NAND2_X1 U9427 ( .A1(n8291), .A2(n9990), .ZN(n7715) );
  OAI211_X1 U9428 ( .C1(n7731), .C2(n8588), .A(n7716), .B(n7715), .ZN(n7717)
         );
  AOI21_X1 U9429 ( .B1(n7718), .B2(n10009), .A(n7717), .ZN(n7719) );
  OAI21_X1 U9430 ( .B1(n7738), .B2(n8592), .A(n7719), .ZN(P2_U3281) );
  AND2_X1 U9431 ( .A1(n10120), .A2(n10097), .ZN(n8639) );
  AOI211_X1 U9432 ( .C1(n7722), .C2(n10069), .A(n7721), .B(n7720), .ZN(n7724)
         );
  MUX2_X1 U9433 ( .A(n8326), .B(n7724), .S(n10120), .Z(n7723) );
  OAI21_X1 U9434 ( .B1(n7727), .B2(n8672), .A(n7723), .ZN(P2_U3534) );
  AND2_X1 U9435 ( .A1(n10101), .A2(n10097), .ZN(n8716) );
  INV_X1 U9436 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7725) );
  MUX2_X1 U9437 ( .A(n7725), .B(n7724), .S(n10101), .Z(n7726) );
  OAI21_X1 U9438 ( .B1(n7727), .B2(n8750), .A(n7726), .ZN(P2_U3493) );
  INV_X1 U9439 ( .A(n7728), .ZN(n7729) );
  OAI222_X1 U9440 ( .A1(n4268), .A2(n7730), .B1(n8768), .B2(n7729), .C1(n6125), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  NAND2_X1 U9441 ( .A1(n7732), .A2(n7731), .ZN(n7735) );
  MUX2_X1 U9442 ( .A(n7735), .B(P2_REG1_REG_15__SCAN_IN), .S(n10117), .Z(n7733) );
  AOI21_X1 U9443 ( .B1(n8670), .B2(n8291), .A(n7733), .ZN(n7734) );
  OAI21_X1 U9444 ( .B1(n7738), .B2(n8672), .A(n7734), .ZN(P2_U3535) );
  MUX2_X1 U9445 ( .A(n7735), .B(P2_REG0_REG_15__SCAN_IN), .S(n10099), .Z(n7736) );
  AOI21_X1 U9446 ( .B1(n8748), .B2(n8291), .A(n7736), .ZN(n7737) );
  OAI21_X1 U9447 ( .B1(n7738), .B2(n8750), .A(n7737), .ZN(P2_U3496) );
  NAND2_X1 U9448 ( .A1(n7743), .A2(n7739), .ZN(n7741) );
  OAI211_X1 U9449 ( .C1(n4268), .C2(n7742), .A(n7741), .B(n7740), .ZN(P2_U3330) );
  INV_X1 U9450 ( .A(n7743), .ZN(n7746) );
  OAI222_X1 U9451 ( .A1(n9645), .A2(n7746), .B1(n7745), .B2(P1_U3084), .C1(
        n7744), .C2(n9641), .ZN(P1_U3325) );
  OAI21_X1 U9452 ( .B1(n7748), .B2(n7968), .A(n7747), .ZN(n7749) );
  INV_X1 U9453 ( .A(n7749), .ZN(n8751) );
  NAND2_X1 U9454 ( .A1(n7767), .A2(n7766), .ZN(n7752) );
  NAND2_X1 U9455 ( .A1(n7752), .A2(n7882), .ZN(n7750) );
  AOI21_X1 U9456 ( .B1(n7750), .B2(n7968), .A(n10000), .ZN(n7756) );
  NAND2_X1 U9457 ( .A1(n7752), .A2(n7751), .ZN(n7755) );
  NAND2_X1 U9458 ( .A1(n8307), .A2(n8269), .ZN(n7754) );
  NAND2_X1 U9459 ( .A1(n8309), .A2(n8251), .ZN(n7753) );
  NAND2_X1 U9460 ( .A1(n7754), .A2(n7753), .ZN(n8215) );
  AOI21_X1 U9461 ( .B1(n7756), .B2(n7755), .A(n8215), .ZN(n8668) );
  INV_X1 U9462 ( .A(n8668), .ZN(n7761) );
  INV_X1 U9463 ( .A(n8747), .ZN(n8221) );
  INV_X1 U9464 ( .A(n7757), .ZN(n7771) );
  OAI211_X1 U9465 ( .C1(n8221), .C2(n7771), .A(n8580), .B(n10049), .ZN(n8667)
         );
  AOI22_X1 U9466 ( .A1(n10011), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8218), .B2(
        n10001), .ZN(n7759) );
  NAND2_X1 U9467 ( .A1(n8747), .A2(n9990), .ZN(n7758) );
  OAI211_X1 U9468 ( .C1(n8667), .C2(n8588), .A(n7759), .B(n7758), .ZN(n7760)
         );
  AOI21_X1 U9469 ( .B1(n7761), .B2(n10009), .A(n7760), .ZN(n7762) );
  OAI21_X1 U9470 ( .B1(n8751), .B2(n8592), .A(n7762), .ZN(P2_U3279) );
  NOR2_X1 U9471 ( .A1(n7763), .A2(n7967), .ZN(n7764) );
  OR2_X1 U9472 ( .A1(n7765), .A2(n7764), .ZN(n8673) );
  XNOR2_X1 U9473 ( .A(n7767), .B(n7766), .ZN(n7769) );
  OAI22_X1 U9474 ( .A1(n7768), .A2(n8267), .B1(n8268), .B2(n8249), .ZN(n8139)
         );
  AOI21_X1 U9475 ( .B1(n7769), .B2(n9968), .A(n8139), .ZN(n7770) );
  OAI21_X1 U9476 ( .B1(n8673), .B2(n9955), .A(n7770), .ZN(n8674) );
  NAND2_X1 U9477 ( .A1(n8674), .A2(n10009), .ZN(n7775) );
  AOI211_X1 U9478 ( .C1(n8143), .C2(n4271), .A(n10086), .B(n7771), .ZN(n8675)
         );
  INV_X1 U9479 ( .A(n8143), .ZN(n8756) );
  AOI22_X1 U9480 ( .A1(n10011), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8138), .B2(
        n10001), .ZN(n7772) );
  OAI21_X1 U9481 ( .B1(n8756), .B2(n10004), .A(n7772), .ZN(n7773) );
  AOI21_X1 U9482 ( .B1(n8675), .B2(n9993), .A(n7773), .ZN(n7774) );
  OAI211_X1 U9483 ( .C1(n8673), .C2(n7776), .A(n7775), .B(n7774), .ZN(P2_U3280) );
  INV_X1 U9484 ( .A(n7777), .ZN(n8134) );
  OAI222_X1 U9485 ( .A1(n9641), .A2(n7778), .B1(n9645), .B2(n8134), .C1(n6414), 
        .C2(P1_U3084), .ZN(P1_U3331) );
  NAND2_X1 U9486 ( .A1(n7779), .A2(n7925), .ZN(n7780) );
  NAND2_X1 U9487 ( .A1(n7780), .A2(n7926), .ZN(n7789) );
  NAND2_X1 U9488 ( .A1(n7782), .A2(n7781), .ZN(n7784) );
  NAND2_X1 U9489 ( .A1(n7784), .A2(n7783), .ZN(n7785) );
  MUX2_X1 U9490 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n7794), .Z(n7791) );
  NAND2_X1 U9491 ( .A1(n8763), .A2(n5706), .ZN(n7788) );
  OR2_X1 U9492 ( .A1(n7798), .A2(n8765), .ZN(n7787) );
  NOR2_X1 U9493 ( .A1(n8420), .A2(n7800), .ZN(n7934) );
  NAND2_X1 U9494 ( .A1(n7792), .A2(n7791), .ZN(n7793) );
  MUX2_X1 U9495 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7794), .Z(n7795) );
  XNOR2_X1 U9496 ( .A(n7795), .B(SI_31_), .ZN(n7796) );
  NOR2_X1 U9497 ( .A1(n7798), .A2(n6250), .ZN(n7799) );
  NAND2_X1 U9498 ( .A1(n8420), .A2(n7800), .ZN(n7930) );
  NOR2_X1 U9499 ( .A1(n8689), .A2(n8414), .ZN(n7941) );
  NAND2_X1 U9500 ( .A1(n5643), .A2(n7801), .ZN(n7987) );
  NAND2_X1 U9501 ( .A1(n7980), .A2(n8480), .ZN(n7802) );
  INV_X1 U9502 ( .A(n7807), .ZN(n7904) );
  NOR2_X1 U9503 ( .A1(n8300), .A2(n7807), .ZN(n7911) );
  INV_X1 U9504 ( .A(n7803), .ZN(n7804) );
  MUX2_X1 U9505 ( .A(n7805), .B(n7804), .S(n7807), .Z(n7879) );
  NAND2_X1 U9506 ( .A1(n7811), .A2(n7806), .ZN(n7808) );
  MUX2_X1 U9507 ( .A(n7808), .B(n7829), .S(n7807), .Z(n7817) );
  INV_X1 U9508 ( .A(n7808), .ZN(n7810) );
  AOI22_X1 U9509 ( .A1(n7817), .A2(n7811), .B1(n7810), .B2(n7809), .ZN(n7813)
         );
  OAI21_X1 U9510 ( .B1(n7813), .B2(n7812), .A(n7807), .ZN(n7827) );
  AOI21_X1 U9511 ( .B1(n7980), .B2(n7949), .A(n7814), .ZN(n7816) );
  NAND2_X1 U9512 ( .A1(n6093), .A2(n7819), .ZN(n7815) );
  OAI211_X1 U9513 ( .C1(n7816), .C2(n7815), .A(n7821), .B(n7807), .ZN(n7818)
         );
  INV_X1 U9514 ( .A(n7817), .ZN(n7835) );
  NAND3_X1 U9515 ( .A1(n7818), .A2(n7835), .A3(n6862), .ZN(n7826) );
  INV_X1 U9516 ( .A(n7819), .ZN(n7820) );
  NOR2_X1 U9517 ( .A1(n7820), .A2(n7807), .ZN(n7825) );
  INV_X1 U9518 ( .A(n6093), .ZN(n7823) );
  OAI211_X1 U9519 ( .C1(n7823), .C2(n7822), .A(n7821), .B(n6092), .ZN(n7824)
         );
  AOI22_X1 U9520 ( .A1(n7827), .A2(n7826), .B1(n7825), .B2(n7824), .ZN(n7840)
         );
  INV_X1 U9521 ( .A(n7828), .ZN(n7834) );
  OAI21_X1 U9522 ( .B1(n7832), .B2(n7831), .A(n7830), .ZN(n7833) );
  OAI21_X1 U9523 ( .B1(n7835), .B2(n7834), .A(n7833), .ZN(n7836) );
  AOI21_X1 U9524 ( .B1(n7836), .B2(n7837), .A(n7807), .ZN(n7839) );
  MUX2_X1 U9525 ( .A(n9965), .B(n7837), .S(n7807), .Z(n7838) );
  MUX2_X1 U9526 ( .A(n7842), .B(n7841), .S(n7807), .Z(n7843) );
  MUX2_X1 U9527 ( .A(n7845), .B(n7844), .S(n7807), .Z(n7846) );
  NAND3_X1 U9528 ( .A1(n7850), .A2(n7904), .A3(n7852), .ZN(n7848) );
  OAI21_X1 U9529 ( .B1(n7959), .B2(n6062), .A(n7848), .ZN(n7857) );
  NAND2_X1 U9530 ( .A1(n7859), .A2(n7849), .ZN(n7855) );
  INV_X1 U9531 ( .A(n7849), .ZN(n7853) );
  OAI211_X1 U9532 ( .C1(n7853), .C2(n7852), .A(n7851), .B(n7850), .ZN(n7854)
         );
  MUX2_X1 U9533 ( .A(n7855), .B(n7854), .S(n7807), .Z(n7856) );
  INV_X1 U9534 ( .A(n7858), .ZN(n7861) );
  NAND2_X1 U9535 ( .A1(n7863), .A2(n7859), .ZN(n7860) );
  MUX2_X1 U9536 ( .A(n7861), .B(n7860), .S(n7807), .Z(n7865) );
  MUX2_X1 U9537 ( .A(n7863), .B(n7862), .S(n7807), .Z(n7864) );
  OAI211_X1 U9538 ( .C1(n7866), .C2(n7865), .A(n7962), .B(n7864), .ZN(n7878)
         );
  NOR2_X1 U9539 ( .A1(n8680), .A2(n7807), .ZN(n7870) );
  NOR2_X1 U9540 ( .A1(n7867), .A2(n7904), .ZN(n7869) );
  MUX2_X1 U9541 ( .A(n7870), .B(n7869), .S(n7868), .Z(n7871) );
  NOR2_X1 U9542 ( .A1(n7946), .A2(n7871), .ZN(n7877) );
  INV_X1 U9543 ( .A(n7872), .ZN(n7875) );
  INV_X1 U9544 ( .A(n7873), .ZN(n7874) );
  MUX2_X1 U9545 ( .A(n7875), .B(n7874), .S(n7807), .Z(n7876) );
  OAI211_X1 U9546 ( .C1(n7968), .C2(n7882), .A(n7887), .B(n7881), .ZN(n7884)
         );
  MUX2_X1 U9547 ( .A(n7884), .B(n7883), .S(n7807), .Z(n7885) );
  OAI21_X1 U9548 ( .B1(n7895), .B2(n4561), .A(n7896), .ZN(n7888) );
  NAND3_X1 U9549 ( .A1(n7888), .A2(n7900), .A3(n8545), .ZN(n7889) );
  NAND2_X1 U9550 ( .A1(n8533), .A2(n8304), .ZN(n7902) );
  NAND3_X1 U9551 ( .A1(n7889), .A2(n7897), .A3(n7902), .ZN(n7891) );
  AOI21_X1 U9552 ( .B1(n7892), .B2(n7807), .A(n8500), .ZN(n7894) );
  NAND3_X1 U9553 ( .A1(n7898), .A2(n7897), .A3(n7896), .ZN(n7901) );
  NAND3_X1 U9554 ( .A1(n7901), .A2(n7900), .A3(n7899), .ZN(n7903) );
  AOI21_X1 U9555 ( .B1(n7908), .B2(n7906), .A(n7807), .ZN(n7907) );
  AOI211_X1 U9556 ( .C1(n7911), .C2(n8636), .A(n7910), .B(n7909), .ZN(n7919)
         );
  NAND2_X1 U9557 ( .A1(n7915), .A2(n8457), .ZN(n7914) );
  NAND2_X1 U9558 ( .A1(n8456), .A2(n7912), .ZN(n7913) );
  MUX2_X1 U9559 ( .A(n7914), .B(n7913), .S(n7807), .Z(n7918) );
  INV_X1 U9560 ( .A(n8439), .ZN(n8437) );
  MUX2_X1 U9561 ( .A(n7916), .B(n7915), .S(n7807), .Z(n7917) );
  OAI211_X1 U9562 ( .C1(n7919), .C2(n7918), .A(n8437), .B(n7917), .ZN(n7924)
         );
  AOI22_X1 U9563 ( .A1(n8616), .A2(n7927), .B1(n8162), .B2(n8699), .ZN(n7920)
         );
  MUX2_X1 U9564 ( .A(n7921), .B(n7920), .S(n7807), .Z(n7923) );
  AND3_X1 U9565 ( .A1(n7924), .A2(n7923), .A3(n7922), .ZN(n7929) );
  MUX2_X1 U9566 ( .A(n7807), .B(n7927), .S(n8616), .Z(n7928) );
  NOR2_X1 U9567 ( .A1(n7974), .A2(n7928), .ZN(n7933) );
  INV_X1 U9568 ( .A(n7929), .ZN(n7932) );
  INV_X1 U9569 ( .A(n7930), .ZN(n7931) );
  AOI211_X1 U9570 ( .C1(n7933), .C2(n7932), .A(n7931), .B(n7934), .ZN(n7938)
         );
  INV_X1 U9571 ( .A(n7934), .ZN(n7935) );
  NAND2_X1 U9572 ( .A1(n4578), .A2(n7935), .ZN(n7944) );
  INV_X1 U9573 ( .A(n7939), .ZN(n7940) );
  MUX2_X1 U9574 ( .A(n7941), .B(n7940), .S(n7807), .Z(n7942) );
  OAI21_X1 U9575 ( .B1(n7943), .B2(n7942), .A(n7947), .ZN(n7985) );
  INV_X1 U9576 ( .A(n7944), .ZN(n7977) );
  INV_X1 U9577 ( .A(n8427), .ZN(n8424) );
  INV_X1 U9578 ( .A(n7945), .ZN(n8544) );
  INV_X1 U9579 ( .A(n8561), .ZN(n7970) );
  NOR2_X1 U9580 ( .A1(n8558), .A2(n4561), .ZN(n8575) );
  NOR3_X1 U9581 ( .A1(n7948), .A2(n6097), .A3(n7947), .ZN(n7952) );
  INV_X1 U9582 ( .A(n7092), .ZN(n7951) );
  AND2_X1 U9583 ( .A1(n7950), .A2(n7949), .ZN(n10002) );
  NAND3_X1 U9584 ( .A1(n7952), .A2(n7951), .A3(n10002), .ZN(n7955) );
  NOR3_X1 U9585 ( .A1(n7955), .A2(n7954), .A3(n7953), .ZN(n7958) );
  NAND4_X1 U9586 ( .A1(n7958), .A2(n7957), .A3(n7956), .A4(n8600), .ZN(n7961)
         );
  NOR4_X1 U9587 ( .A1(n7961), .A2(n7960), .A3(n7959), .A4(n6062), .ZN(n7963)
         );
  NAND4_X1 U9588 ( .A1(n4516), .A2(n7964), .A3(n7963), .A4(n7962), .ZN(n7965)
         );
  NOR4_X1 U9589 ( .A1(n7968), .A2(n7967), .A3(n7966), .A4(n7965), .ZN(n7969)
         );
  NAND4_X1 U9590 ( .A1(n8544), .A2(n7970), .A3(n8575), .A4(n7969), .ZN(n7971)
         );
  NOR4_X1 U9591 ( .A1(n8500), .A2(n8528), .A3(n8514), .A4(n7971), .ZN(n7972)
         );
  NAND4_X1 U9592 ( .A1(n8456), .A2(n8471), .A3(n8489), .A4(n7972), .ZN(n7973)
         );
  NOR4_X1 U9593 ( .A1(n7974), .A2(n8424), .A3(n8439), .A4(n7973), .ZN(n7975)
         );
  NAND3_X1 U9594 ( .A1(n7977), .A2(n7976), .A3(n7975), .ZN(n7978) );
  XNOR2_X1 U9595 ( .A(n7978), .B(n8405), .ZN(n7981) );
  OAI22_X1 U9596 ( .A1(n7981), .A2(n7980), .B1(n7979), .B2(n7983), .ZN(n7982)
         );
  INV_X1 U9597 ( .A(n7983), .ZN(n7984) );
  NOR3_X1 U9598 ( .A1(n7985), .A2(n7984), .A3(n4415), .ZN(n7986) );
  NAND4_X1 U9599 ( .A1(n10013), .A2(n7989), .A3(n8251), .A4(n7988), .ZN(n7990)
         );
  OAI211_X1 U9600 ( .C1(n7991), .C2(n7993), .A(n7990), .B(P2_B_REG_SCAN_IN), 
        .ZN(n7992) );
  OAI21_X1 U9601 ( .B1(n7994), .B2(n7993), .A(n7992), .ZN(P2_U3244) );
  INV_X1 U9602 ( .A(n7997), .ZN(n7999) );
  NAND2_X1 U9603 ( .A1(n7999), .A2(n7998), .ZN(n8000) );
  NAND2_X1 U9604 ( .A1(n8001), .A2(n8000), .ZN(n8840) );
  INV_X1 U9605 ( .A(n8840), .ZN(n8013) );
  NAND2_X1 U9606 ( .A1(n9594), .A2(n8098), .ZN(n8003) );
  NAND2_X1 U9607 ( .A1(n4269), .A2(n9498), .ZN(n8002) );
  NAND2_X1 U9608 ( .A1(n8003), .A2(n8002), .ZN(n8004) );
  XNOR2_X1 U9609 ( .A(n8004), .B(n8063), .ZN(n8007) );
  NOR2_X1 U9610 ( .A1(n6660), .A2(n8005), .ZN(n8006) );
  AOI21_X1 U9611 ( .B1(n9594), .B2(n4269), .A(n8006), .ZN(n8008) );
  NAND2_X1 U9612 ( .A1(n8007), .A2(n8008), .ZN(n8014) );
  INV_X1 U9613 ( .A(n8007), .ZN(n8010) );
  INV_X1 U9614 ( .A(n8008), .ZN(n8009) );
  NAND2_X1 U9615 ( .A1(n8010), .A2(n8009), .ZN(n8011) );
  NAND2_X1 U9616 ( .A1(n8014), .A2(n8011), .ZN(n8843) );
  NAND2_X1 U9617 ( .A1(n9587), .A2(n8098), .ZN(n8016) );
  NAND2_X1 U9618 ( .A1(n4269), .A2(n9471), .ZN(n8015) );
  NAND2_X1 U9619 ( .A1(n8016), .A2(n8015), .ZN(n8017) );
  XNOR2_X1 U9620 ( .A(n8017), .B(n8096), .ZN(n8019) );
  NOR2_X1 U9621 ( .A1(n6660), .A2(n9512), .ZN(n8018) );
  AOI21_X1 U9622 ( .B1(n9587), .B2(n4269), .A(n8018), .ZN(n8020) );
  XNOR2_X1 U9623 ( .A(n8019), .B(n8020), .ZN(n8851) );
  INV_X1 U9624 ( .A(n8019), .ZN(n8021) );
  NAND2_X1 U9625 ( .A1(n8021), .A2(n8020), .ZN(n8022) );
  NAND2_X1 U9626 ( .A1(n9575), .A2(n8098), .ZN(n8024) );
  NAND2_X1 U9627 ( .A1(n9472), .A2(n4269), .ZN(n8023) );
  NAND2_X1 U9628 ( .A1(n8024), .A2(n8023), .ZN(n8025) );
  XNOR2_X1 U9629 ( .A(n8025), .B(n8096), .ZN(n8034) );
  NAND2_X1 U9630 ( .A1(n9575), .A2(n4269), .ZN(n8027) );
  NAND2_X1 U9631 ( .A1(n9472), .A2(n8073), .ZN(n8026) );
  NAND2_X1 U9632 ( .A1(n8027), .A2(n8026), .ZN(n8035) );
  NAND2_X1 U9633 ( .A1(n8034), .A2(n8035), .ZN(n8800) );
  NAND2_X1 U9634 ( .A1(n9582), .A2(n8098), .ZN(n8029) );
  NAND2_X1 U9635 ( .A1(n9500), .A2(n4269), .ZN(n8028) );
  NAND2_X1 U9636 ( .A1(n8029), .A2(n8028), .ZN(n8030) );
  XNOR2_X1 U9637 ( .A(n8030), .B(n8063), .ZN(n8798) );
  INV_X1 U9638 ( .A(n8798), .ZN(n8796) );
  AND2_X1 U9639 ( .A1(n8073), .A2(n9500), .ZN(n8031) );
  AOI21_X1 U9640 ( .B1(n9582), .B2(n4269), .A(n8031), .ZN(n8917) );
  INV_X1 U9641 ( .A(n8917), .ZN(n8032) );
  NAND2_X1 U9642 ( .A1(n8796), .A2(n8032), .ZN(n8033) );
  AND2_X1 U9643 ( .A1(n8800), .A2(n8033), .ZN(n8039) );
  NAND3_X1 U9644 ( .A1(n8800), .A2(n8917), .A3(n8798), .ZN(n8038) );
  INV_X1 U9645 ( .A(n8034), .ZN(n8037) );
  INV_X1 U9646 ( .A(n8035), .ZN(n8036) );
  NAND2_X1 U9647 ( .A1(n8037), .A2(n8036), .ZN(n8866) );
  NAND2_X1 U9648 ( .A1(n9570), .A2(n8098), .ZN(n8041) );
  NAND2_X1 U9649 ( .A1(n9463), .A2(n4269), .ZN(n8040) );
  NAND2_X1 U9650 ( .A1(n8041), .A2(n8040), .ZN(n8042) );
  XNOR2_X1 U9651 ( .A(n8042), .B(n8063), .ZN(n8044) );
  AND2_X1 U9652 ( .A1(n9463), .A2(n8073), .ZN(n8043) );
  AOI21_X1 U9653 ( .B1(n9570), .B2(n4269), .A(n8043), .ZN(n8045) );
  NAND2_X1 U9654 ( .A1(n8044), .A2(n8045), .ZN(n8051) );
  INV_X1 U9655 ( .A(n8044), .ZN(n8047) );
  INV_X1 U9656 ( .A(n8045), .ZN(n8046) );
  NAND2_X1 U9657 ( .A1(n8047), .A2(n8046), .ZN(n8048) );
  NAND2_X1 U9658 ( .A1(n8051), .A2(n8048), .ZN(n8867) );
  INV_X1 U9659 ( .A(n8867), .ZN(n8049) );
  NAND2_X1 U9660 ( .A1(n8050), .A2(n8049), .ZN(n8868) );
  NAND2_X1 U9661 ( .A1(n8868), .A2(n8051), .ZN(n8809) );
  NAND2_X1 U9662 ( .A1(n9429), .A2(n8098), .ZN(n8053) );
  NAND2_X1 U9663 ( .A1(n9447), .A2(n4269), .ZN(n8052) );
  NAND2_X1 U9664 ( .A1(n8053), .A2(n8052), .ZN(n8054) );
  XNOR2_X1 U9665 ( .A(n8054), .B(n8096), .ZN(n8056) );
  AND2_X1 U9666 ( .A1(n9447), .A2(n8073), .ZN(n8055) );
  AOI21_X1 U9667 ( .B1(n9429), .B2(n4269), .A(n8055), .ZN(n8057) );
  XNOR2_X1 U9668 ( .A(n8056), .B(n8057), .ZN(n8810) );
  NAND2_X1 U9669 ( .A1(n8809), .A2(n8810), .ZN(n8808) );
  INV_X1 U9670 ( .A(n8056), .ZN(n8058) );
  NAND2_X1 U9671 ( .A1(n8058), .A2(n8057), .ZN(n8059) );
  AND2_X1 U9672 ( .A1(n9426), .A2(n8073), .ZN(n8060) );
  AOI21_X1 U9673 ( .B1(n9560), .B2(n4269), .A(n8060), .ZN(n8066) );
  NAND2_X1 U9674 ( .A1(n9560), .A2(n8098), .ZN(n8062) );
  NAND2_X1 U9675 ( .A1(n9426), .A2(n4269), .ZN(n8061) );
  NAND2_X1 U9676 ( .A1(n8062), .A2(n8061), .ZN(n8064) );
  XNOR2_X1 U9677 ( .A(n8064), .B(n8063), .ZN(n8892) );
  INV_X1 U9678 ( .A(n8066), .ZN(n8067) );
  NAND2_X1 U9679 ( .A1(n9555), .A2(n8098), .ZN(n8069) );
  NAND2_X1 U9680 ( .A1(n9246), .A2(n4269), .ZN(n8068) );
  NAND2_X1 U9681 ( .A1(n8069), .A2(n8068), .ZN(n8070) );
  XNOR2_X1 U9682 ( .A(n8070), .B(n8096), .ZN(n8071) );
  AOI22_X1 U9683 ( .A1(n9555), .A2(n4269), .B1(n8073), .B2(n9246), .ZN(n8789)
         );
  AOI22_X1 U9684 ( .A1(n9550), .A2(n8098), .B1(n4269), .B2(n9394), .ZN(n8072)
         );
  XNOR2_X1 U9685 ( .A(n8072), .B(n8096), .ZN(n8075) );
  AOI22_X1 U9686 ( .A1(n9550), .A2(n4269), .B1(n8073), .B2(n9394), .ZN(n8074)
         );
  NAND2_X1 U9687 ( .A1(n8075), .A2(n8074), .ZN(n8076) );
  OAI21_X1 U9688 ( .B1(n8075), .B2(n8074), .A(n8076), .ZN(n8860) );
  INV_X1 U9689 ( .A(n8076), .ZN(n8077) );
  AOI22_X1 U9690 ( .A1(n9543), .A2(n4269), .B1(n8073), .B2(n9355), .ZN(n8081)
         );
  NAND2_X1 U9691 ( .A1(n9543), .A2(n8098), .ZN(n8079) );
  NAND2_X1 U9692 ( .A1(n9355), .A2(n4269), .ZN(n8078) );
  NAND2_X1 U9693 ( .A1(n8079), .A2(n8078), .ZN(n8080) );
  XNOR2_X1 U9694 ( .A(n8080), .B(n8096), .ZN(n8083) );
  XOR2_X1 U9695 ( .A(n8081), .B(n8083), .Z(n8833) );
  INV_X1 U9696 ( .A(n8081), .ZN(n8082) );
  AND2_X1 U9697 ( .A1(n9372), .A2(n8073), .ZN(n8084) );
  AOI21_X1 U9698 ( .B1(n9538), .B2(n4269), .A(n8084), .ZN(n8088) );
  NAND2_X1 U9699 ( .A1(n9538), .A2(n8098), .ZN(n8086) );
  NAND2_X1 U9700 ( .A1(n9372), .A2(n4269), .ZN(n8085) );
  NAND2_X1 U9701 ( .A1(n8086), .A2(n8085), .ZN(n8087) );
  XNOR2_X1 U9702 ( .A(n8087), .B(n8096), .ZN(n8090) );
  XOR2_X1 U9703 ( .A(n8088), .B(n8090), .Z(n8931) );
  INV_X1 U9704 ( .A(n8088), .ZN(n8089) );
  AOI22_X1 U9705 ( .A1(n9535), .A2(n8098), .B1(n4269), .B2(n9356), .ZN(n8091)
         );
  XNOR2_X1 U9706 ( .A(n8091), .B(n8096), .ZN(n8093) );
  AOI22_X1 U9707 ( .A1(n9535), .A2(n4269), .B1(n8073), .B2(n9356), .ZN(n8092)
         );
  NAND2_X1 U9708 ( .A1(n8093), .A2(n8092), .ZN(n8105) );
  OAI21_X1 U9709 ( .B1(n8093), .B2(n8092), .A(n8105), .ZN(n8150) );
  NAND2_X1 U9710 ( .A1(n9530), .A2(n4269), .ZN(n8095) );
  NAND2_X1 U9711 ( .A1(n9245), .A2(n8073), .ZN(n8094) );
  NAND2_X1 U9712 ( .A1(n8095), .A2(n8094), .ZN(n8097) );
  XNOR2_X1 U9713 ( .A(n8097), .B(n8096), .ZN(n8100) );
  AOI22_X1 U9714 ( .A1(n9530), .A2(n8098), .B1(n4269), .B2(n9245), .ZN(n8099)
         );
  XNOR2_X1 U9715 ( .A(n8100), .B(n8099), .ZN(n8101) );
  INV_X1 U9716 ( .A(n8101), .ZN(n8106) );
  NAND3_X1 U9717 ( .A1(n8106), .A2(n8935), .A3(n8105), .ZN(n8111) );
  NAND3_X1 U9718 ( .A1(n4290), .A2(n8935), .A3(n8101), .ZN(n8110) );
  INV_X1 U9719 ( .A(n8102), .ZN(n9323) );
  AOI22_X1 U9720 ( .A1(n9323), .A2(n8937), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8104) );
  NAND2_X1 U9721 ( .A1(n9356), .A2(n8936), .ZN(n8103) );
  OAI211_X1 U9722 ( .C1(n9321), .C2(n8923), .A(n8104), .B(n8103), .ZN(n8108)
         );
  NOR3_X1 U9723 ( .A1(n8106), .A2(n4653), .A3(n8105), .ZN(n8107) );
  AOI211_X1 U9724 ( .C1(n8928), .C2(n9530), .A(n8108), .B(n8107), .ZN(n8109)
         );
  OAI211_X1 U9725 ( .C1(n4290), .C2(n8111), .A(n8110), .B(n8109), .ZN(P1_U3218) );
  NAND2_X1 U9726 ( .A1(n8758), .A2(n8114), .ZN(n8113) );
  OR2_X1 U9727 ( .A1(n8115), .A2(n6369), .ZN(n8112) );
  NAND2_X1 U9728 ( .A1(n8763), .A2(n8114), .ZN(n8117) );
  INV_X1 U9729 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9640) );
  OR2_X1 U9730 ( .A1(n8115), .A2(n9640), .ZN(n8116) );
  NAND2_X1 U9731 ( .A1(n8119), .A2(n8118), .ZN(n9710) );
  NOR2_X1 U9732 ( .A1(n9692), .A2(n9710), .ZN(n9299) );
  AOI21_X1 U9733 ( .B1(n9887), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9299), .ZN(
        n8121) );
  NAND2_X1 U9734 ( .A1(n9525), .A2(n9693), .ZN(n8120) );
  OAI211_X1 U9735 ( .C1(n9527), .C2(n9308), .A(n8121), .B(n8120), .ZN(P1_U3261) );
  NAND2_X1 U9736 ( .A1(n8127), .A2(n8639), .ZN(n8126) );
  NAND2_X1 U9737 ( .A1(n8123), .A2(n8122), .ZN(n8128) );
  NAND2_X1 U9738 ( .A1(n8126), .A2(n8125), .ZN(P2_U3549) );
  NAND2_X1 U9739 ( .A1(n8127), .A2(n8716), .ZN(n8132) );
  NAND2_X1 U9740 ( .A1(n8132), .A2(n8131), .ZN(P2_U3517) );
  OAI222_X1 U9741 ( .A1(n4268), .A2(n8135), .B1(n8768), .B2(n8134), .C1(n4262), 
        .C2(n8133), .ZN(P2_U3336) );
  OAI222_X1 U9742 ( .A1(n4268), .A2(n8137), .B1(n8768), .B2(n8136), .C1(
        P2_U3152), .C2(n8405), .ZN(P2_U3339) );
  INV_X1 U9743 ( .A(n8138), .ZN(n8141) );
  NAND2_X1 U9744 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n8345) );
  NAND2_X1 U9745 ( .A1(n8285), .A2(n8139), .ZN(n8140) );
  OAI211_X1 U9746 ( .C1(n8287), .C2(n8141), .A(n8345), .B(n8140), .ZN(n8142)
         );
  AOI21_X1 U9747 ( .B1(n8143), .B2(n8290), .A(n8142), .ZN(n8148) );
  NAND2_X1 U9748 ( .A1(n8244), .A2(n8310), .ZN(n8294) );
  OAI21_X1 U9749 ( .B1(n8280), .B2(n8259), .A(n8294), .ZN(n8146) );
  INV_X1 U9750 ( .A(n8144), .ZN(n8145) );
  NAND3_X1 U9751 ( .A1(n8146), .A2(n8145), .A3(n8279), .ZN(n8147) );
  OAI211_X1 U9752 ( .C1(n8149), .C2(n8259), .A(n8148), .B(n8147), .ZN(P2_U3228) );
  INV_X1 U9753 ( .A(n9341), .ZN(n8153) );
  AOI22_X1 U9754 ( .A1(n9372), .A2(n8936), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n8152) );
  OAI21_X1 U9755 ( .B1(n8926), .B2(n8153), .A(n8152), .ZN(n8154) );
  AOI21_X1 U9756 ( .B1(n8942), .B2(n9245), .A(n8154), .ZN(n8155) );
  AOI21_X1 U9757 ( .B1(n8156), .B2(n8157), .A(n8259), .ZN(n8161) );
  NOR3_X1 U9758 ( .A1(n8159), .A2(n8158), .A3(n8262), .ZN(n8160) );
  NOR2_X1 U9759 ( .A1(n8161), .A2(n8160), .ZN(n8167) );
  INV_X1 U9760 ( .A(n8162), .ZN(n8297) );
  AOI22_X1 U9761 ( .A1(n8297), .A2(n8269), .B1(n8251), .B2(n8299), .ZN(n8460)
         );
  INV_X1 U9762 ( .A(n8464), .ZN(n8163) );
  AOI22_X1 U9763 ( .A1(n8163), .A2(n8275), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n8164) );
  OAI21_X1 U9764 ( .B1(n8460), .B2(n8273), .A(n8164), .ZN(n8165) );
  AOI21_X1 U9765 ( .B1(n8626), .B2(n8290), .A(n8165), .ZN(n8166) );
  OAI21_X1 U9766 ( .B1(n8167), .B2(n6139), .A(n8166), .ZN(P2_U3242) );
  AOI22_X1 U9767 ( .A1(n8169), .A2(n8282), .B1(n8244), .B2(n8301), .ZN(n8174)
         );
  INV_X1 U9768 ( .A(n8507), .ZN(n8171) );
  OAI22_X1 U9769 ( .A1(n8226), .A2(n8249), .B1(n8196), .B2(n8267), .ZN(n8502)
         );
  AOI22_X1 U9770 ( .A1(n8502), .A2(n8285), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        n4262), .ZN(n8170) );
  OAI21_X1 U9771 ( .B1(n8171), .B2(n8287), .A(n8170), .ZN(n8172) );
  AOI21_X1 U9772 ( .B1(n8715), .B2(n8290), .A(n8172), .ZN(n8173) );
  OAI21_X1 U9773 ( .B1(n8174), .B2(n8223), .A(n8173), .ZN(P2_U3218) );
  INV_X1 U9774 ( .A(n8264), .ZN(n8178) );
  NOR3_X1 U9775 ( .A1(n8176), .A2(n8175), .A3(n8262), .ZN(n8177) );
  AOI21_X1 U9776 ( .B1(n8178), .B2(n8282), .A(n8177), .ZN(n8188) );
  INV_X1 U9777 ( .A(n8568), .ZN(n8182) );
  NAND2_X1 U9778 ( .A1(n4262), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8408) );
  OR2_X1 U9779 ( .A1(n8197), .A2(n8249), .ZN(n8180) );
  NAND2_X1 U9780 ( .A1(n8307), .A2(n8251), .ZN(n8179) );
  NAND2_X1 U9781 ( .A1(n8180), .A2(n8179), .ZN(n8564) );
  NAND2_X1 U9782 ( .A1(n8285), .A2(n8564), .ZN(n8181) );
  OAI211_X1 U9783 ( .C1(n8287), .C2(n8182), .A(n8408), .B(n8181), .ZN(n8185)
         );
  NOR2_X1 U9784 ( .A1(n8183), .A2(n8259), .ZN(n8184) );
  AOI211_X1 U9785 ( .C1(n8290), .C2(n8737), .A(n8185), .B(n8184), .ZN(n8186)
         );
  OAI21_X1 U9786 ( .B1(n8188), .B2(n8187), .A(n8186), .ZN(P2_U3221) );
  OR2_X1 U9787 ( .A1(n8237), .A2(n8236), .ZN(n8238) );
  AOI21_X1 U9788 ( .B1(n8238), .B2(n8189), .A(n8259), .ZN(n8195) );
  NOR3_X1 U9789 ( .A1(n8190), .A2(n8197), .A3(n8262), .ZN(n8194) );
  AND2_X1 U9790 ( .A1(n8192), .A2(n8191), .ZN(n8193) );
  OAI21_X1 U9791 ( .B1(n8195), .B2(n8194), .A(n8193), .ZN(n8203) );
  OR2_X1 U9792 ( .A1(n8196), .A2(n8249), .ZN(n8199) );
  OR2_X1 U9793 ( .A1(n8197), .A2(n8267), .ZN(n8198) );
  NAND2_X1 U9794 ( .A1(n8199), .A2(n8198), .ZN(n8530) );
  AOI22_X1 U9795 ( .A1(n8285), .A2(n8530), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3152), .ZN(n8200) );
  OAI21_X1 U9796 ( .B1(n8534), .B2(n8287), .A(n8200), .ZN(n8201) );
  AOI21_X1 U9797 ( .B1(n8728), .B2(n8290), .A(n8201), .ZN(n8202) );
  NAND2_X1 U9798 ( .A1(n8203), .A2(n8202), .ZN(P2_U3225) );
  OAI211_X1 U9799 ( .C1(n8205), .C2(n8204), .A(n8156), .B(n8282), .ZN(n8210)
         );
  NOR2_X1 U9800 ( .A1(n8226), .A2(n8267), .ZN(n8206) );
  AOI21_X1 U9801 ( .B1(n8298), .B2(n8269), .A(n8206), .ZN(n8472) );
  OAI22_X1 U9802 ( .A1(n8472), .A2(n8273), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8207), .ZN(n8208) );
  AOI21_X1 U9803 ( .B1(n8477), .B2(n8275), .A(n8208), .ZN(n8209) );
  OAI211_X1 U9804 ( .C1(n8211), .C2(n8278), .A(n8210), .B(n8209), .ZN(P2_U3227) );
  AOI21_X1 U9805 ( .B1(n8213), .B2(n8212), .A(n8259), .ZN(n8214) );
  NAND2_X1 U9806 ( .A1(n8214), .A2(n8261), .ZN(n8220) );
  INV_X1 U9807 ( .A(n8215), .ZN(n8216) );
  OAI22_X1 U9808 ( .A1(n8273), .A2(n8216), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8363), .ZN(n8217) );
  AOI21_X1 U9809 ( .B1(n8218), .B2(n8275), .A(n8217), .ZN(n8219) );
  OAI211_X1 U9810 ( .C1(n8221), .C2(n8278), .A(n8220), .B(n8219), .ZN(P2_U3230) );
  XNOR2_X1 U9811 ( .A(n8225), .B(n8224), .ZN(n8229) );
  OAI22_X1 U9812 ( .A1(n8229), .A2(n8259), .B1(n8226), .B2(n8262), .ZN(n8227)
         );
  OAI21_X1 U9813 ( .B1(n8229), .B2(n8228), .A(n8227), .ZN(n8235) );
  INV_X1 U9814 ( .A(n8230), .ZN(n8494) );
  NOR2_X1 U9815 ( .A1(n8250), .A2(n8267), .ZN(n8231) );
  AOI21_X1 U9816 ( .B1(n8299), .B2(n8269), .A(n8231), .ZN(n8491) );
  OAI22_X1 U9817 ( .A1(n8491), .A2(n8273), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8232), .ZN(n8233) );
  AOI21_X1 U9818 ( .B1(n8494), .B2(n8275), .A(n8233), .ZN(n8234) );
  OAI211_X1 U9819 ( .C1(n4506), .C2(n8278), .A(n8235), .B(n8234), .ZN(P2_U3231) );
  INV_X1 U9820 ( .A(n8549), .ZN(n8734) );
  AOI21_X1 U9821 ( .B1(n8237), .B2(n8236), .A(n8259), .ZN(n8239) );
  NAND2_X1 U9822 ( .A1(n8239), .A2(n8238), .ZN(n8243) );
  AOI22_X1 U9823 ( .A1(n8304), .A2(n8269), .B1(n8251), .B2(n8306), .ZN(n8546)
         );
  OAI22_X1 U9824 ( .A1(n8273), .A2(n8546), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8240), .ZN(n8241) );
  AOI21_X1 U9825 ( .B1(n4843), .B2(n8275), .A(n8241), .ZN(n8242) );
  OAI211_X1 U9826 ( .C1(n8734), .C2(n8278), .A(n8243), .B(n8242), .ZN(P2_U3235) );
  NAND2_X1 U9827 ( .A1(n8244), .A2(n8302), .ZN(n8248) );
  NAND2_X1 U9828 ( .A1(n8282), .A2(n8245), .ZN(n8247) );
  MUX2_X1 U9829 ( .A(n8248), .B(n8247), .S(n8246), .Z(n8257) );
  OR2_X1 U9830 ( .A1(n8250), .A2(n8249), .ZN(n8253) );
  NAND2_X1 U9831 ( .A1(n8304), .A2(n8251), .ZN(n8252) );
  AND2_X1 U9832 ( .A1(n8253), .A2(n8252), .ZN(n8518) );
  OAI22_X1 U9833 ( .A1(n8518), .A2(n8273), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8254), .ZN(n8255) );
  AOI21_X1 U9834 ( .B1(n8521), .B2(n8275), .A(n8255), .ZN(n8256) );
  OAI211_X1 U9835 ( .C1(n8524), .C2(n8278), .A(n8257), .B(n8256), .ZN(P2_U3237) );
  INV_X1 U9836 ( .A(n8258), .ZN(n8260) );
  AOI21_X1 U9837 ( .B1(n8261), .B2(n8260), .A(n8259), .ZN(n8266) );
  NOR3_X1 U9838 ( .A1(n8263), .A2(n8268), .A3(n8262), .ZN(n8265) );
  OAI21_X1 U9839 ( .B1(n8266), .B2(n8265), .A(n8264), .ZN(n8277) );
  OR2_X1 U9840 ( .A1(n8268), .A2(n8267), .ZN(n8271) );
  NAND2_X1 U9841 ( .A1(n8306), .A2(n8269), .ZN(n8270) );
  NAND2_X1 U9842 ( .A1(n8271), .A2(n8270), .ZN(n8578) );
  INV_X1 U9843 ( .A(n8578), .ZN(n8272) );
  NAND2_X1 U9844 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8385) );
  OAI21_X1 U9845 ( .B1(n8273), .B2(n8272), .A(n8385), .ZN(n8274) );
  AOI21_X1 U9846 ( .B1(n8585), .B2(n8275), .A(n8274), .ZN(n8276) );
  OAI211_X1 U9847 ( .C1(n8584), .C2(n8278), .A(n8277), .B(n8276), .ZN(P2_U3240) );
  AND2_X1 U9848 ( .A1(n8280), .A2(n8279), .ZN(n8295) );
  NAND3_X1 U9849 ( .A1(n8295), .A2(n8282), .A3(n8281), .ZN(n8293) );
  INV_X1 U9850 ( .A(n8283), .ZN(n8288) );
  AOI22_X1 U9851 ( .A1(n8285), .A2(n8284), .B1(P2_REG3_REG_15__SCAN_IN), .B2(
        n4262), .ZN(n8286) );
  OAI21_X1 U9852 ( .B1(n8288), .B2(n8287), .A(n8286), .ZN(n8289) );
  AOI21_X1 U9853 ( .B1(n8291), .B2(n8290), .A(n8289), .ZN(n8292) );
  OAI211_X1 U9854 ( .C1(n8295), .C2(n8294), .A(n8293), .B(n8292), .ZN(P2_U3243) );
  MUX2_X1 U9855 ( .A(n8296), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8303), .Z(
        P2_U3580) );
  MUX2_X1 U9856 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8297), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U9857 ( .A(n8298), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8303), .Z(
        P2_U3578) );
  MUX2_X1 U9858 ( .A(n8299), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8303), .Z(
        P2_U3577) );
  MUX2_X1 U9859 ( .A(n8300), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8303), .Z(
        P2_U3576) );
  MUX2_X1 U9860 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8301), .S(P2_U3966), .Z(
        P2_U3575) );
  MUX2_X1 U9861 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8302), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U9862 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8304), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U9863 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8305), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U9864 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8306), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U9865 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8307), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U9866 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8308), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9867 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8309), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9868 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8310), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9869 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8311), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9870 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8312), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9871 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8313), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U9872 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8314), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U9873 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8315), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U9874 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8316), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U9875 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8317), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U9876 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8318), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U9877 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8319), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U9878 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8320), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U9879 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8321), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U9880 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8322), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U9881 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n8323), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U9882 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n8324), .S(P2_U3966), .Z(
        P2_U3553) );
  AOI21_X1 U9883 ( .B1(n8327), .B2(n8326), .A(n8325), .ZN(n8339) );
  XNOR2_X1 U9884 ( .A(n8339), .B(n8349), .ZN(n8328) );
  NAND2_X1 U9885 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n8328), .ZN(n8341) );
  OAI211_X1 U9886 ( .C1(n8328), .C2(P2_REG1_REG_15__SCAN_IN), .A(n9936), .B(
        n8341), .ZN(n8338) );
  XNOR2_X1 U9887 ( .A(n8348), .B(n8340), .ZN(n8332) );
  INV_X1 U9888 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8331) );
  NAND2_X1 U9889 ( .A1(n8332), .A2(n8331), .ZN(n8350) );
  OAI21_X1 U9890 ( .B1(n8332), .B2(n8331), .A(n8350), .ZN(n8333) );
  NAND2_X1 U9891 ( .A1(n8333), .A2(n9937), .ZN(n8337) );
  AND2_X1 U9892 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8334) );
  AOI21_X1 U9893 ( .B1(n9943), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n8334), .ZN(
        n8336) );
  NAND2_X1 U9894 ( .A1(n9668), .A2(n8340), .ZN(n8335) );
  NAND4_X1 U9895 ( .A1(n8338), .A2(n8337), .A3(n8336), .A4(n8335), .ZN(
        P2_U3260) );
  NAND2_X1 U9896 ( .A1(n8340), .A2(n8339), .ZN(n8342) );
  NAND2_X1 U9897 ( .A1(n8342), .A2(n8341), .ZN(n8344) );
  XNOR2_X1 U9898 ( .A(n8365), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8343) );
  NOR2_X1 U9899 ( .A1(n8343), .A2(n8344), .ZN(n8366) );
  AOI21_X1 U9900 ( .B1(n8344), .B2(n8343), .A(n8366), .ZN(n8358) );
  INV_X1 U9901 ( .A(n8345), .ZN(n8346) );
  AOI21_X1 U9902 ( .B1(n9943), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8346), .ZN(
        n8347) );
  INV_X1 U9903 ( .A(n8347), .ZN(n8356) );
  NAND2_X1 U9904 ( .A1(n8349), .A2(n8348), .ZN(n8351) );
  NAND2_X1 U9905 ( .A1(n8351), .A2(n8350), .ZN(n8354) );
  NAND2_X1 U9906 ( .A1(n8365), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8352) );
  OAI21_X1 U9907 ( .B1(n8365), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8352), .ZN(
        n8353) );
  NOR2_X1 U9908 ( .A1(n8353), .A2(n8354), .ZN(n8359) );
  AOI211_X1 U9909 ( .C1(n8354), .C2(n8353), .A(n8359), .B(n9662), .ZN(n8355)
         );
  AOI211_X1 U9910 ( .C1(n9668), .C2(n8365), .A(n8356), .B(n8355), .ZN(n8357)
         );
  OAI21_X1 U9911 ( .B1(n8358), .B2(n9941), .A(n8357), .ZN(P2_U3261) );
  NAND2_X1 U9912 ( .A1(n8381), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8360) );
  OAI21_X1 U9913 ( .B1(n8381), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8360), .ZN(
        n8361) );
  AOI211_X1 U9914 ( .C1(n8362), .C2(n8361), .A(n8380), .B(n9662), .ZN(n8374)
         );
  NOR2_X1 U9915 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8363), .ZN(n8364) );
  AOI21_X1 U9916 ( .B1(n9943), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8364), .ZN(
        n8372) );
  XNOR2_X1 U9917 ( .A(n8376), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8370) );
  OR2_X1 U9918 ( .A1(n8365), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8368) );
  INV_X1 U9919 ( .A(n8366), .ZN(n8367) );
  AND2_X1 U9920 ( .A1(n8368), .A2(n8367), .ZN(n8369) );
  NAND2_X1 U9921 ( .A1(n8370), .A2(n8369), .ZN(n8375) );
  OAI211_X1 U9922 ( .C1(n8370), .C2(n8369), .A(n9936), .B(n8375), .ZN(n8371)
         );
  OAI211_X1 U9923 ( .C1(n9939), .C2(n8376), .A(n8372), .B(n8371), .ZN(n8373)
         );
  OR2_X1 U9924 ( .A1(n8374), .A2(n8373), .ZN(P2_U3262) );
  INV_X1 U9925 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8377) );
  OAI21_X1 U9926 ( .B1(n8377), .B2(n8376), .A(n8375), .ZN(n8379) );
  INV_X1 U9927 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8397) );
  AOI22_X1 U9928 ( .A1(n8387), .A2(n8397), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n8396), .ZN(n8378) );
  NOR2_X1 U9929 ( .A1(n8379), .A2(n8378), .ZN(n8395) );
  AOI21_X1 U9930 ( .B1(n8379), .B2(n8378), .A(n8395), .ZN(n8390) );
  INV_X1 U9931 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8382) );
  NAND2_X1 U9932 ( .A1(n8383), .A2(n8382), .ZN(n8393) );
  OAI21_X1 U9933 ( .B1(n8383), .B2(n8382), .A(n8393), .ZN(n8384) );
  NAND2_X1 U9934 ( .A1(n8384), .A2(n9937), .ZN(n8389) );
  OAI21_X1 U9935 ( .B1(n9650), .B2(n10158), .A(n8385), .ZN(n8386) );
  AOI21_X1 U9936 ( .B1(n9668), .B2(n8387), .A(n8386), .ZN(n8388) );
  OAI211_X1 U9937 ( .C1(n8390), .C2(n9941), .A(n8389), .B(n8388), .ZN(P2_U3263) );
  INV_X1 U9938 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8410) );
  NAND2_X1 U9939 ( .A1(n8391), .A2(n8396), .ZN(n8392) );
  NAND2_X1 U9940 ( .A1(n8393), .A2(n8392), .ZN(n8394) );
  XNOR2_X1 U9941 ( .A(n8394), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8404) );
  AOI21_X1 U9942 ( .B1(n8397), .B2(n8396), .A(n8395), .ZN(n8399) );
  INV_X1 U9943 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8398) );
  XOR2_X1 U9944 ( .A(n8399), .B(n8398), .Z(n8402) );
  AOI21_X1 U9945 ( .B1(n8402), .B2(n9936), .A(n9668), .ZN(n8400) );
  OAI21_X1 U9946 ( .B1(n8404), .B2(n9662), .A(n8400), .ZN(n8401) );
  INV_X1 U9947 ( .A(n8401), .ZN(n8407) );
  INV_X1 U9948 ( .A(n8402), .ZN(n8403) );
  AOI22_X1 U9949 ( .A1(n8404), .A2(n9937), .B1(n9936), .B2(n8403), .ZN(n8406)
         );
  OAI211_X1 U9950 ( .C1(n8410), .C2(n9650), .A(n8409), .B(n8408), .ZN(P2_U3264) );
  XNOR2_X1 U9951 ( .A(n8418), .B(n8689), .ZN(n8411) );
  NAND2_X1 U9952 ( .A1(n8607), .A2(n9993), .ZN(n8417) );
  INV_X1 U9953 ( .A(n8412), .ZN(n8413) );
  AND2_X1 U9954 ( .A1(n8414), .A2(n8413), .ZN(n8610) );
  INV_X1 U9955 ( .A(n8610), .ZN(n8415) );
  NOR2_X1 U9956 ( .A1(n10011), .A2(n8415), .ZN(n8421) );
  AOI21_X1 U9957 ( .B1(n10011), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8421), .ZN(
        n8416) );
  OAI211_X1 U9958 ( .C1(n8689), .C2(n10004), .A(n8417), .B(n8416), .ZN(
        P2_U3265) );
  AOI211_X1 U9959 ( .C1(n8420), .C2(n8419), .A(n10086), .B(n8418), .ZN(n8611)
         );
  NAND2_X1 U9960 ( .A1(n8611), .A2(n9993), .ZN(n8423) );
  AOI21_X1 U9961 ( .B1(n10011), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8421), .ZN(
        n8422) );
  OAI211_X1 U9962 ( .C1(n4579), .C2(n10004), .A(n8423), .B(n8422), .ZN(
        P2_U3266) );
  OAI211_X1 U9963 ( .C1(n8428), .C2(n8427), .A(n8426), .B(n9968), .ZN(n8430)
         );
  NAND2_X1 U9964 ( .A1(n8430), .A2(n8429), .ZN(n8614) );
  AOI211_X1 U9965 ( .C1(n8616), .C2(n8445), .A(n10086), .B(n8431), .ZN(n8615)
         );
  NAND2_X1 U9966 ( .A1(n8615), .A2(n9993), .ZN(n8434) );
  AOI22_X1 U9967 ( .A1(n8432), .A2(n10001), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n10011), .ZN(n8433) );
  OAI211_X1 U9968 ( .C1(n4481), .C2(n10004), .A(n8434), .B(n8433), .ZN(n8435)
         );
  AOI21_X1 U9969 ( .B1(n8614), .B2(n10009), .A(n8435), .ZN(n8436) );
  OAI21_X1 U9970 ( .B1(n8696), .B2(n8592), .A(n8436), .ZN(P2_U3268) );
  NAND2_X1 U9971 ( .A1(n8440), .A2(n8439), .ZN(n8441) );
  NAND3_X1 U9972 ( .A1(n8442), .A2(n9968), .A3(n8441), .ZN(n8444) );
  AND2_X1 U9973 ( .A1(n8444), .A2(n8443), .ZN(n8620) );
  INV_X1 U9974 ( .A(n8620), .ZN(n8451) );
  OAI211_X1 U9975 ( .C1(n8446), .C2(n8463), .A(n10049), .B(n8445), .ZN(n8619)
         );
  AOI22_X1 U9976 ( .A1(n8447), .A2(n10001), .B1(n10011), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n8449) );
  NAND2_X1 U9977 ( .A1(n8699), .A2(n9990), .ZN(n8448) );
  OAI211_X1 U9978 ( .C1(n8619), .C2(n8588), .A(n8449), .B(n8448), .ZN(n8450)
         );
  AOI21_X1 U9979 ( .B1(n8451), .B2(n10009), .A(n8450), .ZN(n8452) );
  OAI21_X1 U9980 ( .B1(n8701), .B2(n8592), .A(n8452), .ZN(P2_U3269) );
  XNOR2_X1 U9981 ( .A(n8454), .B(n8453), .ZN(n8705) );
  AOI22_X1 U9982 ( .A1(n8626), .A2(n9990), .B1(n10011), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8467) );
  INV_X1 U9983 ( .A(n8455), .ZN(n8459) );
  AOI21_X1 U9984 ( .B1(n8469), .B2(n8457), .A(n8456), .ZN(n8458) );
  OAI21_X1 U9985 ( .B1(n8459), .B2(n8458), .A(n9968), .ZN(n8461) );
  NAND2_X1 U9986 ( .A1(n8461), .A2(n8460), .ZN(n8624) );
  OAI21_X1 U9987 ( .B1(n4504), .B2(n8475), .A(n10049), .ZN(n8462) );
  OR2_X1 U9988 ( .A1(n8463), .A2(n8462), .ZN(n8623) );
  OAI22_X1 U9989 ( .A1(n8623), .A2(n8480), .B1(n8479), .B2(n8464), .ZN(n8465)
         );
  OAI21_X1 U9990 ( .B1(n8624), .B2(n8465), .A(n10009), .ZN(n8466) );
  OAI211_X1 U9991 ( .C1(n8705), .C2(n8592), .A(n8467), .B(n8466), .ZN(P2_U3270) );
  XNOR2_X1 U9992 ( .A(n8468), .B(n8471), .ZN(n8710) );
  AOI22_X1 U9993 ( .A1(n8708), .A2(n9990), .B1(n10011), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n8483) );
  OAI211_X1 U9994 ( .C1(n8471), .C2(n8470), .A(n8469), .B(n9968), .ZN(n8473)
         );
  NAND2_X1 U9995 ( .A1(n8473), .A2(n8472), .ZN(n8629) );
  NAND2_X1 U9996 ( .A1(n8493), .A2(n8708), .ZN(n8474) );
  NAND2_X1 U9997 ( .A1(n8474), .A2(n10049), .ZN(n8476) );
  OR2_X1 U9998 ( .A1(n8476), .A2(n8475), .ZN(n8630) );
  INV_X1 U9999 ( .A(n8477), .ZN(n8478) );
  OAI22_X1 U10000 ( .A1(n8630), .A2(n8480), .B1(n8479), .B2(n8478), .ZN(n8481)
         );
  OAI21_X1 U10001 ( .B1(n8629), .B2(n8481), .A(n10009), .ZN(n8482) );
  OAI211_X1 U10002 ( .C1(n8710), .C2(n8592), .A(n8483), .B(n8482), .ZN(
        P2_U3271) );
  OAI21_X1 U10003 ( .B1(n8486), .B2(n8485), .A(n8484), .ZN(n8487) );
  INV_X1 U10004 ( .A(n8487), .ZN(n8714) );
  OAI211_X1 U10005 ( .C1(n8490), .C2(n8489), .A(n8488), .B(n9968), .ZN(n8492)
         );
  NAND2_X1 U10006 ( .A1(n8492), .A2(n8491), .ZN(n8634) );
  AOI211_X1 U10007 ( .C1(n8636), .C2(n4276), .A(n10086), .B(n4470), .ZN(n8635)
         );
  NAND2_X1 U10008 ( .A1(n8635), .A2(n9993), .ZN(n8496) );
  AOI22_X1 U10009 ( .A1(n10011), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8494), 
        .B2(n10001), .ZN(n8495) );
  OAI211_X1 U10010 ( .C1(n4506), .C2(n10004), .A(n8496), .B(n8495), .ZN(n8497)
         );
  AOI21_X1 U10011 ( .B1(n8634), .B2(n10009), .A(n8497), .ZN(n8498) );
  OAI21_X1 U10012 ( .B1(n8714), .B2(n8592), .A(n8498), .ZN(P2_U3272) );
  NAND2_X1 U10013 ( .A1(n8516), .A2(n8499), .ZN(n8501) );
  XNOR2_X1 U10014 ( .A(n8501), .B(n8500), .ZN(n8503) );
  AOI21_X1 U10015 ( .B1(n8503), .B2(n9968), .A(n8502), .ZN(n8641) );
  AOI21_X1 U10016 ( .B1(n8506), .B2(n8505), .A(n8504), .ZN(n8717) );
  NAND2_X1 U10017 ( .A1(n8717), .A2(n10006), .ZN(n8513) );
  OAI211_X1 U10018 ( .C1(n8509), .C2(n8520), .A(n4276), .B(n10049), .ZN(n8640)
         );
  INV_X1 U10019 ( .A(n8640), .ZN(n8511) );
  AOI22_X1 U10020 ( .A1(n10011), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8507), 
        .B2(n10001), .ZN(n8508) );
  OAI21_X1 U10021 ( .B1(n8509), .B2(n10004), .A(n8508), .ZN(n8510) );
  AOI21_X1 U10022 ( .B1(n8511), .B2(n9993), .A(n8510), .ZN(n8512) );
  OAI211_X1 U10023 ( .C1(n10011), .C2(n8641), .A(n8513), .B(n8512), .ZN(
        P2_U3273) );
  XNOR2_X1 U10024 ( .A(n8515), .B(n8514), .ZN(n8725) );
  OAI211_X1 U10025 ( .C1(n4308), .C2(n8517), .A(n9968), .B(n8516), .ZN(n8519)
         );
  NAND2_X1 U10026 ( .A1(n8519), .A2(n8518), .ZN(n8645) );
  AOI211_X1 U10027 ( .C1(n8647), .C2(n4340), .A(n10086), .B(n8520), .ZN(n8646)
         );
  NAND2_X1 U10028 ( .A1(n8646), .A2(n9993), .ZN(n8523) );
  AOI22_X1 U10029 ( .A1(n10011), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8521), 
        .B2(n10001), .ZN(n8522) );
  OAI211_X1 U10030 ( .C1(n8524), .C2(n10004), .A(n8523), .B(n8522), .ZN(n8525)
         );
  AOI21_X1 U10031 ( .B1(n8645), .B2(n10009), .A(n8525), .ZN(n8526) );
  OAI21_X1 U10032 ( .B1(n8725), .B2(n8592), .A(n8526), .ZN(P2_U3274) );
  XOR2_X1 U10033 ( .A(n8528), .B(n8527), .Z(n8730) );
  XNOR2_X1 U10034 ( .A(n8529), .B(n8528), .ZN(n8531) );
  AOI21_X1 U10035 ( .B1(n8531), .B2(n9968), .A(n8530), .ZN(n8651) );
  INV_X1 U10036 ( .A(n8651), .ZN(n8539) );
  INV_X1 U10037 ( .A(n8550), .ZN(n8532) );
  OAI211_X1 U10038 ( .C1(n8533), .C2(n8532), .A(n4340), .B(n10049), .ZN(n8650)
         );
  INV_X1 U10039 ( .A(n8534), .ZN(n8535) );
  AOI22_X1 U10040 ( .A1(n10011), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8535), 
        .B2(n10001), .ZN(n8537) );
  NAND2_X1 U10041 ( .A1(n8728), .A2(n9990), .ZN(n8536) );
  OAI211_X1 U10042 ( .C1(n8650), .C2(n8588), .A(n8537), .B(n8536), .ZN(n8538)
         );
  AOI21_X1 U10043 ( .B1(n8539), .B2(n10009), .A(n8538), .ZN(n8540) );
  OAI21_X1 U10044 ( .B1(n8730), .B2(n8592), .A(n8540), .ZN(P2_U3275) );
  XNOR2_X1 U10045 ( .A(n8541), .B(n8544), .ZN(n8656) );
  INV_X1 U10046 ( .A(n8656), .ZN(n8556) );
  NAND2_X1 U10047 ( .A1(n8542), .A2(n9968), .ZN(n8548) );
  AOI21_X1 U10048 ( .B1(n8543), .B2(n8545), .A(n8544), .ZN(n8547) );
  OAI21_X1 U10049 ( .B1(n8548), .B2(n8547), .A(n8546), .ZN(n8654) );
  AOI21_X1 U10050 ( .B1(n8566), .B2(n8549), .A(n10086), .ZN(n8551) );
  AND2_X1 U10051 ( .A1(n8551), .A2(n8550), .ZN(n8655) );
  NAND2_X1 U10052 ( .A1(n8655), .A2(n9993), .ZN(n8553) );
  AOI22_X1 U10053 ( .A1(n10011), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n4843), 
        .B2(n10001), .ZN(n8552) );
  OAI211_X1 U10054 ( .C1(n8734), .C2(n10004), .A(n8553), .B(n8552), .ZN(n8554)
         );
  AOI21_X1 U10055 ( .B1(n8654), .B2(n10009), .A(n8554), .ZN(n8555) );
  OAI21_X1 U10056 ( .B1(n8556), .B2(n8592), .A(n8555), .ZN(P2_U3276) );
  XNOR2_X1 U10057 ( .A(n8557), .B(n8561), .ZN(n8739) );
  INV_X1 U10058 ( .A(n8558), .ZN(n8559) );
  NAND2_X1 U10059 ( .A1(n8560), .A2(n8559), .ZN(n8562) );
  NAND2_X1 U10060 ( .A1(n8562), .A2(n8561), .ZN(n8563) );
  NAND2_X1 U10061 ( .A1(n8563), .A2(n8543), .ZN(n8565) );
  AOI21_X1 U10062 ( .B1(n8565), .B2(n9968), .A(n8564), .ZN(n8660) );
  INV_X1 U10063 ( .A(n8660), .ZN(n8572) );
  OAI211_X1 U10064 ( .C1(n8567), .C2(n8581), .A(n8566), .B(n10049), .ZN(n8659)
         );
  AOI22_X1 U10065 ( .A1(n10011), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8568), 
        .B2(n10001), .ZN(n8570) );
  NAND2_X1 U10066 ( .A1(n8737), .A2(n9990), .ZN(n8569) );
  OAI211_X1 U10067 ( .C1(n8659), .C2(n8588), .A(n8570), .B(n8569), .ZN(n8571)
         );
  AOI21_X1 U10068 ( .B1(n8572), .B2(n10009), .A(n8571), .ZN(n8573) );
  OAI21_X1 U10069 ( .B1(n8739), .B2(n8592), .A(n8573), .ZN(P2_U3277) );
  XNOR2_X1 U10070 ( .A(n8574), .B(n8575), .ZN(n8744) );
  INV_X1 U10071 ( .A(n8575), .ZN(n8576) );
  XNOR2_X1 U10072 ( .A(n8577), .B(n8576), .ZN(n8579) );
  AOI21_X1 U10073 ( .B1(n8579), .B2(n9968), .A(n8578), .ZN(n8664) );
  INV_X1 U10074 ( .A(n8664), .ZN(n8590) );
  INV_X1 U10075 ( .A(n8580), .ZN(n8583) );
  INV_X1 U10076 ( .A(n8581), .ZN(n8582) );
  OAI211_X1 U10077 ( .C1(n8584), .C2(n8583), .A(n8582), .B(n10049), .ZN(n8663)
         );
  AOI22_X1 U10078 ( .A1(n10011), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8585), 
        .B2(n10001), .ZN(n8587) );
  NAND2_X1 U10079 ( .A1(n8742), .A2(n9990), .ZN(n8586) );
  OAI211_X1 U10080 ( .C1(n8663), .C2(n8588), .A(n8587), .B(n8586), .ZN(n8589)
         );
  AOI21_X1 U10081 ( .B1(n8590), .B2(n10009), .A(n8589), .ZN(n8591) );
  OAI21_X1 U10082 ( .B1(n8744), .B2(n8592), .A(n8591), .ZN(P2_U3278) );
  XNOR2_X1 U10083 ( .A(n8593), .B(n8600), .ZN(n8596) );
  INV_X1 U10084 ( .A(n8594), .ZN(n8595) );
  AOI21_X1 U10085 ( .B1(n8596), .B2(n9968), .A(n8595), .ZN(n10052) );
  MUX2_X1 U10086 ( .A(n10052), .B(n6474), .S(n10011), .Z(n8606) );
  AOI22_X1 U10087 ( .A1(n9990), .A2(n10048), .B1(n10001), .B2(n8597), .ZN(
        n8605) );
  NAND2_X1 U10088 ( .A1(n8599), .A2(n8600), .ZN(n10047) );
  NAND3_X1 U10089 ( .A1(n8598), .A2(n10047), .A3(n10006), .ZN(n8604) );
  AOI21_X1 U10090 ( .B1(n10048), .B2(n8601), .A(n9979), .ZN(n10050) );
  NAND2_X1 U10091 ( .A1(n10050), .A2(n8602), .ZN(n8603) );
  NAND4_X1 U10092 ( .A1(n8606), .A2(n8605), .A3(n8604), .A4(n8603), .ZN(
        P2_U3290) );
  INV_X1 U10093 ( .A(n8670), .ZN(n8679) );
  NOR2_X1 U10094 ( .A1(n8607), .A2(n8610), .ZN(n8686) );
  MUX2_X1 U10095 ( .A(n8608), .B(n8686), .S(n10120), .Z(n8609) );
  OAI21_X1 U10096 ( .B1(n8689), .B2(n8679), .A(n8609), .ZN(P2_U3551) );
  INV_X1 U10097 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8612) );
  NOR2_X1 U10098 ( .A1(n8611), .A2(n8610), .ZN(n8690) );
  MUX2_X1 U10099 ( .A(n8612), .B(n8690), .S(n10120), .Z(n8613) );
  OAI21_X1 U10100 ( .B1(n4579), .B2(n8679), .A(n8613), .ZN(P2_U3550) );
  AOI211_X1 U10101 ( .C1(n8616), .C2(n10069), .A(n8615), .B(n8614), .ZN(n8693)
         );
  MUX2_X1 U10102 ( .A(n8617), .B(n8693), .S(n10120), .Z(n8618) );
  OAI21_X1 U10103 ( .B1(n8696), .B2(n8672), .A(n8618), .ZN(P2_U3548) );
  NAND2_X1 U10104 ( .A1(n8620), .A2(n8619), .ZN(n8697) );
  MUX2_X1 U10105 ( .A(n8697), .B(P2_REG1_REG_27__SCAN_IN), .S(n10117), .Z(
        n8621) );
  AOI21_X1 U10106 ( .B1(n8670), .B2(n8699), .A(n8621), .ZN(n8622) );
  OAI21_X1 U10107 ( .B1(n8701), .B2(n8672), .A(n8622), .ZN(P2_U3547) );
  INV_X1 U10108 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8627) );
  INV_X1 U10109 ( .A(n8623), .ZN(n8625) );
  AOI211_X1 U10110 ( .C1(n8626), .C2(n10069), .A(n8625), .B(n8624), .ZN(n8702)
         );
  MUX2_X1 U10111 ( .A(n8627), .B(n8702), .S(n10120), .Z(n8628) );
  OAI21_X1 U10112 ( .B1(n8705), .B2(n8672), .A(n8628), .ZN(P2_U3546) );
  INV_X1 U10113 ( .A(n8629), .ZN(n8631) );
  NAND2_X1 U10114 ( .A1(n8631), .A2(n8630), .ZN(n8706) );
  MUX2_X1 U10115 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8706), .S(n10120), .Z(
        n8632) );
  AOI21_X1 U10116 ( .B1(n8670), .B2(n8708), .A(n8632), .ZN(n8633) );
  OAI21_X1 U10117 ( .B1(n8710), .B2(n8672), .A(n8633), .ZN(P2_U3545) );
  INV_X1 U10118 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8637) );
  AOI211_X1 U10119 ( .C1(n8636), .C2(n10069), .A(n8635), .B(n8634), .ZN(n8711)
         );
  MUX2_X1 U10120 ( .A(n8637), .B(n8711), .S(n10120), .Z(n8638) );
  OAI21_X1 U10121 ( .B1(n8714), .B2(n8672), .A(n8638), .ZN(P2_U3544) );
  AOI22_X1 U10122 ( .A1(n8717), .A2(n8639), .B1(n8670), .B2(n8715), .ZN(n8644)
         );
  AND2_X1 U10123 ( .A1(n8641), .A2(n8640), .ZN(n8719) );
  INV_X1 U10124 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8642) );
  MUX2_X1 U10125 ( .A(n8719), .B(n8642), .S(n10117), .Z(n8643) );
  NAND2_X1 U10126 ( .A1(n8644), .A2(n8643), .ZN(P2_U3543) );
  AOI211_X1 U10127 ( .C1(n8647), .C2(n10069), .A(n8646), .B(n8645), .ZN(n8722)
         );
  MUX2_X1 U10128 ( .A(n8648), .B(n8722), .S(n10120), .Z(n8649) );
  OAI21_X1 U10129 ( .B1(n8725), .B2(n8672), .A(n8649), .ZN(P2_U3542) );
  NAND2_X1 U10130 ( .A1(n8651), .A2(n8650), .ZN(n8726) );
  MUX2_X1 U10131 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8726), .S(n10120), .Z(
        n8652) );
  AOI21_X1 U10132 ( .B1(n8670), .B2(n8728), .A(n8652), .ZN(n8653) );
  OAI21_X1 U10133 ( .B1(n8730), .B2(n8672), .A(n8653), .ZN(P2_U3541) );
  INV_X1 U10134 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8657) );
  AOI211_X1 U10135 ( .C1(n8656), .C2(n10097), .A(n8655), .B(n8654), .ZN(n8731)
         );
  MUX2_X1 U10136 ( .A(n8657), .B(n8731), .S(n10120), .Z(n8658) );
  OAI21_X1 U10137 ( .B1(n8734), .B2(n8679), .A(n8658), .ZN(P2_U3540) );
  NAND2_X1 U10138 ( .A1(n8660), .A2(n8659), .ZN(n8735) );
  MUX2_X1 U10139 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8735), .S(n10120), .Z(
        n8661) );
  AOI21_X1 U10140 ( .B1(n8670), .B2(n8737), .A(n8661), .ZN(n8662) );
  OAI21_X1 U10141 ( .B1(n8739), .B2(n8672), .A(n8662), .ZN(P2_U3539) );
  NAND2_X1 U10142 ( .A1(n8664), .A2(n8663), .ZN(n8740) );
  MUX2_X1 U10143 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8740), .S(n10120), .Z(
        n8665) );
  AOI21_X1 U10144 ( .B1(n8670), .B2(n8742), .A(n8665), .ZN(n8666) );
  OAI21_X1 U10145 ( .B1(n8744), .B2(n8672), .A(n8666), .ZN(P2_U3538) );
  NAND2_X1 U10146 ( .A1(n8668), .A2(n8667), .ZN(n8745) );
  MUX2_X1 U10147 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8745), .S(n10120), .Z(
        n8669) );
  AOI21_X1 U10148 ( .B1(n8670), .B2(n8747), .A(n8669), .ZN(n8671) );
  OAI21_X1 U10149 ( .B1(n8751), .B2(n8672), .A(n8671), .ZN(P2_U3537) );
  INV_X1 U10150 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8677) );
  INV_X1 U10151 ( .A(n8673), .ZN(n8676) );
  INV_X1 U10152 ( .A(n10073), .ZN(n10082) );
  AOI211_X1 U10153 ( .C1(n8676), .C2(n10082), .A(n8675), .B(n8674), .ZN(n8752)
         );
  MUX2_X1 U10154 ( .A(n8677), .B(n8752), .S(n10120), .Z(n8678) );
  OAI21_X1 U10155 ( .B1(n8756), .B2(n8679), .A(n8678), .ZN(P2_U3536) );
  NAND2_X1 U10156 ( .A1(n8680), .A2(n10069), .ZN(n8682) );
  OAI211_X1 U10157 ( .C1(n8683), .C2(n10073), .A(n8682), .B(n8681), .ZN(n8684)
         );
  OR2_X1 U10158 ( .A1(n8685), .A2(n8684), .ZN(n8757) );
  MUX2_X1 U10159 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n8757), .S(n10120), .Z(
        P2_U3533) );
  INV_X1 U10160 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8687) );
  MUX2_X1 U10161 ( .A(n8687), .B(n8686), .S(n10101), .Z(n8688) );
  OAI21_X1 U10162 ( .B1(n8689), .B2(n8755), .A(n8688), .ZN(P2_U3519) );
  MUX2_X1 U10163 ( .A(n8691), .B(n8690), .S(n10101), .Z(n8692) );
  OAI21_X1 U10164 ( .B1(n4579), .B2(n8755), .A(n8692), .ZN(P2_U3518) );
  INV_X1 U10165 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8694) );
  MUX2_X1 U10166 ( .A(n8694), .B(n8693), .S(n10101), .Z(n8695) );
  OAI21_X1 U10167 ( .B1(n8696), .B2(n8750), .A(n8695), .ZN(P2_U3516) );
  MUX2_X1 U10168 ( .A(n8697), .B(P2_REG0_REG_27__SCAN_IN), .S(n10099), .Z(
        n8698) );
  AOI21_X1 U10169 ( .B1(n8748), .B2(n8699), .A(n8698), .ZN(n8700) );
  OAI21_X1 U10170 ( .B1(n8701), .B2(n8750), .A(n8700), .ZN(P2_U3515) );
  MUX2_X1 U10171 ( .A(n8703), .B(n8702), .S(n10101), .Z(n8704) );
  OAI21_X1 U10172 ( .B1(n8705), .B2(n8750), .A(n8704), .ZN(P2_U3514) );
  MUX2_X1 U10173 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8706), .S(n10101), .Z(
        n8707) );
  AOI21_X1 U10174 ( .B1(n8748), .B2(n8708), .A(n8707), .ZN(n8709) );
  OAI21_X1 U10175 ( .B1(n8710), .B2(n8750), .A(n8709), .ZN(P2_U3513) );
  MUX2_X1 U10176 ( .A(n8712), .B(n8711), .S(n10101), .Z(n8713) );
  OAI21_X1 U10177 ( .B1(n8714), .B2(n8750), .A(n8713), .ZN(P2_U3512) );
  AOI22_X1 U10178 ( .A1(n8717), .A2(n8716), .B1(n8748), .B2(n8715), .ZN(n8721)
         );
  INV_X1 U10179 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8718) );
  MUX2_X1 U10180 ( .A(n8719), .B(n8718), .S(n10099), .Z(n8720) );
  NAND2_X1 U10181 ( .A1(n8721), .A2(n8720), .ZN(P2_U3511) );
  INV_X1 U10182 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8723) );
  MUX2_X1 U10183 ( .A(n8723), .B(n8722), .S(n10101), .Z(n8724) );
  OAI21_X1 U10184 ( .B1(n8725), .B2(n8750), .A(n8724), .ZN(P2_U3510) );
  MUX2_X1 U10185 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8726), .S(n10101), .Z(
        n8727) );
  AOI21_X1 U10186 ( .B1(n8748), .B2(n8728), .A(n8727), .ZN(n8729) );
  OAI21_X1 U10187 ( .B1(n8730), .B2(n8750), .A(n8729), .ZN(P2_U3509) );
  INV_X1 U10188 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8732) );
  MUX2_X1 U10189 ( .A(n8732), .B(n8731), .S(n10101), .Z(n8733) );
  OAI21_X1 U10190 ( .B1(n8734), .B2(n8755), .A(n8733), .ZN(P2_U3508) );
  MUX2_X1 U10191 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8735), .S(n10101), .Z(
        n8736) );
  AOI21_X1 U10192 ( .B1(n8748), .B2(n8737), .A(n8736), .ZN(n8738) );
  OAI21_X1 U10193 ( .B1(n8739), .B2(n8750), .A(n8738), .ZN(P2_U3507) );
  MUX2_X1 U10194 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8740), .S(n10101), .Z(
        n8741) );
  AOI21_X1 U10195 ( .B1(n8748), .B2(n8742), .A(n8741), .ZN(n8743) );
  OAI21_X1 U10196 ( .B1(n8744), .B2(n8750), .A(n8743), .ZN(P2_U3505) );
  MUX2_X1 U10197 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8745), .S(n10101), .Z(
        n8746) );
  AOI21_X1 U10198 ( .B1(n8748), .B2(n8747), .A(n8746), .ZN(n8749) );
  OAI21_X1 U10199 ( .B1(n8751), .B2(n8750), .A(n8749), .ZN(P2_U3502) );
  INV_X1 U10200 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8753) );
  MUX2_X1 U10201 ( .A(n8753), .B(n8752), .S(n10101), .Z(n8754) );
  OAI21_X1 U10202 ( .B1(n8756), .B2(n8755), .A(n8754), .ZN(P2_U3499) );
  MUX2_X1 U10203 ( .A(n8757), .B(P2_REG0_REG_13__SCAN_IN), .S(n10099), .Z(
        P2_U3490) );
  INV_X1 U10204 ( .A(n8758), .ZN(n9636) );
  INV_X1 U10205 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8759) );
  NAND3_X1 U10206 ( .A1(n8759), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n8760) );
  OAI22_X1 U10207 ( .A1(n5555), .A2(n8760), .B1(n6250), .B2(n4268), .ZN(n8761)
         );
  INV_X1 U10208 ( .A(n8761), .ZN(n8762) );
  OAI21_X1 U10209 ( .B1(n9636), .B2(n8768), .A(n8762), .ZN(P2_U3327) );
  INV_X1 U10210 ( .A(n8763), .ZN(n9638) );
  OAI222_X1 U10211 ( .A1(n4268), .A2(n8765), .B1(n8768), .B2(n9638), .C1(n4262), .C2(n8764), .ZN(P2_U3328) );
  INV_X1 U10212 ( .A(n8766), .ZN(n9644) );
  OAI222_X1 U10213 ( .A1(n4268), .A2(n8769), .B1(n8768), .B2(n9644), .C1(n8767), .C2(n4262), .ZN(P2_U3329) );
  MUX2_X1 U10214 ( .A(n8770), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  NAND2_X1 U10215 ( .A1(n8818), .A2(n8771), .ZN(n8773) );
  NAND2_X1 U10216 ( .A1(n8773), .A2(n8772), .ZN(n8775) );
  AND2_X1 U10217 ( .A1(n8775), .A2(n8774), .ZN(n8781) );
  AOI21_X1 U10218 ( .B1(n8777), .B2(n4352), .A(n8776), .ZN(n8778) );
  NOR2_X1 U10219 ( .A1(n8778), .A2(n4653), .ZN(n8779) );
  OAI21_X1 U10220 ( .B1(n8781), .B2(n8780), .A(n8779), .ZN(n8787) );
  NOR2_X1 U10221 ( .A1(n8926), .A2(n8782), .ZN(n8785) );
  OAI21_X1 U10222 ( .B1(n8897), .B2(n8825), .A(n8783), .ZN(n8784) );
  AOI211_X1 U10223 ( .C1(n8942), .C2(n9247), .A(n8785), .B(n8784), .ZN(n8786)
         );
  OAI211_X1 U10224 ( .C1(n9718), .C2(n8945), .A(n8787), .B(n8786), .ZN(
        P1_U3213) );
  NAND2_X1 U10225 ( .A1(n4318), .A2(n8788), .ZN(n8790) );
  XNOR2_X1 U10226 ( .A(n8790), .B(n8789), .ZN(n8795) );
  NAND2_X1 U10227 ( .A1(n9394), .A2(n8942), .ZN(n8792) );
  AOI22_X1 U10228 ( .A1(n9426), .A2(n8936), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8791) );
  OAI211_X1 U10229 ( .C1(n8926), .C2(n9400), .A(n8792), .B(n8791), .ZN(n8793)
         );
  AOI21_X1 U10230 ( .B1(n9555), .B2(n8928), .A(n8793), .ZN(n8794) );
  OAI21_X1 U10231 ( .B1(n8795), .B2(n4653), .A(n8794), .ZN(P1_U3214) );
  INV_X1 U10232 ( .A(n8799), .ZN(n8797) );
  NAND2_X1 U10233 ( .A1(n8797), .A2(n8796), .ZN(n8918) );
  NAND2_X1 U10234 ( .A1(n8918), .A2(n8917), .ZN(n8916) );
  NAND2_X1 U10235 ( .A1(n8799), .A2(n8798), .ZN(n8920) );
  NAND2_X1 U10236 ( .A1(n8800), .A2(n8866), .ZN(n8801) );
  AOI21_X1 U10237 ( .B1(n8916), .B2(n8920), .A(n8801), .ZN(n8870) );
  AND3_X1 U10238 ( .A1(n8916), .A2(n8920), .A3(n8801), .ZN(n8802) );
  OAI21_X1 U10239 ( .B1(n8870), .B2(n8802), .A(n8935), .ZN(n8807) );
  NAND2_X1 U10240 ( .A1(n8942), .A2(n9463), .ZN(n8803) );
  NAND2_X1 U10241 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9293) );
  NAND2_X1 U10242 ( .A1(n8803), .A2(n9293), .ZN(n8805) );
  NOR2_X1 U10243 ( .A1(n8926), .A2(n9454), .ZN(n8804) );
  AOI211_X1 U10244 ( .C1(n8936), .C2(n9500), .A(n8805), .B(n8804), .ZN(n8806)
         );
  OAI211_X1 U10245 ( .C1(n4546), .C2(n8945), .A(n8807), .B(n8806), .ZN(
        P1_U3217) );
  OAI21_X1 U10246 ( .B1(n8810), .B2(n8809), .A(n8808), .ZN(n8811) );
  NAND2_X1 U10247 ( .A1(n8811), .A2(n8935), .ZN(n8816) );
  AOI22_X1 U10248 ( .A1(n8936), .A2(n9463), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8812) );
  OAI21_X1 U10249 ( .B1(n8813), .B2(n8923), .A(n8812), .ZN(n8814) );
  AOI21_X1 U10250 ( .B1(n9432), .B2(n8937), .A(n8814), .ZN(n8815) );
  OAI211_X1 U10251 ( .C1(n9565), .C2(n8945), .A(n8816), .B(n8815), .ZN(
        P1_U3221) );
  NAND2_X1 U10252 ( .A1(n8818), .A2(n8817), .ZN(n8910) );
  OR2_X1 U10253 ( .A1(n8910), .A2(n8911), .ZN(n8908) );
  NAND2_X1 U10254 ( .A1(n8908), .A2(n8819), .ZN(n8823) );
  XNOR2_X1 U10255 ( .A(n8821), .B(n8820), .ZN(n8822) );
  XNOR2_X1 U10256 ( .A(n8823), .B(n8822), .ZN(n8832) );
  NOR2_X1 U10257 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8824), .ZN(n9785) );
  NOR2_X1 U10258 ( .A1(n8923), .A2(n8825), .ZN(n8826) );
  AOI211_X1 U10259 ( .C1(n8936), .C2(n9251), .A(n9785), .B(n8826), .ZN(n8827)
         );
  OAI21_X1 U10260 ( .B1(n8926), .B2(n8828), .A(n8827), .ZN(n8829) );
  AOI21_X1 U10261 ( .B1(n8928), .B2(n8830), .A(n8829), .ZN(n8831) );
  OAI21_X1 U10262 ( .B1(n8832), .B2(n4653), .A(n8831), .ZN(P1_U3222) );
  AOI21_X1 U10263 ( .B1(n8834), .B2(n8833), .A(n8933), .ZN(n8839) );
  NAND2_X1 U10264 ( .A1(n9372), .A2(n8942), .ZN(n8836) );
  AOI22_X1 U10265 ( .A1(n9394), .A2(n8936), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8835) );
  OAI211_X1 U10266 ( .C1(n8926), .C2(n9364), .A(n8836), .B(n8835), .ZN(n8837)
         );
  AOI21_X1 U10267 ( .B1(n9543), .B2(n8928), .A(n8837), .ZN(n8838) );
  OAI21_X1 U10268 ( .B1(n8839), .B2(n4653), .A(n8838), .ZN(P1_U3223) );
  INV_X1 U10269 ( .A(n8841), .ZN(n8842) );
  AOI21_X1 U10270 ( .B1(n8840), .B2(n8843), .A(n8842), .ZN(n8848) );
  NAND2_X1 U10271 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9825) );
  OAI21_X1 U10272 ( .B1(n8897), .B2(n9511), .A(n9825), .ZN(n8844) );
  AOI21_X1 U10273 ( .B1(n8942), .B2(n9471), .A(n8844), .ZN(n8845) );
  OAI21_X1 U10274 ( .B1(n8926), .B2(n9513), .A(n8845), .ZN(n8846) );
  AOI21_X1 U10275 ( .B1(n9594), .B2(n8928), .A(n8846), .ZN(n8847) );
  OAI21_X1 U10276 ( .B1(n8848), .B2(n4653), .A(n8847), .ZN(P1_U3224) );
  OAI21_X1 U10277 ( .B1(n8851), .B2(n8850), .A(n8849), .ZN(n8852) );
  NAND2_X1 U10278 ( .A1(n8852), .A2(n8935), .ZN(n8857) );
  NOR2_X1 U10279 ( .A1(n8926), .A2(n9491), .ZN(n8855) );
  NAND2_X1 U10280 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9843) );
  OAI21_X1 U10281 ( .B1(n8923), .B2(n8853), .A(n9843), .ZN(n8854) );
  AOI211_X1 U10282 ( .C1(n8936), .C2(n9498), .A(n8855), .B(n8854), .ZN(n8856)
         );
  OAI211_X1 U10283 ( .C1(n9494), .C2(n8945), .A(n8857), .B(n8856), .ZN(
        P1_U3226) );
  AOI21_X1 U10284 ( .B1(n8860), .B2(n8859), .A(n8858), .ZN(n8865) );
  AOI22_X1 U10285 ( .A1(n9246), .A2(n8936), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8862) );
  NAND2_X1 U10286 ( .A1(n8937), .A2(n9384), .ZN(n8861) );
  OAI211_X1 U10287 ( .C1(n9382), .C2(n8923), .A(n8862), .B(n8861), .ZN(n8863)
         );
  AOI21_X1 U10288 ( .B1(n9550), .B2(n8928), .A(n8863), .ZN(n8864) );
  OAI21_X1 U10289 ( .B1(n8865), .B2(n4653), .A(n8864), .ZN(P1_U3227) );
  NAND2_X1 U10290 ( .A1(n8867), .A2(n8866), .ZN(n8869) );
  OAI21_X1 U10291 ( .B1(n8870), .B2(n8869), .A(n8868), .ZN(n8871) );
  NAND2_X1 U10292 ( .A1(n8871), .A2(n8935), .ZN(n8876) );
  NOR2_X1 U10293 ( .A1(n8926), .A2(n9441), .ZN(n8874) );
  OAI22_X1 U10294 ( .A1(n8923), .A2(n9411), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8872), .ZN(n8873) );
  AOI211_X1 U10295 ( .C1(n8936), .C2(n9472), .A(n8874), .B(n8873), .ZN(n8875)
         );
  OAI211_X1 U10296 ( .C1(n9444), .C2(n8945), .A(n8876), .B(n8875), .ZN(
        P1_U3231) );
  OR2_X1 U10297 ( .A1(n8910), .A2(n8877), .ZN(n8880) );
  AND2_X1 U10298 ( .A1(n8880), .A2(n8878), .ZN(n8884) );
  NAND2_X1 U10299 ( .A1(n8880), .A2(n8879), .ZN(n8882) );
  NAND2_X1 U10300 ( .A1(n4293), .A2(n8883), .ZN(n8881) );
  AOI22_X1 U10301 ( .A1(n8884), .A2(n8883), .B1(n8882), .B2(n8881), .ZN(n8891)
         );
  AND2_X1 U10302 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9800) );
  NOR2_X1 U10303 ( .A1(n8897), .A2(n8885), .ZN(n8886) );
  AOI211_X1 U10304 ( .C1(n8942), .C2(n9248), .A(n9800), .B(n8886), .ZN(n8887)
         );
  OAI21_X1 U10305 ( .B1(n8926), .B2(n8888), .A(n8887), .ZN(n8889) );
  AOI21_X1 U10306 ( .B1(n8928), .B2(n9605), .A(n8889), .ZN(n8890) );
  OAI21_X1 U10307 ( .B1(n8891), .B2(n4653), .A(n8890), .ZN(P1_U3232) );
  OAI21_X1 U10308 ( .B1(n8895), .B2(n8893), .A(n8892), .ZN(n8894) );
  OAI211_X1 U10309 ( .C1(n4298), .C2(n8895), .A(n8935), .B(n8894), .ZN(n8901)
         );
  NOR2_X1 U10310 ( .A1(n8926), .A2(n9414), .ZN(n8899) );
  OAI22_X1 U10311 ( .A1(n8897), .A2(n9411), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8896), .ZN(n8898) );
  AOI211_X1 U10312 ( .C1(n8942), .C2(n9246), .A(n8899), .B(n8898), .ZN(n8900)
         );
  OAI211_X1 U10313 ( .C1(n8902), .C2(n8945), .A(n8901), .B(n8900), .ZN(
        P1_U3233) );
  INV_X1 U10314 ( .A(n8903), .ZN(n8904) );
  AOI21_X1 U10315 ( .B1(n8936), .B2(n9252), .A(n8904), .ZN(n8906) );
  NAND2_X1 U10316 ( .A1(n8942), .A2(n9250), .ZN(n8905) );
  OAI211_X1 U10317 ( .C1(n8926), .C2(n8907), .A(n8906), .B(n8905), .ZN(n8913)
         );
  INV_X1 U10318 ( .A(n8908), .ZN(n8909) );
  AOI211_X1 U10319 ( .C1(n8911), .C2(n8910), .A(n4653), .B(n8909), .ZN(n8912)
         );
  AOI211_X1 U10320 ( .C1(n8928), .C2(n8914), .A(n8913), .B(n8912), .ZN(n8915)
         );
  INV_X1 U10321 ( .A(n8915), .ZN(P1_U3234) );
  INV_X1 U10322 ( .A(n8916), .ZN(n8921) );
  AOI21_X1 U10323 ( .B1(n8918), .B2(n8920), .A(n8917), .ZN(n8919) );
  AOI21_X1 U10324 ( .B1(n8921), .B2(n8920), .A(n8919), .ZN(n8930) );
  NAND2_X1 U10325 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9860) );
  OAI21_X1 U10326 ( .B1(n8923), .B2(n8922), .A(n9860), .ZN(n8924) );
  AOI21_X1 U10327 ( .B1(n8936), .B2(n9471), .A(n8924), .ZN(n8925) );
  OAI21_X1 U10328 ( .B1(n8926), .B2(n9477), .A(n8925), .ZN(n8927) );
  AOI21_X1 U10329 ( .B1(n9582), .B2(n8928), .A(n8927), .ZN(n8929) );
  OAI21_X1 U10330 ( .B1(n8930), .B2(n4653), .A(n8929), .ZN(P1_U3236) );
  OAI21_X1 U10331 ( .B1(n8933), .B2(n8932), .A(n8931), .ZN(n8934) );
  NAND3_X1 U10332 ( .A1(n4656), .A2(n8935), .A3(n8934), .ZN(n8944) );
  NAND2_X1 U10333 ( .A1(n9355), .A2(n8936), .ZN(n8939) );
  NAND2_X1 U10334 ( .A1(n9349), .A2(n8937), .ZN(n8938) );
  OAI211_X1 U10335 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n8940), .A(n8939), .B(
        n8938), .ZN(n8941) );
  AOI21_X1 U10336 ( .B1(n9356), .B2(n8942), .A(n8941), .ZN(n8943) );
  OAI211_X1 U10337 ( .C1(n4553), .C2(n8945), .A(n8944), .B(n8943), .ZN(
        P1_U3238) );
  INV_X1 U10338 ( .A(n9214), .ZN(n9159) );
  NAND2_X1 U10339 ( .A1(n8946), .A2(n9159), .ZN(n8947) );
  NAND2_X1 U10340 ( .A1(n9219), .A2(n8947), .ZN(n8950) );
  INV_X1 U10341 ( .A(n9368), .ZN(n8948) );
  OAI21_X1 U10342 ( .B1(n9217), .B2(n8948), .A(n9351), .ZN(n8949) );
  MUX2_X1 U10343 ( .A(n8950), .B(n8949), .S(n9068), .Z(n9048) );
  AND2_X1 U10344 ( .A1(n9023), .A2(n8951), .ZN(n9021) );
  INV_X1 U10345 ( .A(n9121), .ZN(n8953) );
  AND2_X1 U10346 ( .A1(n9458), .A2(n8953), .ZN(n8952) );
  MUX2_X1 U10347 ( .A(n8952), .B(n9151), .S(n9068), .Z(n9019) );
  AND2_X1 U10348 ( .A1(n8953), .A2(n9468), .ZN(n9495) );
  MUX2_X1 U10349 ( .A(n9141), .B(n9120), .S(n9068), .Z(n9017) );
  INV_X1 U10350 ( .A(n9508), .ZN(n9015) );
  NAND4_X1 U10351 ( .A1(n8954), .A2(n9196), .A3(n9192), .A4(n9202), .ZN(n8961)
         );
  NAND2_X1 U10352 ( .A1(n9199), .A2(n9193), .ZN(n8956) );
  NAND3_X1 U10353 ( .A1(n8956), .A2(n8955), .A3(n9196), .ZN(n8957) );
  AND2_X1 U10354 ( .A1(n8957), .A2(n9200), .ZN(n8960) );
  AND2_X1 U10355 ( .A1(n8967), .A2(n8958), .ZN(n9203) );
  INV_X1 U10356 ( .A(n9203), .ZN(n8959) );
  AOI21_X1 U10357 ( .B1(n8961), .B2(n8960), .A(n8959), .ZN(n9145) );
  INV_X1 U10358 ( .A(n9145), .ZN(n8962) );
  NAND2_X1 U10359 ( .A1(n8962), .A2(n9122), .ZN(n8970) );
  INV_X1 U10360 ( .A(n9095), .ZN(n8963) );
  NAND2_X1 U10361 ( .A1(n8964), .A2(n8963), .ZN(n8966) );
  NAND3_X1 U10362 ( .A1(n8966), .A2(n9122), .A3(n8965), .ZN(n8968) );
  NAND2_X1 U10363 ( .A1(n8968), .A2(n8967), .ZN(n8969) );
  INV_X1 U10364 ( .A(n8971), .ZN(n8973) );
  OAI211_X1 U10365 ( .C1(n8982), .C2(n8973), .A(n8972), .B(n9123), .ZN(n8975)
         );
  NAND3_X1 U10366 ( .A1(n8975), .A2(n9130), .A3(n8974), .ZN(n8980) );
  NAND2_X1 U10367 ( .A1(n8977), .A2(n8976), .ZN(n8996) );
  AND2_X1 U10368 ( .A1(n8996), .A2(n9000), .ZN(n9124) );
  AND4_X1 U10369 ( .A1(n9125), .A2(n9103), .A3(n8978), .A4(n9068), .ZN(n8979)
         );
  NAND3_X1 U10370 ( .A1(n8980), .A2(n9124), .A3(n8979), .ZN(n9011) );
  OAI21_X1 U10371 ( .B1(n8982), .B2(n8981), .A(n9129), .ZN(n8985) );
  INV_X1 U10372 ( .A(n8983), .ZN(n8984) );
  NAND2_X1 U10373 ( .A1(n8985), .A2(n8984), .ZN(n8988) );
  AND2_X1 U10374 ( .A1(n9135), .A2(n8992), .ZN(n8999) );
  INV_X1 U10375 ( .A(n9068), .ZN(n9074) );
  NAND2_X1 U10376 ( .A1(n8990), .A2(n9074), .ZN(n9001) );
  INV_X1 U10377 ( .A(n9130), .ZN(n8986) );
  NOR2_X1 U10378 ( .A1(n9001), .A2(n8986), .ZN(n8987) );
  NAND4_X1 U10379 ( .A1(n8988), .A2(n8999), .A3(n8987), .A4(n9103), .ZN(n9010)
         );
  NAND2_X1 U10380 ( .A1(n8990), .A2(n8989), .ZN(n8991) );
  NAND2_X1 U10381 ( .A1(n8991), .A2(n9125), .ZN(n8993) );
  NAND2_X1 U10382 ( .A1(n8993), .A2(n8992), .ZN(n9131) );
  NAND3_X1 U10383 ( .A1(n9131), .A2(n9000), .A3(n9068), .ZN(n8994) );
  NAND2_X1 U10384 ( .A1(n8996), .A2(n8994), .ZN(n8995) );
  OAI21_X1 U10385 ( .B1(n8996), .B2(n9074), .A(n8995), .ZN(n8998) );
  OR2_X1 U10386 ( .A1(n9135), .A2(n9074), .ZN(n8997) );
  AND2_X1 U10387 ( .A1(n8998), .A2(n8997), .ZN(n9009) );
  INV_X1 U10388 ( .A(n8999), .ZN(n9007) );
  INV_X1 U10389 ( .A(n9000), .ZN(n9005) );
  INV_X1 U10390 ( .A(n9001), .ZN(n9004) );
  NAND2_X1 U10391 ( .A1(n9125), .A2(n9002), .ZN(n9003) );
  AOI22_X1 U10392 ( .A1(n9005), .A2(n9074), .B1(n9004), .B2(n9003), .ZN(n9006)
         );
  OR2_X1 U10393 ( .A1(n9007), .A2(n9006), .ZN(n9008) );
  NAND4_X1 U10394 ( .A1(n9011), .A2(n9010), .A3(n9009), .A4(n9008), .ZN(n9012)
         );
  NAND2_X1 U10395 ( .A1(n9012), .A2(n9105), .ZN(n9014) );
  MUX2_X1 U10396 ( .A(n9138), .B(n9140), .S(n9068), .Z(n9013) );
  NAND3_X1 U10397 ( .A1(n9015), .A2(n9014), .A3(n9013), .ZN(n9016) );
  NAND3_X1 U10398 ( .A1(n9495), .A2(n9017), .A3(n9016), .ZN(n9018) );
  NAND2_X1 U10399 ( .A1(n9019), .A2(n9018), .ZN(n9024) );
  INV_X1 U10400 ( .A(n9022), .ZN(n9119) );
  OR2_X1 U10401 ( .A1(n9084), .A2(n9119), .ZN(n9020) );
  AOI21_X1 U10402 ( .B1(n9021), .B2(n9024), .A(n9020), .ZN(n9026) );
  AND2_X1 U10403 ( .A1(n9022), .A2(n9458), .ZN(n9146) );
  NAND2_X1 U10404 ( .A1(n9085), .A2(n9023), .ZN(n9147) );
  AOI21_X1 U10405 ( .B1(n9146), .B2(n9024), .A(n9147), .ZN(n9025) );
  MUX2_X1 U10406 ( .A(n9026), .B(n9025), .S(n9068), .Z(n9030) );
  INV_X1 U10407 ( .A(n9085), .ZN(n9027) );
  OAI21_X1 U10408 ( .B1(n9030), .B2(n9027), .A(n9031), .ZN(n9029) );
  AND2_X1 U10409 ( .A1(n9155), .A2(n9149), .ZN(n9028) );
  AOI21_X1 U10410 ( .B1(n9029), .B2(n9028), .A(n4805), .ZN(n9038) );
  NAND2_X1 U10411 ( .A1(n9030), .A2(n9149), .ZN(n9036) );
  NAND2_X1 U10412 ( .A1(n9149), .A2(n9084), .ZN(n9032) );
  AND2_X1 U10413 ( .A1(n9032), .A2(n9031), .ZN(n9034) );
  AND2_X1 U10414 ( .A1(n9034), .A2(n9033), .ZN(n9118) );
  INV_X1 U10415 ( .A(n9155), .ZN(n9035) );
  AOI21_X1 U10416 ( .B1(n9036), .B2(n9118), .A(n9035), .ZN(n9037) );
  MUX2_X1 U10417 ( .A(n9038), .B(n9037), .S(n9068), .Z(n9040) );
  NAND3_X1 U10418 ( .A1(n9217), .A2(n9214), .A3(n9368), .ZN(n9039) );
  NOR2_X1 U10419 ( .A1(n9040), .A2(n9039), .ZN(n9047) );
  INV_X1 U10420 ( .A(n9169), .ZN(n9042) );
  NAND2_X1 U10421 ( .A1(n9041), .A2(n9068), .ZN(n9049) );
  NAND2_X1 U10422 ( .A1(n9042), .A2(n9049), .ZN(n9046) );
  OR2_X1 U10423 ( .A1(n9043), .A2(n9074), .ZN(n9044) );
  AND2_X1 U10424 ( .A1(n9162), .A2(n9044), .ZN(n9045) );
  OAI211_X1 U10425 ( .C1(n9048), .C2(n9047), .A(n9046), .B(n9045), .ZN(n9054)
         );
  INV_X1 U10426 ( .A(n9049), .ZN(n9050) );
  NAND2_X1 U10427 ( .A1(n9316), .A2(n9050), .ZN(n9052) );
  NAND2_X1 U10428 ( .A1(n9162), .A2(n9074), .ZN(n9051) );
  NAND2_X1 U10429 ( .A1(n9052), .A2(n9051), .ZN(n9053) );
  AND2_X1 U10430 ( .A1(n9054), .A2(n9053), .ZN(n9058) );
  NAND2_X1 U10431 ( .A1(n9058), .A2(n9059), .ZN(n9057) );
  AOI21_X1 U10432 ( .B1(n9057), .B2(n9056), .A(n9055), .ZN(n9064) );
  INV_X1 U10433 ( .A(n9058), .ZN(n9062) );
  AND2_X1 U10434 ( .A1(n9060), .A2(n9059), .ZN(n9161) );
  INV_X1 U10435 ( .A(n9167), .ZN(n9061) );
  AOI21_X1 U10436 ( .B1(n9062), .B2(n9161), .A(n9061), .ZN(n9063) );
  MUX2_X1 U10437 ( .A(n9064), .B(n9063), .S(n9068), .Z(n9067) );
  NAND2_X1 U10438 ( .A1(n9525), .A2(n9075), .ZN(n9069) );
  INV_X1 U10439 ( .A(n9244), .ZN(n9070) );
  OR2_X1 U10440 ( .A1(n9298), .A2(n9070), .ZN(n9065) );
  NAND2_X1 U10441 ( .A1(n9229), .A2(n9525), .ZN(n9175) );
  MUX2_X1 U10442 ( .A(n9223), .B(n9168), .S(n9068), .Z(n9066) );
  OAI211_X1 U10443 ( .C1(n9067), .C2(n9114), .A(n9175), .B(n9066), .ZN(n9073)
         );
  NAND2_X1 U10444 ( .A1(n9069), .A2(n9068), .ZN(n9072) );
  NAND2_X1 U10445 ( .A1(n9298), .A2(n9070), .ZN(n9224) );
  NAND2_X1 U10446 ( .A1(n9298), .A2(n9075), .ZN(n9071) );
  NAND2_X1 U10447 ( .A1(n9224), .A2(n9071), .ZN(n9170) );
  MUX2_X1 U10448 ( .A(n9073), .B(n9072), .S(n9170), .Z(n9078) );
  NAND3_X1 U10449 ( .A1(n9229), .A2(n9074), .A3(n9525), .ZN(n9076) );
  AND2_X1 U10450 ( .A1(n9076), .A2(n9230), .ZN(n9077) );
  AND2_X2 U10451 ( .A1(n9078), .A2(n9077), .ZN(n9180) );
  INV_X1 U10452 ( .A(n9079), .ZN(n9117) );
  INV_X1 U10453 ( .A(n9229), .ZN(n9116) );
  INV_X1 U10454 ( .A(n9317), .ZN(n9113) );
  INV_X1 U10455 ( .A(n9080), .ZN(n9081) );
  INV_X1 U10456 ( .A(n9083), .ZN(n9408) );
  INV_X1 U10457 ( .A(n9424), .ZN(n9110) );
  INV_X1 U10458 ( .A(n9084), .ZN(n9086) );
  AND2_X1 U10459 ( .A1(n9086), .A2(n9085), .ZN(n9445) );
  INV_X1 U10460 ( .A(n9495), .ZN(n9486) );
  INV_X1 U10461 ( .A(n9087), .ZN(n9102) );
  INV_X1 U10462 ( .A(n9089), .ZN(n9092) );
  NAND4_X1 U10463 ( .A1(n9093), .A2(n9092), .A3(n9091), .A4(n9090), .ZN(n9096)
         );
  NOR4_X1 U10464 ( .A1(n9096), .A2(n6844), .A3(n9095), .A4(n9094), .ZN(n9097)
         );
  NAND4_X1 U10465 ( .A1(n9099), .A2(n9098), .A3(n4829), .A4(n9097), .ZN(n9100)
         );
  NOR4_X1 U10466 ( .A1(n9102), .A2(n9101), .A3(n9676), .A4(n9100), .ZN(n9104)
         );
  NAND3_X1 U10467 ( .A1(n9105), .A2(n9104), .A3(n9103), .ZN(n9106) );
  NOR4_X1 U10468 ( .A1(n9486), .A2(n9107), .A3(n9508), .A4(n9106), .ZN(n9108)
         );
  NAND4_X1 U10469 ( .A1(n9445), .A2(n9457), .A3(n9481), .A4(n9108), .ZN(n9109)
         );
  NOR4_X1 U10470 ( .A1(n9391), .A2(n9408), .A3(n9110), .A4(n9109), .ZN(n9111)
         );
  XNOR2_X1 U10471 ( .A(n9550), .B(n9394), .ZN(n9379) );
  NAND4_X1 U10472 ( .A1(n9354), .A2(n9370), .A3(n9111), .A4(n9379), .ZN(n9112)
         );
  NOR4_X1 U10473 ( .A1(n9114), .A2(n9113), .A3(n9112), .A4(n9329), .ZN(n9115)
         );
  NAND4_X1 U10474 ( .A1(n9116), .A2(n9115), .A3(n9224), .A4(n9230), .ZN(n9177)
         );
  INV_X1 U10475 ( .A(n9118), .ZN(n9154) );
  NOR2_X1 U10476 ( .A1(n9154), .A2(n9119), .ZN(n9209) );
  NOR2_X1 U10477 ( .A1(n9121), .A2(n4819), .ZN(n9144) );
  NAND3_X1 U10478 ( .A1(n9138), .A2(n9123), .A3(n9122), .ZN(n9127) );
  INV_X1 U10479 ( .A(n9124), .ZN(n9133) );
  INV_X1 U10480 ( .A(n9125), .ZN(n9126) );
  OR3_X1 U10481 ( .A1(n9133), .A2(n9126), .A3(n4351), .ZN(n9137) );
  NOR2_X1 U10482 ( .A1(n9127), .A2(n9137), .ZN(n9128) );
  NAND3_X1 U10483 ( .A1(n9144), .A2(n9128), .A3(n9458), .ZN(n9207) );
  AND2_X1 U10484 ( .A1(n9130), .A2(n9129), .ZN(n9136) );
  INV_X1 U10485 ( .A(n9131), .ZN(n9132) );
  OR2_X1 U10486 ( .A1(n9133), .A2(n9132), .ZN(n9134) );
  OAI211_X1 U10487 ( .C1(n9137), .C2(n9136), .A(n9135), .B(n9134), .ZN(n9139)
         );
  NAND2_X1 U10488 ( .A1(n9139), .A2(n9138), .ZN(n9142) );
  NAND3_X1 U10489 ( .A1(n9142), .A2(n9141), .A3(n9140), .ZN(n9143) );
  NAND3_X1 U10490 ( .A1(n9144), .A2(n9458), .A3(n9143), .ZN(n9205) );
  OAI21_X1 U10491 ( .B1(n9207), .B2(n9145), .A(n9205), .ZN(n9157) );
  INV_X1 U10492 ( .A(n9146), .ZN(n9150) );
  INV_X1 U10493 ( .A(n9147), .ZN(n9148) );
  OAI211_X1 U10494 ( .C1(n9151), .C2(n9150), .A(n9149), .B(n9148), .ZN(n9152)
         );
  INV_X1 U10495 ( .A(n9152), .ZN(n9153) );
  OR2_X1 U10496 ( .A1(n9154), .A2(n9153), .ZN(n9156) );
  NAND2_X1 U10497 ( .A1(n9156), .A2(n9155), .ZN(n9210) );
  AOI21_X1 U10498 ( .B1(n9209), .B2(n9157), .A(n9210), .ZN(n9158) );
  OAI21_X1 U10499 ( .B1(n9159), .B2(n9158), .A(n9217), .ZN(n9160) );
  NAND2_X1 U10500 ( .A1(n9219), .A2(n9160), .ZN(n9166) );
  INV_X1 U10501 ( .A(n9161), .ZN(n9165) );
  INV_X1 U10502 ( .A(n9162), .ZN(n9163) );
  AND2_X1 U10503 ( .A1(n9316), .A2(n9163), .ZN(n9164) );
  OR2_X1 U10504 ( .A1(n9165), .A2(n9164), .ZN(n9222) );
  AOI21_X1 U10505 ( .B1(n9316), .B2(n9166), .A(n9222), .ZN(n9172) );
  OAI211_X1 U10506 ( .C1(n9222), .C2(n9169), .A(n9168), .B(n9167), .ZN(n9225)
         );
  INV_X1 U10507 ( .A(n9170), .ZN(n9171) );
  OAI211_X1 U10508 ( .C1(n9172), .C2(n9225), .A(n9171), .B(n9223), .ZN(n9174)
         );
  INV_X1 U10509 ( .A(n9230), .ZN(n9173) );
  AOI21_X1 U10510 ( .B1(n9175), .B2(n9174), .A(n9173), .ZN(n9176) );
  MUX2_X1 U10511 ( .A(n9177), .B(n9176), .S(n9186), .Z(n9178) );
  MUX2_X1 U10512 ( .A(n9179), .B(n9178), .S(n9878), .Z(n9184) );
  INV_X1 U10513 ( .A(n9180), .ZN(n9181) );
  NAND4_X1 U10514 ( .A1(n9181), .A2(n9186), .A3(n6414), .A4(n9230), .ZN(n9182)
         );
  AND3_X1 U10515 ( .A1(n9184), .A2(n9183), .A3(n9182), .ZN(n9243) );
  NAND2_X1 U10516 ( .A1(n9262), .A2(n6556), .ZN(n9188) );
  INV_X1 U10517 ( .A(n9185), .ZN(n9187) );
  NAND3_X1 U10518 ( .A1(n9188), .A2(n9187), .A3(n9186), .ZN(n9190) );
  NAND3_X1 U10519 ( .A1(n9190), .A2(n9193), .A3(n9189), .ZN(n9197) );
  NAND2_X1 U10520 ( .A1(n9192), .A2(n9191), .ZN(n9194) );
  NAND2_X1 U10521 ( .A1(n9194), .A2(n9193), .ZN(n9195) );
  OAI211_X1 U10522 ( .C1(n9198), .C2(n9197), .A(n9196), .B(n9195), .ZN(n9201)
         );
  NAND3_X1 U10523 ( .A1(n9201), .A2(n9200), .A3(n9199), .ZN(n9204) );
  AND3_X1 U10524 ( .A1(n9204), .A2(n9203), .A3(n9202), .ZN(n9206) );
  OAI21_X1 U10525 ( .B1(n9207), .B2(n9206), .A(n9205), .ZN(n9208) );
  INV_X1 U10526 ( .A(n9208), .ZN(n9213) );
  INV_X1 U10527 ( .A(n9209), .ZN(n9212) );
  INV_X1 U10528 ( .A(n9210), .ZN(n9211) );
  OAI21_X1 U10529 ( .B1(n9213), .B2(n9212), .A(n9211), .ZN(n9215) );
  NAND2_X1 U10530 ( .A1(n9215), .A2(n9214), .ZN(n9216) );
  NAND2_X1 U10531 ( .A1(n9217), .A2(n9216), .ZN(n9218) );
  NAND2_X1 U10532 ( .A1(n9219), .A2(n9218), .ZN(n9220) );
  AND2_X1 U10533 ( .A1(n9333), .A2(n9220), .ZN(n9221) );
  NOR2_X1 U10534 ( .A1(n9222), .A2(n9221), .ZN(n9226) );
  OAI211_X1 U10535 ( .C1(n9226), .C2(n9225), .A(n9224), .B(n9223), .ZN(n9227)
         );
  INV_X1 U10536 ( .A(n9227), .ZN(n9228) );
  OR2_X1 U10537 ( .A1(n9229), .A2(n9228), .ZN(n9231) );
  NAND2_X1 U10538 ( .A1(n9231), .A2(n9230), .ZN(n9236) );
  NAND3_X1 U10539 ( .A1(n9236), .A2(n9434), .A3(n9232), .ZN(n9234) );
  OAI211_X1 U10540 ( .C1(n9236), .C2(n9235), .A(n9234), .B(n9233), .ZN(n9242)
         );
  NOR3_X1 U10541 ( .A1(n9238), .A2(n9629), .A3(n9237), .ZN(n9241) );
  OAI21_X1 U10542 ( .B1(n5488), .B2(n9239), .A(P1_B_REG_SCAN_IN), .ZN(n9240)
         );
  OAI22_X1 U10543 ( .A1(n9243), .A2(n9242), .B1(n9241), .B2(n9240), .ZN(
        P1_U3240) );
  MUX2_X1 U10544 ( .A(n9244), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9261), .Z(
        P1_U3585) );
  MUX2_X1 U10545 ( .A(n9245), .B(P1_DATAO_REG_28__SCAN_IN), .S(n9261), .Z(
        P1_U3583) );
  MUX2_X1 U10546 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9356), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10547 ( .A(n9372), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9261), .Z(
        P1_U3581) );
  MUX2_X1 U10548 ( .A(n9355), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9261), .Z(
        P1_U3580) );
  MUX2_X1 U10549 ( .A(n9394), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9261), .Z(
        P1_U3579) );
  MUX2_X1 U10550 ( .A(n9246), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9261), .Z(
        P1_U3578) );
  MUX2_X1 U10551 ( .A(n9426), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9261), .Z(
        P1_U3577) );
  MUX2_X1 U10552 ( .A(n9447), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9261), .Z(
        P1_U3576) );
  MUX2_X1 U10553 ( .A(n9463), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9261), .Z(
        P1_U3575) );
  MUX2_X1 U10554 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9472), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10555 ( .A(n9500), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9261), .Z(
        P1_U3573) );
  MUX2_X1 U10556 ( .A(n9471), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9261), .Z(
        P1_U3572) );
  MUX2_X1 U10557 ( .A(n9498), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9261), .Z(
        P1_U3571) );
  MUX2_X1 U10558 ( .A(n9247), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9261), .Z(
        P1_U3570) );
  MUX2_X1 U10559 ( .A(n9248), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9261), .Z(
        P1_U3569) );
  MUX2_X1 U10560 ( .A(n9249), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9261), .Z(
        P1_U3568) );
  MUX2_X1 U10561 ( .A(n9250), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9261), .Z(
        P1_U3567) );
  MUX2_X1 U10562 ( .A(n9251), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9261), .Z(
        P1_U3566) );
  MUX2_X1 U10563 ( .A(n9252), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9261), .Z(
        P1_U3565) );
  MUX2_X1 U10564 ( .A(n9253), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9261), .Z(
        P1_U3564) );
  MUX2_X1 U10565 ( .A(n9254), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9261), .Z(
        P1_U3563) );
  MUX2_X1 U10566 ( .A(n9255), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9261), .Z(
        P1_U3562) );
  MUX2_X1 U10567 ( .A(n9256), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9261), .Z(
        P1_U3561) );
  MUX2_X1 U10568 ( .A(n9257), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9261), .Z(
        P1_U3560) );
  MUX2_X1 U10569 ( .A(n9258), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9261), .Z(
        P1_U3559) );
  MUX2_X1 U10570 ( .A(n9259), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9261), .Z(
        P1_U3558) );
  MUX2_X1 U10571 ( .A(n9260), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9261), .Z(
        P1_U3557) );
  MUX2_X1 U10572 ( .A(n9262), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9261), .Z(
        P1_U3556) );
  INV_X1 U10573 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9295) );
  NOR2_X1 U10574 ( .A1(n9263), .A2(n9275), .ZN(n9265) );
  NOR2_X1 U10575 ( .A1(n9265), .A2(n9264), .ZN(n9266) );
  NOR2_X1 U10576 ( .A1(n9266), .A2(n9276), .ZN(n9267) );
  NAND2_X1 U10577 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9831), .ZN(n9268) );
  OAI21_X1 U10578 ( .B1(n9831), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9268), .ZN(
        n9828) );
  AOI21_X1 U10579 ( .B1(n9831), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9827), .ZN(
        n9839) );
  OR2_X1 U10580 ( .A1(n9842), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9270) );
  NAND2_X1 U10581 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9842), .ZN(n9269) );
  NAND2_X1 U10582 ( .A1(n9270), .A2(n9269), .ZN(n9840) );
  NOR2_X1 U10583 ( .A1(n9839), .A2(n9840), .ZN(n9838) );
  AOI21_X1 U10584 ( .B1(n9842), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9838), .ZN(
        n9854) );
  OR2_X1 U10585 ( .A1(n9858), .A2(n9478), .ZN(n9272) );
  NAND2_X1 U10586 ( .A1(n9858), .A2(n9478), .ZN(n9271) );
  AND2_X1 U10587 ( .A1(n9272), .A2(n9271), .ZN(n9855) );
  NOR2_X1 U10588 ( .A1(n9854), .A2(n9855), .ZN(n9853) );
  AOI21_X1 U10589 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n9858), .A(n9853), .ZN(
        n9273) );
  XNOR2_X1 U10590 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9273), .ZN(n9291) );
  INV_X1 U10591 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9284) );
  XNOR2_X1 U10592 ( .A(n9858), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9865) );
  INV_X1 U10593 ( .A(n9842), .ZN(n9282) );
  XOR2_X1 U10594 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9842), .Z(n9849) );
  INV_X1 U10595 ( .A(n9831), .ZN(n9280) );
  INV_X1 U10596 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9279) );
  XOR2_X1 U10597 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9831), .Z(n9833) );
  NAND2_X1 U10598 ( .A1(n9819), .A2(n9277), .ZN(n9278) );
  XNOR2_X1 U10599 ( .A(n9277), .B(n9276), .ZN(n9821) );
  NAND2_X1 U10600 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n9821), .ZN(n9820) );
  NAND2_X1 U10601 ( .A1(n9833), .A2(n9834), .ZN(n9832) );
  NAND2_X1 U10602 ( .A1(n9849), .A2(n9848), .ZN(n9846) );
  OAI21_X1 U10603 ( .B1(n9282), .B2(n9281), .A(n9846), .ZN(n9864) );
  NOR2_X1 U10604 ( .A1(n9865), .A2(n9864), .ZN(n9863) );
  XOR2_X1 U10605 ( .A(n9286), .B(n9285), .Z(n9289) );
  AOI21_X1 U10606 ( .B1(n9289), .B2(n9847), .A(n9859), .ZN(n9287) );
  INV_X1 U10607 ( .A(n9289), .ZN(n9290) );
  AOI22_X1 U10608 ( .A1(n9291), .A2(n9857), .B1(n9290), .B2(n9847), .ZN(n9292)
         );
  OAI211_X1 U10609 ( .C1(n9295), .C2(n9870), .A(n9294), .B(n9293), .ZN(
        P1_U3260) );
  INV_X1 U10610 ( .A(n9298), .ZN(n9711) );
  AOI21_X1 U10611 ( .B1(n9298), .B2(n9297), .A(n9296), .ZN(n9714) );
  NAND2_X1 U10612 ( .A1(n9714), .A2(n9504), .ZN(n9301) );
  AOI21_X1 U10613 ( .B1(n9887), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9299), .ZN(
        n9300) );
  OAI211_X1 U10614 ( .C1(n9711), .C2(n9519), .A(n9301), .B(n9300), .ZN(
        P1_U3262) );
  INV_X1 U10615 ( .A(n9302), .ZN(n9313) );
  INV_X1 U10616 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9303) );
  OAI22_X1 U10617 ( .A1(n9304), .A2(n9876), .B1(n9303), .B2(n9885), .ZN(n9305)
         );
  AOI21_X1 U10618 ( .B1(n9306), .B2(n9693), .A(n9305), .ZN(n9307) );
  OAI21_X1 U10619 ( .B1(n9309), .B2(n9308), .A(n9307), .ZN(n9310) );
  AOI21_X1 U10620 ( .B1(n9311), .B2(n9885), .A(n9310), .ZN(n9312) );
  OAI21_X1 U10621 ( .B1(n9313), .B2(n9524), .A(n9312), .ZN(P1_U3355) );
  AOI21_X1 U10622 ( .B1(n9317), .B2(n9314), .A(n4336), .ZN(n9315) );
  INV_X1 U10623 ( .A(n9315), .ZN(n9532) );
  NAND2_X1 U10624 ( .A1(n9332), .A2(n9316), .ZN(n9318) );
  XNOR2_X1 U10625 ( .A(n9318), .B(n9317), .ZN(n9319) );
  OAI222_X1 U10626 ( .A1(n9681), .A2(n9321), .B1(n9682), .B2(n9320), .C1(n9510), .C2(n9319), .ZN(n9528) );
  INV_X1 U10627 ( .A(n9530), .ZN(n9326) );
  AOI211_X1 U10628 ( .C1(n9530), .C2(n9338), .A(n9921), .B(n4551), .ZN(n9529)
         );
  NAND2_X1 U10629 ( .A1(n9529), .A2(n9698), .ZN(n9325) );
  AOI22_X1 U10630 ( .A1(n9323), .A2(n9690), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9692), .ZN(n9324) );
  OAI211_X1 U10631 ( .C1(n9326), .C2(n9519), .A(n9325), .B(n9324), .ZN(n9327)
         );
  AOI21_X1 U10632 ( .B1(n9528), .B2(n9885), .A(n9327), .ZN(n9328) );
  OAI21_X1 U10633 ( .B1(n9532), .B2(n9524), .A(n9328), .ZN(P1_U3263) );
  XNOR2_X1 U10634 ( .A(n9330), .B(n9329), .ZN(n9537) );
  INV_X1 U10635 ( .A(n9331), .ZN(n9334) );
  OAI211_X1 U10636 ( .C1(n9334), .C2(n9333), .A(n9332), .B(n9685), .ZN(n9336)
         );
  NAND2_X1 U10637 ( .A1(n9372), .A2(n9497), .ZN(n9335) );
  OAI211_X1 U10638 ( .C1(n9337), .C2(n9681), .A(n9336), .B(n9335), .ZN(n9533)
         );
  INV_X1 U10639 ( .A(n9348), .ZN(n9340) );
  INV_X1 U10640 ( .A(n9338), .ZN(n9339) );
  AOI211_X1 U10641 ( .C1(n9535), .C2(n9340), .A(n9921), .B(n9339), .ZN(n9534)
         );
  NAND2_X1 U10642 ( .A1(n9534), .A2(n9698), .ZN(n9343) );
  AOI22_X1 U10643 ( .A1(n9341), .A2(n9690), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9692), .ZN(n9342) );
  OAI211_X1 U10644 ( .C1(n9344), .C2(n9519), .A(n9343), .B(n9342), .ZN(n9345)
         );
  AOI21_X1 U10645 ( .B1(n9533), .B2(n9885), .A(n9345), .ZN(n9346) );
  OAI21_X1 U10646 ( .B1(n9537), .B2(n9524), .A(n9346), .ZN(P1_U3264) );
  XNOR2_X1 U10647 ( .A(n9347), .B(n9354), .ZN(n9542) );
  AOI21_X1 U10648 ( .B1(n9538), .B2(n9362), .A(n9348), .ZN(n9539) );
  AOI22_X1 U10649 ( .A1(n9349), .A2(n9690), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9887), .ZN(n9350) );
  OAI21_X1 U10650 ( .B1(n4553), .B2(n9519), .A(n9350), .ZN(n9359) );
  NAND2_X1 U10651 ( .A1(n9352), .A2(n9351), .ZN(n9353) );
  XOR2_X1 U10652 ( .A(n9354), .B(n9353), .Z(n9357) );
  AOI222_X1 U10653 ( .A1(n9685), .A2(n9357), .B1(n9356), .B2(n9499), .C1(n9355), .C2(n9497), .ZN(n9541) );
  NOR2_X1 U10654 ( .A1(n9541), .A2(n9887), .ZN(n9358) );
  AOI211_X1 U10655 ( .C1(n9539), .C2(n9504), .A(n9359), .B(n9358), .ZN(n9360)
         );
  OAI21_X1 U10656 ( .B1(n9542), .B2(n9524), .A(n9360), .ZN(P1_U3265) );
  XOR2_X1 U10657 ( .A(n9370), .B(n9361), .Z(n9547) );
  INV_X1 U10658 ( .A(n9362), .ZN(n9363) );
  AOI21_X1 U10659 ( .B1(n9543), .B2(n4557), .A(n9363), .ZN(n9544) );
  INV_X1 U10660 ( .A(n9364), .ZN(n9365) );
  AOI22_X1 U10661 ( .A1(n9365), .A2(n9690), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9887), .ZN(n9366) );
  OAI21_X1 U10662 ( .B1(n9367), .B2(n9519), .A(n9366), .ZN(n9375) );
  NAND2_X1 U10663 ( .A1(n9369), .A2(n9368), .ZN(n9371) );
  XNOR2_X1 U10664 ( .A(n9371), .B(n9370), .ZN(n9373) );
  AOI222_X1 U10665 ( .A1(n9685), .A2(n9373), .B1(n9372), .B2(n9499), .C1(n9394), .C2(n9497), .ZN(n9546) );
  NOR2_X1 U10666 ( .A1(n9546), .A2(n9692), .ZN(n9374) );
  AOI211_X1 U10667 ( .C1(n9544), .C2(n9504), .A(n9375), .B(n9374), .ZN(n9376)
         );
  OAI21_X1 U10668 ( .B1(n9547), .B2(n9524), .A(n9376), .ZN(P1_U3266) );
  XOR2_X1 U10669 ( .A(n9379), .B(n9377), .Z(n9552) );
  NAND2_X1 U10670 ( .A1(n9392), .A2(n9378), .ZN(n9380) );
  XNOR2_X1 U10671 ( .A(n9380), .B(n9379), .ZN(n9381) );
  OAI222_X1 U10672 ( .A1(n9681), .A2(n9382), .B1(n9682), .B2(n9412), .C1(n9381), .C2(n9510), .ZN(n9548) );
  AOI211_X1 U10673 ( .C1(n9550), .C2(n9397), .A(n9921), .B(n9383), .ZN(n9549)
         );
  NAND2_X1 U10674 ( .A1(n9549), .A2(n9698), .ZN(n9386) );
  AOI22_X1 U10675 ( .A1(n9384), .A2(n9690), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9692), .ZN(n9385) );
  OAI211_X1 U10676 ( .C1(n9387), .C2(n9519), .A(n9386), .B(n9385), .ZN(n9388)
         );
  AOI21_X1 U10677 ( .B1(n9548), .B2(n9885), .A(n9388), .ZN(n9389) );
  OAI21_X1 U10678 ( .B1(n9552), .B2(n9524), .A(n9389), .ZN(P1_U3267) );
  XNOR2_X1 U10679 ( .A(n9390), .B(n9391), .ZN(n9557) );
  INV_X1 U10680 ( .A(n9391), .ZN(n9393) );
  OAI211_X1 U10681 ( .C1(n4304), .C2(n9393), .A(n9392), .B(n9685), .ZN(n9396)
         );
  AOI22_X1 U10682 ( .A1(n9394), .A2(n9499), .B1(n9497), .B2(n9426), .ZN(n9395)
         );
  NAND2_X1 U10683 ( .A1(n9396), .A2(n9395), .ZN(n9553) );
  INV_X1 U10684 ( .A(n9397), .ZN(n9398) );
  AOI211_X1 U10685 ( .C1(n9555), .C2(n9399), .A(n9921), .B(n9398), .ZN(n9554)
         );
  NAND2_X1 U10686 ( .A1(n9554), .A2(n9698), .ZN(n9403) );
  INV_X1 U10687 ( .A(n9400), .ZN(n9401) );
  AOI22_X1 U10688 ( .A1(n9401), .A2(n9690), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9692), .ZN(n9402) );
  OAI211_X1 U10689 ( .C1(n9404), .C2(n9519), .A(n9403), .B(n9402), .ZN(n9405)
         );
  AOI21_X1 U10690 ( .B1(n9553), .B2(n9885), .A(n9405), .ZN(n9406) );
  OAI21_X1 U10691 ( .B1(n9557), .B2(n9524), .A(n9406), .ZN(P1_U3268) );
  XNOR2_X1 U10692 ( .A(n9407), .B(n9408), .ZN(n9562) );
  AOI22_X1 U10693 ( .A1(n9560), .A2(n9693), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9692), .ZN(n9418) );
  XNOR2_X1 U10694 ( .A(n9409), .B(n9408), .ZN(n9410) );
  OAI222_X1 U10695 ( .A1(n9681), .A2(n9412), .B1(n9682), .B2(n9411), .C1(n9410), .C2(n9510), .ZN(n9558) );
  AOI211_X1 U10696 ( .C1(n9560), .C2(n9430), .A(n9921), .B(n9413), .ZN(n9559)
         );
  INV_X1 U10697 ( .A(n9559), .ZN(n9415) );
  OAI22_X1 U10698 ( .A1(n9415), .A2(n9434), .B1(n9876), .B2(n9414), .ZN(n9416)
         );
  OAI21_X1 U10699 ( .B1(n9558), .B2(n9416), .A(n9885), .ZN(n9417) );
  OAI211_X1 U10700 ( .C1(n9562), .C2(n9524), .A(n9418), .B(n9417), .ZN(
        P1_U3269) );
  NAND2_X1 U10701 ( .A1(n9419), .A2(n9424), .ZN(n9420) );
  NAND2_X1 U10702 ( .A1(n9421), .A2(n9420), .ZN(n9563) );
  AOI22_X1 U10703 ( .A1(n9429), .A2(n9693), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9692), .ZN(n9437) );
  OAI21_X1 U10704 ( .B1(n9424), .B2(n9423), .A(n9422), .ZN(n9425) );
  NAND2_X1 U10705 ( .A1(n9425), .A2(n9685), .ZN(n9428) );
  AOI22_X1 U10706 ( .A1(n9426), .A2(n9499), .B1(n9497), .B2(n9463), .ZN(n9427)
         );
  NAND2_X1 U10707 ( .A1(n9428), .A2(n9427), .ZN(n9567) );
  AOI21_X1 U10708 ( .B1(n9439), .B2(n9429), .A(n9921), .ZN(n9431) );
  NAND2_X1 U10709 ( .A1(n9431), .A2(n9430), .ZN(n9564) );
  INV_X1 U10710 ( .A(n9432), .ZN(n9433) );
  OAI22_X1 U10711 ( .A1(n9564), .A2(n9434), .B1(n9876), .B2(n9433), .ZN(n9435)
         );
  OAI21_X1 U10712 ( .B1(n9567), .B2(n9435), .A(n9885), .ZN(n9436) );
  OAI211_X1 U10713 ( .C1(n9563), .C2(n9524), .A(n9437), .B(n9436), .ZN(
        P1_U3270) );
  XOR2_X1 U10714 ( .A(n9445), .B(n9438), .Z(n9574) );
  INV_X1 U10715 ( .A(n9439), .ZN(n9440) );
  AOI21_X1 U10716 ( .B1(n9570), .B2(n4548), .A(n9440), .ZN(n9571) );
  INV_X1 U10717 ( .A(n9441), .ZN(n9442) );
  AOI22_X1 U10718 ( .A1(n9692), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9442), .B2(
        n9690), .ZN(n9443) );
  OAI21_X1 U10719 ( .B1(n9444), .B2(n9519), .A(n9443), .ZN(n9450) );
  XNOR2_X1 U10720 ( .A(n9446), .B(n9445), .ZN(n9448) );
  AOI222_X1 U10721 ( .A1(n9685), .A2(n9448), .B1(n9447), .B2(n9499), .C1(n9472), .C2(n9497), .ZN(n9573) );
  NOR2_X1 U10722 ( .A1(n9573), .A2(n9692), .ZN(n9449) );
  AOI211_X1 U10723 ( .C1(n9571), .C2(n9504), .A(n9450), .B(n9449), .ZN(n9451)
         );
  OAI21_X1 U10724 ( .B1(n9524), .B2(n9574), .A(n9451), .ZN(P1_U3271) );
  XOR2_X1 U10725 ( .A(n9452), .B(n9457), .Z(n9579) );
  AOI21_X1 U10726 ( .B1(n9575), .B2(n9474), .A(n9453), .ZN(n9576) );
  INV_X1 U10727 ( .A(n9454), .ZN(n9455) );
  AOI22_X1 U10728 ( .A1(n9692), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9455), .B2(
        n9690), .ZN(n9456) );
  OAI21_X1 U10729 ( .B1(n4546), .B2(n9519), .A(n9456), .ZN(n9466) );
  INV_X1 U10730 ( .A(n9457), .ZN(n9459) );
  NAND3_X1 U10731 ( .A1(n9460), .A2(n9459), .A3(n9458), .ZN(n9461) );
  NAND2_X1 U10732 ( .A1(n9462), .A2(n9461), .ZN(n9464) );
  AOI222_X1 U10733 ( .A1(n9685), .A2(n9464), .B1(n9463), .B2(n9499), .C1(n9500), .C2(n9497), .ZN(n9578) );
  NOR2_X1 U10734 ( .A1(n9578), .A2(n9692), .ZN(n9465) );
  AOI211_X1 U10735 ( .C1(n9576), .C2(n9504), .A(n9466), .B(n9465), .ZN(n9467)
         );
  OAI21_X1 U10736 ( .B1(n9524), .B2(n9579), .A(n9467), .ZN(P1_U3272) );
  NAND2_X1 U10737 ( .A1(n9469), .A2(n9468), .ZN(n9470) );
  XOR2_X1 U10738 ( .A(n9481), .B(n9470), .Z(n9473) );
  AOI222_X1 U10739 ( .A1(n9685), .A2(n9473), .B1(n9472), .B2(n9499), .C1(n9471), .C2(n9497), .ZN(n9585) );
  INV_X1 U10740 ( .A(n9474), .ZN(n9475) );
  AOI21_X1 U10741 ( .B1(n9582), .B2(n9488), .A(n9475), .ZN(n9583) );
  INV_X1 U10742 ( .A(n9582), .ZN(n9476) );
  NOR2_X1 U10743 ( .A1(n9476), .A2(n9519), .ZN(n9480) );
  OAI22_X1 U10744 ( .A1(n9885), .A2(n9478), .B1(n9477), .B2(n9876), .ZN(n9479)
         );
  AOI211_X1 U10745 ( .C1(n9583), .C2(n9504), .A(n9480), .B(n9479), .ZN(n9485)
         );
  NAND2_X1 U10746 ( .A1(n9482), .A2(n9481), .ZN(n9580) );
  NAND3_X1 U10747 ( .A1(n9581), .A2(n9580), .A3(n9483), .ZN(n9484) );
  OAI211_X1 U10748 ( .C1(n9585), .C2(n9692), .A(n9485), .B(n9484), .ZN(
        P1_U3273) );
  XNOR2_X1 U10749 ( .A(n9487), .B(n9486), .ZN(n9591) );
  INV_X1 U10750 ( .A(n9516), .ZN(n9490) );
  INV_X1 U10751 ( .A(n9488), .ZN(n9489) );
  AOI21_X1 U10752 ( .B1(n9587), .B2(n9490), .A(n9489), .ZN(n9588) );
  INV_X1 U10753 ( .A(n9491), .ZN(n9492) );
  AOI22_X1 U10754 ( .A1(n9692), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9492), .B2(
        n9690), .ZN(n9493) );
  OAI21_X1 U10755 ( .B1(n9494), .B2(n9519), .A(n9493), .ZN(n9503) );
  XNOR2_X1 U10756 ( .A(n9496), .B(n9495), .ZN(n9501) );
  AOI222_X1 U10757 ( .A1(n9685), .A2(n9501), .B1(n9500), .B2(n9499), .C1(n9498), .C2(n9497), .ZN(n9590) );
  NOR2_X1 U10758 ( .A1(n9590), .A2(n9887), .ZN(n9502) );
  AOI211_X1 U10759 ( .C1(n9588), .C2(n9504), .A(n9503), .B(n9502), .ZN(n9505)
         );
  OAI21_X1 U10760 ( .B1(n9524), .B2(n9591), .A(n9505), .ZN(P1_U3274) );
  XNOR2_X1 U10761 ( .A(n9506), .B(n9508), .ZN(n9596) );
  AOI21_X1 U10762 ( .B1(n9508), .B2(n9507), .A(n4345), .ZN(n9509) );
  OAI222_X1 U10763 ( .A1(n9681), .A2(n9512), .B1(n9682), .B2(n9511), .C1(n9510), .C2(n9509), .ZN(n9592) );
  NOR2_X1 U10764 ( .A1(n9876), .A2(n9513), .ZN(n9514) );
  OAI21_X1 U10765 ( .B1(n9592), .B2(n9514), .A(n9885), .ZN(n9523) );
  INV_X1 U10766 ( .A(n9515), .ZN(n9517) );
  AOI211_X1 U10767 ( .C1(n9594), .C2(n9517), .A(n9921), .B(n9516), .ZN(n9593)
         );
  INV_X1 U10768 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9518) );
  OAI22_X1 U10769 ( .A1(n9520), .A2(n9519), .B1(n9518), .B2(n9885), .ZN(n9521)
         );
  AOI21_X1 U10770 ( .B1(n9593), .B2(n9698), .A(n9521), .ZN(n9522) );
  OAI211_X1 U10771 ( .C1(n9596), .C2(n9524), .A(n9523), .B(n9522), .ZN(
        P1_U3275) );
  NAND2_X1 U10772 ( .A1(n9525), .A2(n9606), .ZN(n9526) );
  OAI211_X1 U10773 ( .C1(n9527), .C2(n9921), .A(n9710), .B(n9526), .ZN(n9613)
         );
  MUX2_X1 U10774 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9613), .S(n9935), .Z(
        P1_U3554) );
  AOI211_X1 U10775 ( .C1(n9606), .C2(n9530), .A(n9529), .B(n9528), .ZN(n9531)
         );
  OAI21_X1 U10776 ( .B1(n9532), .B2(n9597), .A(n9531), .ZN(n9614) );
  MUX2_X1 U10777 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9614), .S(n9935), .Z(
        P1_U3551) );
  AOI211_X1 U10778 ( .C1(n9606), .C2(n9535), .A(n9534), .B(n9533), .ZN(n9536)
         );
  OAI21_X1 U10779 ( .B1(n9537), .B2(n9597), .A(n9536), .ZN(n9615) );
  MUX2_X1 U10780 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9615), .S(n9935), .Z(
        P1_U3550) );
  AOI22_X1 U10781 ( .A1(n9539), .A2(n9713), .B1(n9606), .B2(n9538), .ZN(n9540)
         );
  OAI211_X1 U10782 ( .C1(n9542), .C2(n9597), .A(n9541), .B(n9540), .ZN(n9616)
         );
  MUX2_X1 U10783 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9616), .S(n9935), .Z(
        P1_U3549) );
  AOI22_X1 U10784 ( .A1(n9544), .A2(n9713), .B1(n9606), .B2(n9543), .ZN(n9545)
         );
  OAI211_X1 U10785 ( .C1(n9547), .C2(n9597), .A(n9546), .B(n9545), .ZN(n9617)
         );
  MUX2_X1 U10786 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9617), .S(n9935), .Z(
        P1_U3548) );
  AOI211_X1 U10787 ( .C1(n9606), .C2(n9550), .A(n9549), .B(n9548), .ZN(n9551)
         );
  OAI21_X1 U10788 ( .B1(n9552), .B2(n9597), .A(n9551), .ZN(n9618) );
  MUX2_X1 U10789 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9618), .S(n9935), .Z(
        P1_U3547) );
  AOI211_X1 U10790 ( .C1(n9606), .C2(n9555), .A(n9554), .B(n9553), .ZN(n9556)
         );
  OAI21_X1 U10791 ( .B1(n9557), .B2(n9597), .A(n9556), .ZN(n9619) );
  MUX2_X1 U10792 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9619), .S(n9935), .Z(
        P1_U3546) );
  AOI211_X1 U10793 ( .C1(n9606), .C2(n9560), .A(n9559), .B(n9558), .ZN(n9561)
         );
  OAI21_X1 U10794 ( .B1(n9562), .B2(n9597), .A(n9561), .ZN(n9620) );
  MUX2_X1 U10795 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9620), .S(n9935), .Z(
        P1_U3545) );
  OR2_X1 U10796 ( .A1(n9563), .A2(n9597), .ZN(n9569) );
  OAI21_X1 U10797 ( .B1(n9565), .B2(n9911), .A(n9564), .ZN(n9566) );
  NOR2_X1 U10798 ( .A1(n9567), .A2(n9566), .ZN(n9568) );
  NAND2_X1 U10799 ( .A1(n9569), .A2(n9568), .ZN(n9621) );
  MUX2_X1 U10800 ( .A(n9621), .B(P1_REG1_REG_21__SCAN_IN), .S(n9933), .Z(
        P1_U3544) );
  AOI22_X1 U10801 ( .A1(n9571), .A2(n9713), .B1(n9606), .B2(n9570), .ZN(n9572)
         );
  OAI211_X1 U10802 ( .C1(n9574), .C2(n9597), .A(n9573), .B(n9572), .ZN(n9622)
         );
  MUX2_X1 U10803 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9622), .S(n9935), .Z(
        P1_U3543) );
  AOI22_X1 U10804 ( .A1(n9576), .A2(n9713), .B1(n9606), .B2(n9575), .ZN(n9577)
         );
  OAI211_X1 U10805 ( .C1(n9579), .C2(n9597), .A(n9578), .B(n9577), .ZN(n9623)
         );
  MUX2_X1 U10806 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9623), .S(n9935), .Z(
        P1_U3542) );
  NAND3_X1 U10807 ( .A1(n9581), .A2(n9926), .A3(n9580), .ZN(n9586) );
  AOI22_X1 U10808 ( .A1(n9583), .A2(n9713), .B1(n9606), .B2(n9582), .ZN(n9584)
         );
  NAND3_X1 U10809 ( .A1(n9586), .A2(n9585), .A3(n9584), .ZN(n9624) );
  MUX2_X1 U10810 ( .A(n9624), .B(P1_REG1_REG_18__SCAN_IN), .S(n9933), .Z(
        P1_U3541) );
  AOI22_X1 U10811 ( .A1(n9588), .A2(n9713), .B1(n9606), .B2(n9587), .ZN(n9589)
         );
  OAI211_X1 U10812 ( .C1(n9591), .C2(n9597), .A(n9590), .B(n9589), .ZN(n9625)
         );
  MUX2_X1 U10813 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9625), .S(n9935), .Z(
        P1_U3540) );
  AOI211_X1 U10814 ( .C1(n9606), .C2(n9594), .A(n9593), .B(n9592), .ZN(n9595)
         );
  OAI21_X1 U10815 ( .B1(n9597), .B2(n9596), .A(n9595), .ZN(n9626) );
  MUX2_X1 U10816 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9626), .S(n9935), .Z(
        P1_U3539) );
  AND2_X1 U10817 ( .A1(n9598), .A2(n9917), .ZN(n9604) );
  INV_X1 U10818 ( .A(n9599), .ZN(n9600) );
  OAI22_X1 U10819 ( .A1(n9601), .A2(n9921), .B1(n9600), .B2(n9911), .ZN(n9602)
         );
  MUX2_X1 U10820 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9627), .S(n9935), .Z(
        P1_U3538) );
  AOI22_X1 U10821 ( .A1(n9607), .A2(n9713), .B1(n9606), .B2(n9605), .ZN(n9608)
         );
  OAI21_X1 U10822 ( .B1(n9610), .B2(n9609), .A(n9608), .ZN(n9611) );
  OR2_X1 U10823 ( .A1(n9612), .A2(n9611), .ZN(n9628) );
  MUX2_X1 U10824 ( .A(n9628), .B(P1_REG1_REG_13__SCAN_IN), .S(n9933), .Z(
        P1_U3536) );
  MUX2_X1 U10825 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9613), .S(n9929), .Z(
        P1_U3522) );
  MUX2_X1 U10826 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9614), .S(n9929), .Z(
        P1_U3519) );
  MUX2_X1 U10827 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9615), .S(n9929), .Z(
        P1_U3518) );
  MUX2_X1 U10828 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9616), .S(n9929), .Z(
        P1_U3517) );
  MUX2_X1 U10829 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9617), .S(n9929), .Z(
        P1_U3516) );
  MUX2_X1 U10830 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9618), .S(n9929), .Z(
        P1_U3515) );
  MUX2_X1 U10831 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9619), .S(n9929), .Z(
        P1_U3514) );
  MUX2_X1 U10832 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9620), .S(n9929), .Z(
        P1_U3513) );
  MUX2_X1 U10833 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9621), .S(n9929), .Z(
        P1_U3512) );
  MUX2_X1 U10834 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9622), .S(n9929), .Z(
        P1_U3511) );
  MUX2_X1 U10835 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9623), .S(n9929), .Z(
        P1_U3510) );
  MUX2_X1 U10836 ( .A(n9624), .B(P1_REG0_REG_18__SCAN_IN), .S(n9927), .Z(
        P1_U3508) );
  MUX2_X1 U10837 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9625), .S(n9929), .Z(
        P1_U3505) );
  MUX2_X1 U10838 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9626), .S(n9929), .Z(
        P1_U3502) );
  MUX2_X1 U10839 ( .A(n9627), .B(P1_REG0_REG_15__SCAN_IN), .S(n9927), .Z(
        P1_U3499) );
  MUX2_X1 U10840 ( .A(n9628), .B(P1_REG0_REG_13__SCAN_IN), .S(n9927), .Z(
        P1_U3493) );
  MUX2_X1 U10841 ( .A(n9630), .B(P1_D_REG_0__SCAN_IN), .S(n9629), .Z(P1_U3440)
         );
  NOR4_X1 U10842 ( .A1(n9632), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n9631), .ZN(n9633) );
  AOI21_X1 U10843 ( .B1(n9634), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9633), .ZN(
        n9635) );
  OAI21_X1 U10844 ( .B1(n9636), .B2(n9639), .A(n9635), .ZN(P1_U3322) );
  OAI222_X1 U10845 ( .A1(n9641), .A2(n9640), .B1(n9639), .B2(n9638), .C1(
        P1_U3084), .C2(n9637), .ZN(P1_U3323) );
  OAI222_X1 U10846 ( .A1(n9645), .A2(n9644), .B1(n9643), .B2(P1_U3084), .C1(
        n9642), .C2(n9641), .ZN(P1_U3324) );
  MUX2_X1 U10847 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9647), .S(P1_U3084), .Z(
        P1_U3353) );
  OAI22_X1 U10848 ( .A1(n9650), .A2(n9649), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9648), .ZN(n9655) );
  NAND2_X1 U10849 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9653) );
  AOI211_X1 U10850 ( .C1(n9653), .C2(n9652), .A(n9651), .B(n9662), .ZN(n9654)
         );
  AOI211_X1 U10851 ( .C1(n9668), .C2(n9656), .A(n9655), .B(n9654), .ZN(n9661)
         );
  INV_X1 U10852 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10102) );
  NOR2_X1 U10853 ( .A1(n9946), .A2(n10102), .ZN(n9659) );
  OAI211_X1 U10854 ( .C1(n9659), .C2(n9658), .A(n9936), .B(n9657), .ZN(n9660)
         );
  NAND2_X1 U10855 ( .A1(n9661), .A2(n9660), .ZN(P2_U3246) );
  AOI22_X1 U10856 ( .A1(n9943), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9674) );
  AOI211_X1 U10857 ( .C1(n9665), .C2(n9664), .A(n9663), .B(n9662), .ZN(n9666)
         );
  AOI21_X1 U10858 ( .B1(n9668), .B2(n9667), .A(n9666), .ZN(n9673) );
  OAI211_X1 U10859 ( .C1(n9671), .C2(n9670), .A(n9936), .B(n9669), .ZN(n9672)
         );
  NAND3_X1 U10860 ( .A1(n9674), .A2(n9673), .A3(n9672), .ZN(P2_U3247) );
  XNOR2_X1 U10861 ( .A(n9675), .B(n9676), .ZN(n9707) );
  OAI21_X1 U10862 ( .B1(n9679), .B2(n9678), .A(n9677), .ZN(n9686) );
  OAI22_X1 U10863 ( .A1(n9683), .A2(n9682), .B1(n9681), .B2(n9680), .ZN(n9684)
         );
  AOI21_X1 U10864 ( .B1(n9686), .B2(n9685), .A(n9684), .ZN(n9704) );
  INV_X1 U10865 ( .A(n9704), .ZN(n9687) );
  AOI21_X1 U10866 ( .B1(n9707), .B2(n9688), .A(n9687), .ZN(n9702) );
  INV_X1 U10867 ( .A(n9689), .ZN(n9691) );
  AOI222_X1 U10868 ( .A1(n9694), .A2(n9693), .B1(P1_REG2_REG_10__SCAN_IN), 
        .B2(n9692), .C1(n9691), .C2(n9690), .ZN(n9701) );
  INV_X1 U10869 ( .A(n9694), .ZN(n9705) );
  OAI211_X1 U10870 ( .C1(n9696), .C2(n9705), .A(n9713), .B(n9695), .ZN(n9703)
         );
  INV_X1 U10871 ( .A(n9703), .ZN(n9697) );
  AOI22_X1 U10872 ( .A1(n9707), .A2(n9699), .B1(n9698), .B2(n9697), .ZN(n9700)
         );
  OAI211_X1 U10873 ( .C1(n9887), .C2(n9702), .A(n9701), .B(n9700), .ZN(
        P1_U3281) );
  OAI211_X1 U10874 ( .C1(n9705), .C2(n9911), .A(n9704), .B(n9703), .ZN(n9706)
         );
  AOI21_X1 U10875 ( .B1(n9707), .B2(n9926), .A(n9706), .ZN(n9709) );
  INV_X1 U10876 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9708) );
  AOI22_X1 U10877 ( .A1(n9929), .A2(n9709), .B1(n9708), .B2(n9927), .ZN(
        P1_U3484) );
  AOI22_X1 U10878 ( .A1(n9935), .A2(n9709), .B1(n6621), .B2(n9933), .ZN(
        P1_U3533) );
  OAI21_X1 U10879 ( .B1(n9711), .B2(n9911), .A(n9710), .ZN(n9712) );
  AOI21_X1 U10880 ( .B1(n9714), .B2(n9713), .A(n9712), .ZN(n9730) );
  INV_X1 U10881 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9715) );
  AOI22_X1 U10882 ( .A1(n9935), .A2(n9730), .B1(n9715), .B2(n9933), .ZN(
        P1_U3553) );
  OAI211_X1 U10883 ( .C1(n9718), .C2(n9911), .A(n9717), .B(n9716), .ZN(n9719)
         );
  AOI21_X1 U10884 ( .B1(n9720), .B2(n9926), .A(n9719), .ZN(n9732) );
  AOI22_X1 U10885 ( .A1(n9935), .A2(n9732), .B1(n9721), .B2(n9933), .ZN(
        P1_U3537) );
  OAI21_X1 U10886 ( .B1(n9723), .B2(n9911), .A(n9722), .ZN(n9724) );
  AOI21_X1 U10887 ( .B1(n9725), .B2(n9917), .A(n9724), .ZN(n9726) );
  AND2_X1 U10888 ( .A1(n9727), .A2(n9726), .ZN(n9734) );
  AOI22_X1 U10889 ( .A1(n9935), .A2(n9734), .B1(n9728), .B2(n9933), .ZN(
        P1_U3535) );
  INV_X1 U10890 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9729) );
  AOI22_X1 U10891 ( .A1(n9929), .A2(n9730), .B1(n9729), .B2(n9927), .ZN(
        P1_U3521) );
  INV_X1 U10892 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9731) );
  AOI22_X1 U10893 ( .A1(n9929), .A2(n9732), .B1(n9731), .B2(n9927), .ZN(
        P1_U3496) );
  INV_X1 U10894 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9733) );
  AOI22_X1 U10895 ( .A1(n9929), .A2(n9734), .B1(n9733), .B2(n9927), .ZN(
        P1_U3490) );
  XNOR2_X1 U10896 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  INV_X1 U10897 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10125) );
  NAND3_X1 U10898 ( .A1(n9847), .A2(P1_IR_REG_0__SCAN_IN), .A3(n9737), .ZN(
        n9745) );
  INV_X1 U10899 ( .A(n9735), .ZN(n9742) );
  OAI21_X1 U10900 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(n9737), .A(n9736), .ZN(
        n9738) );
  AOI21_X1 U10901 ( .B1(n9740), .B2(n9739), .A(n9738), .ZN(n9741) );
  OAI21_X1 U10902 ( .B1(n9742), .B2(n9741), .A(P1_STATE_REG_SCAN_IN), .ZN(
        n9743) );
  OAI211_X1 U10903 ( .C1(P1_STATE_REG_SCAN_IN), .C2(P1_REG3_REG_0__SCAN_IN), 
        .A(P1_U3083), .B(n9743), .ZN(n9744) );
  OAI211_X1 U10904 ( .C1(n10125), .C2(n9870), .A(n9745), .B(n9744), .ZN(
        P1_U3241) );
  OAI21_X1 U10905 ( .B1(n9748), .B2(n9747), .A(n9746), .ZN(n9749) );
  AOI22_X1 U10906 ( .A1(n9750), .A2(n9859), .B1(n9857), .B2(n9749), .ZN(n9759)
         );
  AOI21_X1 U10907 ( .B1(n9753), .B2(n9752), .A(n9751), .ZN(n9754) );
  NOR2_X1 U10908 ( .A1(n9867), .A2(n9754), .ZN(n9755) );
  AOI211_X1 U10909 ( .C1(P1_ADDR_REG_4__SCAN_IN), .C2(n9773), .A(n9756), .B(
        n9755), .ZN(n9758) );
  NAND3_X1 U10910 ( .A1(n9759), .A2(n9758), .A3(n9757), .ZN(P1_U3245) );
  AOI22_X1 U10911 ( .A1(n9773), .A2(P1_ADDR_REG_5__SCAN_IN), .B1(n9859), .B2(
        n9760), .ZN(n9771) );
  OAI21_X1 U10912 ( .B1(n9763), .B2(n9762), .A(n9761), .ZN(n9764) );
  NAND2_X1 U10913 ( .A1(n9857), .A2(n9764), .ZN(n9769) );
  OAI211_X1 U10914 ( .C1(n9767), .C2(n9766), .A(n9847), .B(n9765), .ZN(n9768)
         );
  NAND4_X1 U10915 ( .A1(n9771), .A2(n9770), .A3(n9769), .A4(n9768), .ZN(
        P1_U3246) );
  AOI22_X1 U10916 ( .A1(n9773), .A2(P1_ADDR_REG_8__SCAN_IN), .B1(n9859), .B2(
        n9772), .ZN(n9784) );
  INV_X1 U10917 ( .A(n9774), .ZN(n9783) );
  XNOR2_X1 U10918 ( .A(n9776), .B(n9775), .ZN(n9777) );
  NAND2_X1 U10919 ( .A1(n9857), .A2(n9777), .ZN(n9782) );
  OAI211_X1 U10920 ( .C1(n9780), .C2(n9779), .A(n9778), .B(n9847), .ZN(n9781)
         );
  NAND4_X1 U10921 ( .A1(n9784), .A2(n9783), .A3(n9782), .A4(n9781), .ZN(
        P1_U3249) );
  INV_X1 U10922 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9799) );
  AOI21_X1 U10923 ( .B1(n9859), .B2(n9786), .A(n9785), .ZN(n9792) );
  AOI21_X1 U10924 ( .B1(n9789), .B2(n9788), .A(n9787), .ZN(n9790) );
  NAND2_X1 U10925 ( .A1(n9857), .A2(n9790), .ZN(n9791) );
  AND2_X1 U10926 ( .A1(n9792), .A2(n9791), .ZN(n9798) );
  AOI21_X1 U10927 ( .B1(n9795), .B2(n9794), .A(n9793), .ZN(n9796) );
  OR2_X1 U10928 ( .A1(n9867), .A2(n9796), .ZN(n9797) );
  OAI211_X1 U10929 ( .C1(n9799), .C2(n9870), .A(n9798), .B(n9797), .ZN(
        P1_U3253) );
  INV_X1 U10930 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9814) );
  AOI21_X1 U10931 ( .B1(n9859), .B2(n9801), .A(n9800), .ZN(n9807) );
  AOI21_X1 U10932 ( .B1(n9804), .B2(n9803), .A(n9802), .ZN(n9805) );
  NAND2_X1 U10933 ( .A1(n9857), .A2(n9805), .ZN(n9806) );
  AND2_X1 U10934 ( .A1(n9807), .A2(n9806), .ZN(n9813) );
  AOI21_X1 U10935 ( .B1(n9810), .B2(n9809), .A(n9808), .ZN(n9811) );
  OR2_X1 U10936 ( .A1(n9867), .A2(n9811), .ZN(n9812) );
  OAI211_X1 U10937 ( .C1(n9814), .C2(n9870), .A(n9813), .B(n9812), .ZN(
        P1_U3254) );
  AOI211_X1 U10938 ( .C1(n9816), .C2(n7599), .A(n9815), .B(n9826), .ZN(n9817)
         );
  AOI211_X1 U10939 ( .C1(n9819), .C2(n9859), .A(n9818), .B(n9817), .ZN(n9823)
         );
  OAI211_X1 U10940 ( .C1(n9821), .C2(P1_REG1_REG_15__SCAN_IN), .A(n9847), .B(
        n9820), .ZN(n9822) );
  OAI211_X1 U10941 ( .C1(n9824), .C2(n9870), .A(n9823), .B(n9822), .ZN(
        P1_U3256) );
  INV_X1 U10942 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9837) );
  INV_X1 U10943 ( .A(n9825), .ZN(n9830) );
  AOI211_X1 U10944 ( .C1(n4344), .C2(n9828), .A(n9827), .B(n9826), .ZN(n9829)
         );
  AOI211_X1 U10945 ( .C1(n9831), .C2(n9859), .A(n9830), .B(n9829), .ZN(n9836)
         );
  OAI211_X1 U10946 ( .C1(n9834), .C2(n9833), .A(n9847), .B(n9832), .ZN(n9835)
         );
  OAI211_X1 U10947 ( .C1(n9837), .C2(n9870), .A(n9836), .B(n9835), .ZN(
        P1_U3257) );
  INV_X1 U10948 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9852) );
  AOI21_X1 U10949 ( .B1(n9840), .B2(n9839), .A(n9838), .ZN(n9841) );
  NAND2_X1 U10950 ( .A1(n9857), .A2(n9841), .ZN(n9845) );
  NAND2_X1 U10951 ( .A1(n9859), .A2(n9842), .ZN(n9844) );
  AND3_X1 U10952 ( .A1(n9845), .A2(n9844), .A3(n9843), .ZN(n9851) );
  OAI211_X1 U10953 ( .C1(n9849), .C2(n9848), .A(n9847), .B(n9846), .ZN(n9850)
         );
  OAI211_X1 U10954 ( .C1(n9852), .C2(n9870), .A(n9851), .B(n9850), .ZN(
        P1_U3258) );
  INV_X1 U10955 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9871) );
  AOI21_X1 U10956 ( .B1(n9855), .B2(n9854), .A(n9853), .ZN(n9856) );
  NAND2_X1 U10957 ( .A1(n9857), .A2(n9856), .ZN(n9862) );
  NAND2_X1 U10958 ( .A1(n9859), .A2(n9858), .ZN(n9861) );
  AND3_X1 U10959 ( .A1(n9862), .A2(n9861), .A3(n9860), .ZN(n9869) );
  AOI21_X1 U10960 ( .B1(n9865), .B2(n9864), .A(n9863), .ZN(n9866) );
  OR2_X1 U10961 ( .A1(n9867), .A2(n9866), .ZN(n9868) );
  OAI211_X1 U10962 ( .C1(n9871), .C2(n9870), .A(n9869), .B(n9868), .ZN(
        P1_U3259) );
  INV_X1 U10963 ( .A(n9872), .ZN(n9882) );
  OAI22_X1 U10964 ( .A1(n9876), .A2(n9875), .B1(n9874), .B2(n9873), .ZN(n9877)
         );
  AOI21_X1 U10965 ( .B1(n9879), .B2(n9878), .A(n9877), .ZN(n9880) );
  OAI211_X1 U10966 ( .C1(n9883), .C2(n9882), .A(n9881), .B(n9880), .ZN(n9884)
         );
  INV_X1 U10967 ( .A(n9884), .ZN(n9886) );
  AOI22_X1 U10968 ( .A1(n9887), .A2(n5055), .B1(n9886), .B2(n9885), .ZN(
        P1_U3286) );
  AND2_X1 U10969 ( .A1(n9895), .A2(n9888), .ZN(n9891) );
  AND2_X1 U10970 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9892), .ZN(P1_U3292) );
  AND2_X1 U10971 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9892), .ZN(P1_U3293) );
  AND2_X1 U10972 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9892), .ZN(P1_U3294) );
  AND2_X1 U10973 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9892), .ZN(P1_U3295) );
  AND2_X1 U10974 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9892), .ZN(P1_U3296) );
  AND2_X1 U10975 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9892), .ZN(P1_U3297) );
  AND2_X1 U10976 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9892), .ZN(P1_U3298) );
  NOR2_X1 U10977 ( .A1(n9891), .A2(n9889), .ZN(P1_U3299) );
  AND2_X1 U10978 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9892), .ZN(P1_U3300) );
  AND2_X1 U10979 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9892), .ZN(P1_U3301) );
  AND2_X1 U10980 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9892), .ZN(P1_U3302) );
  AND2_X1 U10981 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9892), .ZN(P1_U3303) );
  AND2_X1 U10982 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9892), .ZN(P1_U3304) );
  AND2_X1 U10983 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9892), .ZN(P1_U3305) );
  AND2_X1 U10984 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9892), .ZN(P1_U3306) );
  AND2_X1 U10985 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9892), .ZN(P1_U3307) );
  AND2_X1 U10986 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9892), .ZN(P1_U3308) );
  AND2_X1 U10987 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9892), .ZN(P1_U3309) );
  AND2_X1 U10988 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9892), .ZN(P1_U3310) );
  NOR2_X1 U10989 ( .A1(n9891), .A2(n9890), .ZN(P1_U3311) );
  AND2_X1 U10990 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9892), .ZN(P1_U3312) );
  AND2_X1 U10991 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9892), .ZN(P1_U3313) );
  AND2_X1 U10992 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9892), .ZN(P1_U3314) );
  AND2_X1 U10993 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9892), .ZN(P1_U3315) );
  AND2_X1 U10994 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9892), .ZN(P1_U3316) );
  AND2_X1 U10995 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9892), .ZN(P1_U3317) );
  AND2_X1 U10996 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9892), .ZN(P1_U3318) );
  AND2_X1 U10997 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9892), .ZN(P1_U3319) );
  AND2_X1 U10998 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9892), .ZN(P1_U3320) );
  AND2_X1 U10999 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9892), .ZN(P1_U3321) );
  INV_X1 U11000 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9894) );
  OAI21_X1 U11001 ( .B1(n9895), .B2(n9894), .A(n9893), .ZN(P1_U3441) );
  INV_X1 U11002 ( .A(n9896), .ZN(n9898) );
  NAND2_X1 U11003 ( .A1(n9898), .A2(n9897), .ZN(n9900) );
  AOI211_X1 U11004 ( .C1(n9901), .C2(n9926), .A(n9900), .B(n9899), .ZN(n9930)
         );
  INV_X1 U11005 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9902) );
  AOI22_X1 U11006 ( .A1(n9929), .A2(n9930), .B1(n9902), .B2(n9927), .ZN(
        P1_U3457) );
  INV_X1 U11007 ( .A(n9903), .ZN(n9904) );
  OAI21_X1 U11008 ( .B1(n9921), .B2(n9905), .A(n9904), .ZN(n9908) );
  INV_X1 U11009 ( .A(n9906), .ZN(n9907) );
  AOI211_X1 U11010 ( .C1(n9926), .C2(n9909), .A(n9908), .B(n9907), .ZN(n9931)
         );
  INV_X1 U11011 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9910) );
  AOI22_X1 U11012 ( .A1(n9929), .A2(n9931), .B1(n9910), .B2(n9927), .ZN(
        P1_U3460) );
  OAI22_X1 U11013 ( .A1(n9913), .A2(n9921), .B1(n9912), .B2(n9911), .ZN(n9915)
         );
  AOI211_X1 U11014 ( .C1(n9917), .C2(n9916), .A(n9915), .B(n9914), .ZN(n9932)
         );
  INV_X1 U11015 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9918) );
  AOI22_X1 U11016 ( .A1(n9929), .A2(n9932), .B1(n9918), .B2(n9927), .ZN(
        P1_U3466) );
  INV_X1 U11017 ( .A(n9919), .ZN(n9920) );
  OAI21_X1 U11018 ( .B1(n9922), .B2(n9921), .A(n9920), .ZN(n9924) );
  AOI211_X1 U11019 ( .C1(n9926), .C2(n9925), .A(n9924), .B(n9923), .ZN(n9934)
         );
  INV_X1 U11020 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9928) );
  AOI22_X1 U11021 ( .A1(n9929), .A2(n9934), .B1(n9928), .B2(n9927), .ZN(
        P1_U3472) );
  AOI22_X1 U11022 ( .A1(n9935), .A2(n9930), .B1(n6173), .B2(n9933), .ZN(
        P1_U3524) );
  AOI22_X1 U11023 ( .A1(n9935), .A2(n9931), .B1(n6176), .B2(n9933), .ZN(
        P1_U3525) );
  AOI22_X1 U11024 ( .A1(n9935), .A2(n9932), .B1(n6180), .B2(n9933), .ZN(
        P1_U3527) );
  AOI22_X1 U11025 ( .A1(n9935), .A2(n9934), .B1(n5081), .B2(n9933), .ZN(
        P1_U3529) );
  AOI22_X1 U11026 ( .A1(n9937), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9936), .ZN(n9947) );
  NAND2_X1 U11027 ( .A1(n9938), .A2(n10008), .ZN(n9940) );
  OAI211_X1 U11028 ( .C1(n9941), .C2(P2_REG1_REG_0__SCAN_IN), .A(n9940), .B(
        n9939), .ZN(n9942) );
  INV_X1 U11029 ( .A(n9942), .ZN(n9945) );
  AOI22_X1 U11030 ( .A1(n9943), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(n4262), .ZN(n9944) );
  OAI221_X1 U11031 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9947), .C1(n9946), .C2(
        n9945), .A(n9944), .ZN(P2_U3245) );
  XNOR2_X1 U11032 ( .A(n9948), .B(n9954), .ZN(n9958) );
  NAND2_X1 U11033 ( .A1(n9950), .A2(n9949), .ZN(n9953) );
  AOI21_X1 U11034 ( .B1(n9954), .B2(n9953), .A(n4349), .ZN(n10074) );
  NOR2_X1 U11035 ( .A1(n10074), .A2(n9955), .ZN(n9956) );
  AOI211_X1 U11036 ( .C1(n9958), .C2(n9968), .A(n9957), .B(n9956), .ZN(n10072)
         );
  AOI222_X1 U11037 ( .A1(n10070), .A2(n9990), .B1(P2_REG2_REG_9__SCAN_IN), 
        .B2(n10011), .C1(n10001), .C2(n9959), .ZN(n9964) );
  INV_X1 U11038 ( .A(n10074), .ZN(n9962) );
  AOI211_X1 U11039 ( .C1(n10070), .C2(n9960), .A(n10086), .B(n4353), .ZN(
        n10068) );
  AOI22_X1 U11040 ( .A1(n9962), .A2(n9961), .B1(n9993), .B2(n10068), .ZN(n9963) );
  OAI211_X1 U11041 ( .C1(n10011), .C2(n10072), .A(n9964), .B(n9963), .ZN(
        P2_U3287) );
  NAND2_X1 U11042 ( .A1(n9966), .A2(n9965), .ZN(n9967) );
  NAND2_X1 U11043 ( .A1(n9967), .A2(n9977), .ZN(n9970) );
  NAND3_X1 U11044 ( .A1(n9970), .A2(n9969), .A3(n9968), .ZN(n9973) );
  INV_X1 U11045 ( .A(n9971), .ZN(n9972) );
  AND2_X1 U11046 ( .A1(n9973), .A2(n9972), .ZN(n10056) );
  AOI222_X1 U11047 ( .A1(n9975), .A2(n9990), .B1(P2_REG2_REG_7__SCAN_IN), .B2(
        n10011), .C1(n10001), .C2(n9974), .ZN(n9982) );
  OAI21_X1 U11048 ( .B1(n7161), .B2(n9977), .A(n9976), .ZN(n10059) );
  OAI211_X1 U11049 ( .C1(n9979), .C2(n10057), .A(n10049), .B(n9978), .ZN(
        n10055) );
  INV_X1 U11050 ( .A(n10055), .ZN(n9980) );
  AOI22_X1 U11051 ( .A1(n10059), .A2(n10006), .B1(n9993), .B2(n9980), .ZN(
        n9981) );
  OAI211_X1 U11052 ( .C1(n10011), .C2(n10056), .A(n9982), .B(n9981), .ZN(
        P2_U3289) );
  AOI22_X1 U11053 ( .A1(n9983), .A2(n10001), .B1(P2_REG2_REG_4__SCAN_IN), .B2(
        n10011), .ZN(n9988) );
  AOI222_X1 U11054 ( .A1(n9986), .A2(n10006), .B1(n9993), .B2(n9985), .C1(
        n9984), .C2(n9990), .ZN(n9987) );
  OAI211_X1 U11055 ( .C1(n10011), .C2(n9989), .A(n9988), .B(n9987), .ZN(
        P2_U3292) );
  AOI22_X1 U11056 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(n10001), .B1(
        P2_REG2_REG_2__SCAN_IN), .B2(n10011), .ZN(n9996) );
  AOI222_X1 U11057 ( .A1(n9994), .A2(n10006), .B1(n9993), .B2(n9992), .C1(
        n9991), .C2(n9990), .ZN(n9995) );
  OAI211_X1 U11058 ( .C1(n10011), .C2(n9997), .A(n9996), .B(n9995), .ZN(
        P2_U3294) );
  INV_X1 U11059 ( .A(n9998), .ZN(n9999) );
  OAI21_X1 U11060 ( .B1(n10002), .B2(n10000), .A(n9999), .ZN(n10029) );
  AOI21_X1 U11061 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n10001), .A(n10029), .ZN(
        n10010) );
  INV_X1 U11062 ( .A(n10002), .ZN(n10031) );
  AOI21_X1 U11063 ( .B1(n10004), .B2(n10003), .A(n10028), .ZN(n10005) );
  AOI21_X1 U11064 ( .B1(n10006), .B2(n10031), .A(n10005), .ZN(n10007) );
  OAI221_X1 U11065 ( .B1(n10011), .B2(n10010), .C1(n10009), .C2(n10008), .A(
        n10007), .ZN(P2_U3296) );
  INV_X1 U11066 ( .A(n10012), .ZN(n10014) );
  NAND2_X1 U11067 ( .A1(n10014), .A2(n10013), .ZN(n10023) );
  AND2_X1 U11068 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10023), .ZN(P2_U3297) );
  AND2_X1 U11069 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10023), .ZN(P2_U3298) );
  AND2_X1 U11070 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10023), .ZN(P2_U3299) );
  AND2_X1 U11071 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10023), .ZN(P2_U3300) );
  INV_X1 U11072 ( .A(n10023), .ZN(n10020) );
  NOR2_X1 U11073 ( .A1(n10020), .A2(n10015), .ZN(P2_U3301) );
  NOR2_X1 U11074 ( .A1(n10020), .A2(n10016), .ZN(P2_U3302) );
  AND2_X1 U11075 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10023), .ZN(P2_U3303) );
  NOR2_X1 U11076 ( .A1(n10020), .A2(n10017), .ZN(P2_U3304) );
  AND2_X1 U11077 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10023), .ZN(P2_U3305) );
  AND2_X1 U11078 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10023), .ZN(P2_U3306) );
  AND2_X1 U11079 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10023), .ZN(P2_U3307) );
  AND2_X1 U11080 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10023), .ZN(P2_U3308) );
  AND2_X1 U11081 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10023), .ZN(P2_U3309) );
  AND2_X1 U11082 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10023), .ZN(P2_U3310) );
  AND2_X1 U11083 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10023), .ZN(P2_U3311) );
  AND2_X1 U11084 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10023), .ZN(P2_U3312) );
  AND2_X1 U11085 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10023), .ZN(P2_U3313) );
  AND2_X1 U11086 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10023), .ZN(P2_U3314) );
  AND2_X1 U11087 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10023), .ZN(P2_U3315) );
  AND2_X1 U11088 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10023), .ZN(P2_U3316) );
  AND2_X1 U11089 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10023), .ZN(P2_U3317) );
  AND2_X1 U11090 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10023), .ZN(P2_U3318) );
  AND2_X1 U11091 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10023), .ZN(P2_U3319) );
  NOR2_X1 U11092 ( .A1(n10020), .A2(n10018), .ZN(P2_U3320) );
  AND2_X1 U11093 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10023), .ZN(P2_U3321) );
  AND2_X1 U11094 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10023), .ZN(P2_U3322) );
  AND2_X1 U11095 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10023), .ZN(P2_U3323) );
  AND2_X1 U11096 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10023), .ZN(P2_U3324) );
  AND2_X1 U11097 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10023), .ZN(P2_U3325) );
  AND2_X1 U11098 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10023), .ZN(P2_U3326) );
  OAI22_X1 U11099 ( .A1(P2_D_REG_0__SCAN_IN), .A2(n10020), .B1(n10019), .B2(
        n10022), .ZN(n10021) );
  INV_X1 U11100 ( .A(n10021), .ZN(P2_U3437) );
  INV_X1 U11101 ( .A(n10022), .ZN(n10025) );
  AOI22_X1 U11102 ( .A1(n10026), .A2(n10025), .B1(n10024), .B2(n10023), .ZN(
        P2_U3438) );
  NOR2_X1 U11103 ( .A1(n10028), .A2(n10027), .ZN(n10030) );
  AOI211_X1 U11104 ( .C1(n10031), .C2(n10097), .A(n10030), .B(n10029), .ZN(
        n10103) );
  INV_X1 U11105 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10032) );
  AOI22_X1 U11106 ( .A1(n10101), .A2(n10103), .B1(n10032), .B2(n10099), .ZN(
        P2_U3451) );
  INV_X1 U11107 ( .A(n10069), .ZN(n10094) );
  NAND3_X1 U11108 ( .A1(n10034), .A2(n10033), .A3(n10049), .ZN(n10035) );
  OAI21_X1 U11109 ( .B1(n6052), .B2(n10094), .A(n10035), .ZN(n10038) );
  INV_X1 U11110 ( .A(n10036), .ZN(n10037) );
  AOI211_X1 U11111 ( .C1(n10097), .C2(n10039), .A(n10038), .B(n10037), .ZN(
        n10104) );
  INV_X1 U11112 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10040) );
  AOI22_X1 U11113 ( .A1(n10101), .A2(n10104), .B1(n10040), .B2(n10099), .ZN(
        P2_U3454) );
  OAI211_X1 U11114 ( .C1(n10043), .C2(n10094), .A(n10042), .B(n10041), .ZN(
        n10044) );
  AOI21_X1 U11115 ( .B1(n10097), .B2(n10045), .A(n10044), .ZN(n10105) );
  INV_X1 U11116 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10046) );
  AOI22_X1 U11117 ( .A1(n10101), .A2(n10105), .B1(n10046), .B2(n10099), .ZN(
        P2_U3466) );
  NAND3_X1 U11118 ( .A1(n8598), .A2(n10047), .A3(n10097), .ZN(n10053) );
  AOI22_X1 U11119 ( .A1(n10050), .A2(n10049), .B1(n10048), .B2(n10069), .ZN(
        n10051) );
  AND3_X1 U11120 ( .A1(n10053), .A2(n10052), .A3(n10051), .ZN(n10107) );
  INV_X1 U11121 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10054) );
  AOI22_X1 U11122 ( .A1(n10101), .A2(n10107), .B1(n10054), .B2(n10099), .ZN(
        P2_U3469) );
  OAI211_X1 U11123 ( .C1(n10057), .C2(n10094), .A(n10056), .B(n10055), .ZN(
        n10058) );
  AOI21_X1 U11124 ( .B1(n10059), .B2(n10097), .A(n10058), .ZN(n10109) );
  INV_X1 U11125 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10060) );
  AOI22_X1 U11126 ( .A1(n10101), .A2(n10109), .B1(n10060), .B2(n10099), .ZN(
        P2_U3472) );
  INV_X1 U11127 ( .A(n10061), .ZN(n10066) );
  OAI22_X1 U11128 ( .A1(n10063), .A2(n10086), .B1(n10062), .B2(n10094), .ZN(
        n10065) );
  AOI211_X1 U11129 ( .C1(n10082), .C2(n10066), .A(n10065), .B(n10064), .ZN(
        n10111) );
  INV_X1 U11130 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10067) );
  AOI22_X1 U11131 ( .A1(n10101), .A2(n10111), .B1(n10067), .B2(n10099), .ZN(
        P2_U3475) );
  AOI21_X1 U11132 ( .B1(n10070), .B2(n10069), .A(n10068), .ZN(n10071) );
  OAI211_X1 U11133 ( .C1(n10074), .C2(n10073), .A(n10072), .B(n10071), .ZN(
        n10075) );
  INV_X1 U11134 ( .A(n10075), .ZN(n10113) );
  INV_X1 U11135 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10076) );
  AOI22_X1 U11136 ( .A1(n10101), .A2(n10113), .B1(n10076), .B2(n10099), .ZN(
        P2_U3478) );
  OAI21_X1 U11137 ( .B1(n10078), .B2(n10094), .A(n10077), .ZN(n10080) );
  AOI211_X1 U11138 ( .C1(n10082), .C2(n10081), .A(n10080), .B(n10079), .ZN(
        n10114) );
  INV_X1 U11139 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10083) );
  AOI22_X1 U11140 ( .A1(n10101), .A2(n10114), .B1(n10083), .B2(n10099), .ZN(
        P2_U3481) );
  INV_X1 U11141 ( .A(n10084), .ZN(n10090) );
  OAI22_X1 U11142 ( .A1(n10087), .A2(n10086), .B1(n10085), .B2(n10094), .ZN(
        n10088) );
  AOI211_X1 U11143 ( .C1(n10090), .C2(n10097), .A(n10089), .B(n10088), .ZN(
        n10116) );
  INV_X1 U11144 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10091) );
  AOI22_X1 U11145 ( .A1(n10101), .A2(n10116), .B1(n10091), .B2(n10099), .ZN(
        P2_U3484) );
  OAI211_X1 U11146 ( .C1(n10095), .C2(n10094), .A(n10093), .B(n10092), .ZN(
        n10096) );
  AOI21_X1 U11147 ( .B1(n10098), .B2(n10097), .A(n10096), .ZN(n10119) );
  INV_X1 U11148 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10100) );
  AOI22_X1 U11149 ( .A1(n10101), .A2(n10119), .B1(n10100), .B2(n10099), .ZN(
        P2_U3487) );
  AOI22_X1 U11150 ( .A1(n10120), .A2(n10103), .B1(n10102), .B2(n10117), .ZN(
        P2_U3520) );
  AOI22_X1 U11151 ( .A1(n10120), .A2(n10104), .B1(n6435), .B2(n10117), .ZN(
        P2_U3521) );
  AOI22_X1 U11152 ( .A1(n10120), .A2(n10105), .B1(n5634), .B2(n10117), .ZN(
        P2_U3525) );
  AOI22_X1 U11153 ( .A1(n10120), .A2(n10107), .B1(n10106), .B2(n10117), .ZN(
        P2_U3526) );
  AOI22_X1 U11154 ( .A1(n10120), .A2(n10109), .B1(n10108), .B2(n10117), .ZN(
        P2_U3527) );
  AOI22_X1 U11155 ( .A1(n10120), .A2(n10111), .B1(n10110), .B2(n10117), .ZN(
        P2_U3528) );
  AOI22_X1 U11156 ( .A1(n10120), .A2(n10113), .B1(n10112), .B2(n10117), .ZN(
        P2_U3529) );
  AOI22_X1 U11157 ( .A1(n10120), .A2(n10114), .B1(n6919), .B2(n10117), .ZN(
        P2_U3530) );
  AOI22_X1 U11158 ( .A1(n10120), .A2(n10116), .B1(n10115), .B2(n10117), .ZN(
        P2_U3531) );
  AOI22_X1 U11159 ( .A1(n10120), .A2(n10119), .B1(n10118), .B2(n10117), .ZN(
        P2_U3532) );
  INV_X1 U11160 ( .A(n10121), .ZN(n10122) );
  NAND2_X1 U11161 ( .A1(n10123), .A2(n10122), .ZN(n10124) );
  XNOR2_X1 U11162 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10124), .ZN(ADD_1071_U5)
         );
  INV_X1 U11163 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10126) );
  AOI22_X1 U11164 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .B1(n10126), .B2(n10125), .ZN(ADD_1071_U46) );
  OAI21_X1 U11165 ( .B1(n10129), .B2(n10128), .A(n10127), .ZN(ADD_1071_U56) );
  OAI21_X1 U11166 ( .B1(n10132), .B2(n10131), .A(n10130), .ZN(ADD_1071_U57) );
  OAI21_X1 U11167 ( .B1(n10135), .B2(n10134), .A(n10133), .ZN(ADD_1071_U58) );
  OAI21_X1 U11168 ( .B1(n10138), .B2(n10137), .A(n10136), .ZN(ADD_1071_U59) );
  OAI21_X1 U11169 ( .B1(n10141), .B2(n10140), .A(n10139), .ZN(ADD_1071_U60) );
  OAI21_X1 U11170 ( .B1(n10144), .B2(n10143), .A(n10142), .ZN(ADD_1071_U61) );
  AOI21_X1 U11171 ( .B1(n10147), .B2(n10146), .A(n10145), .ZN(ADD_1071_U62) );
  AOI21_X1 U11172 ( .B1(n10150), .B2(n10149), .A(n10148), .ZN(ADD_1071_U63) );
  XOR2_X1 U11173 ( .A(n10151), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11174 ( .A1(n10153), .A2(n10152), .ZN(n10154) );
  XOR2_X1 U11175 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10154), .Z(ADD_1071_U51) );
  XOR2_X1 U11176 ( .A(n10155), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1071_U48) );
  OAI21_X1 U11177 ( .B1(n10158), .B2(n10157), .A(n10156), .ZN(n10159) );
  XNOR2_X1 U11178 ( .A(n10159), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XOR2_X1 U11179 ( .A(n10160), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  AOI21_X1 U11180 ( .B1(n10163), .B2(n10162), .A(n10161), .ZN(ADD_1071_U47) );
  XOR2_X1 U11181 ( .A(n10165), .B(n10164), .Z(ADD_1071_U54) );
  XOR2_X1 U11182 ( .A(n10167), .B(n10166), .Z(ADD_1071_U53) );
  XNOR2_X1 U11183 ( .A(n10169), .B(n10168), .ZN(ADD_1071_U52) );
  OR2_X1 U4772 ( .A1(n6932), .A2(n5470), .ZN(n5471) );
  NAND2_X1 U4786 ( .A1(n5471), .A2(n9196), .ZN(n7152) );
  CLKBUF_X1 U4813 ( .A(n7259), .Z(n8098) );
  CLKBUF_X3 U4863 ( .A(n5062), .Z(n8115) );
  CLKBUF_X2 U6104 ( .A(n5050), .Z(n6244) );
  CLKBUF_X1 U6921 ( .A(n5649), .Z(n6038) );
endmodule

