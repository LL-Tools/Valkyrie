

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput127, keyinput126, keyinput125, keyinput124, keyinput123, 
        keyinput122, keyinput121, keyinput120, keyinput119, keyinput118, 
        keyinput117, keyinput116, keyinput115, keyinput114, keyinput113, 
        keyinput112, keyinput111, keyinput110, keyinput109, keyinput108, 
        keyinput107, keyinput106, keyinput105, keyinput104, keyinput103, 
        keyinput102, keyinput101, keyinput100, keyinput99, keyinput98, 
        keyinput97, keyinput96, keyinput95, keyinput94, keyinput93, keyinput92, 
        keyinput91, keyinput90, keyinput89, keyinput88, keyinput87, keyinput86, 
        keyinput85, keyinput84, keyinput83, keyinput82, keyinput81, keyinput80, 
        keyinput79, keyinput78, keyinput77, keyinput76, keyinput75, keyinput74, 
        keyinput73, keyinput72, keyinput71, keyinput70, keyinput69, keyinput68, 
        keyinput67, keyinput66, keyinput65, keyinput64, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4421, n4422, n4423, n4424, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303;

  XNOR2_X1 U4927 ( .A(n6541), .B(n7237), .ZN(n7242) );
  INV_X1 U4929 ( .A(n5979), .ZN(n9176) );
  CLKBUF_X1 U4930 ( .A(n5931), .Z(n6480) );
  CLKBUF_X2 U4931 ( .A(n5176), .Z(n5177) );
  AND2_X1 U4932 ( .A1(n4588), .A2(n5914), .ZN(n7439) );
  NAND2_X2 U4933 ( .A1(n8222), .A2(n5101), .ZN(n4529) );
  NAND2_X1 U4934 ( .A1(n5031), .A2(n5030), .ZN(n5333) );
  OAI22_X1 U4935 ( .A1(n6566), .A2(n5147), .B1(P2_IR_REG_2__SCAN_IN), .B2(
        P2_IR_REG_31__SCAN_IN), .ZN(n5149) );
  NOR2_X1 U4936 ( .A1(n8284), .A2(n8283), .ZN(n8296) );
  OR2_X1 U4937 ( .A1(n8674), .A2(n4778), .ZN(n4777) );
  OAI22_X1 U4938 ( .A1(n4859), .A2(n10133), .B1(n7242), .B2(n4858), .ZN(n10132) );
  AND2_X2 U4939 ( .A1(n5102), .A2(n8222), .ZN(n5155) );
  INV_X1 U4940 ( .A(n5135), .ZN(n5756) );
  XNOR2_X1 U4941 ( .A(n6215), .B(n6213), .ZN(n9028) );
  NAND2_X1 U4944 ( .A1(n4936), .A2(n4934), .ZN(n7641) );
  CLKBUF_X3 U4945 ( .A(n5122), .Z(n8392) );
  NOR2_X1 U4946 ( .A1(n8178), .A2(n9841), .ZN(n8177) );
  AND2_X1 U4947 ( .A1(n4867), .A2(n4481), .ZN(n8725) );
  AND2_X2 U4948 ( .A1(n5168), .A2(n5192), .ZN(n6708) );
  AND2_X1 U4949 ( .A1(n9608), .A2(n8520), .ZN(n9758) );
  NAND2_X1 U4950 ( .A1(n6217), .A2(n6219), .ZN(n6221) );
  XNOR2_X1 U4951 ( .A(n5187), .B(SI_3_), .ZN(n5209) );
  XNOR2_X1 U4952 ( .A(n5098), .B(n5097), .ZN(n5102) );
  OR2_X2 U4953 ( .A1(n9620), .A2(n9621), .ZN(n4961) );
  INV_X4 U4954 ( .A(n8774), .ZN(n4713) );
  INV_X2 U4955 ( .A(n8468), .ZN(n5925) );
  INV_X2 U4956 ( .A(n6742), .ZN(n9280) );
  OAI21_X2 U4957 ( .B1(n6221), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6269) );
  INV_X4 U4958 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5154) );
  AOI21_X2 U4959 ( .B1(n7154), .B2(n7155), .A(n7156), .ZN(n7153) );
  OR3_X4 U4960 ( .A1(n5333), .A2(P2_REG3_REG_10__SCAN_IN), .A3(
        P2_REG3_REG_11__SCAN_IN), .ZN(n5348) );
  OAI21_X2 U4961 ( .B1(n5505), .B2(n5504), .A(n5503), .ZN(n5518) );
  NAND2_X4 U4962 ( .A1(n7854), .A2(n9584), .ZN(n9285) );
  XNOR2_X2 U4963 ( .A(n6600), .B(n6599), .ZN(n8674) );
  NAND2_X1 U4964 ( .A1(n5134), .A2(n4587), .ZN(n4421) );
  NAND2_X1 U4965 ( .A1(n5134), .A2(n4587), .ZN(n4422) );
  NAND2_X1 U4966 ( .A1(n5906), .A2(n7112), .ZN(n4423) );
  INV_X2 U4967 ( .A(n6439), .ZN(n6418) );
  OAI21_X2 U4968 ( .B1(n5343), .B2(n5342), .A(n5341), .ZN(n5367) );
  OAI21_X4 U4969 ( .B1(n5322), .B2(n5321), .A(n5320), .ZN(n5343) );
  NOR2_X2 U4970 ( .A1(n8047), .A2(n8046), .ZN(n8088) );
  AOI21_X2 U4971 ( .B1(n7602), .B2(n9299), .A(n5016), .ZN(n9929) );
  NAND2_X2 U4972 ( .A1(n7472), .A2(n7471), .ZN(n7602) );
  AND2_X2 U4973 ( .A1(n6284), .A2(n9321), .ZN(n9415) );
  NAND2_X2 U4974 ( .A1(n6467), .A2(n6284), .ZN(n7112) );
  OAI211_X2 U4975 ( .C1(n5296), .C2(n5913), .A(n4897), .B(n4896), .ZN(n5136)
         );
  NOR2_X4 U4976 ( .A1(n5149), .A2(n5165), .ZN(n6632) );
  AND2_X2 U4977 ( .A1(n6566), .A2(n5148), .ZN(n5165) );
  BUF_X4 U4978 ( .A(n6441), .Z(n4424) );
  INV_X1 U4979 ( .A(n6393), .ZN(n6441) );
  AOI21_X2 U4980 ( .B1(n7641), .B2(n7643), .A(n7640), .ZN(n9911) );
  CLKBUF_X1 U4982 ( .A(n7028), .Z(n4426) );
  AOI21_X2 U4983 ( .B1(n6534), .B2(n6708), .A(n6535), .ZN(n7252) );
  NAND2_X2 U4984 ( .A1(n9361), .A2(n9321), .ZN(n7477) );
  XNOR2_X2 U4985 ( .A(n5885), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9361) );
  OAI211_X2 U4986 ( .C1(n4850), .C2(n6533), .A(n4847), .B(n4846), .ZN(n4848)
         );
  OR2_X1 U4987 ( .A1(n8711), .A2(n8933), .ZN(n4867) );
  NOR2_X1 U4988 ( .A1(n8691), .A2(n4868), .ZN(n6559) );
  OAI21_X1 U4989 ( .B1(n8505), .B2(n4951), .A(n4490), .ZN(n4949) );
  NAND2_X1 U4990 ( .A1(n5607), .A2(n5606), .ZN(n5676) );
  NAND2_X1 U4991 ( .A1(n5586), .A2(n5585), .ZN(n5605) );
  INV_X4 U4992 ( .A(n5834), .ZN(n5828) );
  INV_X2 U4993 ( .A(n5762), .ZN(n5834) );
  INV_X1 U4994 ( .A(n9285), .ZN(n9287) );
  INV_X1 U4995 ( .A(n7617), .ZN(n10021) );
  NAND2_X1 U4996 ( .A1(n7114), .A2(n7550), .ZN(n9974) );
  INV_X4 U4997 ( .A(n8399), .ZN(n8383) );
  AND3_X1 U4998 ( .A1(n5984), .A2(n5983), .A3(n5982), .ZN(n10015) );
  BUF_X2 U4999 ( .A(n5986), .Z(n9284) );
  INV_X1 U5000 ( .A(n5986), .ZN(n5931) );
  MUX2_X1 U5001 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5112), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5114) );
  AND3_X1 U5002 ( .A1(n5895), .A2(n4439), .A3(n4502), .ZN(n5922) );
  OR2_X1 U5003 ( .A1(n5233), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5235) );
  CLKBUF_X2 U5004 ( .A(n5105), .Z(n6566) );
  INV_X1 U5005 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5891) );
  OAI21_X1 U5006 ( .B1(n9291), .B2(n9748), .A(n4569), .ZN(n9325) );
  AOI21_X1 U5007 ( .B1(n4553), .B2(n8894), .A(n4556), .ZN(n4844) );
  AOI21_X1 U5008 ( .B1(n4680), .B2(n8399), .A(n4679), .ZN(n4678) );
  MUX2_X1 U5009 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n6698), .S(n10261), .Z(n6694) );
  OAI21_X1 U5010 ( .B1(n9278), .B2(n9601), .A(n9277), .ZN(n9288) );
  NOR2_X1 U5011 ( .A1(n9103), .A2(n6383), .ZN(n9066) );
  AOI21_X1 U5012 ( .B1(n5730), .B2(n8894), .A(n5729), .ZN(n8769) );
  NOR2_X1 U5013 ( .A1(n8743), .A2(n6609), .ZN(n6610) );
  NAND2_X1 U5014 ( .A1(n9179), .A2(n9178), .ZN(n9596) );
  AND2_X1 U5015 ( .A1(n8364), .A2(n8363), .ZN(n4646) );
  AND2_X2 U5016 ( .A1(n6347), .A2(n6346), .ZN(n9125) );
  NOR2_X1 U5017 ( .A1(n8740), .A2(n8739), .ZN(n8743) );
  NAND2_X1 U5018 ( .A1(n4979), .A2(n4977), .ZN(n6347) );
  AOI21_X1 U5019 ( .B1(n4874), .B2(n4875), .A(n4434), .ZN(n4537) );
  OAI21_X1 U5020 ( .B1(n4874), .B2(n4539), .A(n4538), .ZN(n4541) );
  AOI21_X1 U5021 ( .B1(n4431), .B2(n9621), .A(n4478), .ZN(n4960) );
  XNOR2_X1 U5022 ( .A(n8395), .B(n8394), .ZN(n9177) );
  NOR2_X1 U5023 ( .A1(n8718), .A2(n6607), .ZN(n8740) );
  OR2_X1 U5024 ( .A1(n6518), .A2(n8234), .ZN(n8445) );
  AOI21_X1 U5025 ( .B1(n8569), .B2(n4459), .A(n4922), .ZN(n8597) );
  XNOR2_X1 U5026 ( .A(n6559), .B(n6614), .ZN(n8711) );
  NAND2_X1 U5027 ( .A1(n5809), .A2(n5808), .ZN(n8569) );
  NAND2_X1 U5028 ( .A1(n6507), .A2(n6506), .ZN(n6518) );
  INV_X1 U5029 ( .A(n4949), .ZN(n9700) );
  NAND2_X1 U5030 ( .A1(n6268), .A2(n6267), .ZN(n6282) );
  XNOR2_X1 U5031 ( .A(n6501), .B(n6500), .ZN(n8217) );
  NAND2_X1 U5032 ( .A1(n5685), .A2(n5684), .ZN(n8765) );
  NAND2_X1 U5033 ( .A1(n5690), .A2(n5689), .ZN(n6501) );
  AND2_X1 U5034 ( .A1(n4978), .A2(n6336), .ZN(n4977) );
  NAND2_X1 U5035 ( .A1(n6395), .A2(n6394), .ZN(n9771) );
  NAND2_X1 U5036 ( .A1(n5688), .A2(n5687), .ZN(n5690) );
  INV_X1 U5037 ( .A(n9655), .ZN(n9776) );
  NAND2_X1 U5038 ( .A1(n5678), .A2(n5677), .ZN(n5688) );
  NAND2_X1 U5039 ( .A1(n4972), .A2(n4971), .ZN(n6215) );
  XNOR2_X1 U5040 ( .A(n5676), .B(n5675), .ZN(n8082) );
  NAND2_X1 U5041 ( .A1(n6349), .A2(n6348), .ZN(n9785) );
  NAND2_X1 U5042 ( .A1(n6364), .A2(n6363), .ZN(n9780) );
  INV_X1 U5043 ( .A(n9691), .ZN(n9790) );
  NAND2_X1 U5044 ( .A1(n5605), .A2(n5604), .ZN(n5607) );
  NAND2_X1 U5045 ( .A1(n4864), .A2(n4450), .ZN(n4863) );
  INV_X1 U5046 ( .A(n9705), .ZN(n9794) );
  AND2_X1 U5047 ( .A1(n6338), .A2(n6337), .ZN(n9691) );
  AND2_X1 U5048 ( .A1(n6317), .A2(n6316), .ZN(n9705) );
  NAND2_X1 U5049 ( .A1(n6550), .A2(n6549), .ZN(n7998) );
  OAI21_X1 U5050 ( .B1(n5469), .B2(n5468), .A(n5467), .ZN(n5488) );
  NAND2_X1 U5051 ( .A1(n4534), .A2(n4533), .ZN(n4530) );
  OR2_X1 U5052 ( .A1(n10132), .A2(n6543), .ZN(n6544) );
  AND2_X1 U5053 ( .A1(n6067), .A2(n6066), .ZN(n10042) );
  INV_X1 U5054 ( .A(n6430), .ZN(n6391) );
  NAND2_X1 U5055 ( .A1(n7782), .A2(n5785), .ZN(n4536) );
  CLKBUF_X3 U5056 ( .A(n5959), .Z(n6430) );
  NAND2_X1 U5057 ( .A1(n6539), .A2(n6538), .ZN(n7217) );
  NAND2_X1 U5058 ( .A1(n6084), .A2(n6083), .ZN(n10058) );
  NOR2_X1 U5059 ( .A1(n7223), .A2(n7222), .ZN(n7221) );
  AND2_X1 U5060 ( .A1(n6050), .A2(n6049), .ZN(n10035) );
  NAND2_X1 U5061 ( .A1(n5304), .A2(n5303), .ZN(n5322) );
  NAND2_X1 U5062 ( .A1(n5653), .A2(n8251), .ZN(n8408) );
  NAND2_X1 U5063 ( .A1(n6393), .A2(n4423), .ZN(n5959) );
  NAND2_X1 U5064 ( .A1(n6011), .A2(n4946), .ZN(n9451) );
  AND2_X1 U5065 ( .A1(n4775), .A2(n4774), .ZN(n7223) );
  OAI211_X1 U5066 ( .C1(n6753), .C2(n7085), .A(n6027), .B(n6026), .ZN(n9948)
         );
  OAI211_X1 U5067 ( .C1(n8491), .C2(n6753), .A(n6005), .B(n6004), .ZN(n7617)
         );
  INV_X1 U5068 ( .A(n7303), .ZN(n8670) );
  AND4_X1 U5069 ( .A1(n5140), .A2(n5139), .A3(n5141), .A4(n5138), .ZN(n7303)
         );
  INV_X1 U5070 ( .A(n4702), .ZN(n4698) );
  CLKBUF_X1 U5071 ( .A(n6467), .Z(n4429) );
  OR2_X1 U5072 ( .A1(n5943), .A2(n5942), .ZN(n7114) );
  INV_X2 U5073 ( .A(n6006), .ZN(n6482) );
  INV_X2 U5074 ( .A(n4529), .ZN(n5178) );
  OR2_X1 U5075 ( .A1(n5431), .A2(n5430), .ZN(n5433) );
  NAND2_X1 U5076 ( .A1(n5886), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6463) );
  XNOR2_X1 U5077 ( .A(n5073), .B(P2_IR_REG_21__SCAN_IN), .ZN(n5753) );
  OR2_X1 U5078 ( .A1(n5440), .A2(n5439), .ZN(n5443) );
  OR2_X1 U5079 ( .A1(n5411), .A2(n5410), .ZN(n5439) );
  INV_X1 U5080 ( .A(n5930), .ZN(n5929) );
  INV_X1 U5081 ( .A(n5103), .ZN(n8222) );
  NAND2_X4 U5082 ( .A1(n5110), .A2(n8460), .ZN(n5134) );
  AND2_X1 U5083 ( .A1(n5409), .A2(n5006), .ZN(n5410) );
  NAND2_X1 U5084 ( .A1(n5878), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5879) );
  INV_X1 U5085 ( .A(n5362), .ZN(n5366) );
  NOR2_X1 U5086 ( .A1(n4765), .A2(n4768), .ZN(n6571) );
  NAND2_X1 U5087 ( .A1(n4742), .A2(n5916), .ZN(n4741) );
  INV_X1 U5088 ( .A(n5283), .ZN(n5031) );
  NAND2_X1 U5089 ( .A1(n5194), .A2(n5216), .ZN(n7164) );
  XNOR2_X1 U5090 ( .A(n5911), .B(n5920), .ZN(n7028) );
  NAND2_X1 U5091 ( .A1(n4568), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5911) );
  INV_X2 U5092 ( .A(n8392), .ZN(n4587) );
  AND2_X1 U5093 ( .A1(n5900), .A2(n5889), .ZN(n6217) );
  OR2_X1 U5094 ( .A1(n5305), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n5326) );
  INV_X2 U5095 ( .A(n9832), .ZN(n4428) );
  INV_X2 U5096 ( .A(n5122), .ZN(n5186) );
  AND3_X1 U5097 ( .A1(n4564), .A2(n4562), .A3(n4563), .ZN(n5895) );
  AND2_X1 U5098 ( .A1(n5106), .A2(n4763), .ZN(n6564) );
  NAND2_X1 U5099 ( .A1(n5119), .A2(n5118), .ZN(n5122) );
  INV_X1 U5100 ( .A(n5235), .ZN(n4928) );
  AND2_X1 U5101 ( .A1(n4503), .A2(n4930), .ZN(n4929) );
  NAND2_X1 U5102 ( .A1(n5116), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5119) );
  NAND2_X1 U5103 ( .A1(n5915), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5916) );
  NAND4_X1 U5104 ( .A1(n5892), .A2(n6785), .A3(n6219), .A4(n5891), .ZN(n5893)
         );
  OAI21_X1 U5105 ( .B1(P1_RD_REG_SCAN_IN), .B2(P1_ADDR_REG_19__SCAN_IN), .A(
        n5117), .ZN(n5118) );
  INV_X4 U5106 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U5107 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n6121) );
  INV_X1 U5108 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6879) );
  INV_X1 U5109 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n6983) );
  NOR2_X1 U5110 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5874) );
  INV_X1 U5111 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9886) );
  INV_X1 U5112 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6219) );
  INV_X1 U5113 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6887) );
  INV_X1 U5114 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6785) );
  INV_X4 U5115 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U5116 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6937) );
  NOR2_X1 U5117 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5051) );
  NOR2_X1 U5118 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5105) );
  NOR2_X1 U5119 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n5050) );
  INV_X1 U5120 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5276) );
  NAND2_X1 U5121 ( .A1(n4863), .A2(n4861), .ZN(n6555) );
  AND2_X1 U5122 ( .A1(n4862), .A2(n4513), .ZN(n4861) );
  OR2_X2 U5123 ( .A1(n5261), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5283) );
  AOI21_X2 U5124 ( .B1(n7160), .B2(n4848), .A(n7161), .ZN(n7159) );
  NAND2_X2 U5125 ( .A1(n5933), .A2(n5932), .ZN(n7440) );
  NAND2_X1 U5126 ( .A1(n4590), .A2(n4593), .ZN(n4589) );
  OAI21_X1 U5127 ( .B1(n9332), .B2(n9285), .A(n4594), .ZN(n4590) );
  NAND2_X1 U5128 ( .A1(n9337), .A2(n4595), .ZN(n4594) );
  AND2_X1 U5129 ( .A1(n9259), .A2(n9285), .ZN(n4595) );
  NAND2_X1 U5130 ( .A1(n8246), .A2(n5711), .ZN(n8434) );
  OR2_X1 U5131 ( .A1(n8826), .A2(n8835), .ZN(n8341) );
  OAI21_X1 U5132 ( .B1(n5518), .B2(n5517), .A(n5516), .ZN(n5520) );
  NAND2_X2 U5133 ( .A1(n4712), .A2(n4711), .ZN(n8357) );
  NAND2_X1 U5134 ( .A1(n4886), .A2(n4884), .ZN(n8830) );
  AND2_X1 U5135 ( .A1(n4888), .A2(n4885), .ZN(n4884) );
  INV_X1 U5136 ( .A(n8833), .ZN(n4885) );
  OAI21_X1 U5137 ( .B1(n8101), .B2(n4494), .A(n5386), .ZN(n8121) );
  XNOR2_X1 U5138 ( .A(n5100), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5103) );
  NAND2_X1 U5139 ( .A1(n8302), .A2(n8304), .ZN(n4641) );
  OAI211_X1 U5140 ( .C1(n4592), .C2(n4591), .A(n4589), .B(n9260), .ZN(n9263)
         );
  NAND2_X1 U5141 ( .A1(n8765), .A2(n8655), .ZN(n5711) );
  INV_X1 U5142 ( .A(n8960), .ZN(n5603) );
  NOR2_X1 U5143 ( .A1(n4698), .A2(n4696), .ZN(n4695) );
  NOR2_X1 U5144 ( .A1(n4705), .A2(n4700), .ZN(n4699) );
  NAND2_X1 U5145 ( .A1(n5779), .A2(n4905), .ZN(n4904) );
  OR2_X1 U5146 ( .A1(n5786), .A2(n5787), .ZN(n4902) );
  AND2_X1 U5147 ( .A1(n4501), .A2(n5773), .ZN(n4898) );
  AND2_X1 U5148 ( .A1(n7185), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6533) );
  NAND2_X1 U5149 ( .A1(n7217), .A2(n6540), .ZN(n6541) );
  NAND2_X1 U5150 ( .A1(n7216), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6540) );
  INV_X1 U5151 ( .A(n8771), .ZN(n4876) );
  NAND2_X1 U5152 ( .A1(n5603), .A2(n5602), .ZN(n8350) );
  OR2_X1 U5153 ( .A1(n8836), .A2(n8822), .ZN(n8335) );
  OR2_X1 U5154 ( .A1(n8930), .A2(n5806), .ZN(n8329) );
  NAND2_X1 U5155 ( .A1(n4549), .A2(n4928), .ZN(n5094) );
  AND3_X1 U5156 ( .A1(n4551), .A2(n4929), .A3(n4550), .ZN(n4549) );
  NAND2_X1 U5157 ( .A1(n4920), .A2(n5054), .ZN(n4919) );
  INV_X1 U5158 ( .A(n5053), .ZN(n4920) );
  OR2_X1 U5159 ( .A1(n9415), .A2(n5884), .ZN(n5887) );
  NOR2_X1 U5160 ( .A1(n9766), .A2(n4676), .ZN(n4675) );
  INV_X1 U5161 ( .A(n4677), .ZN(n4676) );
  AND2_X1 U5162 ( .A1(n9314), .A2(n4945), .ZN(n4944) );
  NAND2_X1 U5163 ( .A1(n8513), .A2(n8512), .ZN(n4945) );
  OR2_X1 U5164 ( .A1(n4952), .A2(n4458), .ZN(n4950) );
  NAND2_X1 U5165 ( .A1(n4626), .A2(n9392), .ZN(n4623) );
  AND2_X1 U5166 ( .A1(n8164), .A2(n4738), .ZN(n4737) );
  NAND2_X1 U5167 ( .A1(n9308), .A2(n4739), .ZN(n4738) );
  INV_X1 U5168 ( .A(n9225), .ZN(n4739) );
  NAND2_X1 U5169 ( .A1(n8371), .A2(n8370), .ZN(n8389) );
  OR2_X1 U5170 ( .A1(n8367), .A2(SI_29_), .ZN(n8371) );
  NAND2_X1 U5171 ( .A1(n8599), .A2(n5823), .ZN(n5824) );
  OAI21_X1 U5172 ( .B1(n4924), .B2(n4923), .A(n4487), .ZN(n4922) );
  OAI22_X1 U5173 ( .A1(n8587), .A2(n8586), .B1(n5829), .B2(n8783), .ZN(n5832)
         );
  OR2_X1 U5174 ( .A1(n8075), .A2(n8076), .ZN(n5796) );
  AND2_X1 U5175 ( .A1(n4850), .A2(n4849), .ZN(n7189) );
  INV_X1 U5176 ( .A(n7190), .ZN(n4849) );
  XNOR2_X1 U5177 ( .A(n6573), .B(n8483), .ZN(n8477) );
  INV_X1 U5178 ( .A(n6583), .ZN(n6584) );
  OR2_X2 U5179 ( .A1(n8177), .A2(n6556), .ZN(n4852) );
  INV_X1 U5180 ( .A(n6555), .ZN(n6553) );
  NAND2_X1 U5181 ( .A1(n4780), .A2(n4451), .ZN(n4779) );
  INV_X1 U5182 ( .A(n8184), .ZN(n4780) );
  AND4_X1 U5183 ( .A1(n5530), .A2(n5529), .A3(n5528), .A4(n5527), .ZN(n8835)
         );
  NAND2_X1 U5184 ( .A1(n4548), .A2(n4466), .ZN(n4886) );
  INV_X1 U5185 ( .A(n5466), .ZN(n4548) );
  OR2_X1 U5186 ( .A1(n8669), .A2(n7395), .ZN(n5173) );
  AOI21_X1 U5187 ( .B1(n4808), .B2(n4806), .A(n4485), .ZN(n4805) );
  INV_X1 U5188 ( .A(n8357), .ZN(n4806) );
  NAND2_X1 U5189 ( .A1(n5692), .A2(n5691), .ZN(n8378) );
  NAND2_X1 U5190 ( .A1(n8217), .A2(n8396), .ZN(n5692) );
  NAND2_X1 U5191 ( .A1(n5661), .A2(n8350), .ZN(n5710) );
  NAND2_X1 U5192 ( .A1(n4822), .A2(n4821), .ZN(n5661) );
  AND2_X1 U5193 ( .A1(n4823), .A2(n8358), .ZN(n4821) );
  NAND2_X1 U5194 ( .A1(n8793), .A2(n4824), .ZN(n4822) );
  NAND2_X1 U5195 ( .A1(n5845), .A2(n8383), .ZN(n10171) );
  NOR2_X1 U5196 ( .A1(n5482), .A2(n4892), .ZN(n4891) );
  INV_X1 U5197 ( .A(n5465), .ZN(n4892) );
  NOR2_X1 U5198 ( .A1(n8930), .A2(n8879), .ZN(n4890) );
  OAI21_X1 U5199 ( .B1(n8121), .B2(n5403), .A(n5402), .ZN(n8888) );
  INV_X1 U5200 ( .A(n4422), .ZN(n5493) );
  NAND2_X1 U5201 ( .A1(n5134), .A2(n8392), .ZN(n5296) );
  INV_X1 U5202 ( .A(n5094), .ZN(n5096) );
  AND2_X1 U5203 ( .A1(n9101), .A2(n6362), .ZN(n9040) );
  OR2_X1 U5204 ( .A1(n9526), .A2(n9525), .ZN(n9534) );
  OR2_X1 U5205 ( .A1(n9611), .A2(n9754), .ZN(n5012) );
  NOR2_X1 U5206 ( .A1(n9655), .A2(n9104), .ZN(n8514) );
  NAND2_X1 U5207 ( .A1(n8206), .A2(n9846), .ZN(n8205) );
  INV_X1 U5208 ( .A(n6003), .ZN(n6286) );
  INV_X1 U5209 ( .A(n6753), .ZN(n6285) );
  BUF_X1 U5210 ( .A(n5960), .Z(n6753) );
  XNOR2_X1 U5211 ( .A(n7463), .B(n10015), .ZN(n9963) );
  AOI21_X1 U5212 ( .B1(n4691), .B2(n5551), .A(n4689), .ZN(n4688) );
  INV_X1 U5213 ( .A(n5558), .ZN(n4689) );
  INV_X1 U5214 ( .A(n5144), .ZN(n5142) );
  AND3_X1 U5215 ( .A1(n5581), .A2(n5580), .A3(n5579), .ZN(n8797) );
  AND4_X1 U5216 ( .A1(n5401), .A2(n5400), .A3(n5399), .A4(n5398), .ZN(n8200)
         );
  INV_X1 U5217 ( .A(n8971), .ZN(n8801) );
  INV_X1 U5218 ( .A(n5653), .ZN(n4636) );
  OAI21_X1 U5219 ( .B1(n8257), .B2(n8252), .A(n4634), .ZN(n4633) );
  AND2_X1 U5220 ( .A1(n5653), .A2(n8399), .ZN(n4634) );
  AND2_X1 U5221 ( .A1(n8296), .A2(n8285), .ZN(n4660) );
  OAI21_X1 U5222 ( .B1(n8278), .B2(n4815), .A(n8277), .ZN(n4659) );
  NAND2_X1 U5223 ( .A1(n4643), .A2(n8383), .ZN(n4642) );
  NAND2_X1 U5224 ( .A1(n4641), .A2(n8399), .ZN(n4640) );
  NAND2_X1 U5225 ( .A1(n8307), .A2(n8306), .ZN(n4643) );
  AND2_X1 U5226 ( .A1(n8312), .A2(n8311), .ZN(n4638) );
  AND2_X1 U5227 ( .A1(n9188), .A2(n9285), .ZN(n4719) );
  OAI22_X1 U5228 ( .A1(n9199), .A2(n9287), .B1(n9285), .B2(n9189), .ZN(n4717)
         );
  OAI21_X1 U5229 ( .B1(n4432), .B2(n4483), .A(n4725), .ZN(n4584) );
  NOR2_X1 U5230 ( .A1(n9212), .A2(n9285), .ZN(n4725) );
  NOR2_X1 U5231 ( .A1(n9374), .A2(n9287), .ZN(n4585) );
  NOR2_X1 U5232 ( .A1(n4432), .A2(n4580), .ZN(n4579) );
  NOR2_X1 U5233 ( .A1(n9228), .A2(n9287), .ZN(n4729) );
  OAI21_X1 U5234 ( .B1(n9249), .B2(n9388), .A(n4469), .ZN(n9250) );
  INV_X1 U5235 ( .A(n9264), .ZN(n4733) );
  INV_X1 U5236 ( .A(n5373), .ZN(n5374) );
  NAND2_X1 U5237 ( .A1(n5366), .A2(n5365), .ZN(n4706) );
  OR2_X1 U5238 ( .A1(n8765), .A2(n8655), .ZN(n8246) );
  AND2_X1 U5239 ( .A1(n4981), .A2(n4982), .ZN(n4980) );
  AND2_X1 U5240 ( .A1(n5444), .A2(SI_16_), .ZN(n5445) );
  NAND2_X1 U5241 ( .A1(n5755), .A2(n4907), .ZN(n5762) );
  AOI21_X1 U5242 ( .B1(n5754), .B2(n5753), .A(n5752), .ZN(n5755) );
  NAND2_X1 U5243 ( .A1(n5750), .A2(n4908), .ZN(n4907) );
  NOR2_X1 U5244 ( .A1(n4909), .A2(n5754), .ZN(n4908) );
  NOR2_X1 U5245 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5063) );
  INV_X1 U5246 ( .A(n7186), .ZN(n4767) );
  NOR2_X1 U5247 ( .A1(n7153), .A2(n4468), .ZN(n6573) );
  INV_X1 U5248 ( .A(n8133), .ZN(n4866) );
  AND2_X1 U5249 ( .A1(n8129), .A2(n6595), .ZN(n6596) );
  NAND2_X1 U5250 ( .A1(n6604), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4778) );
  NOR2_X1 U5251 ( .A1(n4474), .A2(n4434), .ZN(n4540) );
  NAND2_X1 U5252 ( .A1(n5048), .A2(n5047), .ZN(n5618) );
  INV_X1 U5253 ( .A(n5595), .ZN(n5048) );
  OR2_X1 U5254 ( .A1(n8624), .A2(n7951), .ZN(n8304) );
  OR2_X1 U5255 ( .A1(n8669), .A2(n7869), .ZN(n8264) );
  INV_X1 U5256 ( .A(n6508), .ZN(n4552) );
  NOR2_X1 U5257 ( .A1(n5568), .A2(n4883), .ZN(n4882) );
  INV_X1 U5258 ( .A(n5549), .ZN(n4883) );
  NAND2_X1 U5259 ( .A1(n8846), .A2(n4830), .ZN(n4828) );
  AOI21_X1 U5260 ( .B1(n8318), .B2(n4798), .A(n4797), .ZN(n4796) );
  INV_X1 U5261 ( .A(n8317), .ZN(n4798) );
  INV_X1 U5262 ( .A(n8322), .ZN(n4797) );
  INV_X1 U5263 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5328) );
  NOR2_X1 U5264 ( .A1(n6315), .A2(n4986), .ZN(n4985) );
  INV_X1 U5265 ( .A(n6300), .ZN(n4986) );
  AOI21_X1 U5266 ( .B1(n4974), .B2(n4976), .A(n4475), .ZN(n4971) );
  NAND2_X1 U5267 ( .A1(n4445), .A2(n4970), .ZN(n4967) );
  OR2_X1 U5268 ( .A1(n6063), .A2(n4514), .ZN(n4445) );
  NAND3_X1 U5269 ( .A1(n6043), .A2(n7369), .A3(n4446), .ZN(n4966) );
  NOR2_X1 U5270 ( .A1(n9498), .A2(n4610), .ZN(n9520) );
  AND2_X1 U5271 ( .A1(n9499), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4610) );
  INV_X1 U5272 ( .A(n9536), .ZN(n4601) );
  OR2_X1 U5273 ( .A1(n9766), .A2(n8501), .ZN(n9331) );
  OR2_X1 U5274 ( .A1(n4736), .A2(n4624), .ZN(n4622) );
  NAND2_X1 U5275 ( .A1(n9392), .A2(n9244), .ZN(n4624) );
  AND2_X1 U5276 ( .A1(n4671), .A2(n9742), .ZN(n4670) );
  NOR2_X1 U5277 ( .A1(n9810), .A2(n9097), .ZN(n4671) );
  AND2_X1 U5278 ( .A1(n7449), .A2(n9200), .ZN(n5002) );
  OR2_X1 U5279 ( .A1(n9190), .A2(n9188), .ZN(n7449) );
  OR2_X1 U5280 ( .A1(n10058), .A2(n9446), .ZN(n4937) );
  NOR2_X1 U5281 ( .A1(n4933), .A2(n7497), .ZN(n4932) );
  NAND2_X1 U5282 ( .A1(n7610), .A2(n9367), .ZN(n9183) );
  NAND2_X1 U5283 ( .A1(n9451), .A2(n10021), .ZN(n9367) );
  NAND2_X1 U5284 ( .A1(n9659), .A2(n9655), .ZN(n9649) );
  OR2_X1 U5285 ( .A1(n9285), .A2(n9410), .ZN(n10000) );
  NAND2_X1 U5286 ( .A1(n5676), .A2(n5675), .ZN(n5678) );
  NAND2_X1 U5287 ( .A1(n4692), .A2(n5535), .ZN(n4691) );
  INV_X1 U5288 ( .A(n5552), .ZN(n4692) );
  INV_X1 U5289 ( .A(n5483), .ZN(n5487) );
  NAND2_X1 U5290 ( .A1(n5319), .A2(SI_10_), .ZN(n5320) );
  INV_X1 U5291 ( .A(n5317), .ZN(n5321) );
  INV_X1 U5292 ( .A(n5253), .ZN(n4684) );
  NAND2_X1 U5293 ( .A1(n5207), .A2(SI_4_), .ZN(n5211) );
  OAI21_X1 U5294 ( .B1(n5122), .B2(n5120), .A(n4613), .ZN(n5145) );
  NAND2_X1 U5295 ( .A1(n5122), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4613) );
  NAND2_X1 U5296 ( .A1(n5132), .A2(n5946), .ZN(n5143) );
  INV_X1 U5297 ( .A(n4904), .ZN(n4903) );
  OR2_X1 U5298 ( .A1(n8671), .A2(n7309), .ZN(n8250) );
  XNOR2_X1 U5299 ( .A(n5762), .B(n7869), .ZN(n5765) );
  NAND2_X1 U5300 ( .A1(n4910), .A2(n7388), .ZN(n7320) );
  AND2_X1 U5301 ( .A1(n5767), .A2(n5766), .ZN(n4910) );
  INV_X1 U5302 ( .A(n7323), .ZN(n5767) );
  OR2_X1 U5303 ( .A1(n8569), .A2(n5812), .ZN(n4927) );
  NOR2_X1 U5304 ( .A1(n7932), .A2(n8660), .ZN(n4914) );
  NAND2_X1 U5305 ( .A1(n7932), .A2(n8660), .ZN(n4916) );
  NOR2_X1 U5306 ( .A1(n5789), .A2(n4914), .ZN(n4913) );
  NOR2_X1 U5307 ( .A1(n5816), .A2(n4926), .ZN(n4925) );
  INV_X1 U5308 ( .A(n5811), .ZN(n4926) );
  XNOR2_X1 U5309 ( .A(n5762), .B(n5136), .ZN(n5758) );
  AND4_X1 U5310 ( .A1(n5481), .A2(n5480), .A3(n5479), .A4(n5478), .ZN(n5806)
         );
  INV_X1 U5311 ( .A(n7983), .ZN(n5088) );
  NAND2_X1 U5312 ( .A1(n6564), .A2(n4761), .ZN(n6567) );
  NAND2_X1 U5313 ( .A1(n4762), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n4761) );
  NOR2_X1 U5314 ( .A1(n7173), .A2(n7385), .ZN(n7172) );
  NOR2_X1 U5315 ( .A1(n7189), .A2(n6533), .ZN(n6534) );
  OR2_X1 U5316 ( .A1(n8477), .A2(n8478), .ZN(n4775) );
  NAND2_X1 U5317 ( .A1(n4860), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4858) );
  INV_X1 U5318 ( .A(n5014), .ZN(n4859) );
  NOR2_X1 U5319 ( .A1(n7699), .A2(n10254), .ZN(n4856) );
  OR2_X1 U5320 ( .A1(n7998), .A2(n10258), .ZN(n4865) );
  XNOR2_X1 U5321 ( .A(n6596), .B(n8186), .ZN(n8184) );
  INV_X1 U5322 ( .A(n10145), .ZN(n4851) );
  OR2_X1 U5323 ( .A1(n8184), .A2(n8183), .ZN(n4784) );
  NAND2_X1 U5324 ( .A1(n4781), .A2(n4779), .ZN(n6600) );
  AND2_X1 U5325 ( .A1(n4782), .A2(n4522), .ZN(n4781) );
  INV_X1 U5326 ( .A(n4799), .ZN(n8446) );
  OAI21_X1 U5327 ( .B1(n5710), .B2(n4803), .A(n4800), .ZN(n4799) );
  NAND2_X1 U5328 ( .A1(n4808), .A2(n6510), .ZN(n4803) );
  INV_X1 U5329 ( .A(n4801), .ZN(n4800) );
  NAND2_X1 U5330 ( .A1(n5044), .A2(n5043), .ZN(n5577) );
  INV_X1 U5331 ( .A(n5563), .ZN(n5044) );
  NAND2_X1 U5332 ( .A1(n5040), .A2(n5039), .ZN(n5524) );
  INV_X1 U5333 ( .A(n5509), .ZN(n5040) );
  INV_X1 U5334 ( .A(n4889), .ZN(n4888) );
  OAI21_X1 U5335 ( .B1(n8844), .B2(n4476), .A(n5502), .ZN(n4889) );
  NAND2_X1 U5336 ( .A1(n5038), .A2(n6842), .ZN(n5476) );
  INV_X1 U5337 ( .A(n5459), .ZN(n5038) );
  OAI21_X1 U5338 ( .B1(n7950), .B2(n5355), .A(n5354), .ZN(n7975) );
  OR2_X1 U5339 ( .A1(n10232), .A2(n8660), .ZN(n5354) );
  AOI21_X1 U5340 ( .B1(n4839), .B2(n8281), .A(n4838), .ZN(n4837) );
  INV_X1 U5341 ( .A(n8288), .ZN(n4838) );
  NAND2_X1 U5342 ( .A1(n7742), .A2(n5654), .ZN(n7624) );
  NAND2_X1 U5343 ( .A1(n7718), .A2(n5198), .ZN(n7717) );
  NAND2_X1 U5344 ( .A1(n5154), .A2(n5025), .ZN(n5199) );
  INV_X1 U5345 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5025) );
  NAND2_X1 U5346 ( .A1(n4547), .A2(n4546), .ZN(n4545) );
  AND2_X1 U5347 ( .A1(n4437), .A2(n5137), .ZN(n4546) );
  NAND2_X1 U5348 ( .A1(n7582), .A2(n8671), .ZN(n7377) );
  NAND2_X1 U5349 ( .A1(n8082), .A2(n8396), .ZN(n4712) );
  OR2_X1 U5350 ( .A1(n4881), .A2(n5582), .ZN(n4880) );
  AND2_X1 U5351 ( .A1(n8966), .A2(n8656), .ZN(n5582) );
  INV_X1 U5352 ( .A(n5567), .ZN(n4881) );
  INV_X1 U5353 ( .A(n4879), .ZN(n4878) );
  OAI22_X1 U5354 ( .A1(n4880), .A2(n4882), .B1(n8966), .B2(n8656), .ZN(n4879)
         );
  NAND2_X1 U5355 ( .A1(n8358), .A2(n8350), .ZN(n8771) );
  AOI21_X1 U5356 ( .B1(n4824), .B2(n8406), .A(n8403), .ZN(n4823) );
  OR2_X1 U5357 ( .A1(n8403), .A2(n8402), .ZN(n8780) );
  OR2_X1 U5358 ( .A1(n8977), .A2(n8657), .ZN(n5549) );
  NAND2_X1 U5359 ( .A1(n5660), .A2(n8346), .ZN(n8793) );
  OR2_X1 U5360 ( .A1(n8826), .A2(n8807), .ZN(n5531) );
  NAND2_X1 U5361 ( .A1(n8346), .A2(n8345), .ZN(n8806) );
  AND2_X1 U5362 ( .A1(n8335), .A2(n8334), .ZN(n4830) );
  NAND2_X1 U5363 ( .A1(n8877), .A2(n8878), .ZN(n5466) );
  NAND2_X1 U5364 ( .A1(n8845), .A2(n8844), .ZN(n8843) );
  OR2_X1 U5365 ( .A1(n9010), .A2(n8227), .ZN(n8874) );
  AND2_X1 U5366 ( .A1(n5847), .A2(n8383), .ZN(n8891) );
  INV_X1 U5367 ( .A(n10171), .ZN(n8889) );
  AND3_X1 U5368 ( .A1(n5260), .A2(n5259), .A3(n5258), .ZN(n10204) );
  AND3_X1 U5369 ( .A1(n5197), .A2(n5196), .A3(n5195), .ZN(n10189) );
  AOI21_X1 U5370 ( .B1(n5633), .B2(n8058), .A(n5632), .ZN(n6724) );
  NOR2_X1 U5371 ( .A1(n4792), .A2(n5076), .ZN(n5081) );
  NAND2_X1 U5372 ( .A1(n5057), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5071) );
  NAND2_X1 U5373 ( .A1(n5255), .A2(n5276), .ZN(n5297) );
  OR2_X1 U5374 ( .A1(n5167), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n5192) );
  NAND2_X1 U5375 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5147) );
  INV_X1 U5376 ( .A(n9451), .ZN(n7467) );
  INV_X1 U5377 ( .A(n7444), .ZN(n7443) );
  NOR2_X1 U5378 ( .A1(n4992), .A2(n4993), .ZN(n4991) );
  INV_X1 U5379 ( .A(n9029), .ZN(n4993) );
  INV_X1 U5380 ( .A(n9122), .ZN(n4998) );
  INV_X1 U5381 ( .A(n9100), .ZN(n4999) );
  INV_X1 U5382 ( .A(n9101), .ZN(n4996) );
  OR2_X1 U5383 ( .A1(n9147), .A2(n9148), .ZN(n6408) );
  OR2_X1 U5384 ( .A1(n9596), .A2(n9290), .ZN(n9408) );
  NAND2_X1 U5385 ( .A1(n4573), .A2(n4571), .ZN(n4570) );
  NOR2_X1 U5386 ( .A1(n9324), .A2(n4572), .ZN(n4571) );
  NAND2_X1 U5387 ( .A1(n9288), .A2(n9751), .ZN(n4573) );
  AND2_X1 U5388 ( .A1(n9354), .A2(n9287), .ZN(n4572) );
  OR2_X1 U5389 ( .A1(n6009), .A2(n7026), .ZN(n4948) );
  OR2_X1 U5390 ( .A1(n9468), .A2(n9467), .ZN(n4607) );
  AOI21_X1 U5391 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n7093), .A(n7088), .ZN(
        n7092) );
  NOR2_X1 U5392 ( .A1(n7564), .A2(n4515), .ZN(n7568) );
  NOR2_X1 U5393 ( .A1(n7568), .A2(n7567), .ZN(n7665) );
  XNOR2_X1 U5394 ( .A(n9520), .B(n4609), .ZN(n9500) );
  NOR2_X1 U5395 ( .A1(n9500), .A2(n8050), .ZN(n9521) );
  AND2_X1 U5396 ( .A1(n9534), .A2(n9533), .ZN(n9535) );
  NAND2_X1 U5397 ( .A1(n9535), .A2(n9536), .ZN(n9553) );
  NOR2_X1 U5398 ( .A1(n9759), .A2(n4674), .ZN(n4673) );
  INV_X1 U5399 ( .A(n4675), .ZN(n4674) );
  OR2_X1 U5400 ( .A1(n4444), .A2(n9394), .ZN(n4751) );
  NAND2_X1 U5401 ( .A1(n4753), .A2(n4731), .ZN(n4752) );
  NOR2_X1 U5402 ( .A1(n9664), .A2(n8500), .ZN(n9644) );
  NAND2_X1 U5403 ( .A1(n4940), .A2(n4939), .ZN(n9642) );
  AOI21_X1 U5404 ( .B1(n4493), .B2(n4941), .A(n4443), .ZN(n4939) );
  NOR2_X1 U5405 ( .A1(n9665), .A2(n9666), .ZN(n9664) );
  AND2_X1 U5406 ( .A1(n9663), .A2(n9673), .ZN(n9659) );
  OR2_X1 U5407 ( .A1(n9719), .A2(n9794), .ZN(n9701) );
  NAND2_X1 U5408 ( .A1(n4498), .A2(n4433), .ZN(n4952) );
  NAND2_X1 U5409 ( .A1(n4433), .A2(n4954), .ZN(n4953) );
  INV_X1 U5410 ( .A(n4956), .ZN(n4954) );
  NAND2_X1 U5411 ( .A1(n4737), .A2(n4740), .ZN(n4735) );
  AND2_X1 U5412 ( .A1(n9390), .A2(n9392), .ZN(n9731) );
  NAND2_X1 U5413 ( .A1(n9083), .A2(n9439), .ZN(n4957) );
  OR2_X1 U5414 ( .A1(n8040), .A2(n8048), .ZN(n8084) );
  INV_X1 U5415 ( .A(n10092), .ZN(n8045) );
  OR2_X1 U5416 ( .A1(n7947), .A2(n8068), .ZN(n9894) );
  NOR2_X1 U5417 ( .A1(n9915), .A2(n4580), .ZN(n4721) );
  OR2_X1 U5418 ( .A1(n9920), .A2(n7642), .ZN(n9209) );
  NAND2_X1 U5419 ( .A1(n4723), .A2(n9371), .ZN(n4722) );
  AND2_X1 U5420 ( .A1(n9369), .A2(n9302), .ZN(n4723) );
  AND2_X1 U5421 ( .A1(n9209), .A2(n9210), .ZN(n9910) );
  NAND2_X1 U5422 ( .A1(n7450), .A2(n5002), .ZN(n9371) );
  INV_X1 U5423 ( .A(n7496), .ZN(n7450) );
  NAND2_X1 U5424 ( .A1(n9183), .A2(n9185), .ZN(n9942) );
  NAND2_X1 U5425 ( .A1(n7593), .A2(n9297), .ZN(n7592) );
  NAND2_X1 U5426 ( .A1(n8541), .A2(n8540), .ZN(n9754) );
  NAND2_X1 U5427 ( .A1(n8082), .A2(n9176), .ZN(n6395) );
  AND2_X1 U5428 ( .A1(n6238), .A2(n6237), .ZN(n9859) );
  OR2_X1 U5429 ( .A1(n6723), .A2(n5979), .ZN(n6067) );
  AND2_X1 U5430 ( .A1(n7552), .A2(n7111), .ZN(n10059) );
  NAND2_X1 U5431 ( .A1(n8391), .A2(n8390), .ZN(n8395) );
  XNOR2_X1 U5432 ( .A(n8389), .B(n8388), .ZN(n8535) );
  NOR2_X1 U5433 ( .A1(n4559), .A2(n5893), .ZN(n4565) );
  XNOR2_X1 U5434 ( .A(n5688), .B(n5687), .ZN(n8126) );
  XNOR2_X1 U5435 ( .A(n5605), .B(n5604), .ZN(n8056) );
  INV_X1 U5436 ( .A(n4691), .ZN(n4687) );
  NAND2_X1 U5437 ( .A1(n4693), .A2(n5535), .ZN(n5553) );
  XNOR2_X1 U5438 ( .A(n5414), .B(n5413), .ZN(n7305) );
  AND2_X1 U5439 ( .A1(n5412), .A2(n5439), .ZN(n5414) );
  NOR2_X1 U5440 ( .A1(n5877), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n4563) );
  NOR2_X1 U5441 ( .A1(n4620), .A2(n4619), .ZN(n4618) );
  INV_X1 U5442 ( .A(n5271), .ZN(n4620) );
  INV_X1 U5443 ( .A(n5231), .ZN(n4619) );
  NAND2_X1 U5444 ( .A1(n4683), .A2(n5271), .ZN(n4617) );
  OAI21_X1 U5445 ( .B1(n5249), .B2(n4684), .A(n5267), .ZN(n4683) );
  XNOR2_X1 U5446 ( .A(n5269), .B(SI_7_), .ZN(n5267) );
  XNOR2_X1 U5447 ( .A(n5251), .B(SI_6_), .ZN(n5249) );
  NAND2_X1 U5448 ( .A1(n5232), .A2(n5231), .ZN(n5250) );
  AOI21_X1 U5449 ( .B1(n8639), .B2(n8774), .A(n5833), .ZN(n8555) );
  AND4_X1 U5450 ( .A1(n5514), .A2(n5513), .A3(n5512), .A4(n5511), .ZN(n8822)
         );
  NOR2_X1 U5451 ( .A1(n5822), .A2(n5022), .ZN(n5826) );
  NAND2_X1 U5452 ( .A1(n8151), .A2(n5800), .ZN(n8196) );
  NAND2_X1 U5453 ( .A1(n7390), .A2(n7389), .ZN(n7388) );
  AND4_X1 U5454 ( .A1(n5501), .A2(n5500), .A3(n5499), .A4(n5498), .ZN(n8865)
         );
  AND4_X1 U5455 ( .A1(n5385), .A2(n5384), .A3(n5383), .A4(n5382), .ZN(n8123)
         );
  AND4_X1 U5456 ( .A1(n5464), .A2(n5463), .A3(n5462), .A4(n5461), .ZN(n8866)
         );
  NAND2_X1 U5457 ( .A1(n5111), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5112) );
  NOR2_X1 U5458 ( .A1(n8444), .A2(n4480), .ZN(n4710) );
  NAND2_X1 U5459 ( .A1(n8387), .A2(n4471), .ZN(n4709) );
  INV_X1 U5460 ( .A(n5806), .ZN(n8879) );
  XNOR2_X1 U5461 ( .A(n5217), .B(P2_IR_REG_5__SCAN_IN), .ZN(n8483) );
  XNOR2_X1 U5462 ( .A(n6605), .B(n8720), .ZN(n8716) );
  OAI21_X1 U5463 ( .B1(n8722), .B2(n10147), .A(n4477), .ZN(n4787) );
  NOR2_X1 U5464 ( .A1(n8716), .A2(n8882), .ZN(n8718) );
  NOR2_X1 U5465 ( .A1(n5707), .A2(n5706), .ZN(n5708) );
  OR2_X1 U5466 ( .A1(n8958), .A2(n8901), .ZN(n5672) );
  NAND2_X1 U5467 ( .A1(n5475), .A2(n5474), .ZN(n8930) );
  NAND2_X1 U5468 ( .A1(n5395), .A2(n5394), .ZN(n8941) );
  AND3_X1 U5469 ( .A1(n5280), .A2(n5279), .A3(n5278), .ZN(n10210) );
  INV_X1 U5470 ( .A(n8839), .ZN(n8898) );
  INV_X1 U5471 ( .A(n4843), .ZN(n6693) );
  OAI21_X1 U5472 ( .B1(n8761), .B2(n4841), .A(n4844), .ZN(n4843) );
  NOR2_X1 U5473 ( .A1(n4842), .A2(n10216), .ZN(n4841) );
  OAI21_X1 U5474 ( .B1(n5710), .B2(n4807), .A(n4805), .ZN(n6511) );
  XOR2_X1 U5475 ( .A(n8436), .B(n5710), .Z(n8958) );
  INV_X1 U5476 ( .A(n4537), .ZN(n5674) );
  AND2_X1 U5477 ( .A1(n5562), .A2(n5561), .ZN(n8971) );
  INV_X1 U5478 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4644) );
  OR3_X1 U5479 ( .A1(n8100), .A2(n8061), .A3(n8027), .ZN(n6705) );
  AND2_X1 U5480 ( .A1(n6469), .A2(n9150), .ZN(n6470) );
  NAND2_X1 U5481 ( .A1(n6100), .A2(n6099), .ZN(n7866) );
  NAND2_X1 U5482 ( .A1(n4586), .A2(n5960), .ZN(n4588) );
  OAI22_X1 U5483 ( .A1(n6722), .A2(n8392), .B1(n4587), .B2(n5120), .ZN(n4586)
         );
  OR2_X1 U5484 ( .A1(n5990), .A2(n5989), .ZN(n7463) );
  OR2_X1 U5485 ( .A1(n7078), .A2(n7077), .ZN(n4605) );
  AND2_X1 U5486 ( .A1(n4607), .A2(n4606), .ZN(n7078) );
  NAND2_X1 U5487 ( .A1(n9473), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4606) );
  NAND2_X1 U5488 ( .A1(n4961), .A2(n8517), .ZN(n8519) );
  OAI21_X1 U5489 ( .B1(n4629), .B2(n9913), .A(n9633), .ZN(n9769) );
  XNOR2_X1 U5490 ( .A(n4754), .B(n9632), .ZN(n4629) );
  NAND2_X1 U5491 ( .A1(n4755), .A2(n9336), .ZN(n4754) );
  AOI21_X1 U5492 ( .B1(n4632), .B2(n4631), .A(n8410), .ZN(n8275) );
  INV_X1 U5493 ( .A(n8262), .ZN(n4631) );
  NAND2_X1 U5494 ( .A1(n4636), .A2(n8383), .ZN(n4635) );
  OAI211_X1 U5495 ( .C1(n8280), .C2(n8399), .A(n4660), .B(n4658), .ZN(n8300)
         );
  NAND2_X1 U5496 ( .A1(n4639), .A2(n4638), .ZN(n4637) );
  INV_X1 U5497 ( .A(n4717), .ZN(n4716) );
  OAI21_X1 U5498 ( .B1(n4479), .B2(n8383), .A(n4652), .ZN(n4651) );
  NOR2_X1 U5499 ( .A1(n8873), .A2(n4653), .ZN(n4652) );
  NOR2_X1 U5500 ( .A1(n8322), .A2(n8399), .ZN(n4653) );
  INV_X1 U5501 ( .A(n4584), .ZN(n4583) );
  INV_X1 U5502 ( .A(n9310), .ZN(n4730) );
  INV_X1 U5503 ( .A(n9057), .ZN(n4981) );
  INV_X1 U5504 ( .A(n5341), .ZN(n4700) );
  AOI21_X1 U5505 ( .B1(n4704), .B2(n4703), .A(n4496), .ZN(n4702) );
  INV_X1 U5506 ( .A(n5365), .ZN(n4703) );
  NOR2_X1 U5507 ( .A1(n4705), .A2(n4697), .ZN(n4696) );
  NAND2_X1 U5508 ( .A1(n5342), .A2(n5341), .ZN(n4697) );
  INV_X1 U5509 ( .A(n5751), .ZN(n4909) );
  NAND2_X1 U5510 ( .A1(n8364), .A2(n8385), .ZN(n4645) );
  AND2_X1 U5511 ( .A1(n5754), .A2(n7409), .ZN(n5752) );
  INV_X1 U5512 ( .A(n4792), .ZN(n4551) );
  NOR2_X1 U5513 ( .A1(n5076), .A2(n4489), .ZN(n4550) );
  AND2_X1 U5514 ( .A1(n8019), .A2(n4975), .ZN(n4974) );
  OR2_X1 U5515 ( .A1(n7941), .A2(n4976), .ZN(n4975) );
  INV_X1 U5516 ( .A(n6183), .ZN(n4976) );
  NAND2_X1 U5517 ( .A1(n4732), .A2(n4731), .ZN(n9265) );
  NOR2_X1 U5518 ( .A1(n9771), .A2(n9776), .ZN(n4677) );
  NAND2_X1 U5519 ( .A1(n6505), .A2(n6504), .ZN(n8369) );
  NAND2_X1 U5520 ( .A1(n6501), .A2(n6500), .ZN(n6505) );
  INV_X1 U5521 ( .A(n5404), .ZN(n5408) );
  INV_X1 U5522 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5115) );
  INV_X1 U5523 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5117) );
  INV_X1 U5524 ( .A(n5821), .ZN(n4923) );
  INV_X1 U5525 ( .A(n8366), .ZN(n8382) );
  OAI21_X1 U5526 ( .B1(n7186), .B2(n6568), .A(n4769), .ZN(n4768) );
  AND2_X1 U5527 ( .A1(n4767), .A2(n7172), .ZN(n4765) );
  NAND2_X1 U5528 ( .A1(n7185), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4769) );
  NAND2_X1 U5529 ( .A1(n6577), .A2(n6576), .ZN(n6578) );
  NAND2_X1 U5530 ( .A1(n7216), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6576) );
  INV_X1 U5531 ( .A(n6579), .ZN(n4771) );
  OR2_X1 U5532 ( .A1(n10130), .A2(n6581), .ZN(n6583) );
  INV_X1 U5533 ( .A(n4760), .ZN(n4759) );
  NAND2_X1 U5534 ( .A1(n6592), .A2(n6593), .ZN(n7990) );
  NAND2_X1 U5535 ( .A1(n6592), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4760) );
  INV_X1 U5536 ( .A(n10143), .ZN(n4785) );
  OAI21_X1 U5537 ( .B1(n4805), .B2(n4802), .A(n4495), .ZN(n4801) );
  INV_X1 U5538 ( .A(n6510), .ZN(n4802) );
  NOR2_X1 U5539 ( .A1(n4895), .A2(n5301), .ZN(n4533) );
  NAND2_X1 U5540 ( .A1(n7627), .A2(n5281), .ZN(n4535) );
  NAND2_X1 U5541 ( .A1(n5281), .A2(n8285), .ZN(n4534) );
  OAI21_X1 U5542 ( .B1(n5198), .B2(n4873), .A(n7755), .ZN(n4872) );
  NAND2_X1 U5543 ( .A1(n5178), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5140) );
  INV_X1 U5544 ( .A(n8439), .ZN(n4554) );
  OR2_X1 U5545 ( .A1(n9003), .A2(n8866), .ZN(n8327) );
  INV_X1 U5546 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5090) );
  INV_X1 U5547 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n4930) );
  INV_X1 U5548 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n4931) );
  NOR2_X1 U5549 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n4764) );
  NOR2_X1 U5550 ( .A1(n4967), .A2(n4965), .ZN(n4964) );
  INV_X1 U5551 ( .A(n6113), .ZN(n4965) );
  INV_X1 U5552 ( .A(n9605), .ZN(n9606) );
  OR2_X1 U5553 ( .A1(n9754), .A2(n9276), .ZN(n9329) );
  OR2_X1 U5554 ( .A1(n9759), .A2(n9606), .ZN(n9328) );
  INV_X1 U5555 ( .A(n9308), .ZN(n4740) );
  NAND2_X1 U5556 ( .A1(n4627), .A2(n9442), .ZN(n9222) );
  NAND2_X1 U5557 ( .A1(n4667), .A2(n10042), .ZN(n4666) );
  INV_X1 U5558 ( .A(n4668), .ZN(n4667) );
  NAND2_X1 U5559 ( .A1(n10035), .A2(n10028), .ZN(n4668) );
  NAND2_X1 U5560 ( .A1(n9366), .A2(n4576), .ZN(n4575) );
  INV_X1 U5561 ( .A(n7445), .ZN(n4576) );
  NAND2_X1 U5562 ( .A1(n9659), .A2(n4677), .ZN(n9634) );
  XNOR2_X1 U5563 ( .A(n8369), .B(n8368), .ZN(n8367) );
  NOR2_X1 U5564 ( .A1(n4440), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n4962) );
  AND2_X1 U5565 ( .A1(n4566), .A2(n5903), .ZN(n4557) );
  INV_X1 U5566 ( .A(n5877), .ZN(n4558) );
  INV_X1 U5567 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n4566) );
  NOR2_X1 U5568 ( .A1(n5893), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n4561) );
  OAI21_X2 U5569 ( .B1(n5883), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5885) );
  OR2_X1 U5570 ( .A1(n5436), .A2(n5435), .ZN(n5437) );
  AND2_X1 U5571 ( .A1(n5405), .A2(n5407), .ZN(n5444) );
  INV_X1 U5572 ( .A(n6044), .ZN(n4564) );
  XNOR2_X1 U5573 ( .A(n5318), .B(SI_10_), .ZN(n5317) );
  OAI211_X1 U5574 ( .C1(n4617), .C2(n5290), .A(n5289), .B(n4615), .ZN(n5302)
         );
  NAND2_X1 U5575 ( .A1(n5208), .A2(n5211), .ZN(n5213) );
  OAI21_X1 U5576 ( .B1(n5186), .B2(P1_DATAO_REG_4__SCAN_IN), .A(n5185), .ZN(
        n5206) );
  OR2_X1 U5577 ( .A1(n5122), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5185) );
  OAI21_X1 U5578 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(P1_IR_REG_1__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6001) );
  INV_X1 U5579 ( .A(SI_1_), .ZN(n4612) );
  OAI21_X1 U5580 ( .B1(n4906), .B2(n4901), .A(n4900), .ZN(n7791) );
  AOI21_X1 U5581 ( .B1(n4904), .B2(n4902), .A(n8662), .ZN(n4900) );
  NAND2_X1 U5582 ( .A1(n5033), .A2(n5032), .ZN(n5356) );
  INV_X1 U5583 ( .A(n5348), .ZN(n5033) );
  NAND2_X1 U5584 ( .A1(n4906), .A2(n5779), .ZN(n7765) );
  AOI21_X1 U5585 ( .B1(n4925), .B2(n5812), .A(n4492), .ZN(n4924) );
  NAND2_X1 U5586 ( .A1(n8615), .A2(n8618), .ZN(n8617) );
  NAND2_X1 U5587 ( .A1(n5774), .A2(n5773), .ZN(n7412) );
  NAND3_X1 U5588 ( .A1(n4430), .A2(n5077), .A3(n5078), .ZN(n5111) );
  INV_X1 U5589 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5078) );
  OR2_X1 U5590 ( .A1(n7172), .A2(n6569), .ZN(n4766) );
  NAND2_X1 U5591 ( .A1(n4845), .A2(n7190), .ZN(n4847) );
  INV_X1 U5592 ( .A(n6533), .ZN(n4845) );
  CLKBUF_X1 U5593 ( .A(n7160), .Z(n7253) );
  NAND2_X1 U5594 ( .A1(n6574), .A2(n6714), .ZN(n4774) );
  INV_X1 U5595 ( .A(n7219), .ZN(n6538) );
  XNOR2_X1 U5596 ( .A(n6578), .B(n7237), .ZN(n7239) );
  AND2_X1 U5597 ( .A1(n6578), .A2(n7237), .ZN(n6579) );
  NOR2_X1 U5598 ( .A1(n4770), .A2(n4772), .ZN(n10130) );
  OAI21_X1 U5599 ( .B1(n6579), .B2(P2_REG2_REG_7__SCAN_IN), .A(n4773), .ZN(
        n4772) );
  AND2_X1 U5600 ( .A1(n4771), .A2(n7239), .ZN(n4770) );
  INV_X1 U5601 ( .A(n10131), .ZN(n4773) );
  NOR2_X1 U5602 ( .A1(n7239), .A2(n7240), .ZN(n7238) );
  NOR2_X1 U5603 ( .A1(n7242), .A2(n10250), .ZN(n7241) );
  XNOR2_X1 U5604 ( .A(n6583), .B(n6582), .ZN(n7530) );
  INV_X1 U5605 ( .A(n7708), .ZN(n6587) );
  INV_X1 U5606 ( .A(n4784), .ZN(n8182) );
  INV_X1 U5607 ( .A(n6600), .ZN(n6601) );
  NAND2_X1 U5608 ( .A1(n4777), .A2(n4776), .ZN(n8702) );
  OR2_X1 U5609 ( .A1(n10162), .A2(n8720), .ZN(n4789) );
  NAND2_X1 U5610 ( .A1(n10141), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n4790) );
  INV_X1 U5611 ( .A(n4867), .ZN(n8710) );
  AND2_X1 U5612 ( .A1(n7307), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4868) );
  INV_X1 U5613 ( .A(n6605), .ZN(n6606) );
  NAND2_X1 U5614 ( .A1(n8445), .A2(n8381), .ZN(n8439) );
  NOR2_X1 U5615 ( .A1(n8646), .A2(n5626), .ZN(n5707) );
  INV_X1 U5616 ( .A(n4540), .ZN(n4539) );
  AOI21_X1 U5617 ( .B1(n4542), .B2(n4540), .A(n4497), .ZN(n4538) );
  NAND2_X1 U5618 ( .A1(n5046), .A2(n5045), .ZN(n5593) );
  INV_X1 U5619 ( .A(n5577), .ZN(n5046) );
  NAND2_X1 U5620 ( .A1(n5042), .A2(n5041), .ZN(n5543) );
  INV_X1 U5621 ( .A(n5524), .ZN(n5042) );
  NAND2_X1 U5622 ( .A1(n5037), .A2(n5036), .ZN(n5421) );
  INV_X1 U5623 ( .A(n5396), .ZN(n5037) );
  AND4_X1 U5624 ( .A1(n5426), .A2(n5425), .A3(n5424), .A4(n5423), .ZN(n8227)
         );
  NAND2_X1 U5625 ( .A1(n5035), .A2(n5034), .ZN(n5380) );
  INV_X1 U5626 ( .A(n5356), .ZN(n5035) );
  AND2_X1 U5627 ( .A1(n7895), .A2(n8306), .ZN(n7956) );
  AND4_X1 U5628 ( .A1(n5353), .A2(n5352), .A3(n5351), .A4(n5350), .ZN(n8621)
         );
  OAI21_X2 U5629 ( .B1(n7901), .B2(n5316), .A(n5315), .ZN(n7893) );
  INV_X1 U5630 ( .A(n8419), .ZN(n7892) );
  AND2_X1 U5631 ( .A1(n8304), .A2(n8306), .ZN(n8419) );
  OAI21_X1 U5632 ( .B1(n7730), .B2(n4834), .A(n4831), .ZN(n7896) );
  AOI21_X1 U5633 ( .B1(n4833), .B2(n4840), .A(n4832), .ZN(n4831) );
  INV_X1 U5634 ( .A(n8301), .ZN(n4832) );
  NAND2_X1 U5635 ( .A1(n4535), .A2(n4532), .ZN(n7778) );
  AND2_X1 U5636 ( .A1(n4534), .A2(n5282), .ZN(n4532) );
  NAND2_X1 U5637 ( .A1(n7733), .A2(n5281), .ZN(n7731) );
  OR2_X1 U5638 ( .A1(n7627), .A2(n8285), .ZN(n7733) );
  NAND2_X1 U5639 ( .A1(n5029), .A2(n5028), .ZN(n5261) );
  INV_X1 U5640 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5028) );
  INV_X1 U5641 ( .A(n5243), .ZN(n5029) );
  AOI21_X1 U5642 ( .B1(n4817), .B2(n4816), .A(n4815), .ZN(n4814) );
  INV_X1 U5643 ( .A(n8265), .ZN(n4816) );
  NAND2_X1 U5644 ( .A1(n4812), .A2(n4817), .ZN(n4813) );
  NAND2_X1 U5645 ( .A1(n4813), .A2(n4811), .ZN(n7742) );
  AND2_X1 U5646 ( .A1(n4814), .A2(n4820), .ZN(n4811) );
  OR2_X1 U5647 ( .A1(n5221), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5243) );
  NAND2_X1 U5648 ( .A1(n5027), .A2(n5026), .ZN(n5221) );
  INV_X1 U5649 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5026) );
  INV_X1 U5650 ( .A(n5199), .ZN(n5027) );
  NAND2_X1 U5651 ( .A1(n8352), .A2(n8357), .ZN(n4809) );
  XNOR2_X1 U5652 ( .A(n8378), .B(n8654), .ZN(n8437) );
  AND2_X1 U5653 ( .A1(n4810), .A2(n8357), .ZN(n8436) );
  NAND2_X1 U5654 ( .A1(n4877), .A2(n5567), .ZN(n8782) );
  NAND2_X1 U5655 ( .A1(n5550), .A2(n4882), .ZN(n4877) );
  OAI21_X1 U5656 ( .B1(n8845), .B2(n4829), .A(n4484), .ZN(n5659) );
  INV_X1 U5657 ( .A(n4830), .ZN(n4829) );
  OR2_X1 U5658 ( .A1(n8836), .A2(n8848), .ZN(n5515) );
  AND4_X1 U5659 ( .A1(n5548), .A2(n5547), .A3(n5546), .A4(n5545), .ZN(n8821)
         );
  NAND2_X1 U5660 ( .A1(n4794), .A2(n4793), .ZN(n8859) );
  AND2_X1 U5661 ( .A1(n4463), .A2(n4796), .ZN(n4793) );
  NAND2_X1 U5662 ( .A1(n4794), .A2(n4796), .ZN(n8854) );
  NOR2_X1 U5663 ( .A1(n9840), .A2(n5372), .ZN(n4893) );
  AND3_X1 U5664 ( .A1(n5239), .A2(n5238), .A3(n5237), .ZN(n10198) );
  AND3_X1 U5665 ( .A1(n5220), .A2(n5219), .A3(n5218), .ZN(n10194) );
  NAND2_X1 U5666 ( .A1(n5072), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5073) );
  INV_X1 U5667 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5070) );
  INV_X1 U5668 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5064) );
  NOR3_X2 U5669 ( .A1(n5326), .A2(n4917), .A3(n4919), .ZN(n5058) );
  NAND2_X1 U5670 ( .A1(n4918), .A2(n5056), .ZN(n4917) );
  INV_X1 U5671 ( .A(n5055), .ZN(n4918) );
  OR2_X1 U5672 ( .A1(n6205), .A2(n9032), .ZN(n6239) );
  NAND2_X1 U5673 ( .A1(n9028), .A2(n9029), .ZN(n9027) );
  AND2_X1 U5674 ( .A1(n6350), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6365) );
  AOI21_X1 U5675 ( .B1(n4985), .B2(n4983), .A(n4491), .ZN(n4982) );
  INV_X1 U5676 ( .A(n9050), .ZN(n4983) );
  INV_X1 U5677 ( .A(n4985), .ZN(n4984) );
  OAI21_X1 U5678 ( .B1(n9039), .B2(n9125), .A(n9040), .ZN(n9038) );
  INV_X1 U5679 ( .A(n4967), .ZN(n4963) );
  OR2_X1 U5680 ( .A1(n6103), .A2(n7278), .ZN(n6144) );
  NOR2_X1 U5681 ( .A1(n6339), .A2(n9132), .ZN(n6350) );
  NOR2_X1 U5682 ( .A1(n9123), .A2(n9122), .ZN(n9039) );
  AND2_X1 U5683 ( .A1(n6146), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6171) );
  AND2_X1 U5684 ( .A1(n6328), .A2(n6327), .ZN(n9116) );
  AND3_X1 U5685 ( .A1(n6293), .A2(n6292), .A3(n6291), .ZN(n9115) );
  AND3_X1 U5686 ( .A1(n6229), .A2(n6228), .A3(n6227), .ZN(n8169) );
  NAND2_X1 U5687 ( .A1(n5930), .A2(n8468), .ZN(n5987) );
  AOI21_X1 U5688 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(n7035), .A(n7055), .ZN(
        n9458) );
  AND2_X1 U5689 ( .A1(n4605), .A2(n4604), .ZN(n7030) );
  NAND2_X1 U5690 ( .A1(n7031), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4604) );
  NOR2_X1 U5691 ( .A1(n7273), .A2(n4608), .ZN(n7275) );
  AND2_X1 U5692 ( .A1(n7274), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4608) );
  NAND2_X1 U5693 ( .A1(n7275), .A2(n7276), .ZN(n7333) );
  NOR2_X1 U5694 ( .A1(n7665), .A2(n4516), .ZN(n7667) );
  NAND2_X1 U5695 ( .A1(n7667), .A2(n7668), .ZN(n7917) );
  NOR2_X1 U5696 ( .A1(n9522), .A2(n9521), .ZN(n9526) );
  OAI21_X1 U5697 ( .B1(n9535), .B2(n4603), .A(n4600), .ZN(n9573) );
  AOI21_X1 U5698 ( .B1(n4602), .B2(n4601), .A(n4523), .ZN(n4600) );
  NOR2_X1 U5699 ( .A1(n5012), .A2(n9354), .ZN(n9591) );
  AND2_X1 U5700 ( .A1(n6752), .A2(n7064), .ZN(n9604) );
  AND2_X1 U5701 ( .A1(n9328), .A2(n9598), .ZN(n9317) );
  NOR2_X1 U5702 ( .A1(n6931), .A2(n6386), .ZN(n6396) );
  OR2_X1 U5703 ( .A1(n9644), .A2(n9643), .ZN(n4755) );
  OAI21_X1 U5704 ( .B1(n9692), .B2(n8498), .A(n9258), .ZN(n9665) );
  INV_X1 U5705 ( .A(n4944), .ZN(n4943) );
  AOI21_X1 U5706 ( .B1(n4944), .B2(n4942), .A(n4457), .ZN(n4941) );
  INV_X1 U5707 ( .A(n8512), .ZN(n4942) );
  AND2_X1 U5708 ( .A1(n9677), .A2(n9688), .ZN(n9673) );
  NAND2_X1 U5709 ( .A1(n4621), .A2(n9338), .ZN(n9693) );
  NOR2_X1 U5710 ( .A1(n9693), .A2(n9694), .ZN(n9692) );
  NOR2_X1 U5711 ( .A1(n9790), .A2(n9701), .ZN(n9688) );
  OR2_X1 U5712 ( .A1(n4953), .A2(n4458), .ZN(n4951) );
  NAND2_X1 U5713 ( .A1(n4622), .A2(n4623), .ZN(n9724) );
  NAND2_X1 U5714 ( .A1(n8170), .A2(n4442), .ZN(n9719) );
  NAND2_X1 U5715 ( .A1(n8170), .A2(n4670), .ZN(n9735) );
  AND2_X1 U5716 ( .A1(n9091), .A2(n6272), .ZN(n6289) );
  OAI21_X1 U5717 ( .B1(n8084), .B2(n4740), .A(n4737), .ZN(n8495) );
  AND2_X1 U5718 ( .A1(n8093), .A2(n9853), .ZN(n8170) );
  NAND2_X1 U5719 ( .A1(n8170), .A2(n9846), .ZN(n8209) );
  NOR2_X1 U5720 ( .A1(n6239), .A2(n9502), .ZN(n6241) );
  AND2_X1 U5721 ( .A1(n6241), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9091) );
  NAND2_X1 U5722 ( .A1(n8084), .A2(n9225), .ZN(n8085) );
  OAI21_X1 U5723 ( .B1(n8090), .B2(n9440), .A(n8089), .ZN(n8091) );
  AND2_X1 U5724 ( .A1(n9380), .A2(n9383), .ZN(n9308) );
  OR2_X1 U5725 ( .A1(n10000), .A2(n9361), .ZN(n7107) );
  NOR2_X1 U5726 ( .A1(n9906), .A2(n8045), .ZN(n8051) );
  AOI21_X1 U5727 ( .B1(n9895), .B2(n7879), .A(n9220), .ZN(n7880) );
  NOR2_X1 U5728 ( .A1(n9896), .A2(n9212), .ZN(n7879) );
  AND2_X1 U5729 ( .A1(n9224), .A2(n9219), .ZN(n9306) );
  NAND2_X1 U5730 ( .A1(n9213), .A2(n9222), .ZN(n9896) );
  NAND2_X1 U5731 ( .A1(n4662), .A2(n4627), .ZN(n9906) );
  OR2_X1 U5732 ( .A1(n6188), .A2(n8020), .ZN(n6205) );
  NAND2_X1 U5733 ( .A1(n6171), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6188) );
  INV_X1 U5734 ( .A(n9896), .ZN(n9902) );
  NAND2_X1 U5735 ( .A1(n4724), .A2(n5002), .ZN(n9369) );
  AND2_X1 U5736 ( .A1(n7491), .A2(n10068), .ZN(n9921) );
  INV_X1 U5737 ( .A(n4935), .ZN(n4934) );
  OAI21_X1 U5738 ( .B1(n7497), .B2(n4938), .A(n4937), .ZN(n4935) );
  NOR2_X1 U5739 ( .A1(n7682), .A2(n10058), .ZN(n7491) );
  NAND2_X1 U5740 ( .A1(n4665), .A2(n4664), .ZN(n7682) );
  NOR2_X1 U5741 ( .A1(n4666), .A2(n7866), .ZN(n4664) );
  NAND2_X1 U5742 ( .A1(n4665), .A2(n4663), .ZN(n9936) );
  INV_X1 U5743 ( .A(n4666), .ZN(n4663) );
  NOR2_X1 U5744 ( .A1(n6068), .A2(n7545), .ZN(n6101) );
  NAND2_X1 U5745 ( .A1(n6051), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6068) );
  NOR2_X1 U5746 ( .A1(n9951), .A2(n4668), .ZN(n9937) );
  NAND2_X1 U5747 ( .A1(n4747), .A2(n9365), .ZN(n7599) );
  NAND2_X1 U5748 ( .A1(n9183), .A2(n4745), .ZN(n4747) );
  NOR2_X1 U5749 ( .A1(n9192), .A2(n4746), .ZN(n4745) );
  INV_X1 U5750 ( .A(n9185), .ZN(n4746) );
  NOR2_X1 U5751 ( .A1(n9951), .A2(n9948), .ZN(n9952) );
  AND2_X1 U5752 ( .A1(n6028), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6051) );
  NAND2_X1 U5753 ( .A1(n9184), .A2(n9365), .ZN(n9950) );
  OR2_X1 U5754 ( .A1(n5979), .A2(n8490), .ZN(n6005) );
  NOR2_X1 U5755 ( .A1(n7442), .A2(n9984), .ZN(n9965) );
  NAND2_X1 U5756 ( .A1(n9976), .A2(n9974), .ZN(n7458) );
  NAND2_X1 U5757 ( .A1(n7439), .A2(n9986), .ZN(n9984) );
  NAND2_X1 U5758 ( .A1(n6410), .A2(n6409), .ZN(n9766) );
  NAND2_X1 U5759 ( .A1(n8126), .A2(n9176), .ZN(n6410) );
  INV_X1 U5760 ( .A(n7480), .ZN(n10068) );
  NOR2_X1 U5761 ( .A1(n4744), .A2(n5917), .ZN(n4743) );
  NAND2_X1 U5762 ( .A1(n5010), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n5917) );
  INV_X1 U5763 ( .A(n5910), .ZN(n4744) );
  INV_X1 U5764 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5920) );
  XNOR2_X1 U5765 ( .A(n5391), .B(n5390), .ZN(n7312) );
  XNOR2_X1 U5766 ( .A(n4630), .B(n5373), .ZN(n7138) );
  XNOR2_X1 U5767 ( .A(n5206), .B(SI_4_), .ZN(n5205) );
  NAND2_X1 U5768 ( .A1(n5188), .A2(SI_3_), .ZN(n5212) );
  XNOR2_X1 U5769 ( .A(n5161), .B(SI_2_), .ZN(n5160) );
  AND4_X1 U5770 ( .A1(n5338), .A2(n5337), .A3(n5336), .A4(n5335), .ZN(n7951)
         );
  NAND2_X1 U5771 ( .A1(n8555), .A2(n8554), .ZN(n8553) );
  NAND2_X1 U5772 ( .A1(n4927), .A2(n4925), .ZN(n8580) );
  NAND2_X1 U5773 ( .A1(n8617), .A2(n5790), .ZN(n7934) );
  NAND2_X1 U5774 ( .A1(n4927), .A2(n5811), .ZN(n8528) );
  NAND2_X1 U5775 ( .A1(n4912), .A2(n4911), .ZN(n8030) );
  OR2_X1 U5776 ( .A1(n4915), .A2(n4914), .ZN(n4911) );
  AND2_X1 U5777 ( .A1(n5790), .A2(n4916), .ZN(n4915) );
  NAND2_X1 U5778 ( .A1(n4921), .A2(n4924), .ZN(n8607) );
  NAND2_X1 U5779 ( .A1(n8569), .A2(n4925), .ZN(n4921) );
  NAND2_X1 U5780 ( .A1(n5332), .A2(n5331), .ZN(n8624) );
  NAND2_X1 U5781 ( .A1(n5761), .A2(n5760), .ZN(n7357) );
  OAI21_X1 U5782 ( .B1(n8225), .B2(n5805), .A(n5804), .ZN(n8630) );
  OR2_X1 U5783 ( .A1(n5849), .A2(n5848), .ZN(n8645) );
  INV_X1 U5784 ( .A(n5831), .ZN(n5830) );
  INV_X1 U5785 ( .A(n8149), .ZN(n5797) );
  NAND2_X1 U5786 ( .A1(n5796), .A2(n5795), .ZN(n8150) );
  INV_X1 U5787 ( .A(n8797), .ZN(n8656) );
  OAI211_X1 U5788 ( .C1(n4529), .C2(n8799), .A(n5566), .B(n5565), .ZN(n8808)
         );
  INV_X1 U5789 ( .A(n8835), .ZN(n8807) );
  INV_X1 U5790 ( .A(n8621), .ZN(n8660) );
  INV_X1 U5791 ( .A(n4766), .ZN(n7187) );
  INV_X1 U5792 ( .A(n4775), .ZN(n8476) );
  NOR2_X1 U5793 ( .A1(n7525), .A2(n10254), .ZN(n7524) );
  NAND2_X1 U5794 ( .A1(n6546), .A2(n4857), .ZN(n4855) );
  INV_X1 U5795 ( .A(n4865), .ZN(n7997) );
  NAND2_X1 U5796 ( .A1(n4863), .A2(n4862), .ZN(n8132) );
  INV_X1 U5797 ( .A(n4852), .ZN(n10146) );
  NAND2_X1 U5798 ( .A1(n4779), .A2(n4782), .ZN(n10142) );
  INV_X1 U5799 ( .A(n6597), .ZN(n4783) );
  NOR2_X1 U5800 ( .A1(n8674), .A2(n8673), .ZN(n8672) );
  NAND2_X1 U5801 ( .A1(n8377), .A2(n8376), .ZN(n8751) );
  XNOR2_X1 U5802 ( .A(n8446), .B(n8439), .ZN(n8761) );
  NAND2_X1 U5803 ( .A1(n4844), .A2(n4555), .ZN(n8755) );
  OR2_X1 U5804 ( .A1(n8761), .A2(n7777), .ZN(n4555) );
  OAI21_X1 U5805 ( .B1(n5710), .B2(n8352), .A(n8357), .ZN(n5731) );
  NAND2_X1 U5806 ( .A1(n4804), .A2(n4808), .ZN(n5733) );
  NAND2_X1 U5807 ( .A1(n5710), .A2(n8357), .ZN(n4804) );
  NAND2_X1 U5808 ( .A1(n8126), .A2(n8396), .ZN(n5685) );
  NAND2_X1 U5809 ( .A1(n5523), .A2(n5522), .ZN(n8826) );
  AND2_X1 U5810 ( .A1(n8843), .A2(n8334), .ZN(n8829) );
  NAND2_X1 U5811 ( .A1(n4886), .A2(n4888), .ZN(n8832) );
  NAND2_X1 U5812 ( .A1(n5466), .A2(n5465), .ZN(n8863) );
  NAND2_X1 U5813 ( .A1(n5347), .A2(n5346), .ZN(n10232) );
  NAND2_X1 U5814 ( .A1(n4836), .A2(n4837), .ZN(n7903) );
  NAND2_X1 U5815 ( .A1(n7730), .A2(n4839), .ZN(n4836) );
  OAI21_X1 U5816 ( .B1(n7730), .B2(n8281), .A(n8292), .ZN(n7776) );
  NAND2_X1 U5817 ( .A1(n7717), .A2(n7720), .ZN(n7757) );
  NAND2_X1 U5818 ( .A1(n4819), .A2(n8272), .ZN(n7756) );
  NAND2_X1 U5819 ( .A1(n7716), .A2(n8265), .ZN(n4819) );
  INV_X1 U5820 ( .A(n5153), .ZN(n10182) );
  NAND2_X1 U5821 ( .A1(n4547), .A2(n5137), .ZN(n10168) );
  OR2_X1 U5822 ( .A1(n5134), .A2(n6564), .ZN(n4896) );
  INV_X1 U5823 ( .A(n10165), .ZN(n8897) );
  NAND2_X1 U5824 ( .A1(n8398), .A2(n8397), .ZN(n8946) );
  INV_X1 U5825 ( .A(n8751), .ZN(n8952) );
  INV_X1 U5826 ( .A(n8378), .ZN(n6700) );
  AND2_X1 U5827 ( .A1(n5592), .A2(n5591), .ZN(n8960) );
  OAI21_X1 U5828 ( .B1(n5550), .B2(n4880), .A(n4878), .ZN(n8772) );
  NAND2_X1 U5829 ( .A1(n4822), .A2(n4823), .ZN(n8770) );
  NAND2_X1 U5830 ( .A1(n5576), .A2(n5575), .ZN(n8966) );
  NAND2_X1 U5831 ( .A1(n4825), .A2(n8404), .ZN(n8779) );
  NAND2_X1 U5832 ( .A1(n4827), .A2(n4826), .ZN(n4825) );
  INV_X1 U5833 ( .A(n8793), .ZN(n4827) );
  NAND2_X1 U5834 ( .A1(n5542), .A2(n5541), .ZN(n8977) );
  NAND2_X1 U5835 ( .A1(n8843), .A2(n4830), .ZN(n8815) );
  NAND2_X1 U5836 ( .A1(n5495), .A2(n5494), .ZN(n8993) );
  INV_X1 U5837 ( .A(n4887), .ZN(n8847) );
  AOI21_X1 U5838 ( .B1(n5466), .B2(n4891), .A(n4890), .ZN(n4887) );
  NAND2_X1 U5839 ( .A1(n5420), .A2(n5419), .ZN(n9010) );
  NAND2_X1 U5840 ( .A1(n5655), .A2(n8317), .ZN(n8118) );
  NAND2_X1 U5841 ( .A1(n5379), .A2(n5378), .ZN(n8114) );
  AND3_X1 U5842 ( .A1(n5172), .A2(n5171), .A3(n5170), .ZN(n7869) );
  NAND2_X1 U5843 ( .A1(n9019), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5098) );
  NAND2_X1 U5844 ( .A1(n5087), .A2(n5086), .ZN(n7983) );
  NOR2_X1 U5845 ( .A1(n5326), .A2(n5053), .ZN(n5368) );
  INV_X1 U5846 ( .A(n6064), .ZN(n4969) );
  AND2_X1 U5847 ( .A1(n6204), .A2(n6203), .ZN(n10092) );
  OR2_X1 U5848 ( .A1(n6678), .A2(n6677), .ZN(n6427) );
  OAI21_X1 U5849 ( .B1(n9051), .B2(n4984), .A(n4982), .ZN(n9056) );
  NAND2_X1 U5850 ( .A1(n6169), .A2(n6168), .ZN(n7947) );
  NAND2_X1 U5851 ( .A1(n4989), .A2(n6249), .ZN(n4988) );
  NAND2_X1 U5852 ( .A1(n4999), .A2(n4996), .ZN(n4995) );
  NAND2_X1 U5853 ( .A1(n4999), .A2(n4470), .ZN(n4997) );
  INV_X1 U5854 ( .A(n7284), .ZN(n6022) );
  NAND2_X1 U5855 ( .A1(n5000), .A2(n5999), .ZN(n7285) );
  NAND2_X1 U5856 ( .A1(n4987), .A2(n6300), .ZN(n9113) );
  NAND2_X1 U5857 ( .A1(n9051), .A2(n9050), .ZN(n4987) );
  NAND2_X1 U5858 ( .A1(n7940), .A2(n7941), .ZN(n4973) );
  AND2_X1 U5859 ( .A1(n9089), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9158) );
  INV_X1 U5860 ( .A(n6676), .ZN(n9151) );
  AND2_X1 U5861 ( .A1(n6479), .A2(n6468), .ZN(n9150) );
  INV_X1 U5862 ( .A(n9150), .ZN(n9174) );
  INV_X1 U5863 ( .A(n9161), .ZN(n9171) );
  NAND2_X1 U5864 ( .A1(n4570), .A2(n4472), .ZN(n4569) );
  INV_X1 U5865 ( .A(n4947), .ZN(n4946) );
  OAI211_X1 U5866 ( .C1(n9284), .C2(n10103), .A(n6010), .B(n4948), .ZN(n4947)
         );
  XNOR2_X1 U5867 ( .A(n5912), .B(P1_IR_REG_1__SCAN_IN), .ZN(n9884) );
  INV_X1 U5868 ( .A(n4607), .ZN(n9466) );
  NOR2_X1 U5869 ( .A1(n7204), .A2(n4508), .ZN(n7208) );
  NOR2_X1 U5870 ( .A1(n7208), .A2(n7207), .ZN(n7273) );
  NAND2_X1 U5871 ( .A1(n9553), .A2(n4602), .ZN(n9571) );
  AND2_X1 U5872 ( .A1(n9553), .A2(n9552), .ZN(n9558) );
  AND2_X1 U5873 ( .A1(n9612), .A2(n5012), .ZN(n9753) );
  AND2_X1 U5874 ( .A1(n4757), .A2(n4756), .ZN(n9756) );
  AOI22_X1 U5875 ( .A1(n9605), .A2(n9604), .B1(n9602), .B2(n9603), .ZN(n4756)
         );
  NAND2_X1 U5876 ( .A1(n4758), .A2(n9980), .ZN(n4757) );
  XNOR2_X1 U5877 ( .A(n9600), .B(n9609), .ZN(n4758) );
  NAND2_X1 U5878 ( .A1(n4750), .A2(n4751), .ZN(n9622) );
  OR2_X1 U5879 ( .A1(n9644), .A2(n4752), .ZN(n4750) );
  INV_X1 U5880 ( .A(n9785), .ZN(n9677) );
  OAI21_X1 U5881 ( .B1(n9687), .B2(n8513), .A(n8512), .ZN(n9672) );
  OAI21_X1 U5882 ( .B1(n8505), .B2(n4953), .A(n4952), .ZN(n9718) );
  NAND2_X1 U5883 ( .A1(n4625), .A2(n9244), .ZN(n9730) );
  NAND2_X1 U5884 ( .A1(n4736), .A2(n4435), .ZN(n4625) );
  OR2_X1 U5885 ( .A1(n8505), .A2(n4956), .ZN(n4955) );
  INV_X1 U5886 ( .A(n4958), .ZN(n9850) );
  NAND2_X1 U5887 ( .A1(n6224), .A2(n6223), .ZN(n9083) );
  INV_X1 U5888 ( .A(n9859), .ZN(n9172) );
  NAND2_X1 U5889 ( .A1(n4722), .A2(n9206), .ZN(n9914) );
  NAND2_X1 U5890 ( .A1(n6127), .A2(n6126), .ZN(n9920) );
  OR2_X1 U5891 ( .A1(n9992), .A2(n7483), .ZN(n9741) );
  AOI21_X1 U5892 ( .B1(n7674), .B2(n7676), .A(n5008), .ZN(n7489) );
  NAND2_X1 U5893 ( .A1(n7592), .A2(n7445), .ZN(n9957) );
  INV_X1 U5894 ( .A(n7439), .ZN(n9982) );
  NAND2_X1 U5895 ( .A1(n9758), .A2(n10095), .ZN(n9763) );
  NOR3_X1 U5896 ( .A1(n9769), .A2(n9770), .A3(n4628), .ZN(n9772) );
  AND2_X1 U5897 ( .A1(n9771), .A2(n10059), .ZN(n4628) );
  INV_X1 U5898 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5921) );
  NAND2_X1 U5899 ( .A1(n5911), .A2(n5910), .ZN(n5918) );
  NOR2_X1 U5900 ( .A1(n5894), .A2(n5893), .ZN(n5901) );
  INV_X1 U5901 ( .A(n4686), .ZN(n5559) );
  AOI21_X1 U5902 ( .B1(n4693), .B2(n4687), .A(n4690), .ZN(n4686) );
  NAND2_X1 U5903 ( .A1(n6269), .A2(n5880), .ZN(n5878) );
  AND2_X1 U5904 ( .A1(n4617), .A2(n4614), .ZN(n5291) );
  INV_X1 U5905 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6964) );
  NAND2_X1 U5906 ( .A1(n4682), .A2(n5253), .ZN(n5268) );
  NAND2_X1 U5907 ( .A1(n5250), .A2(n5249), .ZN(n4682) );
  INV_X1 U5908 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n8492) );
  INV_X1 U5909 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6711) );
  INV_X1 U5910 ( .A(n7035), .ZN(n7054) );
  NAND2_X1 U5911 ( .A1(n7388), .A2(n5766), .ZN(n7322) );
  INV_X1 U5912 ( .A(n4787), .ZN(n4786) );
  AOI21_X1 U5913 ( .B1(n5716), .B2(n5715), .A(n5714), .ZN(n5717) );
  NAND2_X1 U5914 ( .A1(n5713), .A2(n5003), .ZN(n5714) );
  NAND2_X1 U5915 ( .A1(n5673), .A2(n4467), .ZN(P2_U3207) );
  NOR2_X1 U5916 ( .A1(n6519), .A2(n6521), .ZN(n6522) );
  NOR2_X1 U5917 ( .A1(n10238), .A2(n6520), .ZN(n6521) );
  INV_X1 U5918 ( .A(n4605), .ZN(n7076) );
  AND2_X1 U5919 ( .A1(n4551), .A2(n4550), .ZN(n4430) );
  INV_X2 U5920 ( .A(n5937), .ZN(n6093) );
  INV_X1 U5921 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5148) );
  AND4_X1 U5922 ( .A1(n5314), .A2(n5313), .A3(n5312), .A4(n5311), .ZN(n8620)
         );
  AND2_X1 U5923 ( .A1(n5102), .A2(n5103), .ZN(n5176) );
  AND2_X1 U5924 ( .A1(n8518), .A2(n8517), .ZN(n4431) );
  NAND2_X1 U5925 ( .A1(n9211), .A2(n9210), .ZN(n4432) );
  NAND2_X1 U5926 ( .A1(n9806), .A2(n9436), .ZN(n4433) );
  NOR2_X1 U5927 ( .A1(n5603), .A2(n8783), .ZN(n4434) );
  AND2_X1 U5928 ( .A1(n8494), .A2(n4735), .ZN(n4435) );
  INV_X1 U5929 ( .A(n9643), .ZN(n4753) );
  AND4_X1 U5930 ( .A1(n5065), .A2(n5376), .A3(n5064), .A4(n5070), .ZN(n4436)
         );
  OR2_X1 U5931 ( .A1(n8670), .A2(n5153), .ZN(n4437) );
  OR2_X1 U5932 ( .A1(n8234), .A2(n8399), .ZN(n4438) );
  AND2_X1 U5933 ( .A1(n4561), .A2(n4560), .ZN(n4439) );
  NAND2_X1 U5934 ( .A1(n5909), .A2(n5908), .ZN(n4440) );
  OR2_X1 U5935 ( .A1(n4894), .A2(n7952), .ZN(n4441) );
  AND2_X1 U5936 ( .A1(n4670), .A2(n4669), .ZN(n4442) );
  AND2_X1 U5937 ( .A1(n9780), .A2(n9432), .ZN(n4443) );
  INV_X1 U5938 ( .A(n7782), .ZN(n10215) );
  AND2_X1 U5939 ( .A1(n5300), .A2(n5299), .ZN(n7782) );
  AND2_X1 U5940 ( .A1(n9336), .A2(n9632), .ZN(n4444) );
  NOR2_X1 U5941 ( .A1(n6064), .A2(n4514), .ZN(n4446) );
  AND2_X1 U5942 ( .A1(n6288), .A2(n6287), .ZN(n9742) );
  INV_X1 U5943 ( .A(n9742), .ZN(n9806) );
  AND2_X1 U5944 ( .A1(n5095), .A2(n4644), .ZN(n4447) );
  OR2_X1 U5945 ( .A1(n5534), .A2(SI_21_), .ZN(n4448) );
  AND2_X1 U5946 ( .A1(n4865), .A2(n6550), .ZN(n4449) );
  AND2_X1 U5947 ( .A1(n4866), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4450) );
  NAND2_X1 U5948 ( .A1(n6187), .A2(n6186), .ZN(n9905) );
  INV_X1 U5949 ( .A(n9905), .ZN(n4627) );
  INV_X1 U5950 ( .A(n8414), .ZN(n4820) );
  AND2_X1 U5951 ( .A1(n4785), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4451) );
  INV_X1 U5952 ( .A(n7777), .ZN(n4842) );
  INV_X1 U5953 ( .A(n5179), .ZN(n5699) );
  AND2_X1 U5954 ( .A1(n5101), .A2(n5103), .ZN(n5179) );
  NAND2_X2 U5955 ( .A1(n5960), .A2(n8392), .ZN(n6003) );
  NOR2_X1 U5956 ( .A1(n6044), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n6046) );
  OR2_X1 U5957 ( .A1(n9776), .A2(n9104), .ZN(n9336) );
  OAI211_X2 U5958 ( .C1(n6753), .C2(n7054), .A(n5962), .B(n5961), .ZN(n7442)
         );
  NOR2_X1 U5959 ( .A1(n8528), .A2(n8529), .ZN(n4452) );
  OR2_X1 U5960 ( .A1(n9780), .A2(n9432), .ZN(n4453) );
  INV_X1 U5961 ( .A(n9621), .ZN(n9619) );
  AND2_X1 U5962 ( .A1(n9331), .A2(n9267), .ZN(n9621) );
  INV_X1 U5963 ( .A(n4705), .ZN(n4704) );
  NAND2_X1 U5964 ( .A1(n4706), .A2(n5374), .ZN(n4705) );
  AND2_X1 U5965 ( .A1(n9659), .A2(n4675), .ZN(n4454) );
  INV_X2 U5966 ( .A(n5134), .ZN(n5169) );
  AND2_X1 U5967 ( .A1(n5697), .A2(n5696), .ZN(n6509) );
  NAND2_X1 U5968 ( .A1(n6271), .A2(n6270), .ZN(n9810) );
  OR2_X1 U5969 ( .A1(n9810), .A2(n9437), .ZN(n4455) );
  NOR2_X1 U5970 ( .A1(n5235), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5255) );
  INV_X1 U5971 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9020) );
  AND2_X1 U5972 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4456) );
  NAND2_X1 U5973 ( .A1(n6257), .A2(n6256), .ZN(n9097) );
  INV_X1 U5974 ( .A(n9206), .ZN(n4580) );
  INV_X1 U5975 ( .A(n8271), .ZN(n4818) );
  OAI21_X1 U5976 ( .B1(n9687), .B2(n4943), .A(n4941), .ZN(n9658) );
  INV_X1 U5977 ( .A(n9666), .ZN(n4593) );
  INV_X1 U5978 ( .A(n8276), .ZN(n4815) );
  NAND2_X1 U5979 ( .A1(n5341), .A2(n5325), .ZN(n5342) );
  INV_X1 U5980 ( .A(n8418), .ZN(n4835) );
  AND2_X1 U5981 ( .A1(n9677), .A2(n9129), .ZN(n4457) );
  NAND2_X1 U5982 ( .A1(n8538), .A2(n8537), .ZN(n9354) );
  INV_X1 U5983 ( .A(n9354), .ZN(n9751) );
  AND2_X1 U5984 ( .A1(n9329), .A2(n9402), .ZN(n9609) );
  INV_X1 U5985 ( .A(n9341), .ZN(n4734) );
  AND2_X1 U5986 ( .A1(n9800), .A2(n9435), .ZN(n4458) );
  AND2_X1 U5987 ( .A1(n4925), .A2(n5821), .ZN(n4459) );
  OR3_X1 U5988 ( .A1(n8387), .A2(n8441), .A3(n8453), .ZN(n4460) );
  INV_X1 U5989 ( .A(n8352), .ZN(n4810) );
  OR2_X1 U5990 ( .A1(n9800), .A2(n9435), .ZN(n4461) );
  AND4_X1 U5991 ( .A1(n5063), .A2(n5062), .A3(n5061), .A4(n5328), .ZN(n4462)
         );
  AND2_X1 U5992 ( .A1(n8960), .A2(n8783), .ZN(n8236) );
  NOR2_X1 U5993 ( .A1(n8855), .A2(n8862), .ZN(n4463) );
  AND3_X1 U5994 ( .A1(n5920), .A2(n5919), .A3(n5915), .ZN(n4464) );
  INV_X1 U5995 ( .A(n6249), .ZN(n4992) );
  INV_X1 U5996 ( .A(n4875), .ZN(n4542) );
  AOI21_X1 U5997 ( .B1(n4878), .B2(n4880), .A(n4876), .ZN(n4875) );
  NOR2_X1 U5998 ( .A1(n6602), .A2(n8672), .ZN(n4465) );
  NOR2_X1 U5999 ( .A1(n8844), .A2(n4890), .ZN(n4466) );
  AND2_X1 U6000 ( .A1(n5672), .A2(n5671), .ZN(n4467) );
  INV_X1 U6001 ( .A(n9394), .ZN(n4731) );
  AND2_X1 U6002 ( .A1(n7164), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4468) );
  INV_X1 U6003 ( .A(n9759), .ZN(n9607) );
  NAND2_X1 U6004 ( .A1(n6429), .A2(n6428), .ZN(n9759) );
  AND2_X1 U6005 ( .A1(n9248), .A2(n9247), .ZN(n4469) );
  AND2_X1 U6006 ( .A1(n9040), .A2(n4998), .ZN(n4470) );
  NOR2_X1 U6007 ( .A1(n8402), .A2(n8405), .ZN(n4824) );
  AND2_X1 U6008 ( .A1(n8442), .A2(n5019), .ZN(n4471) );
  INV_X1 U6009 ( .A(n4840), .ZN(n4839) );
  OR2_X1 U6010 ( .A1(n8283), .A2(n8282), .ZN(n4840) );
  AND2_X1 U6011 ( .A1(n9408), .A2(n9355), .ZN(n4472) );
  OR2_X1 U6012 ( .A1(n5326), .A2(n4792), .ZN(n4473) );
  NOR2_X1 U6013 ( .A1(n8955), .A2(n4713), .ZN(n4474) );
  AND2_X1 U6014 ( .A1(n8971), .A2(n8808), .ZN(n8406) );
  INV_X1 U6015 ( .A(n8406), .ZN(n4826) );
  AND2_X1 U6016 ( .A1(n6200), .A2(n6199), .ZN(n4475) );
  AND2_X1 U6017 ( .A1(n6385), .A2(n6384), .ZN(n9655) );
  OR2_X1 U6018 ( .A1(n8966), .A2(n8797), .ZN(n8401) );
  OR2_X1 U6019 ( .A1(n4891), .A2(n4890), .ZN(n4476) );
  NOR2_X1 U6020 ( .A1(n8721), .A2(n4788), .ZN(n4477) );
  NOR2_X1 U6021 ( .A1(n9607), .A2(n9606), .ZN(n4478) );
  AND2_X1 U6022 ( .A1(n8318), .A2(n8874), .ZN(n4479) );
  NAND2_X1 U6023 ( .A1(n8459), .A2(n8458), .ZN(n4480) );
  OR2_X1 U6024 ( .A1(n6614), .A2(n6559), .ZN(n4481) );
  NAND2_X1 U6025 ( .A1(n5077), .A2(n5081), .ZN(n4482) );
  AND2_X1 U6026 ( .A1(n9209), .A2(n9208), .ZN(n4483) );
  AND2_X1 U6027 ( .A1(n8337), .A2(n4828), .ZN(n4484) );
  NOR2_X1 U6028 ( .A1(n8765), .A2(n8646), .ZN(n4485) );
  AND2_X1 U6029 ( .A1(n4899), .A2(n4902), .ZN(n4486) );
  INV_X1 U6030 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6866) );
  NAND2_X1 U6031 ( .A1(n8608), .A2(n8821), .ZN(n4487) );
  AND2_X1 U6032 ( .A1(n8334), .A2(n8332), .ZN(n8844) );
  NAND2_X1 U6033 ( .A1(n8580), .A2(n8579), .ZN(n4488) );
  OR2_X1 U6034 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n4489) );
  AND2_X1 U6035 ( .A1(n4950), .A2(n4461), .ZN(n4490) );
  AND2_X1 U6036 ( .A1(n6314), .A2(n6313), .ZN(n4491) );
  NAND2_X1 U6037 ( .A1(n5819), .A2(n8579), .ZN(n4492) );
  AND2_X1 U6038 ( .A1(n4943), .A2(n4453), .ZN(n4493) );
  INV_X1 U6039 ( .A(n4834), .ZN(n4833) );
  NAND2_X1 U6040 ( .A1(n4837), .A2(n4835), .ZN(n4834) );
  AND2_X1 U6041 ( .A1(n8114), .A2(n8659), .ZN(n4494) );
  INV_X1 U6042 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5888) );
  NAND2_X1 U6043 ( .A1(n6700), .A2(n8654), .ZN(n4495) );
  NAND2_X1 U6044 ( .A1(n5441), .A2(n5443), .ZN(n4496) );
  INV_X1 U6045 ( .A(n4808), .ZN(n4807) );
  AND2_X1 U6046 ( .A1(n4809), .A2(n8434), .ZN(n4808) );
  OAI21_X1 U6047 ( .B1(n4435), .B2(n9245), .A(n9731), .ZN(n4626) );
  AND2_X1 U6048 ( .A1(n8955), .A2(n4713), .ZN(n4497) );
  NAND2_X1 U6049 ( .A1(n4455), .A2(n8508), .ZN(n4498) );
  NAND2_X1 U6050 ( .A1(n5550), .A2(n5549), .ZN(n8794) );
  AND2_X1 U6051 ( .A1(n4941), .A2(n4453), .ZN(n4499) );
  AND2_X1 U6052 ( .A1(n4955), .A2(n4455), .ZN(n4500) );
  NAND2_X1 U6053 ( .A1(n5289), .A2(n5275), .ZN(n5290) );
  INV_X1 U6054 ( .A(n5290), .ZN(n4616) );
  NOR2_X1 U6055 ( .A1(n7411), .A2(n5778), .ZN(n4501) );
  INV_X1 U6056 ( .A(n9197), .ZN(n4720) );
  OR2_X1 U6057 ( .A1(n9083), .A2(n8169), .ZN(n9380) );
  AND2_X1 U6058 ( .A1(n4962), .A2(n4464), .ZN(n4502) );
  NAND2_X1 U6059 ( .A1(n8259), .A2(n8258), .ZN(n8255) );
  INV_X1 U6060 ( .A(n8255), .ZN(n4543) );
  AND2_X1 U6061 ( .A1(n9771), .A2(n9261), .ZN(n9394) );
  AND2_X1 U6062 ( .A1(n5276), .A2(n4931), .ZN(n4503) );
  AND2_X1 U6063 ( .A1(n4818), .A2(n8272), .ZN(n4817) );
  AND2_X1 U6064 ( .A1(n5797), .A2(n5795), .ZN(n4504) );
  AND2_X1 U6065 ( .A1(n6022), .A2(n5999), .ZN(n4505) );
  AND2_X1 U6066 ( .A1(n4999), .A2(n9040), .ZN(n4506) );
  AND2_X1 U6067 ( .A1(n7446), .A2(n4575), .ZN(n4507) );
  XNOR2_X1 U6068 ( .A(n5060), .B(n5064), .ZN(n7409) );
  AND2_X1 U6069 ( .A1(n4966), .A2(n4963), .ZN(n7858) );
  NAND2_X1 U6070 ( .A1(n9027), .A2(n6216), .ZN(n9072) );
  NAND2_X1 U6071 ( .A1(n8085), .A2(n9308), .ZN(n8165) );
  INV_X1 U6072 ( .A(n5753), .ZN(n5750) );
  NAND2_X1 U6073 ( .A1(n4722), .A2(n4721), .ZN(n7645) );
  INV_X1 U6074 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4762) );
  OAI21_X1 U6075 ( .B1(n7974), .B2(n8314), .A(n7973), .ZN(n8106) );
  AND2_X1 U6076 ( .A1(n7205), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4508) );
  NAND2_X1 U6077 ( .A1(n5429), .A2(n5428), .ZN(n8877) );
  NAND2_X1 U6078 ( .A1(n4973), .A2(n6183), .ZN(n8018) );
  INV_X1 U6079 ( .A(n5305), .ZN(n5077) );
  NAND2_X1 U6080 ( .A1(n4759), .A2(n6593), .ZN(n7988) );
  INV_X1 U6081 ( .A(n7699), .ZN(n4857) );
  INV_X1 U6082 ( .A(n10133), .ZN(n4860) );
  OR2_X1 U6083 ( .A1(n5326), .A2(n4919), .ZN(n4509) );
  NAND2_X1 U6084 ( .A1(n8170), .A2(n4671), .ZN(n4672) );
  OR3_X1 U6085 ( .A1(n5326), .A2(n4919), .A3(n5055), .ZN(n4510) );
  AND2_X1 U6086 ( .A1(n4784), .A2(n4783), .ZN(n4511) );
  NAND2_X1 U6087 ( .A1(n6548), .A2(n7073), .ZN(n6550) );
  NOR2_X1 U6088 ( .A1(n9190), .A2(n9197), .ZN(n4512) );
  INV_X1 U6089 ( .A(n5551), .ZN(n4690) );
  NAND2_X1 U6090 ( .A1(n5774), .A2(n4898), .ZN(n4906) );
  INV_X1 U6091 ( .A(n10176), .ZN(n10174) );
  INV_X1 U6092 ( .A(n8895), .ZN(n10176) );
  INV_X1 U6093 ( .A(n7676), .ZN(n4933) );
  NAND2_X1 U6094 ( .A1(n6302), .A2(n6301), .ZN(n9800) );
  INV_X1 U6095 ( .A(n9800), .ZN(n4669) );
  OR2_X1 U6096 ( .A1(n6622), .A2(n6552), .ZN(n4513) );
  AND2_X1 U6097 ( .A1(n6078), .A2(n6077), .ZN(n4514) );
  AND2_X1 U6098 ( .A1(n7565), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4515) );
  INV_X1 U6099 ( .A(n5155), .ZN(n5310) );
  AND2_X1 U6100 ( .A1(n7666), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4516) );
  NOR2_X1 U6101 ( .A1(n7524), .A2(n6546), .ZN(n4517) );
  NOR2_X1 U6102 ( .A1(n7238), .A2(n6579), .ZN(n4518) );
  NOR2_X1 U6103 ( .A1(n7241), .A2(n5014), .ZN(n4519) );
  AND2_X1 U6104 ( .A1(n10161), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4520) );
  INV_X1 U6105 ( .A(n4662), .ZN(n9904) );
  NOR2_X1 U6106 ( .A1(n7651), .A2(n7947), .ZN(n4662) );
  INV_X1 U6107 ( .A(n4661), .ZN(n8093) );
  NAND2_X1 U6108 ( .A1(n8051), .A2(n9859), .ZN(n4661) );
  AND2_X1 U6109 ( .A1(n7369), .A2(n4969), .ZN(n4521) );
  INV_X1 U6110 ( .A(n5282), .ZN(n4895) );
  NAND2_X1 U6111 ( .A1(n10161), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4522) );
  INV_X1 U6112 ( .A(n9513), .ZN(n4609) );
  AND2_X1 U6113 ( .A1(n9575), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4523) );
  NAND2_X1 U6114 ( .A1(n5371), .A2(n5370), .ZN(n9840) );
  OR2_X1 U6115 ( .A1(n9964), .A2(n7617), .ZN(n9951) );
  INV_X1 U6116 ( .A(n9951), .ZN(n4665) );
  OR2_X1 U6117 ( .A1(n5666), .A2(n8464), .ZN(n10205) );
  INV_X1 U6118 ( .A(n4603), .ZN(n4602) );
  NAND2_X1 U6119 ( .A1(n9557), .A2(n9552), .ZN(n4603) );
  NAND2_X1 U6120 ( .A1(n7307), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4524) );
  INV_X1 U6121 ( .A(n6564), .ZN(n6707) );
  INV_X1 U6122 ( .A(n4850), .ZN(n7188) );
  OR2_X1 U6123 ( .A1(n7175), .A2(n6531), .ZN(n4850) );
  AND2_X1 U6124 ( .A1(n4766), .A2(n4767), .ZN(n4525) );
  INV_X1 U6125 ( .A(n4848), .ZN(n6535) );
  INV_X1 U6126 ( .A(n7998), .ZN(n4864) );
  OR2_X1 U6127 ( .A1(n8723), .A2(n6561), .ZN(n6562) );
  NOR2_X1 U6128 ( .A1(n7174), .A2(n10241), .ZN(n7175) );
  NAND2_X1 U6129 ( .A1(n6547), .A2(n5013), .ZN(n6548) );
  NAND2_X2 U6130 ( .A1(n9137), .A2(n6283), .ZN(n9051) );
  NAND2_X1 U6131 ( .A1(n7230), .A2(n7231), .ZN(n5000) );
  NAND2_X1 U6132 ( .A1(n4966), .A2(n4964), .ZN(n6119) );
  NAND2_X1 U6133 ( .A1(n8384), .A2(n4645), .ZN(n8366) );
  NAND2_X1 U6134 ( .A1(n8386), .A2(n4678), .ZN(n8387) );
  XNOR2_X1 U6135 ( .A(n4708), .B(n7409), .ZN(n8467) );
  NAND2_X1 U6136 ( .A1(n5367), .A2(n5365), .ZN(n4701) );
  NAND2_X1 U6137 ( .A1(n4701), .A2(n4704), .ZN(n5442) );
  NAND3_X1 U6138 ( .A1(n5210), .A2(n5213), .A3(n5209), .ZN(n5215) );
  NAND3_X1 U6139 ( .A1(n4527), .A2(n5104), .A3(n4526), .ZN(n5135) );
  NAND2_X1 U6140 ( .A1(n5155), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n4526) );
  AOI21_X1 U6141 ( .B1(n5176), .B2(P2_REG1_REG_1__SCAN_IN), .A(n4528), .ZN(
        n4527) );
  NOR2_X1 U6142 ( .A1(n4529), .A2(n7385), .ZN(n4528) );
  OAI21_X2 U6143 ( .B1(n4531), .B2(n4530), .A(n4536), .ZN(n7901) );
  INV_X1 U6144 ( .A(n4535), .ZN(n4531) );
  INV_X1 U6145 ( .A(n4541), .ZN(n5728) );
  NAND2_X1 U6146 ( .A1(n4543), .A2(n4437), .ZN(n4544) );
  NAND2_X1 U6147 ( .A1(n4545), .A2(n4544), .ZN(n7301) );
  NAND2_X1 U6148 ( .A1(n8408), .A2(n7377), .ZN(n4547) );
  NAND2_X1 U6149 ( .A1(n4928), .A2(n4929), .ZN(n5305) );
  XNOR2_X1 U6150 ( .A(n4552), .B(n4554), .ZN(n4553) );
  INV_X1 U6151 ( .A(n6517), .ZN(n4556) );
  OAI21_X2 U6152 ( .B1(n7975), .B2(n4893), .A(n4441), .ZN(n8101) );
  NAND2_X1 U6153 ( .A1(n4558), .A2(n4557), .ZN(n4559) );
  INV_X1 U6154 ( .A(n5894), .ZN(n4560) );
  INV_X1 U6155 ( .A(n6767), .ZN(n4562) );
  NOR2_X1 U6156 ( .A1(n5894), .A2(n6767), .ZN(n4567) );
  NAND4_X1 U6157 ( .A1(n4962), .A2(n4567), .A3(n4565), .A4(n4564), .ZN(n4568)
         );
  NAND2_X1 U6158 ( .A1(n4574), .A2(n4507), .ZN(n7610) );
  NAND3_X1 U6159 ( .A1(n7593), .A2(n9366), .A3(n9297), .ZN(n4574) );
  NAND2_X1 U6160 ( .A1(n4577), .A2(n4583), .ZN(n4581) );
  NAND2_X1 U6161 ( .A1(n9207), .A2(n4579), .ZN(n4577) );
  NAND2_X1 U6162 ( .A1(n4578), .A2(n4585), .ZN(n4582) );
  NAND2_X1 U6163 ( .A1(n9203), .A2(n9375), .ZN(n4578) );
  INV_X1 U6164 ( .A(n9218), .ZN(n9223) );
  NAND2_X1 U6165 ( .A1(n4582), .A2(n4581), .ZN(n9218) );
  NAND2_X1 U6166 ( .A1(n5960), .A2(n4587), .ZN(n5979) );
  XNOR2_X2 U6167 ( .A(n7440), .B(n7439), .ZN(n9976) );
  NAND3_X1 U6168 ( .A1(n4593), .A2(n9680), .A3(n9254), .ZN(n4591) );
  INV_X1 U6169 ( .A(n4596), .ZN(n4592) );
  NAND2_X1 U6170 ( .A1(n9255), .A2(n9258), .ZN(n9332) );
  OAI211_X1 U6171 ( .C1(n9253), .C2(n9252), .A(n9250), .B(n9251), .ZN(n4596)
         );
  NAND2_X1 U6172 ( .A1(n4597), .A2(n4719), .ZN(n4718) );
  NAND2_X1 U6173 ( .A1(n4598), .A2(n4720), .ZN(n4597) );
  NAND2_X1 U6174 ( .A1(n4599), .A2(n9194), .ZN(n4598) );
  NAND2_X1 U6175 ( .A1(n9187), .A2(n9191), .ZN(n4599) );
  NAND2_X1 U6176 ( .A1(n4611), .A2(n5160), .ZN(n5164) );
  XNOR2_X1 U6177 ( .A(n4611), .B(n5160), .ZN(n6710) );
  NAND2_X1 U6178 ( .A1(n4707), .A2(n5146), .ZN(n4611) );
  XNOR2_X1 U6179 ( .A(n5145), .B(n4612), .ZN(n5144) );
  NAND3_X1 U6180 ( .A1(n5232), .A2(n5253), .A3(n4618), .ZN(n4614) );
  NAND4_X1 U6181 ( .A1(n5232), .A2(n5253), .A3(n4618), .A4(n4616), .ZN(n4615)
         );
  NAND3_X1 U6182 ( .A1(n4622), .A2(n4623), .A3(n9232), .ZN(n4621) );
  NAND2_X1 U6183 ( .A1(n7138), .A2(n9176), .ZN(n6187) );
  OAI21_X1 U6184 ( .B1(n5367), .B2(n5366), .A(n5365), .ZN(n4630) );
  NAND3_X1 U6185 ( .A1(n8263), .A2(n4635), .A3(n4633), .ZN(n4632) );
  NAND2_X1 U6186 ( .A1(n4637), .A2(n8316), .ZN(n8321) );
  NAND3_X1 U6187 ( .A1(n4642), .A2(n4640), .A3(n8308), .ZN(n4639) );
  NAND2_X1 U6188 ( .A1(n5096), .A2(n4447), .ZN(n9019) );
  NAND2_X1 U6189 ( .A1(n5096), .A2(n5095), .ZN(n5099) );
  NAND3_X1 U6190 ( .A1(n8361), .A2(n8362), .A3(n4646), .ZN(n8384) );
  NAND2_X1 U6191 ( .A1(n4647), .A2(n8326), .ZN(n4654) );
  NAND3_X1 U6192 ( .A1(n4649), .A2(n4648), .A3(n4650), .ZN(n4647) );
  OR2_X1 U6193 ( .A1(n8323), .A2(n8399), .ZN(n4648) );
  OR2_X1 U6194 ( .A1(n8319), .A2(n8383), .ZN(n4649) );
  INV_X1 U6195 ( .A(n4651), .ZN(n4650) );
  NAND2_X1 U6196 ( .A1(n4654), .A2(n8328), .ZN(n8333) );
  NAND3_X1 U6197 ( .A1(n4657), .A2(n8344), .A3(n4655), .ZN(n8349) );
  NAND4_X1 U6198 ( .A1(n4656), .A2(n8341), .A3(n8335), .A4(n8383), .ZN(n4655)
         );
  NAND3_X1 U6199 ( .A1(n8331), .A2(n8332), .A3(n8814), .ZN(n4656) );
  OR2_X1 U6200 ( .A1(n8339), .A2(n8383), .ZN(n4657) );
  NAND3_X1 U6201 ( .A1(n4659), .A2(n8399), .A3(n8279), .ZN(n4658) );
  INV_X1 U6202 ( .A(n4672), .ZN(n9734) );
  NAND2_X1 U6203 ( .A1(n9659), .A2(n4673), .ZN(n9611) );
  NOR2_X1 U6204 ( .A1(n8384), .A2(n8365), .ZN(n4679) );
  NAND2_X1 U6205 ( .A1(n4681), .A2(n8451), .ZN(n4680) );
  NAND2_X1 U6206 ( .A1(n8366), .A2(n6509), .ZN(n4681) );
  NAND2_X1 U6207 ( .A1(n4685), .A2(n4688), .ZN(n5570) );
  NAND4_X1 U6208 ( .A1(n5519), .A2(n5520), .A3(n5551), .A4(n4448), .ZN(n4685)
         );
  NAND2_X1 U6209 ( .A1(n5520), .A2(n5519), .ZN(n5536) );
  NAND3_X1 U6210 ( .A1(n5520), .A2(n5519), .A3(n4448), .ZN(n4693) );
  NAND2_X1 U6211 ( .A1(n4694), .A2(n4695), .ZN(n5448) );
  NAND2_X1 U6212 ( .A1(n5343), .A2(n4699), .ZN(n4694) );
  MUX2_X1 U6213 ( .A(n6711), .B(n6784), .S(n5122), .Z(n5161) );
  NAND2_X1 U6214 ( .A1(n5144), .A2(n5143), .ZN(n4707) );
  NAND3_X1 U6215 ( .A1(n4460), .A2(n4710), .A3(n4709), .ZN(n4708) );
  NAND2_X1 U6216 ( .A1(n4712), .A2(n5611), .ZN(n8955) );
  AND2_X2 U6217 ( .A1(n4713), .A2(n5611), .ZN(n4711) );
  OR2_X1 U6218 ( .A1(n8357), .A2(n8383), .ZN(n8237) );
  NAND3_X1 U6219 ( .A1(n4718), .A2(n4716), .A3(n4714), .ZN(n9205) );
  NAND4_X1 U6220 ( .A1(n4715), .A2(n9198), .A3(n9287), .A4(n4720), .ZN(n4714)
         );
  NAND3_X1 U6221 ( .A1(n9196), .A2(n9194), .A3(n9195), .ZN(n4715) );
  NAND2_X1 U6222 ( .A1(n4512), .A2(n9186), .ZN(n4724) );
  AND3_X1 U6223 ( .A1(n4728), .A2(n4730), .A3(n4726), .ZN(n9249) );
  OAI21_X1 U6224 ( .B1(n4727), .B2(n9216), .A(n4729), .ZN(n4726) );
  INV_X1 U6225 ( .A(n9229), .ZN(n4727) );
  NAND2_X1 U6226 ( .A1(n9230), .A2(n9287), .ZN(n4728) );
  OAI21_X1 U6227 ( .B1(n9263), .B2(n4734), .A(n4733), .ZN(n4732) );
  NAND2_X1 U6228 ( .A1(n8084), .A2(n4737), .ZN(n4736) );
  NAND2_X2 U6229 ( .A1(n4741), .A2(n9830), .ZN(n5930) );
  NAND2_X1 U6230 ( .A1(n5911), .A2(n4743), .ZN(n4742) );
  NAND3_X1 U6231 ( .A1(n4749), .A2(n9267), .A3(n4748), .ZN(n8502) );
  NAND3_X1 U6232 ( .A1(n9621), .A2(n4752), .A3(n4751), .ZN(n4748) );
  NAND3_X1 U6233 ( .A1(n9644), .A2(n4751), .A3(n9621), .ZN(n4749) );
  INV_X1 U6234 ( .A(n4755), .ZN(n9647) );
  NAND3_X1 U6235 ( .A1(n9755), .A2(n9756), .A3(n9757), .ZN(n9816) );
  NAND2_X1 U6236 ( .A1(n4760), .A2(n6593), .ZN(n8130) );
  AOI21_X1 U6237 ( .B1(n4456), .B2(P2_IR_REG_1__SCAN_IN), .A(n4764), .ZN(n4763) );
  NAND2_X1 U6238 ( .A1(n6602), .A2(n6604), .ZN(n4776) );
  NAND3_X1 U6239 ( .A1(n4777), .A2(n4776), .A3(n4524), .ZN(n6605) );
  NAND2_X1 U6240 ( .A1(n6597), .A2(n4785), .ZN(n4782) );
  NAND2_X1 U6241 ( .A1(n4791), .A2(n4786), .ZN(P2_U3199) );
  NAND3_X1 U6242 ( .A1(n4790), .A2(n8719), .A3(n4789), .ZN(n4788) );
  OAI21_X1 U6243 ( .B1(n8717), .B2(n8718), .A(n8741), .ZN(n4791) );
  NOR2_X1 U6244 ( .A1(n6571), .A2(n6708), .ZN(n6572) );
  NAND2_X1 U6245 ( .A1(n7706), .A2(n6589), .ZN(n6591) );
  NOR2_X1 U6246 ( .A1(n7529), .A2(n6585), .ZN(n7709) );
  NAND2_X1 U6247 ( .A1(n7254), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7154) );
  NOR2_X1 U6248 ( .A1(n7530), .A2(n7785), .ZN(n7529) );
  NAND2_X1 U6249 ( .A1(n6567), .A2(n6568), .ZN(n7173) );
  NAND2_X1 U6250 ( .A1(n6588), .A2(n6587), .ZN(n7706) );
  NOR2_X1 U6251 ( .A1(n4792), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n5067) );
  NAND2_X1 U6252 ( .A1(n4462), .A2(n4436), .ZN(n4792) );
  NAND2_X1 U6253 ( .A1(n5153), .A2(n7303), .ZN(n8258) );
  NAND3_X1 U6254 ( .A1(n5150), .A2(n5151), .A3(n5152), .ZN(n5153) );
  NAND2_X1 U6255 ( .A1(n5113), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5109) );
  NAND3_X1 U6256 ( .A1(n4430), .A2(n5077), .A3(n5107), .ZN(n5113) );
  NAND2_X1 U6257 ( .A1(n4795), .A2(n8318), .ZN(n4794) );
  INV_X1 U6258 ( .A(n5655), .ZN(n4795) );
  INV_X1 U6259 ( .A(n7716), .ZN(n4812) );
  NAND2_X1 U6260 ( .A1(n4813), .A2(n4814), .ZN(n7744) );
  INV_X1 U6261 ( .A(n6708), .ZN(n4846) );
  NOR2_X2 U6262 ( .A1(n10144), .A2(n4520), .ZN(n6557) );
  AND2_X2 U6263 ( .A1(n4852), .A2(n4851), .ZN(n10144) );
  NAND2_X1 U6264 ( .A1(n4855), .A2(n4853), .ZN(n7698) );
  NAND2_X1 U6265 ( .A1(n4854), .A2(n4856), .ZN(n4853) );
  INV_X1 U6266 ( .A(n7525), .ZN(n4854) );
  XNOR2_X2 U6267 ( .A(n6544), .B(n6582), .ZN(n7525) );
  NAND2_X1 U6268 ( .A1(n6551), .A2(n4866), .ZN(n4862) );
  INV_X1 U6269 ( .A(n7720), .ZN(n4873) );
  NAND3_X1 U6270 ( .A1(n4870), .A2(n7754), .A3(n4869), .ZN(n7747) );
  OR2_X1 U6271 ( .A1(n4872), .A2(n7720), .ZN(n4869) );
  NAND2_X1 U6272 ( .A1(n4871), .A2(n7718), .ZN(n4870) );
  INV_X1 U6273 ( .A(n4872), .ZN(n4871) );
  NAND2_X1 U6274 ( .A1(n5550), .A2(n4878), .ZN(n4874) );
  NAND3_X1 U6275 ( .A1(n5105), .A2(n5050), .A3(n5051), .ZN(n5233) );
  INV_X1 U6276 ( .A(n9840), .ZN(n4894) );
  OR2_X1 U6277 ( .A1(n4421), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4897) );
  XNOR2_X1 U6278 ( .A(n5674), .B(n8436), .ZN(n5627) );
  NAND2_X1 U6279 ( .A1(n4906), .A2(n4903), .ZN(n4899) );
  INV_X1 U6280 ( .A(n4902), .ZN(n4901) );
  INV_X1 U6281 ( .A(n5786), .ZN(n4905) );
  NAND2_X1 U6282 ( .A1(n8615), .A2(n4913), .ZN(n4912) );
  NAND2_X1 U6283 ( .A1(n5796), .A2(n4504), .ZN(n8151) );
  OAI22_X2 U6284 ( .A1(n9929), .A2(n4427), .B1(n9448), .B2(n9934), .ZN(n7674)
         );
  NAND2_X1 U6285 ( .A1(n7674), .A2(n4932), .ZN(n4936) );
  INV_X1 U6286 ( .A(n5008), .ZN(n4938) );
  NAND2_X1 U6287 ( .A1(n9687), .A2(n4499), .ZN(n4940) );
  INV_X2 U6288 ( .A(n6009), .ZN(n9279) );
  AND2_X1 U6289 ( .A1(n9810), .A2(n9437), .ZN(n4956) );
  AND2_X2 U6290 ( .A1(n4958), .A2(n4957), .ZN(n8206) );
  OR2_X2 U6291 ( .A1(n8091), .A2(n9308), .ZN(n4958) );
  NAND2_X1 U6292 ( .A1(n4959), .A2(n4960), .ZN(n9610) );
  NAND2_X1 U6293 ( .A1(n9620), .A2(n4431), .ZN(n4959) );
  NAND2_X1 U6294 ( .A1(n4961), .A2(n4431), .ZN(n9608) );
  NAND3_X1 U6295 ( .A1(n5895), .A2(n4439), .A3(n6866), .ZN(n5907) );
  NAND2_X1 U6296 ( .A1(n6043), .A2(n7369), .ZN(n7424) );
  NAND2_X1 U6297 ( .A1(n4968), .A2(n6063), .ZN(n7542) );
  NAND2_X1 U6298 ( .A1(n4521), .A2(n6043), .ZN(n4968) );
  INV_X1 U6299 ( .A(n7540), .ZN(n4970) );
  NAND2_X1 U6300 ( .A1(n7940), .A2(n4974), .ZN(n4972) );
  NAND2_X1 U6301 ( .A1(n6221), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6255) );
  NAND2_X1 U6302 ( .A1(n9051), .A2(n4980), .ZN(n4979) );
  NAND3_X1 U6303 ( .A1(n4981), .A2(n4982), .A3(n4984), .ZN(n4978) );
  NAND2_X1 U6304 ( .A1(n9028), .A2(n4991), .ZN(n4990) );
  INV_X1 U6305 ( .A(n6216), .ZN(n4989) );
  NAND3_X1 U6306 ( .A1(n4990), .A2(n6254), .A3(n4988), .ZN(n9087) );
  OAI211_X1 U6307 ( .C1(n9123), .C2(n4997), .A(n4994), .B(n4995), .ZN(n9103)
         );
  NAND2_X1 U6308 ( .A1(n9125), .A2(n4506), .ZN(n4994) );
  NAND2_X1 U6309 ( .A1(n5000), .A2(n4505), .ZN(n7286) );
  NAND2_X1 U6310 ( .A1(n9763), .A2(n5023), .ZN(n9817) );
  OAI21_X1 U6311 ( .B1(n5728), .B2(n5686), .A(n5711), .ZN(n6499) );
  NAND2_X1 U6312 ( .A1(n7460), .A2(n7444), .ZN(n9364) );
  OAI21_X2 U6313 ( .B1(n9631), .B2(n8516), .A(n8515), .ZN(n9620) );
  OAI22_X1 U6314 ( .A1(n5987), .A2(n5941), .B1(n5986), .B2(n5953), .ZN(n5942)
         );
  NAND2_X1 U6315 ( .A1(n8468), .A2(n5929), .ZN(n5986) );
  NAND2_X1 U6316 ( .A1(n5340), .A2(n5339), .ZN(n7950) );
  NAND2_X1 U6317 ( .A1(n5756), .A2(n5125), .ZN(n5653) );
  NAND2_X1 U6318 ( .A1(n9138), .A2(n9139), .ZN(n9137) );
  OAI222_X1 U6319 ( .A1(n5628), .A2(n5627), .B1(n8646), .B2(n10171), .C1(n5602), .C2(n5626), .ZN(n5629) );
  OAI22_X2 U6320 ( .A1(n9642), .A2(n8514), .B1(n9431), .B2(n9776), .ZN(n9631)
         );
  NOR2_X2 U6321 ( .A1(n9066), .A2(n9065), .ZN(n9064) );
  NAND2_X4 U6322 ( .A1(n5114), .A2(n5113), .ZN(n8460) );
  OR2_X1 U6323 ( .A1(n10261), .A2(n6821), .ZN(n5001) );
  INV_X1 U6324 ( .A(n10261), .ZN(n6692) );
  OR2_X1 U6325 ( .A1(n10174), .A2(n5712), .ZN(n5003) );
  AND4_X1 U6326 ( .A1(n5361), .A2(n5360), .A3(n5359), .A4(n5358), .ZN(n7952)
         );
  OR2_X1 U6327 ( .A1(n10238), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5004) );
  AND2_X1 U6328 ( .A1(n5074), .A2(n5090), .ZN(n5005) );
  OR2_X1 U6329 ( .A1(n5408), .A2(n6808), .ZN(n5006) );
  AND2_X1 U6330 ( .A1(n6537), .A2(n6714), .ZN(n5007) );
  AND2_X1 U6331 ( .A1(n10052), .A2(n7475), .ZN(n5008) );
  AND3_X1 U6332 ( .A1(n5888), .A2(n5880), .A3(n5891), .ZN(n5009) );
  INV_X1 U6333 ( .A(n5900), .ZN(n6235) );
  INV_X1 U6334 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5121) );
  NAND2_X1 U6335 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n5010) );
  AND2_X1 U6336 ( .A1(n5303), .A2(n5295), .ZN(n5011) );
  INV_X1 U6337 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6718) );
  INV_X1 U6338 ( .A(n8901), .ZN(n5715) );
  INV_X1 U6339 ( .A(n6625), .ZN(n6582) );
  INV_X1 U6340 ( .A(n6518), .ZN(n8233) );
  INV_X1 U6341 ( .A(n8946), .ZN(n8448) );
  NAND2_X1 U6342 ( .A1(n7020), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5013) );
  NOR2_X1 U6343 ( .A1(n8946), .A2(n8455), .ZN(n8441) );
  AND2_X1 U6344 ( .A1(n6541), .A2(n7237), .ZN(n5014) );
  NOR2_X1 U6345 ( .A1(n8233), .A2(n8989), .ZN(n6519) );
  NAND2_X1 U6346 ( .A1(n8857), .A2(n8856), .ZN(n5015) );
  INV_X1 U6347 ( .A(n9097), .ZN(n9846) );
  AND2_X1 U6348 ( .A1(n7473), .A2(n10035), .ZN(n5016) );
  NAND2_X1 U6349 ( .A1(n5624), .A2(n5623), .ZN(n8655) );
  NAND2_X1 U6350 ( .A1(n5601), .A2(n5600), .ZN(n8783) );
  AND2_X1 U6351 ( .A1(n7164), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5017) );
  OR2_X1 U6352 ( .A1(n8751), .A2(n8748), .ZN(n5018) );
  AND4_X1 U6353 ( .A1(n8400), .A2(n5753), .A3(n8464), .A4(n5754), .ZN(n5019)
         );
  AND3_X1 U6354 ( .A1(n8451), .A2(n8450), .A3(n8449), .ZN(n5020) );
  OR3_X1 U6355 ( .A1(n8596), .A2(n8656), .A3(n8808), .ZN(n5021) );
  AND2_X1 U6356 ( .A1(n8596), .A2(n8808), .ZN(n5022) );
  AND3_X1 U6357 ( .A1(n9762), .A2(n9761), .A3(n9760), .ZN(n5023) );
  NAND2_X1 U6358 ( .A1(n5212), .A2(n5211), .ZN(n5024) );
  NAND2_X1 U6359 ( .A1(n8448), .A2(n5018), .ZN(n8449) );
  NAND2_X1 U6360 ( .A1(n8379), .A2(n8383), .ZN(n8386) );
  AND2_X1 U6361 ( .A1(n5439), .A2(n5440), .ZN(n5430) );
  INV_X1 U6362 ( .A(n6580), .ZN(n6581) );
  NAND2_X1 U6363 ( .A1(n5005), .A2(n5075), .ZN(n5076) );
  INV_X1 U6364 ( .A(n9438), .ZN(n8204) );
  AND2_X1 U6365 ( .A1(n5441), .A2(n5433), .ZN(n5432) );
  OR2_X1 U6366 ( .A1(n8529), .A2(n5818), .ZN(n5816) );
  AND2_X1 U6367 ( .A1(n7477), .A2(n6705), .ZN(n5906) );
  AOI22_X1 U6368 ( .A1(n5931), .A2(P1_REG1_REG_1__SCAN_IN), .B1(n6008), .B2(
        P1_REG0_REG_1__SCAN_IN), .ZN(n5932) );
  OR2_X1 U6369 ( .A1(n9766), .A2(n9429), .ZN(n8517) );
  OR2_X1 U6370 ( .A1(n6321), .A2(n6320), .ZN(n6339) );
  INV_X1 U6371 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5915) );
  OR2_X1 U6372 ( .A1(n5446), .A2(n5445), .ZN(n5447) );
  INV_X1 U6373 ( .A(n5387), .ZN(n5405) );
  NAND2_X1 U6374 ( .A1(n5824), .A2(n5021), .ZN(n5825) );
  INV_X1 U6375 ( .A(n8635), .ZN(n8640) );
  INV_X1 U6376 ( .A(n7706), .ZN(n7707) );
  OR2_X1 U6377 ( .A1(n10205), .A2(n5753), .ZN(n5719) );
  AND2_X1 U6378 ( .A1(n5635), .A2(n6730), .ZN(n5751) );
  AND2_X1 U6379 ( .A1(n8955), .A2(n8774), .ZN(n8352) );
  AND2_X1 U6380 ( .A1(n9010), .A2(n8227), .ZN(n8873) );
  INV_X1 U6381 ( .A(n5634), .ZN(n5632) );
  INV_X1 U6382 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5376) );
  INV_X1 U6383 ( .A(n5165), .ZN(n5167) );
  NOR2_X1 U6384 ( .A1(n6988), .A2(n6411), .ZN(n6481) );
  NAND2_X1 U6385 ( .A1(n6365), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6386) );
  NAND2_X1 U6386 ( .A1(n6289), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6321) );
  NAND2_X1 U6387 ( .A1(n8088), .A2(n9859), .ZN(n8089) );
  NAND2_X1 U6388 ( .A1(n7443), .A2(n7442), .ZN(n7445) );
  AND2_X1 U6389 ( .A1(n8045), .A2(n9441), .ZN(n8046) );
  NOR2_X1 U6390 ( .A1(n7947), .A2(n9443), .ZN(n7875) );
  NOR2_X1 U6391 ( .A1(n7480), .A2(n9445), .ZN(n7640) );
  INV_X1 U6392 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5923) );
  NAND2_X1 U6393 ( .A1(n5323), .A2(n6846), .ZN(n5341) );
  NAND2_X1 U6394 ( .A1(n5293), .A2(n5292), .ZN(n5303) );
  AND2_X1 U6395 ( .A1(n5832), .A2(n5831), .ZN(n5833) );
  XNOR2_X1 U6396 ( .A(n8971), .B(n5828), .ZN(n8596) );
  INV_X1 U6397 ( .A(n8655), .ZN(n8646) );
  INV_X1 U6398 ( .A(n8186), .ZN(n6554) );
  INV_X1 U6399 ( .A(n8679), .ZN(n6599) );
  OR2_X1 U6400 ( .A1(n5618), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8749) );
  AND2_X1 U6401 ( .A1(n8335), .A2(n8814), .ZN(n8833) );
  AND2_X1 U6402 ( .A1(n8309), .A2(n8310), .ZN(n8308) );
  AND2_X1 U6403 ( .A1(n8966), .A2(n8797), .ZN(n8402) );
  OR2_X1 U6404 ( .A1(n8977), .A2(n8821), .ZN(n8346) );
  OR2_X1 U6405 ( .A1(n8993), .A2(n8865), .ZN(n8334) );
  NOR2_X1 U6406 ( .A1(n6144), .A2(n7966), .ZN(n6146) );
  AND2_X1 U6407 ( .A1(n6426), .A2(n6425), .ZN(n6677) );
  OR2_X1 U6408 ( .A1(n5960), .A2(n7036), .ZN(n5914) );
  INV_X1 U6409 ( .A(n9431), .ZN(n9104) );
  AND2_X1 U6410 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6028) );
  INV_X1 U6411 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7545) );
  INV_X1 U6412 ( .A(n9609), .ZN(n9601) );
  NAND2_X1 U6413 ( .A1(n5570), .A2(n5569), .ZN(n5584) );
  XNOR2_X1 U6414 ( .A(n5363), .B(SI_12_), .ZN(n5362) );
  NAND2_X1 U6415 ( .A1(n5230), .A2(SI_5_), .ZN(n5231) );
  INV_X1 U6416 ( .A(n8645), .ZN(n8632) );
  AND2_X1 U6417 ( .A1(n7521), .A2(n5705), .ZN(n8234) );
  NAND2_X1 U6418 ( .A1(n5092), .A2(n6726), .ZN(n10165) );
  NAND2_X1 U6419 ( .A1(n7298), .A2(n8264), .ZN(n7716) );
  OAI21_X1 U6420 ( .B1(n8233), .B2(n8925), .A(n5001), .ZN(n6690) );
  INV_X1 U6421 ( .A(n8925), .ZN(n8937) );
  NAND2_X1 U6422 ( .A1(n5508), .A2(n5507), .ZN(n8836) );
  NAND2_X1 U6423 ( .A1(n5458), .A2(n5457), .ZN(n9003) );
  INV_X1 U6424 ( .A(n8989), .ZN(n9009) );
  AND2_X1 U6425 ( .A1(n6524), .A2(n6732), .ZN(n6726) );
  AND2_X1 U6426 ( .A1(n5069), .A2(n5089), .ZN(n8464) );
  INV_X1 U6427 ( .A(n9987), .ZN(n9967) );
  INV_X1 U6428 ( .A(n9741), .ZN(n9981) );
  NAND2_X1 U6429 ( .A1(n10048), .A2(n10000), .ZN(n10095) );
  INV_X1 U6430 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5903) );
  XNOR2_X1 U6431 ( .A(n5229), .B(SI_5_), .ZN(n5227) );
  AND2_X1 U6432 ( .A1(n5867), .A2(n5866), .ZN(n5872) );
  INV_X1 U6433 ( .A(n8616), .ZN(n8650) );
  INV_X1 U6434 ( .A(n6509), .ZN(n8654) );
  INV_X1 U6435 ( .A(n8200), .ZN(n8892) );
  AND2_X1 U6436 ( .A1(n6668), .A2(n6667), .ZN(n10162) );
  OR2_X1 U6437 ( .A1(n6563), .A2(n6611), .ZN(n10147) );
  NAND2_X1 U6438 ( .A1(n5668), .A2(n10165), .ZN(n8895) );
  NAND2_X1 U6439 ( .A1(n10174), .A2(n10173), .ZN(n8901) );
  INV_X1 U6440 ( .A(n6690), .ZN(n6691) );
  AND2_X1 U6441 ( .A1(n5745), .A2(n5744), .ZN(n10240) );
  INV_X1 U6442 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6809) );
  INV_X1 U6443 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6784) );
  INV_X1 U6444 ( .A(n6687), .ZN(n6688) );
  AND2_X1 U6445 ( .A1(n6473), .A2(n8523), .ZN(n9161) );
  OR2_X1 U6446 ( .A1(n6435), .A2(n6434), .ZN(n9605) );
  INV_X1 U6447 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9590) );
  INV_X1 U6448 ( .A(n9968), .ZN(n9746) );
  NAND2_X1 U6449 ( .A1(n7438), .A2(n8523), .ZN(n9744) );
  INV_X1 U6450 ( .A(n10120), .ZN(n10118) );
  INV_X1 U6451 ( .A(n10098), .ZN(n10097) );
  INV_X1 U6452 ( .A(n9998), .ZN(n9999) );
  AND2_X1 U6453 ( .A1(n7910), .A2(n6466), .ZN(n9828) );
  INV_X1 U6454 ( .A(n4429), .ZN(n7854) );
  OAI21_X1 U6455 ( .B1(n5718), .B2(n10176), .A(n5717), .ZN(P2_U3205) );
  OAI21_X1 U6456 ( .B1(n8925), .B2(n5749), .A(n5736), .ZN(P2_U3486) );
  OAI21_X1 U6457 ( .B1(n8989), .B2(n5749), .A(n5748), .ZN(P2_U3454) );
  AND2_X1 U6458 ( .A1(n7910), .A2(n6706), .ZN(P1_U3973) );
  INV_X1 U6459 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5030) );
  INV_X1 U6460 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5032) );
  INV_X1 U6461 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5034) );
  OR2_X2 U6462 ( .A1(n5380), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5396) );
  INV_X1 U6463 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5036) );
  OR2_X2 U6464 ( .A1(n5421), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5459) );
  INV_X1 U6465 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6842) );
  OR2_X2 U6466 ( .A1(n5476), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5496) );
  OR2_X2 U6467 ( .A1(n5496), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5509) );
  INV_X1 U6468 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n5039) );
  INV_X1 U6469 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5041) );
  OR2_X2 U6470 ( .A1(n5543), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5563) );
  INV_X1 U6471 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n5043) );
  INV_X1 U6472 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5045) );
  OR2_X2 U6473 ( .A1(n5593), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5595) );
  INV_X1 U6474 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n5047) );
  NAND2_X1 U6475 ( .A1(n5595), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5049) );
  NAND2_X1 U6476 ( .A1(n5618), .A2(n5049), .ZN(n8642) );
  INV_X1 U6477 ( .A(n8642), .ZN(n5630) );
  INV_X1 U6478 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5052) );
  NAND2_X1 U6479 ( .A1(n5052), .A2(n5328), .ZN(n5053) );
  INV_X1 U6480 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5054) );
  INV_X1 U6481 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5065) );
  NAND3_X1 U6482 ( .A1(n5063), .A2(n5065), .A3(n5376), .ZN(n5055) );
  INV_X1 U6483 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5056) );
  NAND2_X1 U6484 ( .A1(n5058), .A2(n5064), .ZN(n5057) );
  XNOR2_X1 U6485 ( .A(n5071), .B(n5070), .ZN(n5754) );
  INV_X1 U6486 ( .A(n5058), .ZN(n5059) );
  NAND2_X1 U6487 ( .A1(n5059), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5060) );
  INV_X1 U6488 ( .A(n7409), .ZN(n5637) );
  NAND2_X1 U6489 ( .A1(n5754), .A2(n5637), .ZN(n5666) );
  NOR2_X1 U6490 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5062) );
  NOR2_X1 U6491 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5061) );
  NAND2_X1 U6492 ( .A1(n4473), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5066) );
  MUX2_X1 U6493 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5066), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n5069) );
  INV_X1 U6494 ( .A(n5326), .ZN(n5068) );
  NAND2_X1 U6495 ( .A1(n5068), .A2(n5067), .ZN(n5089) );
  NAND2_X1 U6496 ( .A1(n5071), .A2(n5070), .ZN(n5072) );
  INV_X1 U6497 ( .A(n5719), .ZN(n5092) );
  INV_X1 U6498 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5074) );
  INV_X1 U6499 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5075) );
  NAND2_X1 U6500 ( .A1(n5094), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5079) );
  MUX2_X1 U6501 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5079), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5080) );
  AND2_X1 U6502 ( .A1(n5111), .A2(n5080), .ZN(n5634) );
  NAND2_X1 U6503 ( .A1(n4482), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5084) );
  INV_X1 U6504 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5082) );
  NAND2_X1 U6505 ( .A1(n5084), .A2(n5082), .ZN(n5086) );
  NAND2_X1 U6506 ( .A1(n5086), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5083) );
  XNOR2_X1 U6507 ( .A(n5083), .B(P2_IR_REG_25__SCAN_IN), .ZN(n5631) );
  INV_X1 U6508 ( .A(n5084), .ZN(n5085) );
  NAND2_X1 U6509 ( .A1(n5085), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n5087) );
  NAND3_X1 U6510 ( .A1(n5634), .A2(n5631), .A3(n5088), .ZN(n6524) );
  NAND2_X1 U6511 ( .A1(n5089), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5091) );
  XNOR2_X1 U6512 ( .A(n5091), .B(n5090), .ZN(n6525) );
  AND2_X1 U6513 ( .A1(n6525), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6732) );
  INV_X1 U6514 ( .A(n5754), .ZN(n5093) );
  NAND2_X1 U6515 ( .A1(n5753), .A2(n5093), .ZN(n8447) );
  NAND2_X1 U6516 ( .A1(n5637), .A2(n8464), .ZN(n5739) );
  NAND2_X1 U6517 ( .A1(n8447), .A2(n5739), .ZN(n8894) );
  INV_X1 U6518 ( .A(n8894), .ZN(n5628) );
  INV_X1 U6519 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5108) );
  NOR2_X1 U6520 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n5107) );
  AND2_X1 U6521 ( .A1(n5108), .A2(n5107), .ZN(n5095) );
  INV_X1 U6522 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5097) );
  INV_X1 U6523 ( .A(n5102), .ZN(n5101) );
  NAND2_X1 U6524 ( .A1(n5099), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5100) );
  NAND2_X1 U6525 ( .A1(n5179), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5104) );
  INV_X1 U6526 ( .A(n6566), .ZN(n5106) );
  XNOR2_X1 U6527 ( .A(n5109), .B(n5108), .ZN(n5110) );
  NAND2_X1 U6528 ( .A1(n5115), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n5116) );
  INV_X1 U6529 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5120) );
  AND2_X1 U6530 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5123) );
  NAND2_X1 U6531 ( .A1(n5186), .A2(n5123), .ZN(n5946) );
  AND2_X1 U6532 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5124) );
  NAND2_X1 U6533 ( .A1(n8392), .A2(n5124), .ZN(n5132) );
  XNOR2_X1 U6534 ( .A(n5142), .B(n5143), .ZN(n5913) );
  INV_X1 U6535 ( .A(n5136), .ZN(n5125) );
  NAND2_X1 U6536 ( .A1(n5135), .A2(n5136), .ZN(n8251) );
  NAND2_X1 U6537 ( .A1(n5179), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5129) );
  NAND2_X1 U6538 ( .A1(n5178), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5128) );
  NAND2_X1 U6539 ( .A1(n5155), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5127) );
  NAND2_X1 U6540 ( .A1(n5176), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5126) );
  NAND4_X1 U6541 ( .A1(n5129), .A2(n5128), .A3(n5127), .A4(n5126), .ZN(n8671)
         );
  NAND2_X1 U6542 ( .A1(n8392), .A2(SI_0_), .ZN(n5131) );
  INV_X1 U6543 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5130) );
  NAND2_X1 U6544 ( .A1(n5131), .A2(n5130), .ZN(n5133) );
  NAND2_X1 U6545 ( .A1(n5133), .A2(n5132), .ZN(n9025) );
  MUX2_X1 U6546 ( .A(n4762), .B(n9025), .S(n5134), .Z(n7309) );
  INV_X1 U6547 ( .A(n7309), .ZN(n7582) );
  NAND2_X1 U6548 ( .A1(n5756), .A2(n5136), .ZN(n5137) );
  NAND2_X1 U6549 ( .A1(n5179), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5141) );
  NAND2_X1 U6550 ( .A1(n5155), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5139) );
  NAND2_X1 U6551 ( .A1(n5176), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5138) );
  OR2_X1 U6552 ( .A1(n4422), .A2(n6784), .ZN(n5152) );
  NAND2_X1 U6553 ( .A1(n5145), .A2(SI_1_), .ZN(n5146) );
  OR2_X1 U6554 ( .A1(n5296), .A2(n6710), .ZN(n5151) );
  NAND2_X1 U6555 ( .A1(n5169), .A2(n6632), .ZN(n5150) );
  NAND2_X1 U6556 ( .A1(n8670), .A2(n10182), .ZN(n8259) );
  NAND2_X1 U6557 ( .A1(n5177), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5159) );
  NAND2_X1 U6558 ( .A1(n5179), .A2(n5154), .ZN(n5158) );
  NAND2_X1 U6559 ( .A1(n5178), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5157) );
  NAND2_X1 U6560 ( .A1(n5155), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5156) );
  NAND4_X1 U6561 ( .A1(n5159), .A2(n5158), .A3(n5157), .A4(n5156), .ZN(n8669)
         );
  INV_X1 U6562 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6709) );
  OR2_X1 U6563 ( .A1(n4422), .A2(n6709), .ZN(n5172) );
  INV_X1 U6564 ( .A(n5161), .ZN(n5162) );
  NAND2_X1 U6565 ( .A1(n5162), .A2(SI_2_), .ZN(n5163) );
  NAND2_X1 U6566 ( .A1(n5164), .A2(n5163), .ZN(n5210) );
  INV_X1 U6567 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6713) );
  MUX2_X1 U6568 ( .A(n6709), .B(n6713), .S(n5186), .Z(n5187) );
  XNOR2_X1 U6569 ( .A(n5210), .B(n5209), .ZN(n6712) );
  OR2_X1 U6570 ( .A1(n5296), .A2(n6712), .ZN(n5171) );
  NAND2_X1 U6571 ( .A1(n5167), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5166) );
  MUX2_X1 U6572 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5166), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5168) );
  NAND2_X1 U6573 ( .A1(n5169), .A2(n6708), .ZN(n5170) );
  INV_X1 U6574 ( .A(n7869), .ZN(n7395) );
  NAND2_X1 U6575 ( .A1(n7301), .A2(n5173), .ZN(n5175) );
  NAND2_X1 U6576 ( .A1(n8669), .A2(n7395), .ZN(n5174) );
  NAND2_X1 U6577 ( .A1(n5175), .A2(n5174), .ZN(n7718) );
  NAND2_X1 U6578 ( .A1(n5177), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5184) );
  NAND2_X1 U6579 ( .A1(n5178), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5183) );
  NAND2_X1 U6580 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5180) );
  NAND2_X1 U6581 ( .A1(n5199), .A2(n5180), .ZN(n7726) );
  NAND2_X1 U6582 ( .A1(n5179), .A2(n7726), .ZN(n5182) );
  NAND2_X1 U6583 ( .A1(n5155), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5181) );
  NAND4_X1 U6584 ( .A1(n5184), .A2(n5183), .A3(n5182), .A4(n5181), .ZN(n8668)
         );
  NAND2_X1 U6585 ( .A1(n5210), .A2(n5209), .ZN(n5189) );
  INV_X1 U6586 ( .A(n5187), .ZN(n5188) );
  NAND2_X1 U6587 ( .A1(n5189), .A2(n5212), .ZN(n5190) );
  XNOR2_X1 U6588 ( .A(n5205), .B(n5190), .ZN(n8490) );
  OR2_X1 U6589 ( .A1(n5296), .A2(n8490), .ZN(n5197) );
  OR2_X1 U6590 ( .A1(n4422), .A2(n6718), .ZN(n5196) );
  NAND2_X1 U6591 ( .A1(n5192), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5191) );
  MUX2_X1 U6592 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5191), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5194) );
  INV_X1 U6593 ( .A(n5192), .ZN(n5193) );
  INV_X1 U6594 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6782) );
  NAND2_X1 U6595 ( .A1(n5193), .A2(n6782), .ZN(n5216) );
  OR2_X1 U6596 ( .A1(n5134), .A2(n7164), .ZN(n5195) );
  INV_X1 U6597 ( .A(n10189), .ZN(n7727) );
  OR2_X1 U6598 ( .A1(n8668), .A2(n7727), .ZN(n5198) );
  NAND2_X1 U6599 ( .A1(n8668), .A2(n7727), .ZN(n7720) );
  NAND2_X1 U6600 ( .A1(n5155), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5204) );
  NAND2_X1 U6601 ( .A1(n5177), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5203) );
  INV_X2 U6602 ( .A(n5699), .ZN(n5526) );
  NAND2_X1 U6603 ( .A1(n5199), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5200) );
  NAND2_X1 U6604 ( .A1(n5221), .A2(n5200), .ZN(n7759) );
  NAND2_X1 U6605 ( .A1(n5526), .A2(n7759), .ZN(n5202) );
  NAND2_X1 U6606 ( .A1(n5178), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5201) );
  NAND4_X1 U6607 ( .A1(n5204), .A2(n5203), .A3(n5202), .A4(n5201), .ZN(n8667)
         );
  INV_X1 U6608 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6715) );
  INV_X1 U6609 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6717) );
  MUX2_X1 U6610 ( .A(n6715), .B(n6717), .S(n5186), .Z(n5229) );
  INV_X1 U6611 ( .A(n5205), .ZN(n5208) );
  INV_X1 U6612 ( .A(n5206), .ZN(n5207) );
  NAND2_X1 U6613 ( .A1(n5213), .A2(n5024), .ZN(n5214) );
  NAND2_X1 U6614 ( .A1(n5215), .A2(n5214), .ZN(n5228) );
  XNOR2_X1 U6615 ( .A(n5227), .B(n5228), .ZN(n6716) );
  OR2_X1 U6616 ( .A1(n5296), .A2(n6716), .ZN(n5220) );
  OR2_X1 U6617 ( .A1(n4422), .A2(n6715), .ZN(n5219) );
  NAND2_X1 U6618 ( .A1(n5216), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5217) );
  NAND2_X1 U6619 ( .A1(n5169), .A2(n8483), .ZN(n5218) );
  INV_X1 U6620 ( .A(n10194), .ZN(n7760) );
  OR2_X1 U6621 ( .A1(n8667), .A2(n7760), .ZN(n7755) );
  NAND2_X1 U6622 ( .A1(n8667), .A2(n7760), .ZN(n7754) );
  NAND2_X1 U6623 ( .A1(n5155), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5226) );
  NAND2_X1 U6624 ( .A1(n5177), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5225) );
  NAND2_X1 U6625 ( .A1(n5221), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5222) );
  NAND2_X1 U6626 ( .A1(n5243), .A2(n5222), .ZN(n7745) );
  NAND2_X1 U6627 ( .A1(n5526), .A2(n7745), .ZN(n5224) );
  NAND2_X1 U6628 ( .A1(n5178), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5223) );
  NAND4_X1 U6629 ( .A1(n5226), .A2(n5225), .A3(n5224), .A4(n5223), .ZN(n8666)
         );
  NAND2_X1 U6630 ( .A1(n5228), .A2(n5227), .ZN(n5232) );
  INV_X1 U6631 ( .A(n5229), .ZN(n5230) );
  INV_X1 U6632 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6721) );
  INV_X1 U6633 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6719) );
  MUX2_X1 U6634 ( .A(n6721), .B(n6719), .S(n5186), .Z(n5251) );
  XNOR2_X1 U6635 ( .A(n5250), .B(n5249), .ZN(n6720) );
  OR2_X1 U6636 ( .A1(n5296), .A2(n6720), .ZN(n5239) );
  OR2_X1 U6637 ( .A1(n4422), .A2(n6721), .ZN(n5238) );
  NAND2_X1 U6638 ( .A1(n5233), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5234) );
  MUX2_X1 U6639 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5234), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n5236) );
  AND2_X1 U6640 ( .A1(n5236), .A2(n5235), .ZN(n6642) );
  NAND2_X1 U6641 ( .A1(n5169), .A2(n6642), .ZN(n5237) );
  INV_X1 U6642 ( .A(n10198), .ZN(n7746) );
  OR2_X1 U6643 ( .A1(n8666), .A2(n7746), .ZN(n5240) );
  NAND2_X1 U6644 ( .A1(n7747), .A2(n5240), .ZN(n5242) );
  NAND2_X1 U6645 ( .A1(n8666), .A2(n7746), .ZN(n5241) );
  NAND2_X1 U6646 ( .A1(n5242), .A2(n5241), .ZN(n7627) );
  NAND2_X1 U6647 ( .A1(n5177), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5248) );
  NAND2_X1 U6648 ( .A1(n5155), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5247) );
  NAND2_X1 U6649 ( .A1(n5243), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5244) );
  NAND2_X1 U6650 ( .A1(n5261), .A2(n5244), .ZN(n7636) );
  NAND2_X1 U6651 ( .A1(n5526), .A2(n7636), .ZN(n5246) );
  NAND2_X1 U6652 ( .A1(n5178), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5245) );
  NAND4_X1 U6653 ( .A1(n5248), .A2(n5247), .A3(n5246), .A4(n5245), .ZN(n8665)
         );
  INV_X1 U6654 ( .A(n5251), .ZN(n5252) );
  NAND2_X1 U6655 ( .A1(n5252), .A2(SI_6_), .ZN(n5253) );
  MUX2_X1 U6656 ( .A(n6809), .B(n6964), .S(n5186), .Z(n5269) );
  XNOR2_X1 U6657 ( .A(n5268), .B(n5267), .ZN(n6723) );
  OR2_X1 U6658 ( .A1(n5296), .A2(n6723), .ZN(n5260) );
  OR2_X1 U6659 ( .A1(n4421), .A2(n6809), .ZN(n5259) );
  NAND2_X1 U6660 ( .A1(n5235), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5254) );
  MUX2_X1 U6661 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5254), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n5257) );
  INV_X1 U6662 ( .A(n5255), .ZN(n5256) );
  NAND2_X1 U6663 ( .A1(n5257), .A2(n5256), .ZN(n7237) );
  OR2_X1 U6664 ( .A1(n5134), .A2(n7237), .ZN(n5258) );
  OR2_X1 U6665 ( .A1(n8665), .A2(n10204), .ZN(n8291) );
  NAND2_X1 U6666 ( .A1(n8665), .A2(n10204), .ZN(n8286) );
  NAND2_X1 U6667 ( .A1(n8291), .A2(n8286), .ZN(n8416) );
  INV_X1 U6668 ( .A(n8416), .ZN(n8285) );
  NAND2_X1 U6669 ( .A1(n5155), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5266) );
  NAND2_X1 U6670 ( .A1(n5177), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5265) );
  NAND2_X1 U6671 ( .A1(n5261), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5262) );
  NAND2_X1 U6672 ( .A1(n5283), .A2(n5262), .ZN(n7737) );
  NAND2_X1 U6673 ( .A1(n5526), .A2(n7737), .ZN(n5264) );
  NAND2_X1 U6674 ( .A1(n5178), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5263) );
  NAND4_X1 U6675 ( .A1(n5266), .A2(n5265), .A3(n5264), .A4(n5263), .ZN(n8664)
         );
  INV_X1 U6676 ( .A(n5269), .ZN(n5270) );
  NAND2_X1 U6677 ( .A1(n5270), .A2(SI_7_), .ZN(n5271) );
  INV_X1 U6678 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6740) );
  INV_X1 U6679 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6939) );
  MUX2_X1 U6680 ( .A(n6740), .B(n6939), .S(n5186), .Z(n5273) );
  INV_X1 U6681 ( .A(SI_8_), .ZN(n5272) );
  NAND2_X1 U6682 ( .A1(n5273), .A2(n5272), .ZN(n5289) );
  INV_X1 U6683 ( .A(n5273), .ZN(n5274) );
  NAND2_X1 U6684 ( .A1(n5274), .A2(SI_8_), .ZN(n5275) );
  XNOR2_X1 U6685 ( .A(n5291), .B(n4616), .ZN(n6739) );
  OR2_X1 U6686 ( .A1(n6739), .A2(n5296), .ZN(n5280) );
  OR2_X1 U6687 ( .A1(n5255), .A2(n9020), .ZN(n5277) );
  XNOR2_X1 U6688 ( .A(n5277), .B(n5276), .ZN(n10140) );
  INV_X1 U6689 ( .A(n10140), .ZN(n6644) );
  NAND2_X1 U6690 ( .A1(n5169), .A2(n6644), .ZN(n5279) );
  OR2_X1 U6691 ( .A1(n4422), .A2(n6740), .ZN(n5278) );
  OR2_X1 U6692 ( .A1(n8664), .A2(n10210), .ZN(n8292) );
  AND2_X1 U6693 ( .A1(n8664), .A2(n10210), .ZN(n8281) );
  INV_X1 U6694 ( .A(n8281), .ZN(n8287) );
  NAND2_X1 U6695 ( .A1(n8292), .A2(n8287), .ZN(n8415) );
  INV_X1 U6696 ( .A(n10204), .ZN(n7637) );
  OR2_X1 U6697 ( .A1(n8665), .A2(n7637), .ZN(n7732) );
  AND2_X1 U6698 ( .A1(n8415), .A2(n7732), .ZN(n5281) );
  INV_X1 U6699 ( .A(n10210), .ZN(n7695) );
  NAND2_X1 U6700 ( .A1(n8664), .A2(n7695), .ZN(n5282) );
  NAND2_X1 U6701 ( .A1(n5155), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5288) );
  NAND2_X1 U6702 ( .A1(n5177), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5287) );
  NAND2_X1 U6703 ( .A1(n5283), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5284) );
  NAND2_X1 U6704 ( .A1(n5333), .A2(n5284), .ZN(n7783) );
  NAND2_X1 U6705 ( .A1(n5526), .A2(n7783), .ZN(n5286) );
  NAND2_X1 U6706 ( .A1(n5178), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5285) );
  NAND4_X1 U6707 ( .A1(n5288), .A2(n5287), .A3(n5286), .A4(n5285), .ZN(n8663)
         );
  INV_X1 U6708 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n7015) );
  INV_X1 U6709 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n7017) );
  MUX2_X1 U6710 ( .A(n7015), .B(n7017), .S(n4587), .Z(n5293) );
  INV_X1 U6711 ( .A(SI_9_), .ZN(n5292) );
  INV_X1 U6712 ( .A(n5293), .ZN(n5294) );
  NAND2_X1 U6713 ( .A1(n5294), .A2(SI_9_), .ZN(n5295) );
  XNOR2_X1 U6714 ( .A(n5302), .B(n5011), .ZN(n7014) );
  NAND2_X1 U6715 ( .A1(n7014), .A2(n8396), .ZN(n5300) );
  NAND2_X1 U6716 ( .A1(n5297), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5298) );
  XNOR2_X1 U6717 ( .A(n5298), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6625) );
  AOI22_X1 U6718 ( .A1(n5493), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5169), .B2(
        n6625), .ZN(n5299) );
  AND2_X1 U6719 ( .A1(n8663), .A2(n10215), .ZN(n5301) );
  NAND2_X1 U6720 ( .A1(n5302), .A2(n5011), .ZN(n5304) );
  INV_X1 U6721 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n7019) );
  INV_X1 U6722 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n7022) );
  MUX2_X1 U6723 ( .A(n7019), .B(n7022), .S(n4587), .Z(n5318) );
  XNOR2_X1 U6724 ( .A(n5322), .B(n5317), .ZN(n7018) );
  NAND2_X1 U6725 ( .A1(n7018), .A2(n8396), .ZN(n5309) );
  NAND2_X1 U6726 ( .A1(n5305), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5306) );
  MUX2_X1 U6727 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5306), .S(
        P2_IR_REG_10__SCAN_IN), .Z(n5307) );
  NAND2_X1 U6728 ( .A1(n5307), .A2(n5326), .ZN(n7020) );
  INV_X1 U6729 ( .A(n7020), .ZN(n7704) );
  AOI22_X1 U6730 ( .A1(n5493), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5169), .B2(
        n7704), .ZN(n5308) );
  NAND2_X1 U6731 ( .A1(n5309), .A2(n5308), .ZN(n7797) );
  NAND2_X1 U6732 ( .A1(n5155), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5314) );
  NAND2_X1 U6733 ( .A1(n5177), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5313) );
  XNOR2_X1 U6734 ( .A(n5333), .B(P2_REG3_REG_10__SCAN_IN), .ZN(n7904) );
  NAND2_X1 U6735 ( .A1(n5526), .A2(n7904), .ZN(n5312) );
  NAND2_X1 U6736 ( .A1(n5178), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5311) );
  INV_X1 U6737 ( .A(n8620), .ZN(n8662) );
  NOR2_X1 U6738 ( .A1(n7797), .A2(n8662), .ZN(n5316) );
  NAND2_X1 U6739 ( .A1(n7797), .A2(n8662), .ZN(n5315) );
  INV_X1 U6740 ( .A(n5318), .ZN(n5319) );
  INV_X1 U6741 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7075) );
  INV_X1 U6742 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n7072) );
  MUX2_X1 U6743 ( .A(n7075), .B(n7072), .S(n4587), .Z(n5323) );
  INV_X1 U6744 ( .A(SI_11_), .ZN(n6846) );
  INV_X1 U6745 ( .A(n5323), .ZN(n5324) );
  NAND2_X1 U6746 ( .A1(n5324), .A2(SI_11_), .ZN(n5325) );
  XNOR2_X1 U6747 ( .A(n5343), .B(n5342), .ZN(n7071) );
  NAND2_X1 U6748 ( .A1(n7071), .A2(n8396), .ZN(n5332) );
  NAND2_X1 U6749 ( .A1(n5326), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5329) );
  INV_X1 U6750 ( .A(n5329), .ZN(n5327) );
  NAND2_X1 U6751 ( .A1(n5327), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n5330) );
  NAND2_X1 U6752 ( .A1(n5329), .A2(n5328), .ZN(n5344) );
  AND2_X1 U6753 ( .A1(n5330), .A2(n5344), .ZN(n7993) );
  AOI22_X1 U6754 ( .A1(n5493), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5169), .B2(
        n7993), .ZN(n5331) );
  NAND2_X1 U6755 ( .A1(n5155), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5338) );
  NAND2_X1 U6756 ( .A1(n5177), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5337) );
  OAI21_X1 U6757 ( .B1(n5333), .B2(P2_REG3_REG_10__SCAN_IN), .A(
        P2_REG3_REG_11__SCAN_IN), .ZN(n5334) );
  NAND2_X1 U6758 ( .A1(n5334), .A2(n5348), .ZN(n8625) );
  NAND2_X1 U6759 ( .A1(n5526), .A2(n8625), .ZN(n5336) );
  NAND2_X1 U6760 ( .A1(n5178), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5335) );
  NAND2_X1 U6761 ( .A1(n8624), .A2(n7951), .ZN(n8306) );
  NAND2_X1 U6762 ( .A1(n7893), .A2(n7892), .ZN(n5340) );
  INV_X1 U6763 ( .A(n7951), .ZN(n8661) );
  NAND2_X1 U6764 ( .A1(n8624), .A2(n8661), .ZN(n5339) );
  INV_X1 U6765 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7131) );
  INV_X1 U6766 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7137) );
  MUX2_X1 U6767 ( .A(n7131), .B(n7137), .S(n4587), .Z(n5363) );
  XNOR2_X1 U6768 ( .A(n5367), .B(n5362), .ZN(n7130) );
  NAND2_X1 U6769 ( .A1(n7130), .A2(n8396), .ZN(n5347) );
  NAND2_X1 U6770 ( .A1(n5344), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5345) );
  XNOR2_X1 U6771 ( .A(n5345), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6622) );
  AOI22_X1 U6772 ( .A1(n5493), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5169), .B2(
        n6622), .ZN(n5346) );
  NAND2_X1 U6773 ( .A1(n5155), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5353) );
  NAND2_X1 U6774 ( .A1(n5177), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5352) );
  NAND2_X1 U6775 ( .A1(n5348), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5349) );
  NAND2_X1 U6776 ( .A1(n5356), .A2(n5349), .ZN(n7958) );
  NAND2_X1 U6777 ( .A1(n5526), .A2(n7958), .ZN(n5351) );
  NAND2_X1 U6778 ( .A1(n5178), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5350) );
  AND2_X1 U6779 ( .A1(n10232), .A2(n8660), .ZN(n5355) );
  NAND2_X1 U6780 ( .A1(n5177), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U6781 ( .A1(n5178), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5360) );
  NAND2_X1 U6782 ( .A1(n5356), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5357) );
  NAND2_X1 U6783 ( .A1(n5380), .A2(n5357), .ZN(n8032) );
  NAND2_X1 U6784 ( .A1(n5526), .A2(n8032), .ZN(n5359) );
  NAND2_X1 U6785 ( .A1(n5155), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5358) );
  INV_X1 U6786 ( .A(n5363), .ZN(n5364) );
  NAND2_X1 U6787 ( .A1(n5364), .A2(SI_12_), .ZN(n5365) );
  MUX2_X1 U6788 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n4587), .Z(n5375) );
  XNOR2_X1 U6789 ( .A(n5375), .B(SI_13_), .ZN(n5373) );
  NAND2_X1 U6790 ( .A1(n7138), .A2(n8396), .ZN(n5371) );
  OR2_X1 U6791 ( .A1(n5368), .A2(n9020), .ZN(n5369) );
  XNOR2_X1 U6792 ( .A(n5369), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8186) );
  AOI22_X1 U6793 ( .A1(n5493), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5169), .B2(
        n8186), .ZN(n5370) );
  INV_X1 U6794 ( .A(n7952), .ZN(n5372) );
  NAND2_X1 U6795 ( .A1(n5375), .A2(SI_13_), .ZN(n5441) );
  NAND2_X1 U6796 ( .A1(n5442), .A2(n5441), .ZN(n5406) );
  MUX2_X1 U6797 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n4587), .Z(n5388) );
  XNOR2_X1 U6798 ( .A(n5388), .B(SI_14_), .ZN(n5387) );
  XNOR2_X1 U6799 ( .A(n5406), .B(n5387), .ZN(n7262) );
  NAND2_X1 U6800 ( .A1(n7262), .A2(n8396), .ZN(n5379) );
  NAND2_X1 U6801 ( .A1(n4509), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5416) );
  NAND2_X1 U6802 ( .A1(n5416), .A2(n5376), .ZN(n5392) );
  OR2_X1 U6803 ( .A1(n5416), .A2(n5376), .ZN(n5377) );
  AND2_X1 U6804 ( .A1(n5392), .A2(n5377), .ZN(n6618) );
  AOI22_X1 U6805 ( .A1(n5493), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5169), .B2(
        n6618), .ZN(n5378) );
  NAND2_X1 U6806 ( .A1(n5177), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5385) );
  NAND2_X1 U6807 ( .A1(n5380), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5381) );
  NAND2_X1 U6808 ( .A1(n5396), .A2(n5381), .ZN(n8103) );
  NAND2_X1 U6809 ( .A1(n5179), .A2(n8103), .ZN(n5384) );
  NAND2_X1 U6810 ( .A1(n5178), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5383) );
  NAND2_X1 U6811 ( .A1(n5155), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5382) );
  INV_X1 U6812 ( .A(n8123), .ZN(n8659) );
  OR2_X1 U6813 ( .A1(n8114), .A2(n8659), .ZN(n5386) );
  NAND2_X1 U6814 ( .A1(n5406), .A2(n5405), .ZN(n5389) );
  NAND2_X1 U6815 ( .A1(n5388), .A2(SI_14_), .ZN(n5409) );
  NAND2_X1 U6816 ( .A1(n5389), .A2(n5409), .ZN(n5391) );
  MUX2_X1 U6817 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n4587), .Z(n5404) );
  XNOR2_X1 U6818 ( .A(n5404), .B(SI_15_), .ZN(n5390) );
  NAND2_X1 U6819 ( .A1(n7312), .A2(n8396), .ZN(n5395) );
  NAND2_X1 U6820 ( .A1(n5392), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5393) );
  XNOR2_X1 U6821 ( .A(n5393), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8679) );
  AOI22_X1 U6822 ( .A1(n5493), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5169), .B2(
        n8679), .ZN(n5394) );
  NAND2_X1 U6823 ( .A1(n5177), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5401) );
  NAND2_X1 U6824 ( .A1(n5155), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5400) );
  NAND2_X1 U6825 ( .A1(n5396), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U6826 ( .A1(n5421), .A2(n5397), .ZN(n8155) );
  NAND2_X1 U6827 ( .A1(n5526), .A2(n8155), .ZN(n5399) );
  NAND2_X1 U6828 ( .A1(n5178), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5398) );
  NOR2_X1 U6829 ( .A1(n8941), .A2(n8892), .ZN(n5403) );
  NAND2_X1 U6830 ( .A1(n8941), .A2(n8892), .ZN(n5402) );
  INV_X1 U6831 ( .A(SI_15_), .ZN(n6808) );
  NAND2_X1 U6832 ( .A1(n5408), .A2(n6808), .ZN(n5407) );
  NAND2_X1 U6833 ( .A1(n5406), .A2(n5444), .ZN(n5412) );
  INV_X1 U6834 ( .A(n5407), .ZN(n5411) );
  MUX2_X1 U6835 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n4587), .Z(n5434) );
  INV_X1 U6836 ( .A(SI_16_), .ZN(n5440) );
  XNOR2_X1 U6837 ( .A(n5434), .B(n5440), .ZN(n5413) );
  NAND2_X1 U6838 ( .A1(n7305), .A2(n8396), .ZN(n5420) );
  OAI21_X1 U6839 ( .B1(P2_IR_REG_14__SCAN_IN), .B2(P2_IR_REG_15__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5415) );
  NAND2_X1 U6840 ( .A1(n5416), .A2(n5415), .ZN(n5417) );
  OR2_X1 U6841 ( .A1(n5417), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5455) );
  NAND2_X1 U6842 ( .A1(n5417), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5418) );
  AND2_X1 U6843 ( .A1(n5455), .A2(n5418), .ZN(n8698) );
  AOI22_X1 U6844 ( .A1(n5493), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5169), .B2(
        n8698), .ZN(n5419) );
  NAND2_X1 U6845 ( .A1(n5155), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5426) );
  NAND2_X1 U6846 ( .A1(n5176), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5425) );
  NAND2_X1 U6847 ( .A1(n5421), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5422) );
  NAND2_X1 U6848 ( .A1(n5459), .A2(n5422), .ZN(n8896) );
  NAND2_X1 U6849 ( .A1(n5526), .A2(n8896), .ZN(n5424) );
  NAND2_X1 U6850 ( .A1(n5178), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5423) );
  INV_X1 U6851 ( .A(n8873), .ZN(n5427) );
  NAND2_X1 U6852 ( .A1(n8874), .A2(n5427), .ZN(n8886) );
  NAND2_X1 U6853 ( .A1(n8888), .A2(n8886), .ZN(n5429) );
  INV_X1 U6854 ( .A(n8227), .ZN(n8880) );
  NAND2_X1 U6855 ( .A1(n9010), .A2(n8880), .ZN(n5428) );
  INV_X1 U6856 ( .A(n5434), .ZN(n5431) );
  NAND2_X1 U6857 ( .A1(n5442), .A2(n5432), .ZN(n5438) );
  INV_X1 U6858 ( .A(n5433), .ZN(n5436) );
  AND2_X1 U6859 ( .A1(n5444), .A2(n5434), .ZN(n5435) );
  NAND2_X1 U6860 ( .A1(n5438), .A2(n5437), .ZN(n5450) );
  INV_X1 U6861 ( .A(n5443), .ZN(n5446) );
  NAND2_X1 U6862 ( .A1(n5448), .A2(n5447), .ZN(n5449) );
  NAND2_X1 U6863 ( .A1(n5450), .A2(n5449), .ZN(n5469) );
  INV_X1 U6864 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7295) );
  INV_X1 U6865 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7297) );
  MUX2_X1 U6866 ( .A(n7295), .B(n7297), .S(n4587), .Z(n5452) );
  INV_X1 U6867 ( .A(SI_17_), .ZN(n5451) );
  NAND2_X1 U6868 ( .A1(n5452), .A2(n5451), .ZN(n5467) );
  INV_X1 U6869 ( .A(n5452), .ZN(n5453) );
  NAND2_X1 U6870 ( .A1(n5453), .A2(SI_17_), .ZN(n5454) );
  NAND2_X1 U6871 ( .A1(n5467), .A2(n5454), .ZN(n5468) );
  XNOR2_X1 U6872 ( .A(n5469), .B(n5468), .ZN(n7294) );
  NAND2_X1 U6873 ( .A1(n7294), .A2(n8396), .ZN(n5458) );
  NAND2_X1 U6874 ( .A1(n5455), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5456) );
  XNOR2_X1 U6875 ( .A(n5456), .B(P2_IR_REG_17__SCAN_IN), .ZN(n6614) );
  AOI22_X1 U6876 ( .A1(n5493), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5169), .B2(
        n6614), .ZN(n5457) );
  NAND2_X1 U6877 ( .A1(n5177), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5464) );
  NAND2_X1 U6878 ( .A1(n5178), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5463) );
  NAND2_X1 U6879 ( .A1(n5459), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5460) );
  NAND2_X1 U6880 ( .A1(n5476), .A2(n5460), .ZN(n8883) );
  NAND2_X1 U6881 ( .A1(n5526), .A2(n8883), .ZN(n5462) );
  NAND2_X1 U6882 ( .A1(n5155), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5461) );
  NAND2_X1 U6883 ( .A1(n9003), .A2(n8866), .ZN(n8428) );
  NAND2_X1 U6884 ( .A1(n8327), .A2(n8428), .ZN(n8878) );
  INV_X1 U6885 ( .A(n8866), .ZN(n8890) );
  NAND2_X1 U6886 ( .A1(n9003), .A2(n8890), .ZN(n5465) );
  INV_X1 U6887 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7332) );
  INV_X1 U6888 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5470) );
  MUX2_X1 U6889 ( .A(n7332), .B(n5470), .S(n4587), .Z(n5484) );
  XNOR2_X1 U6890 ( .A(n5484), .B(SI_18_), .ZN(n5483) );
  XNOR2_X1 U6891 ( .A(n5488), .B(n5483), .ZN(n7318) );
  NAND2_X1 U6892 ( .A1(n7318), .A2(n8396), .ZN(n5475) );
  NAND2_X1 U6893 ( .A1(n4510), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5471) );
  MUX2_X1 U6894 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5471), .S(
        P2_IR_REG_18__SCAN_IN), .Z(n5472) );
  INV_X1 U6895 ( .A(n5472), .ZN(n5473) );
  NOR2_X1 U6896 ( .A1(n5473), .A2(n5058), .ZN(n8734) );
  AOI22_X1 U6897 ( .A1(n5493), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5169), .B2(
        n8734), .ZN(n5474) );
  NAND2_X1 U6898 ( .A1(n5155), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5481) );
  NAND2_X1 U6899 ( .A1(n5176), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5480) );
  NAND2_X1 U6900 ( .A1(n5476), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5477) );
  NAND2_X1 U6901 ( .A1(n5496), .A2(n5477), .ZN(n8867) );
  NAND2_X1 U6902 ( .A1(n5526), .A2(n8867), .ZN(n5479) );
  NAND2_X1 U6903 ( .A1(n5178), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5478) );
  AND2_X1 U6904 ( .A1(n8930), .A2(n8879), .ZN(n5482) );
  INV_X1 U6905 ( .A(n5484), .ZN(n5485) );
  NAND2_X1 U6906 ( .A1(n5485), .A2(SI_18_), .ZN(n5486) );
  OAI21_X1 U6907 ( .B1(n5488), .B2(n5487), .A(n5486), .ZN(n5505) );
  INV_X1 U6908 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7410) );
  INV_X1 U6909 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8473) );
  MUX2_X1 U6910 ( .A(n7410), .B(n8473), .S(n4587), .Z(n5490) );
  INV_X1 U6911 ( .A(SI_19_), .ZN(n5489) );
  NAND2_X1 U6912 ( .A1(n5490), .A2(n5489), .ZN(n5503) );
  INV_X1 U6913 ( .A(n5490), .ZN(n5491) );
  NAND2_X1 U6914 ( .A1(n5491), .A2(SI_19_), .ZN(n5492) );
  NAND2_X1 U6915 ( .A1(n5503), .A2(n5492), .ZN(n5504) );
  XNOR2_X1 U6916 ( .A(n5505), .B(n5504), .ZN(n7408) );
  NAND2_X1 U6917 ( .A1(n7408), .A2(n8396), .ZN(n5495) );
  AOI22_X1 U6918 ( .A1(n5493), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5637), .B2(
        n5169), .ZN(n5494) );
  NAND2_X1 U6919 ( .A1(n5155), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5501) );
  NAND2_X1 U6920 ( .A1(n5176), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5500) );
  NAND2_X1 U6921 ( .A1(n5496), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5497) );
  NAND2_X1 U6922 ( .A1(n5509), .A2(n5497), .ZN(n8851) );
  NAND2_X1 U6923 ( .A1(n5526), .A2(n8851), .ZN(n5499) );
  NAND2_X1 U6924 ( .A1(n5178), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5498) );
  NAND2_X1 U6925 ( .A1(n8993), .A2(n8865), .ZN(n8332) );
  INV_X1 U6926 ( .A(n8865), .ZN(n8658) );
  NAND2_X1 U6927 ( .A1(n8993), .A2(n8658), .ZN(n5502) );
  INV_X1 U6928 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7433) );
  INV_X1 U6929 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7538) );
  MUX2_X1 U6930 ( .A(n7433), .B(n7538), .S(n4587), .Z(n5516) );
  XNOR2_X1 U6931 ( .A(n5516), .B(SI_20_), .ZN(n5506) );
  XNOR2_X1 U6932 ( .A(n5518), .B(n5506), .ZN(n7432) );
  NAND2_X1 U6933 ( .A1(n7432), .A2(n8396), .ZN(n5508) );
  OR2_X1 U6934 ( .A1(n4422), .A2(n7433), .ZN(n5507) );
  NAND2_X1 U6935 ( .A1(n5155), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5514) );
  NAND2_X1 U6936 ( .A1(n5177), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5513) );
  NAND2_X1 U6937 ( .A1(n5509), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5510) );
  NAND2_X1 U6938 ( .A1(n5524), .A2(n5510), .ZN(n8837) );
  NAND2_X1 U6939 ( .A1(n5179), .A2(n8837), .ZN(n5512) );
  NAND2_X1 U6940 ( .A1(n5178), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5511) );
  NAND2_X1 U6941 ( .A1(n8836), .A2(n8822), .ZN(n8814) );
  INV_X1 U6942 ( .A(n8822), .ZN(n8848) );
  NAND2_X1 U6943 ( .A1(n8830), .A2(n5515), .ZN(n8818) );
  INV_X1 U6944 ( .A(SI_20_), .ZN(n5517) );
  NAND2_X1 U6945 ( .A1(n5518), .A2(n5517), .ZN(n5519) );
  INV_X1 U6946 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n8550) );
  INV_X1 U6947 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7586) );
  MUX2_X1 U6948 ( .A(n8550), .B(n7586), .S(n5186), .Z(n5533) );
  XNOR2_X1 U6949 ( .A(n5533), .B(SI_21_), .ZN(n5521) );
  XNOR2_X1 U6950 ( .A(n5536), .B(n5521), .ZN(n7585) );
  NAND2_X1 U6951 ( .A1(n7585), .A2(n8396), .ZN(n5523) );
  OR2_X1 U6952 ( .A1(n4421), .A2(n8550), .ZN(n5522) );
  NAND2_X1 U6953 ( .A1(n5176), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5530) );
  NAND2_X1 U6954 ( .A1(n5178), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5529) );
  NAND2_X1 U6955 ( .A1(n5524), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5525) );
  NAND2_X1 U6956 ( .A1(n5543), .A2(n5525), .ZN(n8825) );
  NAND2_X1 U6957 ( .A1(n5526), .A2(n8825), .ZN(n5528) );
  NAND2_X1 U6958 ( .A1(n5155), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5527) );
  NAND2_X1 U6959 ( .A1(n8826), .A2(n8835), .ZN(n8340) );
  NAND2_X1 U6960 ( .A1(n8341), .A2(n8340), .ZN(n8816) );
  NAND2_X1 U6961 ( .A1(n8818), .A2(n8816), .ZN(n5532) );
  NAND2_X1 U6962 ( .A1(n5532), .A2(n5531), .ZN(n8805) );
  INV_X1 U6963 ( .A(n5533), .ZN(n5534) );
  NAND2_X1 U6964 ( .A1(n5534), .A2(SI_21_), .ZN(n5535) );
  INV_X1 U6965 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7857) );
  INV_X1 U6966 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7855) );
  MUX2_X1 U6967 ( .A(n7857), .B(n7855), .S(n4587), .Z(n5538) );
  INV_X1 U6968 ( .A(SI_22_), .ZN(n5537) );
  NAND2_X1 U6969 ( .A1(n5538), .A2(n5537), .ZN(n5551) );
  INV_X1 U6970 ( .A(n5538), .ZN(n5539) );
  NAND2_X1 U6971 ( .A1(n5539), .A2(SI_22_), .ZN(n5540) );
  NAND2_X1 U6972 ( .A1(n5551), .A2(n5540), .ZN(n5552) );
  XNOR2_X1 U6973 ( .A(n5553), .B(n5552), .ZN(n7853) );
  NAND2_X1 U6974 ( .A1(n7853), .A2(n8396), .ZN(n5542) );
  OR2_X1 U6975 ( .A1(n4421), .A2(n7857), .ZN(n5541) );
  NAND2_X1 U6976 ( .A1(n5543), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5544) );
  NAND2_X1 U6977 ( .A1(n5563), .A2(n5544), .ZN(n8811) );
  NAND2_X1 U6978 ( .A1(n8811), .A2(n5179), .ZN(n5548) );
  NAND2_X1 U6979 ( .A1(n5177), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5547) );
  NAND2_X1 U6980 ( .A1(n5178), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5546) );
  NAND2_X1 U6981 ( .A1(n5155), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5545) );
  NAND2_X1 U6982 ( .A1(n8977), .A2(n8821), .ZN(n8345) );
  NAND2_X1 U6983 ( .A1(n8805), .A2(n8806), .ZN(n5550) );
  INV_X1 U6984 ( .A(n8821), .ZN(n8657) );
  INV_X1 U6985 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7916) );
  INV_X1 U6986 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7912) );
  MUX2_X1 U6987 ( .A(n7916), .B(n7912), .S(n4587), .Z(n5555) );
  INV_X1 U6988 ( .A(SI_23_), .ZN(n5554) );
  NAND2_X1 U6989 ( .A1(n5555), .A2(n5554), .ZN(n5569) );
  INV_X1 U6990 ( .A(n5555), .ZN(n5556) );
  NAND2_X1 U6991 ( .A1(n5556), .A2(SI_23_), .ZN(n5557) );
  AND2_X1 U6992 ( .A1(n5569), .A2(n5557), .ZN(n5558) );
  OR2_X1 U6993 ( .A1(n5559), .A2(n5558), .ZN(n5560) );
  NAND2_X1 U6994 ( .A1(n5570), .A2(n5560), .ZN(n7913) );
  NAND2_X1 U6995 ( .A1(n7913), .A2(n8396), .ZN(n5562) );
  OR2_X1 U6996 ( .A1(n4421), .A2(n7916), .ZN(n5561) );
  INV_X1 U6997 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8799) );
  NAND2_X1 U6998 ( .A1(n5563), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5564) );
  NAND2_X1 U6999 ( .A1(n5577), .A2(n5564), .ZN(n8800) );
  NAND2_X1 U7000 ( .A1(n8800), .A2(n5179), .ZN(n5566) );
  AOI22_X1 U7001 ( .A1(n5155), .A2(P2_REG0_REG_23__SCAN_IN), .B1(n5176), .B2(
        P2_REG1_REG_23__SCAN_IN), .ZN(n5565) );
  NOR2_X1 U7002 ( .A1(n8801), .A2(n8808), .ZN(n5568) );
  NAND2_X1 U7003 ( .A1(n8801), .A2(n8808), .ZN(n5567) );
  INV_X1 U7004 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7982) );
  INV_X1 U7005 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8025) );
  MUX2_X1 U7006 ( .A(n7982), .B(n8025), .S(n5186), .Z(n5572) );
  INV_X1 U7007 ( .A(SI_24_), .ZN(n5571) );
  NAND2_X1 U7008 ( .A1(n5572), .A2(n5571), .ZN(n5585) );
  INV_X1 U7009 ( .A(n5572), .ZN(n5573) );
  NAND2_X1 U7010 ( .A1(n5573), .A2(SI_24_), .ZN(n5574) );
  AND2_X1 U7011 ( .A1(n5585), .A2(n5574), .ZN(n5583) );
  XNOR2_X1 U7012 ( .A(n5584), .B(n5583), .ZN(n7981) );
  NAND2_X1 U7013 ( .A1(n7981), .A2(n8396), .ZN(n5576) );
  OR2_X1 U7014 ( .A1(n4422), .A2(n7982), .ZN(n5575) );
  NAND2_X1 U7015 ( .A1(n5577), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5578) );
  NAND2_X1 U7016 ( .A1(n5593), .A2(n5578), .ZN(n8790) );
  NAND2_X1 U7017 ( .A1(n8790), .A2(n5179), .ZN(n5581) );
  AOI22_X1 U7018 ( .A1(n5155), .A2(P2_REG0_REG_24__SCAN_IN), .B1(n5177), .B2(
        P2_REG1_REG_24__SCAN_IN), .ZN(n5580) );
  NAND2_X1 U7019 ( .A1(n5178), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5579) );
  NAND2_X1 U7020 ( .A1(n5584), .A2(n5583), .ZN(n5586) );
  INV_X1 U7021 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8057) );
  INV_X1 U7022 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8059) );
  MUX2_X1 U7023 ( .A(n8057), .B(n8059), .S(n5186), .Z(n5588) );
  INV_X1 U7024 ( .A(SI_25_), .ZN(n5587) );
  NAND2_X1 U7025 ( .A1(n5588), .A2(n5587), .ZN(n5606) );
  INV_X1 U7026 ( .A(n5588), .ZN(n5589) );
  NAND2_X1 U7027 ( .A1(n5589), .A2(SI_25_), .ZN(n5590) );
  AND2_X1 U7028 ( .A1(n5606), .A2(n5590), .ZN(n5604) );
  NAND2_X1 U7029 ( .A1(n8056), .A2(n8396), .ZN(n5592) );
  OR2_X1 U7030 ( .A1(n4422), .A2(n8057), .ZN(n5591) );
  NAND2_X1 U7031 ( .A1(n5593), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5594) );
  NAND2_X1 U7032 ( .A1(n5595), .A2(n5594), .ZN(n8776) );
  NAND2_X1 U7033 ( .A1(n8776), .A2(n5179), .ZN(n5601) );
  INV_X1 U7034 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n5598) );
  NAND2_X1 U7035 ( .A1(n5155), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5597) );
  NAND2_X1 U7036 ( .A1(n5176), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5596) );
  OAI211_X1 U7037 ( .C1(n5598), .C2(n4529), .A(n5597), .B(n5596), .ZN(n5599)
         );
  INV_X1 U7038 ( .A(n5599), .ZN(n5600) );
  INV_X1 U7039 ( .A(n8236), .ZN(n8358) );
  INV_X1 U7040 ( .A(n8783), .ZN(n5602) );
  INV_X1 U7041 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8083) );
  INV_X1 U7042 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8098) );
  MUX2_X1 U7043 ( .A(n8083), .B(n8098), .S(n5186), .Z(n5608) );
  INV_X1 U7044 ( .A(SI_26_), .ZN(n6849) );
  NAND2_X1 U7045 ( .A1(n5608), .A2(n6849), .ZN(n5677) );
  INV_X1 U7046 ( .A(n5608), .ZN(n5609) );
  NAND2_X1 U7047 ( .A1(n5609), .A2(SI_26_), .ZN(n5610) );
  AND2_X1 U7048 ( .A1(n5677), .A2(n5610), .ZN(n5675) );
  OR2_X1 U7049 ( .A1(n4422), .A2(n8083), .ZN(n5611) );
  NAND2_X1 U7050 ( .A1(n8642), .A2(n5179), .ZN(n5617) );
  INV_X1 U7051 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n5614) );
  NAND2_X1 U7052 ( .A1(n5176), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U7053 ( .A1(n5155), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5612) );
  OAI211_X1 U7054 ( .C1(n4529), .C2(n5614), .A(n5613), .B(n5612), .ZN(n5615)
         );
  INV_X1 U7055 ( .A(n5615), .ZN(n5616) );
  AND2_X2 U7056 ( .A1(n5617), .A2(n5616), .ZN(n8774) );
  NAND2_X1 U7057 ( .A1(n5618), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5619) );
  NAND2_X1 U7058 ( .A1(n8749), .A2(n5619), .ZN(n8556) );
  NAND2_X1 U7059 ( .A1(n8556), .A2(n5179), .ZN(n5624) );
  INV_X1 U7060 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n6829) );
  NAND2_X1 U7061 ( .A1(n5178), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5621) );
  NAND2_X1 U7062 ( .A1(n5177), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5620) );
  OAI211_X1 U7063 ( .C1(n5310), .C2(n6829), .A(n5621), .B(n5620), .ZN(n5622)
         );
  INV_X1 U7064 ( .A(n5622), .ZN(n5623) );
  INV_X1 U7065 ( .A(n5110), .ZN(n8461) );
  INV_X1 U7066 ( .A(n8460), .ZN(n6611) );
  NAND2_X1 U7067 ( .A1(n8461), .A2(n6611), .ZN(n5625) );
  NAND2_X1 U7068 ( .A1(n5134), .A2(n5625), .ZN(n5845) );
  NAND2_X2 U7069 ( .A1(n5753), .A2(n8464), .ZN(n8399) );
  INV_X1 U7070 ( .A(n5845), .ZN(n5847) );
  INV_X1 U7071 ( .A(n8891), .ZN(n5626) );
  INV_X1 U7072 ( .A(n5629), .ZN(n8953) );
  OAI21_X1 U7073 ( .B1(n5630), .B2(n10165), .A(n8953), .ZN(n5650) );
  XNOR2_X1 U7074 ( .A(n7983), .B(P2_B_REG_SCAN_IN), .ZN(n5633) );
  INV_X1 U7075 ( .A(n5631), .ZN(n8058) );
  INV_X1 U7076 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6733) );
  NAND2_X1 U7077 ( .A1(n6724), .A2(n6733), .ZN(n5635) );
  NAND2_X1 U7078 ( .A1(n5632), .A2(n7983), .ZN(n6730) );
  INV_X1 U7079 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6729) );
  NAND2_X1 U7080 ( .A1(n6724), .A2(n6729), .ZN(n5636) );
  NAND2_X1 U7081 ( .A1(n5632), .A2(n8058), .ZN(n6727) );
  AND2_X1 U7082 ( .A1(n5636), .A2(n6727), .ZN(n5722) );
  NAND2_X1 U7083 ( .A1(n7409), .A2(n8464), .ZN(n5662) );
  OR2_X1 U7084 ( .A1(n5754), .A2(n5662), .ZN(n5638) );
  AND2_X1 U7085 ( .A1(n8399), .A2(n5638), .ZN(n5721) );
  MUX2_X1 U7086 ( .A(n5751), .B(n5722), .S(n5721), .Z(n5649) );
  OR2_X1 U7087 ( .A1(n8399), .A2(n5752), .ZN(n5852) );
  NOR4_X1 U7088 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n6802) );
  NOR2_X1 U7089 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .ZN(
        n5641) );
  NOR4_X1 U7090 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_31__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n5640) );
  NOR4_X1 U7091 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n5639) );
  NAND4_X1 U7092 ( .A1(n6802), .A2(n5641), .A3(n5640), .A4(n5639), .ZN(n5647)
         );
  NOR4_X1 U7093 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n5645) );
  NOR4_X1 U7094 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n5644) );
  NOR4_X1 U7095 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n5643) );
  NOR4_X1 U7096 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n5642) );
  NAND4_X1 U7097 ( .A1(n5645), .A2(n5644), .A3(n5643), .A4(n5642), .ZN(n5646)
         );
  OAI21_X1 U7098 ( .B1(n5647), .B2(n5646), .A(n6724), .ZN(n5737) );
  AND3_X1 U7099 ( .A1(n5852), .A2(n6726), .A3(n5737), .ZN(n5648) );
  NAND2_X1 U7100 ( .A1(n5751), .A2(n5722), .ZN(n5738) );
  AND2_X1 U7101 ( .A1(n5648), .A2(n5738), .ZN(n5727) );
  NAND2_X1 U7102 ( .A1(n5649), .A2(n5727), .ZN(n5668) );
  NAND2_X1 U7103 ( .A1(n5650), .A2(n10174), .ZN(n5673) );
  INV_X1 U7104 ( .A(n8408), .ZN(n5652) );
  INV_X1 U7105 ( .A(n8250), .ZN(n5651) );
  NAND2_X1 U7106 ( .A1(n5652), .A2(n5651), .ZN(n7378) );
  NAND2_X1 U7107 ( .A1(n7378), .A2(n5653), .ZN(n10164) );
  NAND2_X1 U7108 ( .A1(n10164), .A2(n4543), .ZN(n10163) );
  NAND2_X1 U7109 ( .A1(n10163), .A2(n8258), .ZN(n7299) );
  NAND2_X1 U7110 ( .A1(n8669), .A2(n7869), .ZN(n8274) );
  NAND2_X1 U7111 ( .A1(n8264), .A2(n8274), .ZN(n7300) );
  INV_X1 U7112 ( .A(n7300), .ZN(n8412) );
  NAND2_X1 U7113 ( .A1(n7299), .A2(n8412), .ZN(n7298) );
  NAND2_X1 U7114 ( .A1(n8668), .A2(n10189), .ZN(n8265) );
  OR2_X1 U7115 ( .A1(n8668), .A2(n10189), .ZN(n8272) );
  NOR2_X1 U7116 ( .A1(n8667), .A2(n10194), .ZN(n8271) );
  NAND2_X1 U7117 ( .A1(n8667), .A2(n10194), .ZN(n8276) );
  OR2_X1 U7118 ( .A1(n8666), .A2(n10198), .ZN(n8277) );
  NAND2_X1 U7119 ( .A1(n8666), .A2(n10198), .ZN(n8279) );
  NAND2_X1 U7120 ( .A1(n8277), .A2(n8279), .ZN(n8414) );
  INV_X1 U7121 ( .A(n8277), .ZN(n8267) );
  NOR2_X1 U7122 ( .A1(n8416), .A2(n8267), .ZN(n5654) );
  NAND2_X1 U7123 ( .A1(n7624), .A2(n8286), .ZN(n7730) );
  OR2_X1 U7124 ( .A1(n8663), .A2(n7782), .ZN(n8293) );
  NAND2_X1 U7125 ( .A1(n8663), .A2(n7782), .ZN(n8288) );
  NAND2_X1 U7126 ( .A1(n8293), .A2(n8288), .ZN(n8283) );
  OR2_X1 U7127 ( .A1(n8620), .A2(n7797), .ZN(n8303) );
  NAND2_X1 U7128 ( .A1(n8620), .A2(n7797), .ZN(n8301) );
  NAND2_X1 U7129 ( .A1(n8303), .A2(n8301), .ZN(n8418) );
  NAND2_X1 U7130 ( .A1(n7896), .A2(n8419), .ZN(n7895) );
  OR2_X1 U7131 ( .A1(n10232), .A2(n8621), .ZN(n8309) );
  NAND2_X1 U7132 ( .A1(n10232), .A2(n8621), .ZN(n8310) );
  NAND2_X1 U7133 ( .A1(n7956), .A2(n8308), .ZN(n7955) );
  NAND2_X1 U7134 ( .A1(n7955), .A2(n8309), .ZN(n7974) );
  NOR2_X1 U7135 ( .A1(n9840), .A2(n7952), .ZN(n8314) );
  NAND2_X1 U7136 ( .A1(n9840), .A2(n7952), .ZN(n7973) );
  OR2_X1 U7137 ( .A1(n8114), .A2(n8123), .ZN(n8320) );
  NAND2_X1 U7138 ( .A1(n8106), .A2(n8320), .ZN(n5655) );
  NAND2_X1 U7139 ( .A1(n8114), .A2(n8123), .ZN(n8317) );
  OR2_X1 U7140 ( .A1(n8941), .A2(n8200), .ZN(n8318) );
  NAND2_X1 U7141 ( .A1(n8941), .A2(n8200), .ZN(n8322) );
  INV_X1 U7142 ( .A(n8428), .ZN(n5657) );
  OR2_X1 U7143 ( .A1(n8873), .A2(n5657), .ZN(n8855) );
  NAND2_X1 U7144 ( .A1(n8930), .A2(n5806), .ZN(n8407) );
  NAND2_X1 U7145 ( .A1(n8329), .A2(n8407), .ZN(n8862) );
  AND2_X1 U7146 ( .A1(n8327), .A2(n8874), .ZN(n5656) );
  OR2_X1 U7147 ( .A1(n5657), .A2(n5656), .ZN(n8856) );
  OR2_X1 U7148 ( .A1(n8862), .A2(n8856), .ZN(n8858) );
  AND2_X1 U7149 ( .A1(n8329), .A2(n8858), .ZN(n5658) );
  NAND2_X1 U7150 ( .A1(n8859), .A2(n5658), .ZN(n8845) );
  AND2_X1 U7151 ( .A1(n8340), .A2(n8814), .ZN(n8337) );
  NAND2_X1 U7152 ( .A1(n5659), .A2(n8341), .ZN(n8804) );
  NAND2_X1 U7153 ( .A1(n8804), .A2(n8345), .ZN(n5660) );
  INV_X1 U7154 ( .A(n8808), .ZN(n8785) );
  NAND2_X1 U7155 ( .A1(n8801), .A2(n8785), .ZN(n8404) );
  INV_X1 U7156 ( .A(n8464), .ZN(n8248) );
  NAND2_X1 U7157 ( .A1(n5750), .A2(n8248), .ZN(n10226) );
  INV_X1 U7158 ( .A(n5752), .ZN(n5664) );
  NAND2_X1 U7159 ( .A1(n5664), .A2(n5662), .ZN(n5663) );
  AND2_X1 U7160 ( .A1(n10226), .A2(n5663), .ZN(n5665) );
  OR2_X1 U7161 ( .A1(n8399), .A2(n5664), .ZN(n7576) );
  NAND2_X1 U7162 ( .A1(n5665), .A2(n7576), .ZN(n7777) );
  INV_X1 U7163 ( .A(n5666), .ZN(n5669) );
  AND2_X1 U7164 ( .A1(n5669), .A2(n5753), .ZN(n7626) );
  INV_X1 U7165 ( .A(n7626), .ZN(n5667) );
  NAND2_X1 U7166 ( .A1(n7777), .A2(n5667), .ZN(n10173) );
  INV_X1 U7167 ( .A(n5668), .ZN(n5670) );
  OR2_X1 U7168 ( .A1(n10226), .A2(n5669), .ZN(n10167) );
  INV_X1 U7169 ( .A(n10167), .ZN(n8104) );
  NAND2_X1 U7170 ( .A1(n5670), .A2(n8104), .ZN(n8839) );
  AOI22_X1 U7171 ( .A1(n8955), .A2(n8898), .B1(P2_REG2_REG_26__SCAN_IN), .B2(
        n10176), .ZN(n5671) );
  INV_X1 U7172 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5683) );
  INV_X1 U7173 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8148) );
  MUX2_X1 U7174 ( .A(n5683), .B(n8148), .S(n5186), .Z(n5680) );
  INV_X1 U7175 ( .A(SI_27_), .ZN(n5679) );
  NAND2_X1 U7176 ( .A1(n5680), .A2(n5679), .ZN(n5689) );
  INV_X1 U7177 ( .A(n5680), .ZN(n5681) );
  NAND2_X1 U7178 ( .A1(n5681), .A2(SI_27_), .ZN(n5682) );
  AND2_X1 U7179 ( .A1(n5689), .A2(n5682), .ZN(n5687) );
  OR2_X1 U7180 ( .A1(n4421), .A2(n5683), .ZN(n5684) );
  INV_X1 U7181 ( .A(n8246), .ZN(n5686) );
  INV_X1 U7182 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8162) );
  INV_X1 U7183 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8219) );
  MUX2_X1 U7184 ( .A(n8162), .B(n8219), .S(n4587), .Z(n6503) );
  XNOR2_X1 U7185 ( .A(n6503), .B(SI_28_), .ZN(n6500) );
  OR2_X1 U7186 ( .A1(n4422), .A2(n8162), .ZN(n5691) );
  XNOR2_X1 U7187 ( .A(n8749), .B(P2_REG3_REG_28__SCAN_IN), .ZN(n5862) );
  NAND2_X1 U7188 ( .A1(n5862), .A2(n5179), .ZN(n5697) );
  INV_X1 U7189 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n5712) );
  NAND2_X1 U7190 ( .A1(n5177), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5694) );
  NAND2_X1 U7191 ( .A1(n5155), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5693) );
  OAI211_X1 U7192 ( .C1(n5712), .C2(n4529), .A(n5694), .B(n5693), .ZN(n5695)
         );
  INV_X1 U7193 ( .A(n5695), .ZN(n5696) );
  XNOR2_X1 U7194 ( .A(n6499), .B(n8437), .ZN(n5698) );
  NAND2_X1 U7195 ( .A1(n5698), .A2(n8894), .ZN(n5709) );
  INV_X1 U7196 ( .A(n8749), .ZN(n5701) );
  NOR2_X1 U7197 ( .A1(n5699), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5700) );
  NAND2_X1 U7198 ( .A1(n5701), .A2(n5700), .ZN(n7521) );
  INV_X1 U7199 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n6877) );
  NAND2_X1 U7200 ( .A1(n5177), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5703) );
  NAND2_X1 U7201 ( .A1(n5155), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5702) );
  OAI211_X1 U7202 ( .C1(n6877), .C2(n4529), .A(n5703), .B(n5702), .ZN(n5704)
         );
  INV_X1 U7203 ( .A(n5704), .ZN(n5705) );
  NOR2_X1 U7204 ( .A1(n8234), .A2(n10171), .ZN(n5706) );
  NAND2_X1 U7205 ( .A1(n5709), .A2(n5708), .ZN(n6698) );
  INV_X1 U7206 ( .A(n6698), .ZN(n5718) );
  XNOR2_X1 U7207 ( .A(n6511), .B(n8437), .ZN(n6701) );
  INV_X1 U7208 ( .A(n6701), .ZN(n5716) );
  AOI22_X1 U7209 ( .A1(n8378), .A2(n8898), .B1(n5862), .B2(n8897), .ZN(n5713)
         );
  NAND2_X1 U7210 ( .A1(n5751), .A2(n5719), .ZN(n5720) );
  NAND2_X1 U7211 ( .A1(n5720), .A2(n5721), .ZN(n5725) );
  INV_X1 U7212 ( .A(n5721), .ZN(n5723) );
  INV_X1 U7213 ( .A(n5722), .ZN(n5742) );
  NAND2_X1 U7214 ( .A1(n5723), .A2(n5742), .ZN(n5724) );
  AND2_X1 U7215 ( .A1(n5725), .A2(n5724), .ZN(n5726) );
  AND2_X2 U7216 ( .A1(n5727), .A2(n5726), .ZN(n10261) );
  INV_X1 U7217 ( .A(n10226), .ZN(n10233) );
  NAND2_X1 U7218 ( .A1(n10261), .A2(n10233), .ZN(n8925) );
  INV_X1 U7219 ( .A(n8434), .ZN(n8244) );
  XNOR2_X1 U7220 ( .A(n5728), .B(n8244), .ZN(n5730) );
  OAI22_X1 U7221 ( .A1(n6509), .A2(n10171), .B1(n8774), .B2(n5626), .ZN(n5729)
         );
  INV_X1 U7222 ( .A(n5731), .ZN(n5732) );
  NAND2_X1 U7223 ( .A1(n5732), .A2(n8244), .ZN(n8766) );
  NAND2_X1 U7224 ( .A1(n7777), .A2(n10205), .ZN(n10234) );
  NAND3_X1 U7225 ( .A1(n8766), .A2(n5733), .A3(n10234), .ZN(n5734) );
  NAND2_X1 U7226 ( .A1(n8769), .A2(n5734), .ZN(n5746) );
  MUX2_X1 U7227 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n5746), .S(n10261), .Z(n5735) );
  INV_X1 U7228 ( .A(n5735), .ZN(n5736) );
  INV_X1 U7229 ( .A(n5737), .ZN(n5741) );
  NOR2_X1 U7230 ( .A1(n5738), .A2(n5741), .ZN(n5850) );
  NAND2_X1 U7231 ( .A1(n5850), .A2(n6726), .ZN(n5843) );
  OR3_X1 U7232 ( .A1(n5753), .A2(n5754), .A3(n5739), .ZN(n5855) );
  AND2_X1 U7233 ( .A1(n7576), .A2(n5855), .ZN(n5740) );
  OR2_X1 U7234 ( .A1(n5843), .A2(n5740), .ZN(n5745) );
  NOR2_X1 U7235 ( .A1(n5751), .A2(n5741), .ZN(n5743) );
  AND2_X1 U7236 ( .A1(n5743), .A2(n5742), .ZN(n5859) );
  NAND2_X1 U7237 ( .A1(n5859), .A2(n6726), .ZN(n5849) );
  NAND3_X1 U7238 ( .A1(n8399), .A2(n5855), .A3(n10226), .ZN(n5836) );
  AND2_X1 U7239 ( .A1(n5836), .A2(n10167), .ZN(n5851) );
  OR2_X1 U7240 ( .A1(n5849), .A2(n5851), .ZN(n5744) );
  INV_X2 U7241 ( .A(n10240), .ZN(n10238) );
  NAND2_X1 U7242 ( .A1(n10238), .A2(n10233), .ZN(n8989) );
  INV_X1 U7243 ( .A(n8765), .ZN(n5749) );
  MUX2_X1 U7244 ( .A(n5746), .B(P2_REG0_REG_27__SCAN_IN), .S(n10240), .Z(n5747) );
  INV_X1 U7245 ( .A(n5747), .ZN(n5748) );
  XNOR2_X1 U7246 ( .A(n5758), .B(n5756), .ZN(n7351) );
  NAND2_X1 U7247 ( .A1(n5834), .A2(n7309), .ZN(n5757) );
  NAND2_X1 U7248 ( .A1(n8250), .A2(n5757), .ZN(n7352) );
  NAND2_X1 U7249 ( .A1(n7351), .A2(n7352), .ZN(n5761) );
  INV_X1 U7250 ( .A(n5758), .ZN(n5759) );
  NAND2_X1 U7251 ( .A1(n5759), .A2(n5756), .ZN(n5760) );
  XNOR2_X1 U7252 ( .A(n5762), .B(n10182), .ZN(n5763) );
  XNOR2_X1 U7253 ( .A(n5763), .B(n7303), .ZN(n7358) );
  NOR2_X1 U7254 ( .A1(n5763), .A2(n8670), .ZN(n5764) );
  AOI21_X1 U7255 ( .B1(n7357), .B2(n7358), .A(n5764), .ZN(n7390) );
  INV_X1 U7256 ( .A(n8669), .ZN(n10170) );
  XNOR2_X1 U7257 ( .A(n5765), .B(n10170), .ZN(n7389) );
  NAND2_X1 U7258 ( .A1(n5765), .A2(n8669), .ZN(n5766) );
  XNOR2_X1 U7259 ( .A(n5762), .B(n10189), .ZN(n5768) );
  XNOR2_X1 U7260 ( .A(n5768), .B(n8668), .ZN(n7323) );
  INV_X1 U7261 ( .A(n5768), .ZN(n5769) );
  INV_X1 U7262 ( .A(n8668), .ZN(n7402) );
  NAND2_X1 U7263 ( .A1(n5769), .A2(n7402), .ZN(n5770) );
  NAND2_X1 U7264 ( .A1(n7320), .A2(n5770), .ZN(n7399) );
  XNOR2_X1 U7265 ( .A(n5828), .B(n10194), .ZN(n5771) );
  INV_X1 U7266 ( .A(n8667), .ZN(n7722) );
  XNOR2_X1 U7267 ( .A(n5771), .B(n7722), .ZN(n7398) );
  NAND2_X1 U7268 ( .A1(n7399), .A2(n7398), .ZN(n5774) );
  INV_X1 U7269 ( .A(n5771), .ZN(n5772) );
  NAND2_X1 U7270 ( .A1(n5772), .A2(n7722), .ZN(n5773) );
  XNOR2_X1 U7271 ( .A(n5828), .B(n10198), .ZN(n5777) );
  XNOR2_X1 U7272 ( .A(n5777), .B(n8666), .ZN(n7411) );
  XNOR2_X1 U7273 ( .A(n5828), .B(n10204), .ZN(n5776) );
  INV_X1 U7274 ( .A(n5776), .ZN(n5775) );
  INV_X1 U7275 ( .A(n8665), .ZN(n7416) );
  AND2_X1 U7276 ( .A1(n5775), .A2(n7416), .ZN(n5778) );
  XNOR2_X1 U7277 ( .A(n5776), .B(n7416), .ZN(n7506) );
  NAND2_X1 U7278 ( .A1(n5777), .A2(n8666), .ZN(n7502) );
  AND2_X1 U7279 ( .A1(n7506), .A2(n7502), .ZN(n7503) );
  OR2_X1 U7280 ( .A1(n5778), .A2(n7503), .ZN(n5779) );
  INV_X1 U7281 ( .A(n8663), .ZN(n5785) );
  XNOR2_X1 U7282 ( .A(n7782), .B(n5828), .ZN(n7767) );
  INV_X1 U7283 ( .A(n7767), .ZN(n5781) );
  XNOR2_X1 U7284 ( .A(n5828), .B(n10210), .ZN(n7764) );
  INV_X1 U7285 ( .A(n7764), .ZN(n5780) );
  INV_X1 U7286 ( .A(n8664), .ZN(n7689) );
  AOI22_X1 U7287 ( .A1(n5785), .A2(n5781), .B1(n5780), .B2(n7689), .ZN(n5787)
         );
  NAND2_X1 U7288 ( .A1(n7764), .A2(n8664), .ZN(n5784) );
  NAND2_X1 U7289 ( .A1(n5784), .A2(n5785), .ZN(n5782) );
  NAND2_X1 U7290 ( .A1(n5782), .A2(n7767), .ZN(n5783) );
  OAI21_X1 U7291 ( .B1(n5785), .B2(n5784), .A(n5783), .ZN(n5786) );
  XNOR2_X1 U7292 ( .A(n7797), .B(n5834), .ZN(n7793) );
  NAND2_X1 U7293 ( .A1(n7791), .A2(n7793), .ZN(n5788) );
  NAND2_X1 U7294 ( .A1(n4486), .A2(n8662), .ZN(n7790) );
  NAND2_X1 U7295 ( .A1(n5788), .A2(n7790), .ZN(n8615) );
  XNOR2_X1 U7296 ( .A(n8419), .B(n5828), .ZN(n8618) );
  INV_X1 U7297 ( .A(n8618), .ZN(n5789) );
  NAND2_X1 U7298 ( .A1(n5789), .A2(n8661), .ZN(n5790) );
  XNOR2_X1 U7299 ( .A(n10232), .B(n5834), .ZN(n7932) );
  XNOR2_X1 U7300 ( .A(n9840), .B(n5828), .ZN(n5791) );
  NAND2_X1 U7301 ( .A1(n5791), .A2(n7952), .ZN(n8028) );
  NAND2_X1 U7302 ( .A1(n8030), .A2(n8028), .ZN(n5793) );
  INV_X1 U7303 ( .A(n5791), .ZN(n5792) );
  NAND2_X1 U7304 ( .A1(n5792), .A2(n5372), .ZN(n8029) );
  NAND2_X1 U7305 ( .A1(n5793), .A2(n8029), .ZN(n8075) );
  XNOR2_X1 U7306 ( .A(n8114), .B(n5828), .ZN(n5794) );
  XNOR2_X1 U7307 ( .A(n5794), .B(n8123), .ZN(n8076) );
  NAND2_X1 U7308 ( .A1(n5794), .A2(n8123), .ZN(n5795) );
  XNOR2_X1 U7309 ( .A(n8941), .B(n5828), .ZN(n5798) );
  XNOR2_X1 U7310 ( .A(n5798), .B(n8200), .ZN(n8149) );
  INV_X1 U7311 ( .A(n5798), .ZN(n5799) );
  NAND2_X1 U7312 ( .A1(n5799), .A2(n8892), .ZN(n5800) );
  XNOR2_X1 U7313 ( .A(n9010), .B(n5834), .ZN(n8194) );
  OAI21_X1 U7314 ( .B1(n8196), .B2(n8194), .A(n8880), .ZN(n5802) );
  NAND2_X1 U7315 ( .A1(n8196), .A2(n8194), .ZN(n5801) );
  NAND2_X1 U7316 ( .A1(n5802), .A2(n5801), .ZN(n8225) );
  XNOR2_X1 U7317 ( .A(n9003), .B(n5834), .ZN(n8223) );
  AND2_X1 U7318 ( .A1(n8223), .A2(n8890), .ZN(n5805) );
  INV_X1 U7319 ( .A(n8223), .ZN(n5803) );
  NAND2_X1 U7320 ( .A1(n5803), .A2(n8866), .ZN(n5804) );
  XNOR2_X1 U7321 ( .A(n8930), .B(n5828), .ZN(n5807) );
  XNOR2_X1 U7322 ( .A(n5807), .B(n8879), .ZN(n8631) );
  NAND2_X1 U7323 ( .A1(n8630), .A2(n8631), .ZN(n5809) );
  NAND2_X1 U7324 ( .A1(n5807), .A2(n5806), .ZN(n5808) );
  XNOR2_X1 U7325 ( .A(n8993), .B(n5828), .ZN(n8567) );
  AND2_X1 U7326 ( .A1(n8567), .A2(n8865), .ZN(n5812) );
  INV_X1 U7327 ( .A(n8567), .ZN(n5810) );
  NAND2_X1 U7328 ( .A1(n5810), .A2(n8658), .ZN(n5811) );
  XNOR2_X1 U7329 ( .A(n8836), .B(n5828), .ZN(n5813) );
  NAND2_X1 U7330 ( .A1(n5813), .A2(n8822), .ZN(n8576) );
  INV_X1 U7331 ( .A(n5813), .ZN(n5814) );
  NAND2_X1 U7332 ( .A1(n5814), .A2(n8848), .ZN(n5815) );
  NAND2_X1 U7333 ( .A1(n8576), .A2(n5815), .ZN(n8529) );
  XNOR2_X1 U7334 ( .A(n8826), .B(n5828), .ZN(n5817) );
  XNOR2_X1 U7335 ( .A(n5817), .B(n8807), .ZN(n8577) );
  INV_X1 U7336 ( .A(n8577), .ZN(n5818) );
  NAND2_X1 U7337 ( .A1(n5817), .A2(n8835), .ZN(n5819) );
  OR2_X1 U7338 ( .A1(n5818), .A2(n8576), .ZN(n8579) );
  XNOR2_X1 U7339 ( .A(n8977), .B(n5828), .ZN(n8608) );
  INV_X1 U7340 ( .A(n8608), .ZN(n5820) );
  NAND2_X1 U7341 ( .A1(n5820), .A2(n8657), .ZN(n5821) );
  INV_X1 U7342 ( .A(n8597), .ZN(n5827) );
  XNOR2_X1 U7343 ( .A(n8966), .B(n5828), .ZN(n8599) );
  NOR2_X1 U7344 ( .A1(n8599), .A2(n8797), .ZN(n5822) );
  OAI21_X1 U7345 ( .B1(n8596), .B2(n8808), .A(n8656), .ZN(n5823) );
  AOI21_X1 U7346 ( .B1(n5827), .B2(n5826), .A(n5825), .ZN(n8587) );
  XNOR2_X1 U7347 ( .A(n8960), .B(n5828), .ZN(n5829) );
  XNOR2_X1 U7348 ( .A(n5829), .B(n8783), .ZN(n8586) );
  XNOR2_X1 U7349 ( .A(n8955), .B(n5828), .ZN(n5831) );
  XNOR2_X1 U7350 ( .A(n5832), .B(n5830), .ZN(n8639) );
  XNOR2_X1 U7351 ( .A(n8765), .B(n5828), .ZN(n5840) );
  NOR2_X1 U7352 ( .A1(n5840), .A2(n8646), .ZN(n5868) );
  AOI21_X1 U7353 ( .B1(n8646), .B2(n5840), .A(n5868), .ZN(n8554) );
  INV_X1 U7354 ( .A(n8553), .ZN(n5839) );
  XNOR2_X1 U7355 ( .A(n6509), .B(n5834), .ZN(n5835) );
  XNOR2_X1 U7356 ( .A(n8378), .B(n5835), .ZN(n5869) );
  INV_X1 U7357 ( .A(n5869), .ZN(n5842) );
  OR2_X1 U7358 ( .A1(n5843), .A2(n5836), .ZN(n5838) );
  OR2_X1 U7359 ( .A1(n5849), .A2(n5855), .ZN(n5837) );
  NAND2_X1 U7360 ( .A1(n5838), .A2(n5837), .ZN(n8616) );
  NAND3_X1 U7361 ( .A1(n5839), .A2(n5842), .A3(n8616), .ZN(n5873) );
  INV_X1 U7362 ( .A(n5840), .ZN(n5841) );
  NAND4_X1 U7363 ( .A1(n5842), .A2(n5841), .A3(n8655), .A4(n8616), .ZN(n5867)
         );
  OR2_X1 U7364 ( .A1(n5843), .A2(n10226), .ZN(n5844) );
  NAND2_X1 U7365 ( .A1(n5844), .A2(n10165), .ZN(n8648) );
  OR2_X1 U7366 ( .A1(n7576), .A2(n5845), .ZN(n5846) );
  OR2_X1 U7367 ( .A1(n5849), .A2(n5846), .ZN(n8635) );
  INV_X1 U7368 ( .A(n8234), .ZN(n8653) );
  OR2_X1 U7369 ( .A1(n5847), .A2(n7576), .ZN(n5848) );
  AOI22_X1 U7370 ( .A1(n8653), .A2(n8632), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n5864) );
  OR2_X1 U7371 ( .A1(n5851), .A2(n5850), .ZN(n5854) );
  AND3_X1 U7372 ( .A1(n5852), .A2(n6524), .A3(n6525), .ZN(n5853) );
  OAI211_X1 U7373 ( .C1(n5859), .C2(n5855), .A(n5854), .B(n5853), .ZN(n5856)
         );
  NAND2_X1 U7374 ( .A1(n5856), .A2(P2_STATE_REG_SCAN_IN), .ZN(n5861) );
  INV_X1 U7375 ( .A(n6726), .ZN(n5857) );
  NOR2_X1 U7376 ( .A1(n7576), .A2(n5857), .ZN(n8462) );
  INV_X1 U7377 ( .A(n8462), .ZN(n5858) );
  OR2_X1 U7378 ( .A1(n5859), .A2(n5858), .ZN(n5860) );
  NAND2_X1 U7379 ( .A1(n5861), .A2(n5860), .ZN(n8641) );
  NAND2_X1 U7380 ( .A1(n5862), .A2(n8641), .ZN(n5863) );
  OAI211_X1 U7381 ( .C1(n8646), .C2(n8635), .A(n5864), .B(n5863), .ZN(n5865)
         );
  AOI21_X1 U7382 ( .B1(n8378), .B2(n8648), .A(n5865), .ZN(n5866) );
  INV_X1 U7383 ( .A(n5868), .ZN(n5870) );
  NAND4_X1 U7384 ( .A1(n8553), .A2(n5870), .A3(n8616), .A4(n5869), .ZN(n5871)
         );
  NAND3_X1 U7385 ( .A1(n5873), .A2(n5872), .A3(n5871), .ZN(P2_U3160) );
  NOR2_X1 U7386 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5875) );
  NAND4_X1 U7387 ( .A1(n5875), .A2(n5874), .A3(n9886), .A4(n6887), .ZN(n6044)
         );
  INV_X1 U7388 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6165) );
  NAND4_X1 U7389 ( .A1(n6165), .A2(n6879), .A3(n6121), .A4(n6983), .ZN(n6767)
         );
  INV_X1 U7390 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n6123) );
  INV_X1 U7391 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5876) );
  INV_X1 U7392 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n6120) );
  NAND3_X1 U7393 ( .A1(n6123), .A2(n5876), .A3(n6120), .ZN(n5877) );
  AND2_X2 U7394 ( .A1(n5895), .A2(n6866), .ZN(n5900) );
  INV_X1 U7395 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5889) );
  INV_X1 U7396 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5880) );
  XNOR2_X2 U7397 ( .A(n5879), .B(n5891), .ZN(n6284) );
  INV_X1 U7398 ( .A(n6221), .ZN(n5881) );
  NAND2_X1 U7399 ( .A1(n5881), .A2(n5009), .ZN(n5883) );
  NAND2_X1 U7400 ( .A1(n5883), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5882) );
  XNOR2_X1 U7401 ( .A(n5882), .B(n6785), .ZN(n9321) );
  INV_X1 U7402 ( .A(n7477), .ZN(n5884) );
  INV_X1 U7403 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5892) );
  NAND2_X1 U7404 ( .A1(n5885), .A2(n5892), .ZN(n5886) );
  XNOR2_X1 U7405 ( .A(n6463), .B(P1_IR_REG_22__SCAN_IN), .ZN(n6467) );
  NAND2_X1 U7406 ( .A1(n5887), .A2(n7112), .ZN(n5905) );
  NOR2_X1 U7407 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5890) );
  NAND4_X1 U7408 ( .A1(n5890), .A2(n5889), .A3(n5888), .A4(n6937), .ZN(n5894)
         );
  NAND2_X1 U7409 ( .A1(n5907), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5897) );
  INV_X1 U7410 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5909) );
  NAND2_X1 U7411 ( .A1(n5897), .A2(n5909), .ZN(n5899) );
  NAND2_X1 U7412 ( .A1(n5899), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5896) );
  INV_X1 U7413 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5908) );
  XNOR2_X1 U7414 ( .A(n5896), .B(n5908), .ZN(n8100) );
  OR2_X1 U7415 ( .A1(n5897), .A2(n5909), .ZN(n5898) );
  NAND2_X1 U7416 ( .A1(n5899), .A2(n5898), .ZN(n8061) );
  NAND2_X1 U7417 ( .A1(n5900), .A2(n5901), .ZN(n5902) );
  NAND2_X1 U7418 ( .A1(n5902), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5904) );
  XNOR2_X1 U7419 ( .A(n5904), .B(n5903), .ZN(n8027) );
  NAND2_X2 U7420 ( .A1(n5905), .A2(n6705), .ZN(n6393) );
  NAND2_X4 U7421 ( .A1(n5906), .A2(n7112), .ZN(n6439) );
  NAND2_X1 U7422 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n5910) );
  XNOR2_X2 U7423 ( .A(n5918), .B(P1_IR_REG_28__SCAN_IN), .ZN(n6487) );
  NAND2_X2 U7424 ( .A1(n6487), .A2(n7028), .ZN(n5960) );
  NAND2_X1 U7425 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5912) );
  INV_X1 U7426 ( .A(n9884), .ZN(n7036) );
  INV_X1 U7427 ( .A(n5913), .ZN(n6722) );
  NAND2_X1 U7428 ( .A1(n5959), .A2(n9982), .ZN(n5935) );
  INV_X1 U7429 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5919) );
  INV_X1 U7430 ( .A(n5922), .ZN(n9830) );
  OR2_X2 U7431 ( .A1(n5922), .A2(n5921), .ZN(n5924) );
  XNOR2_X2 U7432 ( .A(n5924), .B(n5923), .ZN(n8468) );
  NAND2_X2 U7433 ( .A1(n5929), .A2(n5925), .ZN(n6006) );
  INV_X1 U7434 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n5927) );
  NAND2_X2 U7435 ( .A1(n5930), .A2(n5925), .ZN(n6009) );
  INV_X1 U7436 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5926) );
  OAI22_X1 U7437 ( .A1(n6006), .A2(n5927), .B1(n6009), .B2(n5926), .ZN(n5928)
         );
  INV_X1 U7438 ( .A(n5928), .ZN(n5933) );
  INV_X1 U7439 ( .A(n5987), .ZN(n6008) );
  INV_X1 U7440 ( .A(n6705), .ZN(n6750) );
  NOR2_X1 U7441 ( .A1(n6750), .A2(n7477), .ZN(n5937) );
  NAND2_X1 U7442 ( .A1(n7440), .A2(n5937), .ZN(n5934) );
  NAND2_X1 U7443 ( .A1(n5935), .A2(n5934), .ZN(n5936) );
  XNOR2_X2 U7444 ( .A(n5936), .B(n6418), .ZN(n5955) );
  NAND2_X1 U7445 ( .A1(n7440), .A2(n6441), .ZN(n5939) );
  OR2_X1 U7446 ( .A1(n7439), .A2(n6093), .ZN(n5938) );
  NAND2_X1 U7447 ( .A1(n5939), .A2(n5938), .ZN(n5956) );
  XNOR2_X1 U7448 ( .A(n5955), .B(n5956), .ZN(n7123) );
  INV_X1 U7449 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7554) );
  INV_X1 U7450 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5940) );
  OAI22_X1 U7451 ( .A1(n6006), .A2(n7554), .B1(n6009), .B2(n5940), .ZN(n5943)
         );
  INV_X1 U7452 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5941) );
  INV_X1 U7453 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5953) );
  NAND2_X1 U7454 ( .A1(n7114), .A2(n4424), .ZN(n5950) );
  INV_X1 U7455 ( .A(SI_0_), .ZN(n5945) );
  INV_X1 U7456 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5944) );
  OAI21_X1 U7457 ( .B1(n8392), .B2(n5945), .A(n5944), .ZN(n5947) );
  AND2_X1 U7458 ( .A1(n5947), .A2(n5946), .ZN(n9836) );
  MUX2_X1 U7459 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9836), .S(n5960), .Z(n7550) );
  INV_X2 U7460 ( .A(n6093), .ZN(n6056) );
  NOR2_X1 U7461 ( .A1(n6705), .A2(n9886), .ZN(n5948) );
  AOI21_X1 U7462 ( .B1(n7550), .B2(n6056), .A(n5948), .ZN(n5949) );
  NAND2_X1 U7463 ( .A1(n5950), .A2(n5949), .ZN(n7062) );
  NAND2_X1 U7464 ( .A1(n5959), .A2(n7550), .ZN(n5952) );
  NAND2_X1 U7465 ( .A1(n7114), .A2(n6056), .ZN(n5951) );
  OAI211_X1 U7466 ( .C1(n6705), .C2(n5953), .A(n5952), .B(n5951), .ZN(n7063)
         );
  NAND2_X1 U7467 ( .A1(n7062), .A2(n7063), .ZN(n7061) );
  OR2_X1 U7468 ( .A1(n6439), .A2(n7550), .ZN(n5954) );
  AND2_X1 U7469 ( .A1(n7061), .A2(n5954), .ZN(n7122) );
  NAND2_X1 U7470 ( .A1(n7123), .A2(n7122), .ZN(n7121) );
  INV_X1 U7471 ( .A(n5956), .ZN(n5957) );
  NAND2_X1 U7472 ( .A1(n5955), .A2(n5957), .ZN(n5958) );
  NAND2_X1 U7473 ( .A1(n7121), .A2(n5958), .ZN(n7141) );
  XNOR2_X1 U7474 ( .A(n6001), .B(P1_IR_REG_2__SCAN_IN), .ZN(n7035) );
  OR2_X1 U7475 ( .A1(n6003), .A2(n6711), .ZN(n5962) );
  OR2_X1 U7476 ( .A1(n5979), .A2(n6710), .ZN(n5961) );
  NAND2_X1 U7477 ( .A1(n5959), .A2(n7442), .ZN(n5972) );
  INV_X1 U7478 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n5964) );
  INV_X1 U7479 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5963) );
  OAI22_X1 U7480 ( .A1(n6006), .A2(n5964), .B1(n6009), .B2(n5963), .ZN(n5965)
         );
  INV_X1 U7481 ( .A(n5965), .ZN(n5970) );
  INV_X1 U7482 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n5967) );
  INV_X1 U7483 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5966) );
  OAI22_X1 U7484 ( .A1(n5986), .A2(n5967), .B1(n5987), .B2(n5966), .ZN(n5968)
         );
  INV_X1 U7485 ( .A(n5968), .ZN(n5969) );
  NAND2_X1 U7486 ( .A1(n5970), .A2(n5969), .ZN(n7444) );
  NAND2_X1 U7487 ( .A1(n7444), .A2(n6056), .ZN(n5971) );
  NAND2_X1 U7488 ( .A1(n5972), .A2(n5971), .ZN(n5973) );
  XNOR2_X1 U7489 ( .A(n5973), .B(n6439), .ZN(n5974) );
  AOI22_X1 U7490 ( .A1(n7444), .A2(n4424), .B1(n6056), .B2(n7442), .ZN(n5975)
         );
  XNOR2_X1 U7491 ( .A(n5974), .B(n5975), .ZN(n7140) );
  NAND2_X1 U7492 ( .A1(n7141), .A2(n7140), .ZN(n5978) );
  INV_X1 U7493 ( .A(n5974), .ZN(n5976) );
  NAND2_X1 U7494 ( .A1(n5976), .A2(n5975), .ZN(n5977) );
  NAND2_X1 U7495 ( .A1(n5978), .A2(n5977), .ZN(n7230) );
  OR2_X1 U7496 ( .A1(n5979), .A2(n6712), .ZN(n5984) );
  OR2_X1 U7497 ( .A1(n6003), .A2(n6713), .ZN(n5983) );
  NAND2_X1 U7498 ( .A1(n6001), .A2(n6887), .ZN(n5980) );
  NAND2_X1 U7499 ( .A1(n5980), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5981) );
  XNOR2_X1 U7500 ( .A(n5981), .B(P1_IR_REG_3__SCAN_IN), .ZN(n7033) );
  INV_X1 U7501 ( .A(n7033), .ZN(n9453) );
  OR2_X1 U7502 ( .A1(n6753), .A2(n9453), .ZN(n5982) );
  INV_X1 U7503 ( .A(n10015), .ZN(n9960) );
  NAND2_X1 U7504 ( .A1(n6430), .A2(n9960), .ZN(n5992) );
  INV_X1 U7505 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n5985) );
  OAI22_X1 U7506 ( .A1(n6006), .A2(P1_REG3_REG_3__SCAN_IN), .B1(n6009), .B2(
        n5985), .ZN(n5990) );
  INV_X1 U7507 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7034) );
  INV_X1 U7508 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5988) );
  OAI22_X1 U7509 ( .A1(n9284), .A2(n7034), .B1(n5987), .B2(n5988), .ZN(n5989)
         );
  NAND2_X1 U7510 ( .A1(n7463), .A2(n6056), .ZN(n5991) );
  NAND2_X1 U7511 ( .A1(n5992), .A2(n5991), .ZN(n5993) );
  XNOR2_X1 U7512 ( .A(n5993), .B(n6418), .ZN(n5998) );
  NAND2_X1 U7513 ( .A1(n7463), .A2(n4424), .ZN(n5995) );
  OR2_X1 U7514 ( .A1(n10015), .A2(n6093), .ZN(n5994) );
  NAND2_X1 U7515 ( .A1(n5995), .A2(n5994), .ZN(n5996) );
  XNOR2_X1 U7516 ( .A(n5998), .B(n5996), .ZN(n7231) );
  INV_X1 U7517 ( .A(n5996), .ZN(n5997) );
  NAND2_X1 U7518 ( .A1(n5998), .A2(n5997), .ZN(n5999) );
  OAI21_X1 U7519 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(P1_IR_REG_3__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6000) );
  NAND2_X1 U7520 ( .A1(n6001), .A2(n6000), .ZN(n6024) );
  INV_X1 U7521 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6002) );
  XNOR2_X1 U7522 ( .A(n6024), .B(n6002), .ZN(n9473) );
  INV_X1 U7523 ( .A(n9473), .ZN(n8491) );
  OR2_X1 U7524 ( .A1(n6003), .A2(n8492), .ZN(n6004) );
  NAND2_X1 U7525 ( .A1(n6430), .A2(n7617), .ZN(n6013) );
  NOR2_X1 U7526 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6007) );
  NOR2_X1 U7527 ( .A1(n6028), .A2(n6007), .ZN(n7618) );
  NAND2_X1 U7528 ( .A1(n6482), .A2(n7618), .ZN(n6011) );
  NAND2_X1 U7529 ( .A1(n6008), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6010) );
  NAND2_X1 U7530 ( .A1(n9451), .A2(n6056), .ZN(n6012) );
  NAND2_X1 U7531 ( .A1(n6013), .A2(n6012), .ZN(n6014) );
  XNOR2_X1 U7532 ( .A(n6014), .B(n6439), .ZN(n6017) );
  NAND2_X1 U7533 ( .A1(n9451), .A2(n4424), .ZN(n6016) );
  NAND2_X1 U7534 ( .A1(n7617), .A2(n6056), .ZN(n6015) );
  NAND2_X1 U7535 ( .A1(n6016), .A2(n6015), .ZN(n6018) );
  NAND2_X1 U7536 ( .A1(n6017), .A2(n6018), .ZN(n6023) );
  INV_X1 U7537 ( .A(n6017), .ZN(n6020) );
  INV_X1 U7538 ( .A(n6018), .ZN(n6019) );
  NAND2_X1 U7539 ( .A1(n6020), .A2(n6019), .ZN(n6021) );
  NAND2_X1 U7540 ( .A1(n6023), .A2(n6021), .ZN(n7284) );
  NAND2_X1 U7541 ( .A1(n7286), .A2(n6023), .ZN(n6039) );
  OAI21_X1 U7542 ( .B1(n6024), .B2(P1_IR_REG_4__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6025) );
  XNOR2_X1 U7543 ( .A(n6025), .B(P1_IR_REG_5__SCAN_IN), .ZN(n7031) );
  INV_X1 U7544 ( .A(n7031), .ZN(n7085) );
  OR2_X1 U7545 ( .A1(n6716), .A2(n5979), .ZN(n6027) );
  OR2_X1 U7546 ( .A1(n6003), .A2(n6717), .ZN(n6026) );
  NAND2_X1 U7547 ( .A1(n6430), .A2(n9948), .ZN(n6035) );
  NOR2_X1 U7548 ( .A1(n6028), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6029) );
  NOR2_X1 U7549 ( .A1(n6051), .A2(n6029), .ZN(n9946) );
  NAND2_X1 U7550 ( .A1(n6482), .A2(n9946), .ZN(n6033) );
  NAND2_X1 U7551 ( .A1(n5931), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6032) );
  NAND2_X1 U7552 ( .A1(n9280), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U7553 ( .A1(n9279), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6030) );
  NAND4_X1 U7554 ( .A1(n6033), .A2(n6032), .A3(n6031), .A4(n6030), .ZN(n9450)
         );
  NAND2_X1 U7555 ( .A1(n9450), .A2(n6056), .ZN(n6034) );
  NAND2_X1 U7556 ( .A1(n6035), .A2(n6034), .ZN(n6036) );
  XNOR2_X1 U7557 ( .A(n6036), .B(n6439), .ZN(n6040) );
  NAND2_X1 U7558 ( .A1(n6039), .A2(n6040), .ZN(n7368) );
  NAND2_X1 U7559 ( .A1(n9450), .A2(n4424), .ZN(n6038) );
  NAND2_X1 U7560 ( .A1(n9948), .A2(n6056), .ZN(n6037) );
  AND2_X1 U7561 ( .A1(n6038), .A2(n6037), .ZN(n7370) );
  NAND2_X1 U7562 ( .A1(n7368), .A2(n7370), .ZN(n6043) );
  INV_X1 U7563 ( .A(n6039), .ZN(n6042) );
  INV_X1 U7564 ( .A(n6040), .ZN(n6041) );
  NAND2_X1 U7565 ( .A1(n6042), .A2(n6041), .ZN(n7369) );
  OR2_X1 U7566 ( .A1(n6720), .A2(n5979), .ZN(n6050) );
  NAND2_X1 U7567 ( .A1(n6044), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6045) );
  MUX2_X1 U7568 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6045), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n6048) );
  INV_X1 U7569 ( .A(n6046), .ZN(n6047) );
  AND2_X1 U7570 ( .A1(n6048), .A2(n6047), .ZN(n7093) );
  AOI22_X1 U7571 ( .A1(n6286), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6285), .B2(
        n7093), .ZN(n6049) );
  OAI21_X1 U7572 ( .B1(n6051), .B2(P1_REG3_REG_6__SCAN_IN), .A(n6068), .ZN(
        n7428) );
  INV_X1 U7573 ( .A(n7428), .ZN(n7604) );
  NAND2_X1 U7574 ( .A1(n6482), .A2(n7604), .ZN(n6055) );
  NAND2_X1 U7575 ( .A1(n5931), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6054) );
  NAND2_X1 U7576 ( .A1(n9280), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U7577 ( .A1(n9279), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6052) );
  NAND4_X1 U7578 ( .A1(n6055), .A2(n6054), .A3(n6053), .A4(n6052), .ZN(n9449)
         );
  NAND2_X1 U7579 ( .A1(n9449), .A2(n6056), .ZN(n6057) );
  OAI21_X1 U7580 ( .B1(n10035), .B2(n6391), .A(n6057), .ZN(n6058) );
  XNOR2_X1 U7581 ( .A(n6058), .B(n6418), .ZN(n7422) );
  OR2_X1 U7582 ( .A1(n10035), .A2(n6093), .ZN(n6060) );
  NAND2_X1 U7583 ( .A1(n9449), .A2(n4424), .ZN(n6059) );
  AND2_X1 U7584 ( .A1(n6060), .A2(n6059), .ZN(n7421) );
  AND2_X1 U7585 ( .A1(n7422), .A2(n7421), .ZN(n6064) );
  INV_X1 U7586 ( .A(n7422), .ZN(n6062) );
  INV_X1 U7587 ( .A(n7421), .ZN(n6061) );
  NAND2_X1 U7588 ( .A1(n6062), .A2(n6061), .ZN(n6063) );
  OR2_X1 U7589 ( .A1(n6046), .A2(n5921), .ZN(n6065) );
  XNOR2_X1 U7590 ( .A(n6065), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7205) );
  AOI22_X1 U7591 ( .A1(n6286), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6285), .B2(
        n7205), .ZN(n6066) );
  AND2_X1 U7592 ( .A1(n6068), .A2(n7545), .ZN(n6069) );
  NOR2_X1 U7593 ( .A1(n6101), .A2(n6069), .ZN(n9933) );
  NAND2_X1 U7594 ( .A1(n6482), .A2(n9933), .ZN(n6073) );
  NAND2_X1 U7595 ( .A1(n5931), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6072) );
  NAND2_X1 U7596 ( .A1(n9280), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6071) );
  NAND2_X1 U7597 ( .A1(n9279), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6070) );
  NAND4_X1 U7598 ( .A1(n6073), .A2(n6072), .A3(n6071), .A4(n6070), .ZN(n9448)
         );
  INV_X1 U7599 ( .A(n9448), .ZN(n7447) );
  OAI22_X1 U7600 ( .A1(n10042), .A2(n6391), .B1(n7447), .B2(n6093), .ZN(n6074)
         );
  XNOR2_X1 U7601 ( .A(n6074), .B(n6439), .ZN(n6080) );
  INV_X1 U7602 ( .A(n6080), .ZN(n6078) );
  OR2_X1 U7603 ( .A1(n10042), .A2(n6093), .ZN(n6076) );
  NAND2_X1 U7604 ( .A1(n9448), .A2(n4424), .ZN(n6075) );
  NAND2_X1 U7605 ( .A1(n6076), .A2(n6075), .ZN(n6079) );
  INV_X1 U7606 ( .A(n6079), .ZN(n6077) );
  AND2_X1 U7607 ( .A1(n6080), .A2(n6079), .ZN(n7540) );
  NAND2_X1 U7608 ( .A1(n7014), .A2(n9176), .ZN(n6084) );
  NAND2_X1 U7609 ( .A1(n6046), .A2(n6121), .ZN(n6081) );
  NAND2_X1 U7610 ( .A1(n6081), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6096) );
  NAND2_X1 U7611 ( .A1(n6096), .A2(n6879), .ZN(n6098) );
  NAND2_X1 U7612 ( .A1(n6098), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6082) );
  XNOR2_X1 U7613 ( .A(n6082), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7337) );
  AOI22_X1 U7614 ( .A1(n6286), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6285), .B2(
        n7337), .ZN(n6083) );
  NAND2_X1 U7615 ( .A1(n10058), .A2(n6430), .ZN(n6091) );
  NAND2_X1 U7616 ( .A1(n6101), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6103) );
  INV_X1 U7617 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7278) );
  NAND2_X1 U7618 ( .A1(n6103), .A2(n7278), .ZN(n6085) );
  AND2_X1 U7619 ( .A1(n6144), .A2(n6085), .ZN(n8014) );
  NAND2_X1 U7620 ( .A1(n6482), .A2(n8014), .ZN(n6089) );
  NAND2_X1 U7621 ( .A1(n6480), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6088) );
  NAND2_X1 U7622 ( .A1(n9279), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6087) );
  NAND2_X1 U7623 ( .A1(n9280), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6086) );
  NAND4_X1 U7624 ( .A1(n6089), .A2(n6088), .A3(n6087), .A4(n6086), .ZN(n9446)
         );
  NAND2_X1 U7625 ( .A1(n9446), .A2(n6436), .ZN(n6090) );
  NAND2_X1 U7626 ( .A1(n6091), .A2(n6090), .ZN(n6092) );
  XNOR2_X1 U7627 ( .A(n6092), .B(n6439), .ZN(n6114) );
  NAND2_X1 U7628 ( .A1(n10058), .A2(n6436), .ZN(n6095) );
  NAND2_X1 U7629 ( .A1(n9446), .A2(n4424), .ZN(n6094) );
  NAND2_X1 U7630 ( .A1(n6095), .A2(n6094), .ZN(n8006) );
  OR2_X1 U7631 ( .A1(n6739), .A2(n5979), .ZN(n6100) );
  OR2_X1 U7632 ( .A1(n6096), .A2(n6879), .ZN(n6097) );
  AND2_X1 U7633 ( .A1(n6098), .A2(n6097), .ZN(n7274) );
  AOI22_X1 U7634 ( .A1(n6286), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6285), .B2(
        n7274), .ZN(n6099) );
  NAND2_X1 U7635 ( .A1(n7866), .A2(n6430), .ZN(n6109) );
  OR2_X1 U7636 ( .A1(n6101), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6102) );
  AND2_X1 U7637 ( .A1(n6103), .A2(n6102), .ZN(n7861) );
  NAND2_X1 U7638 ( .A1(n6482), .A2(n7861), .ZN(n6107) );
  NAND2_X1 U7639 ( .A1(n6480), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6106) );
  NAND2_X1 U7640 ( .A1(n9280), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6105) );
  NAND2_X1 U7641 ( .A1(n9279), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6104) );
  NAND4_X1 U7642 ( .A1(n6107), .A2(n6106), .A3(n6105), .A4(n6104), .ZN(n9447)
         );
  NAND2_X1 U7643 ( .A1(n9447), .A2(n6436), .ZN(n6108) );
  NAND2_X1 U7644 ( .A1(n6109), .A2(n6108), .ZN(n6110) );
  XNOR2_X1 U7645 ( .A(n6110), .B(n6439), .ZN(n6115) );
  NAND2_X1 U7646 ( .A1(n7866), .A2(n6436), .ZN(n6112) );
  NAND2_X1 U7647 ( .A1(n9447), .A2(n4424), .ZN(n6111) );
  NAND2_X1 U7648 ( .A1(n6112), .A2(n6111), .ZN(n7860) );
  AOI22_X1 U7649 ( .A1(n6114), .A2(n8006), .B1(n6115), .B2(n7860), .ZN(n6113)
         );
  INV_X1 U7650 ( .A(n6114), .ZN(n8007) );
  OAI21_X1 U7651 ( .B1(n6115), .B2(n7860), .A(n8006), .ZN(n6117) );
  NOR2_X1 U7652 ( .A1(n8006), .A2(n7860), .ZN(n6116) );
  INV_X1 U7653 ( .A(n6115), .ZN(n8005) );
  AOI22_X1 U7654 ( .A1(n8007), .A2(n6117), .B1(n6116), .B2(n8005), .ZN(n6118)
         );
  NAND2_X1 U7655 ( .A1(n6119), .A2(n6118), .ZN(n7963) );
  NAND2_X1 U7656 ( .A1(n7071), .A2(n9176), .ZN(n6127) );
  AND3_X1 U7657 ( .A1(n6879), .A2(n6121), .A3(n6120), .ZN(n6122) );
  NAND2_X1 U7658 ( .A1(n6046), .A2(n6122), .ZN(n6138) );
  OR2_X1 U7659 ( .A1(n6138), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6140) );
  NAND2_X1 U7660 ( .A1(n6140), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6124) );
  MUX2_X1 U7661 ( .A(n6124), .B(P1_IR_REG_31__SCAN_IN), .S(n6123), .Z(n6125)
         );
  OR2_X1 U7662 ( .A1(n6140), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n6163) );
  AND2_X1 U7663 ( .A1(n6125), .A2(n6163), .ZN(n7666) );
  AOI22_X1 U7664 ( .A1(n6286), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6285), .B2(
        n7666), .ZN(n6126) );
  NAND2_X1 U7665 ( .A1(n9920), .A2(n6430), .ZN(n6134) );
  INV_X1 U7666 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7966) );
  NOR2_X1 U7667 ( .A1(n6146), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6128) );
  OR2_X1 U7668 ( .A1(n6171), .A2(n6128), .ZN(n8071) );
  INV_X1 U7669 ( .A(n8071), .ZN(n9919) );
  NAND2_X1 U7670 ( .A1(n6482), .A2(n9919), .ZN(n6132) );
  NAND2_X1 U7671 ( .A1(n6480), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6131) );
  NAND2_X1 U7672 ( .A1(n9280), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6130) );
  NAND2_X1 U7673 ( .A1(n9279), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6129) );
  NAND4_X1 U7674 ( .A1(n6132), .A2(n6131), .A3(n6130), .A4(n6129), .ZN(n9444)
         );
  NAND2_X1 U7675 ( .A1(n9444), .A2(n6436), .ZN(n6133) );
  NAND2_X1 U7676 ( .A1(n6134), .A2(n6133), .ZN(n6135) );
  XNOR2_X1 U7677 ( .A(n6135), .B(n6439), .ZN(n6157) );
  NAND2_X1 U7678 ( .A1(n9920), .A2(n6436), .ZN(n6137) );
  NAND2_X1 U7679 ( .A1(n9444), .A2(n4424), .ZN(n6136) );
  NAND2_X1 U7680 ( .A1(n6137), .A2(n6136), .ZN(n8064) );
  NAND2_X1 U7681 ( .A1(n7018), .A2(n9176), .ZN(n6143) );
  NAND2_X1 U7682 ( .A1(n6138), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6139) );
  MUX2_X1 U7683 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6139), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n6141) );
  AND2_X1 U7684 ( .A1(n6141), .A2(n6140), .ZN(n7565) );
  AOI22_X1 U7685 ( .A1(n6286), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6285), .B2(
        n7565), .ZN(n6142) );
  NAND2_X1 U7686 ( .A1(n6143), .A2(n6142), .ZN(n7480) );
  NAND2_X1 U7687 ( .A1(n7480), .A2(n6430), .ZN(n6152) );
  AND2_X1 U7688 ( .A1(n6144), .A2(n7966), .ZN(n6145) );
  NOR2_X1 U7689 ( .A1(n6146), .A2(n6145), .ZN(n7970) );
  NAND2_X1 U7690 ( .A1(n6482), .A2(n7970), .ZN(n6150) );
  NAND2_X1 U7691 ( .A1(n6480), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6149) );
  NAND2_X1 U7692 ( .A1(n9279), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U7693 ( .A1(n9280), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6147) );
  NAND4_X1 U7694 ( .A1(n6150), .A2(n6149), .A3(n6148), .A4(n6147), .ZN(n9445)
         );
  NAND2_X1 U7695 ( .A1(n9445), .A2(n6436), .ZN(n6151) );
  NAND2_X1 U7696 ( .A1(n6152), .A2(n6151), .ZN(n6153) );
  XNOR2_X1 U7697 ( .A(n6153), .B(n6439), .ZN(n6158) );
  NAND2_X1 U7698 ( .A1(n7480), .A2(n6436), .ZN(n6155) );
  NAND2_X1 U7699 ( .A1(n9445), .A2(n4424), .ZN(n6154) );
  NAND2_X1 U7700 ( .A1(n6155), .A2(n6154), .ZN(n7964) );
  AOI22_X1 U7701 ( .A1(n6157), .A2(n8064), .B1(n6158), .B2(n7964), .ZN(n6156)
         );
  NAND2_X1 U7702 ( .A1(n7963), .A2(n6156), .ZN(n6162) );
  INV_X1 U7703 ( .A(n6157), .ZN(n8065) );
  OAI21_X1 U7704 ( .B1(n6158), .B2(n7964), .A(n8064), .ZN(n6160) );
  NOR2_X1 U7705 ( .A1(n8064), .A2(n7964), .ZN(n6159) );
  INV_X1 U7706 ( .A(n6158), .ZN(n8063) );
  AOI22_X1 U7707 ( .A1(n8065), .A2(n6160), .B1(n6159), .B2(n8063), .ZN(n6161)
         );
  NAND2_X1 U7708 ( .A1(n6162), .A2(n6161), .ZN(n7940) );
  NAND2_X1 U7709 ( .A1(n7130), .A2(n9176), .ZN(n6169) );
  NAND2_X1 U7710 ( .A1(n6163), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6166) );
  INV_X1 U7711 ( .A(n6166), .ZN(n6164) );
  NAND2_X1 U7712 ( .A1(n6164), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n6167) );
  NAND2_X1 U7713 ( .A1(n6166), .A2(n6165), .ZN(n6184) );
  AND2_X1 U7714 ( .A1(n6167), .A2(n6184), .ZN(n7921) );
  AOI22_X1 U7715 ( .A1(n6286), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6285), .B2(
        n7921), .ZN(n6168) );
  NAND2_X1 U7716 ( .A1(n7947), .A2(n6430), .ZN(n6177) );
  INV_X1 U7717 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6170) );
  INV_X1 U7718 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7653) );
  OAI22_X1 U7719 ( .A1(n9284), .A2(n6170), .B1(n6009), .B2(n7653), .ZN(n6175)
         );
  OR2_X1 U7720 ( .A1(n6171), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6172) );
  NAND2_X1 U7721 ( .A1(n6188), .A2(n6172), .ZN(n7945) );
  INV_X1 U7722 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n6173) );
  OAI22_X1 U7723 ( .A1(n6006), .A2(n7945), .B1(n6742), .B2(n6173), .ZN(n6174)
         );
  OR2_X1 U7724 ( .A1(n6175), .A2(n6174), .ZN(n9443) );
  NAND2_X1 U7725 ( .A1(n9443), .A2(n6436), .ZN(n6176) );
  NAND2_X1 U7726 ( .A1(n6177), .A2(n6176), .ZN(n6178) );
  XNOR2_X1 U7727 ( .A(n6178), .B(n6439), .ZN(n6180) );
  AND2_X1 U7728 ( .A1(n9443), .A2(n4424), .ZN(n6179) );
  AOI21_X1 U7729 ( .B1(n7947), .B2(n6436), .A(n6179), .ZN(n6181) );
  XNOR2_X1 U7730 ( .A(n6180), .B(n6181), .ZN(n7941) );
  INV_X1 U7731 ( .A(n6180), .ZN(n6182) );
  NAND2_X1 U7732 ( .A1(n6182), .A2(n6181), .ZN(n6183) );
  NAND2_X1 U7733 ( .A1(n6184), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6185) );
  XNOR2_X1 U7734 ( .A(n6185), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9484) );
  AOI22_X1 U7735 ( .A1(n6286), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6285), .B2(
        n9484), .ZN(n6186) );
  NAND2_X1 U7736 ( .A1(n9905), .A2(n6430), .ZN(n6195) );
  INV_X1 U7737 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8020) );
  NAND2_X1 U7738 ( .A1(n6188), .A2(n8020), .ZN(n6189) );
  AND2_X1 U7739 ( .A1(n6205), .A2(n6189), .ZN(n9901) );
  NAND2_X1 U7740 ( .A1(n6482), .A2(n9901), .ZN(n6193) );
  NAND2_X1 U7741 ( .A1(n6480), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6192) );
  NAND2_X1 U7742 ( .A1(n9280), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6191) );
  NAND2_X1 U7743 ( .A1(n9279), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6190) );
  NAND4_X1 U7744 ( .A1(n6193), .A2(n6192), .A3(n6191), .A4(n6190), .ZN(n9442)
         );
  INV_X2 U7745 ( .A(n6093), .ZN(n6436) );
  NAND2_X1 U7746 ( .A1(n9442), .A2(n6436), .ZN(n6194) );
  NAND2_X1 U7747 ( .A1(n6195), .A2(n6194), .ZN(n6196) );
  XNOR2_X1 U7748 ( .A(n6196), .B(n6439), .ZN(n6198) );
  AND2_X1 U7749 ( .A1(n9442), .A2(n4424), .ZN(n6197) );
  AOI21_X1 U7750 ( .B1(n9905), .B2(n6436), .A(n6197), .ZN(n6199) );
  XNOR2_X1 U7751 ( .A(n6198), .B(n6199), .ZN(n8019) );
  INV_X1 U7752 ( .A(n6198), .ZN(n6200) );
  NAND2_X1 U7753 ( .A1(n7262), .A2(n9176), .ZN(n6204) );
  NOR2_X1 U7754 ( .A1(n5895), .A2(n5921), .ZN(n6201) );
  MUX2_X1 U7755 ( .A(n5921), .B(n6201), .S(P1_IR_REG_14__SCAN_IN), .Z(n6202)
         );
  OR2_X1 U7756 ( .A1(n6202), .A2(n5900), .ZN(n9505) );
  INV_X1 U7757 ( .A(n9505), .ZN(n9499) );
  AOI22_X1 U7758 ( .A1(n6286), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6285), .B2(
        n9499), .ZN(n6203) );
  INV_X1 U7759 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9489) );
  INV_X1 U7760 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7886) );
  OAI22_X1 U7761 ( .A1(n9284), .A2(n9489), .B1(n6009), .B2(n7886), .ZN(n6209)
         );
  INV_X1 U7762 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9032) );
  NAND2_X1 U7763 ( .A1(n6205), .A2(n9032), .ZN(n6206) );
  NAND2_X1 U7764 ( .A1(n6239), .A2(n6206), .ZN(n9031) );
  INV_X1 U7765 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n6207) );
  OAI22_X1 U7766 ( .A1(n6006), .A2(n9031), .B1(n6742), .B2(n6207), .ZN(n6208)
         );
  OR2_X1 U7767 ( .A1(n6209), .A2(n6208), .ZN(n9441) );
  INV_X1 U7768 ( .A(n9441), .ZN(n8044) );
  OAI22_X1 U7769 ( .A1(n10092), .A2(n6391), .B1(n8044), .B2(n6093), .ZN(n6210)
         );
  XNOR2_X1 U7770 ( .A(n6210), .B(n6439), .ZN(n6213) );
  OR2_X1 U7771 ( .A1(n10092), .A2(n6093), .ZN(n6212) );
  NAND2_X1 U7772 ( .A1(n9441), .A2(n4424), .ZN(n6211) );
  AND2_X1 U7773 ( .A1(n6212), .A2(n6211), .ZN(n9029) );
  INV_X1 U7774 ( .A(n6213), .ZN(n6214) );
  NAND2_X1 U7775 ( .A1(n6215), .A2(n6214), .ZN(n6216) );
  NAND2_X1 U7776 ( .A1(n7305), .A2(n9176), .ZN(n6224) );
  INV_X1 U7777 ( .A(n6217), .ZN(n6218) );
  NAND2_X1 U7778 ( .A1(n6218), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6220) );
  MUX2_X1 U7779 ( .A(n6220), .B(P1_IR_REG_31__SCAN_IN), .S(n6219), .Z(n6222)
         );
  NAND2_X1 U7780 ( .A1(n6222), .A2(n6221), .ZN(n9537) );
  INV_X1 U7781 ( .A(n9537), .ZN(n9532) );
  AOI22_X1 U7782 ( .A1(n6286), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6285), .B2(
        n9532), .ZN(n6223) );
  NAND2_X1 U7783 ( .A1(n9083), .A2(n6430), .ZN(n6231) );
  INV_X1 U7784 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9502) );
  NOR2_X1 U7785 ( .A1(n6241), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6225) );
  OR2_X1 U7786 ( .A1(n9091), .A2(n6225), .ZN(n9078) );
  INV_X1 U7787 ( .A(n9078), .ZN(n6226) );
  NAND2_X1 U7788 ( .A1(n6226), .A2(n6482), .ZN(n6229) );
  AOI22_X1 U7789 ( .A1(n6480), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n9280), .B2(
        P1_REG0_REG_16__SCAN_IN), .ZN(n6228) );
  NAND2_X1 U7790 ( .A1(n9279), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6227) );
  OR2_X1 U7791 ( .A1(n8169), .A2(n6093), .ZN(n6230) );
  NAND2_X1 U7792 ( .A1(n6231), .A2(n6230), .ZN(n6232) );
  XNOR2_X1 U7793 ( .A(n6232), .B(n6439), .ZN(n6250) );
  NAND2_X1 U7794 ( .A1(n9083), .A2(n6436), .ZN(n6234) );
  OR2_X1 U7795 ( .A1(n8169), .A2(n6393), .ZN(n6233) );
  NAND2_X1 U7796 ( .A1(n6234), .A2(n6233), .ZN(n9074) );
  NAND2_X1 U7797 ( .A1(n7312), .A2(n9176), .ZN(n6238) );
  NAND2_X1 U7798 ( .A1(n6235), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6236) );
  XNOR2_X1 U7799 ( .A(n6236), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9513) );
  AOI22_X1 U7800 ( .A1(n6286), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6285), .B2(
        n9513), .ZN(n6237) );
  AND2_X1 U7801 ( .A1(n6239), .A2(n9502), .ZN(n6240) );
  NOR2_X1 U7802 ( .A1(n6241), .A2(n6240), .ZN(n8049) );
  NAND2_X1 U7803 ( .A1(n8049), .A2(n6482), .ZN(n6245) );
  NAND2_X1 U7804 ( .A1(n6480), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6244) );
  NAND2_X1 U7805 ( .A1(n9280), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6243) );
  NAND2_X1 U7806 ( .A1(n9279), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6242) );
  NAND4_X1 U7807 ( .A1(n6245), .A2(n6244), .A3(n6243), .A4(n6242), .ZN(n9440)
         );
  INV_X1 U7808 ( .A(n9440), .ZN(n8039) );
  OAI22_X1 U7809 ( .A1(n9859), .A2(n6391), .B1(n8039), .B2(n6093), .ZN(n6246)
         );
  XNOR2_X1 U7810 ( .A(n6246), .B(n6439), .ZN(n6251) );
  OR2_X1 U7811 ( .A1(n9859), .A2(n6093), .ZN(n6248) );
  NAND2_X1 U7812 ( .A1(n9440), .A2(n4424), .ZN(n6247) );
  NAND2_X1 U7813 ( .A1(n6248), .A2(n6247), .ZN(n9163) );
  AOI22_X1 U7814 ( .A1(n6250), .A2(n9074), .B1(n6251), .B2(n9163), .ZN(n6249)
         );
  OAI21_X1 U7815 ( .B1(n6251), .B2(n9163), .A(n9074), .ZN(n6253) );
  INV_X1 U7816 ( .A(n6250), .ZN(n9075) );
  INV_X1 U7817 ( .A(n6251), .ZN(n9073) );
  NOR2_X1 U7818 ( .A1(n9074), .A2(n9163), .ZN(n6252) );
  AOI22_X1 U7819 ( .A1(n6253), .A2(n9075), .B1(n9073), .B2(n6252), .ZN(n6254)
         );
  NAND2_X1 U7820 ( .A1(n7294), .A2(n9176), .ZN(n6257) );
  XNOR2_X1 U7821 ( .A(n6255), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9561) );
  AOI22_X1 U7822 ( .A1(n6286), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6285), .B2(
        n9561), .ZN(n6256) );
  NAND2_X1 U7823 ( .A1(n9097), .A2(n6430), .ZN(n6261) );
  INV_X1 U7824 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9538) );
  INV_X1 U7825 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9094) );
  XNOR2_X1 U7826 ( .A(n9091), .B(n9094), .ZN(n8171) );
  NAND2_X1 U7827 ( .A1(n8171), .A2(n6482), .ZN(n6259) );
  AOI22_X1 U7828 ( .A1(n9279), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9280), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n6258) );
  OAI211_X1 U7829 ( .C1(n9284), .C2(n9538), .A(n6259), .B(n6258), .ZN(n9438)
         );
  NAND2_X1 U7830 ( .A1(n9438), .A2(n6436), .ZN(n6260) );
  NAND2_X1 U7831 ( .A1(n6261), .A2(n6260), .ZN(n6262) );
  XNOR2_X1 U7832 ( .A(n6262), .B(n6439), .ZN(n6264) );
  AND2_X1 U7833 ( .A1(n9438), .A2(n4424), .ZN(n6263) );
  AOI21_X1 U7834 ( .B1(n9097), .B2(n6436), .A(n6263), .ZN(n6265) );
  XNOR2_X1 U7835 ( .A(n6264), .B(n6265), .ZN(n9086) );
  NAND2_X1 U7836 ( .A1(n9087), .A2(n9086), .ZN(n6268) );
  INV_X1 U7837 ( .A(n6264), .ZN(n6266) );
  NAND2_X1 U7838 ( .A1(n6266), .A2(n6265), .ZN(n6267) );
  NAND2_X1 U7839 ( .A1(n7318), .A2(n9176), .ZN(n6271) );
  XNOR2_X1 U7840 ( .A(n6269), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9575) );
  AOI22_X1 U7841 ( .A1(n6286), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6285), .B2(
        n9575), .ZN(n6270) );
  NAND2_X1 U7842 ( .A1(n9810), .A2(n6430), .ZN(n6277) );
  AND2_X1 U7843 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_17__SCAN_IN), 
        .ZN(n6272) );
  AOI21_X1 U7844 ( .B1(n9091), .B2(P1_REG3_REG_17__SCAN_IN), .A(
        P1_REG3_REG_18__SCAN_IN), .ZN(n6273) );
  OR2_X1 U7845 ( .A1(n6289), .A2(n6273), .ZN(n9143) );
  AOI22_X1 U7846 ( .A1(n9279), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9280), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n6275) );
  NAND2_X1 U7847 ( .A1(n6480), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6274) );
  OAI211_X1 U7848 ( .C1(n9143), .C2(n6006), .A(n6275), .B(n6274), .ZN(n9437)
         );
  NAND2_X1 U7849 ( .A1(n9437), .A2(n6436), .ZN(n6276) );
  NAND2_X1 U7850 ( .A1(n6277), .A2(n6276), .ZN(n6278) );
  XNOR2_X1 U7851 ( .A(n6278), .B(n6439), .ZN(n6280) );
  XNOR2_X1 U7852 ( .A(n6282), .B(n6280), .ZN(n9138) );
  AND2_X1 U7853 ( .A1(n9437), .A2(n4424), .ZN(n6279) );
  AOI21_X1 U7854 ( .B1(n9810), .B2(n6436), .A(n6279), .ZN(n9139) );
  INV_X1 U7855 ( .A(n6280), .ZN(n6281) );
  NAND2_X1 U7856 ( .A1(n6282), .A2(n6281), .ZN(n6283) );
  NAND2_X1 U7857 ( .A1(n7408), .A2(n9176), .ZN(n6288) );
  INV_X1 U7858 ( .A(n6284), .ZN(n9584) );
  AOI22_X1 U7859 ( .A1(n6286), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n6285), .B2(
        n9584), .ZN(n6287) );
  OR2_X1 U7860 ( .A1(n6289), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6290) );
  AND2_X1 U7861 ( .A1(n6290), .A2(n6321), .ZN(n9738) );
  NAND2_X1 U7862 ( .A1(n9738), .A2(n6482), .ZN(n6293) );
  AOI22_X1 U7863 ( .A1(n9279), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9280), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n6292) );
  NAND2_X1 U7864 ( .A1(n6480), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6291) );
  OAI22_X1 U7865 ( .A1(n9742), .A2(n6391), .B1(n9115), .B2(n6093), .ZN(n6294)
         );
  XNOR2_X1 U7866 ( .A(n6294), .B(n6418), .ZN(n6299) );
  OR2_X1 U7867 ( .A1(n9742), .A2(n6093), .ZN(n6296) );
  INV_X1 U7868 ( .A(n9115), .ZN(n9436) );
  NAND2_X1 U7869 ( .A1(n9436), .A2(n4424), .ZN(n6295) );
  NAND2_X1 U7870 ( .A1(n6296), .A2(n6295), .ZN(n6297) );
  XNOR2_X1 U7871 ( .A(n6299), .B(n6297), .ZN(n9050) );
  INV_X1 U7872 ( .A(n6297), .ZN(n6298) );
  NAND2_X1 U7873 ( .A1(n6299), .A2(n6298), .ZN(n6300) );
  NAND2_X1 U7874 ( .A1(n7432), .A2(n9176), .ZN(n6302) );
  OR2_X1 U7875 ( .A1(n6003), .A2(n7538), .ZN(n6301) );
  NAND2_X1 U7876 ( .A1(n9800), .A2(n6430), .ZN(n6310) );
  XNOR2_X1 U7877 ( .A(n6321), .B(P1_REG3_REG_20__SCAN_IN), .ZN(n9721) );
  NAND2_X1 U7878 ( .A1(n9721), .A2(n6482), .ZN(n6308) );
  INV_X1 U7879 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n6305) );
  NAND2_X1 U7880 ( .A1(n9279), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6304) );
  NAND2_X1 U7881 ( .A1(n9280), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6303) );
  OAI211_X1 U7882 ( .C1(n9284), .C2(n6305), .A(n6304), .B(n6303), .ZN(n6306)
         );
  INV_X1 U7883 ( .A(n6306), .ZN(n6307) );
  NAND2_X1 U7884 ( .A1(n6308), .A2(n6307), .ZN(n9435) );
  NAND2_X1 U7885 ( .A1(n9435), .A2(n6436), .ZN(n6309) );
  NAND2_X1 U7886 ( .A1(n6310), .A2(n6309), .ZN(n6311) );
  XNOR2_X1 U7887 ( .A(n6311), .B(n6418), .ZN(n9111) );
  AND2_X1 U7888 ( .A1(n9435), .A2(n4424), .ZN(n6312) );
  AOI21_X1 U7889 ( .B1(n9800), .B2(n6436), .A(n6312), .ZN(n9110) );
  AND2_X1 U7890 ( .A1(n9111), .A2(n9110), .ZN(n6315) );
  INV_X1 U7891 ( .A(n9111), .ZN(n6314) );
  INV_X1 U7892 ( .A(n9110), .ZN(n6313) );
  NAND2_X1 U7893 ( .A1(n7585), .A2(n9176), .ZN(n6317) );
  OR2_X1 U7894 ( .A1(n6003), .A2(n7586), .ZN(n6316) );
  INV_X1 U7895 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n6319) );
  INV_X1 U7896 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n6318) );
  OAI21_X1 U7897 ( .B1(n6321), .B2(n6319), .A(n6318), .ZN(n6322) );
  NAND2_X1 U7898 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_21__SCAN_IN), 
        .ZN(n6320) );
  AND2_X1 U7899 ( .A1(n6322), .A2(n6339), .ZN(n9703) );
  NAND2_X1 U7900 ( .A1(n9703), .A2(n6482), .ZN(n6328) );
  INV_X1 U7901 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n6325) );
  NAND2_X1 U7902 ( .A1(n9280), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6324) );
  NAND2_X1 U7903 ( .A1(n9279), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6323) );
  OAI211_X1 U7904 ( .C1(n9284), .C2(n6325), .A(n6324), .B(n6323), .ZN(n6326)
         );
  INV_X1 U7905 ( .A(n6326), .ZN(n6327) );
  OAI22_X1 U7906 ( .A1(n9705), .A2(n6391), .B1(n9116), .B2(n6093), .ZN(n6329)
         );
  XNOR2_X1 U7907 ( .A(n6329), .B(n6439), .ZN(n6332) );
  OR2_X1 U7908 ( .A1(n9705), .A2(n6093), .ZN(n6331) );
  INV_X1 U7909 ( .A(n9116), .ZN(n9434) );
  NAND2_X1 U7910 ( .A1(n9434), .A2(n4424), .ZN(n6330) );
  NAND2_X1 U7911 ( .A1(n6331), .A2(n6330), .ZN(n6333) );
  XNOR2_X1 U7912 ( .A(n6332), .B(n6333), .ZN(n9057) );
  INV_X1 U7913 ( .A(n6332), .ZN(n6335) );
  INV_X1 U7914 ( .A(n6333), .ZN(n6334) );
  NAND2_X1 U7915 ( .A1(n6335), .A2(n6334), .ZN(n6336) );
  NAND2_X1 U7916 ( .A1(n7853), .A2(n9176), .ZN(n6338) );
  OR2_X1 U7917 ( .A1(n6003), .A2(n7855), .ZN(n6337) );
  INV_X1 U7918 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9132) );
  AND2_X1 U7919 ( .A1(n6339), .A2(n9132), .ZN(n6340) );
  OR2_X1 U7920 ( .A1(n6340), .A2(n6350), .ZN(n9133) );
  INV_X1 U7921 ( .A(n9133), .ZN(n9689) );
  INV_X1 U7922 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n6343) );
  NAND2_X1 U7923 ( .A1(n9280), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6342) );
  NAND2_X1 U7924 ( .A1(n9279), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6341) );
  OAI211_X1 U7925 ( .C1(n9284), .C2(n6343), .A(n6342), .B(n6341), .ZN(n6344)
         );
  AOI21_X1 U7926 ( .B1(n9689), .B2(n6482), .A(n6344), .ZN(n9256) );
  OAI22_X1 U7927 ( .A1(n9691), .A2(n6391), .B1(n9256), .B2(n6093), .ZN(n6345)
         );
  XNOR2_X1 U7928 ( .A(n6345), .B(n6418), .ZN(n6346) );
  NOR2_X1 U7929 ( .A1(n6347), .A2(n6346), .ZN(n9123) );
  OAI22_X1 U7930 ( .A1(n9691), .A2(n6093), .B1(n9256), .B2(n6393), .ZN(n9122)
         );
  NAND2_X1 U7931 ( .A1(n7913), .A2(n9176), .ZN(n6349) );
  OR2_X1 U7932 ( .A1(n6003), .A2(n7912), .ZN(n6348) );
  NAND2_X1 U7933 ( .A1(n9785), .A2(n6430), .ZN(n6357) );
  NOR2_X1 U7934 ( .A1(n6350), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6351) );
  OR2_X1 U7935 ( .A1(n6365), .A2(n6351), .ZN(n9046) );
  INV_X1 U7936 ( .A(n9046), .ZN(n9675) );
  INV_X1 U7937 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n6354) );
  NAND2_X1 U7938 ( .A1(n9279), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6353) );
  NAND2_X1 U7939 ( .A1(n9280), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6352) );
  OAI211_X1 U7940 ( .C1(n9284), .C2(n6354), .A(n6353), .B(n6352), .ZN(n6355)
         );
  AOI21_X1 U7941 ( .B1(n9675), .B2(n6482), .A(n6355), .ZN(n9129) );
  OR2_X1 U7942 ( .A1(n9129), .A2(n6093), .ZN(n6356) );
  NAND2_X1 U7943 ( .A1(n6357), .A2(n6356), .ZN(n6358) );
  XNOR2_X1 U7944 ( .A(n6358), .B(n6418), .ZN(n6361) );
  NOR2_X1 U7945 ( .A1(n9129), .A2(n6393), .ZN(n6359) );
  AOI21_X1 U7946 ( .B1(n9785), .B2(n6436), .A(n6359), .ZN(n6360) );
  NAND2_X1 U7947 ( .A1(n6361), .A2(n6360), .ZN(n9101) );
  OR2_X1 U7948 ( .A1(n6361), .A2(n6360), .ZN(n6362) );
  NAND2_X1 U7949 ( .A1(n7981), .A2(n9176), .ZN(n6364) );
  OR2_X1 U7950 ( .A1(n6003), .A2(n8025), .ZN(n6363) );
  NAND2_X1 U7951 ( .A1(n9780), .A2(n6430), .ZN(n6374) );
  OR2_X1 U7952 ( .A1(n6365), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6366) );
  AND2_X1 U7953 ( .A1(n6366), .A2(n6386), .ZN(n9661) );
  NAND2_X1 U7954 ( .A1(n9661), .A2(n6482), .ZN(n6372) );
  INV_X1 U7955 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n6369) );
  NAND2_X1 U7956 ( .A1(n9279), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6368) );
  NAND2_X1 U7957 ( .A1(n9280), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6367) );
  OAI211_X1 U7958 ( .C1(n9284), .C2(n6369), .A(n6368), .B(n6367), .ZN(n6370)
         );
  INV_X1 U7959 ( .A(n6370), .ZN(n6371) );
  NAND2_X1 U7960 ( .A1(n6372), .A2(n6371), .ZN(n9432) );
  NAND2_X1 U7961 ( .A1(n9432), .A2(n6436), .ZN(n6373) );
  NAND2_X1 U7962 ( .A1(n6374), .A2(n6373), .ZN(n6375) );
  XNOR2_X1 U7963 ( .A(n6375), .B(n6418), .ZN(n6377) );
  AND2_X1 U7964 ( .A1(n9432), .A2(n4424), .ZN(n6376) );
  AOI21_X1 U7965 ( .B1(n9780), .B2(n6436), .A(n6376), .ZN(n6378) );
  NAND2_X1 U7966 ( .A1(n6377), .A2(n6378), .ZN(n6382) );
  INV_X1 U7967 ( .A(n6377), .ZN(n6380) );
  INV_X1 U7968 ( .A(n6378), .ZN(n6379) );
  NAND2_X1 U7969 ( .A1(n6380), .A2(n6379), .ZN(n6381) );
  NAND2_X1 U7970 ( .A1(n6382), .A2(n6381), .ZN(n9100) );
  INV_X1 U7971 ( .A(n6382), .ZN(n6383) );
  NAND2_X1 U7972 ( .A1(n8056), .A2(n9176), .ZN(n6385) );
  OR2_X1 U7973 ( .A1(n6003), .A2(n8059), .ZN(n6384) );
  INV_X1 U7974 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6931) );
  AOI21_X1 U7975 ( .B1(n6931), .B2(n6386), .A(n6396), .ZN(n9652) );
  NAND2_X1 U7976 ( .A1(n6482), .A2(n9652), .ZN(n6390) );
  NAND2_X1 U7977 ( .A1(n6480), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6389) );
  NAND2_X1 U7978 ( .A1(n9279), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6388) );
  NAND2_X1 U7979 ( .A1(n9280), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6387) );
  NAND4_X1 U7980 ( .A1(n6390), .A2(n6389), .A3(n6388), .A4(n6387), .ZN(n9431)
         );
  OAI22_X1 U7981 ( .A1(n9655), .A2(n6391), .B1(n9104), .B2(n6093), .ZN(n6392)
         );
  XNOR2_X1 U7982 ( .A(n6392), .B(n6439), .ZN(n6407) );
  OAI22_X1 U7983 ( .A1(n9655), .A2(n6093), .B1(n9104), .B2(n6393), .ZN(n6406)
         );
  XNOR2_X1 U7984 ( .A(n6407), .B(n6406), .ZN(n9065) );
  OR2_X1 U7985 ( .A1(n6003), .A2(n8098), .ZN(n6394) );
  NAND2_X1 U7986 ( .A1(n9771), .A2(n6430), .ZN(n6403) );
  NAND2_X1 U7987 ( .A1(n6396), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6411) );
  OAI21_X1 U7988 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n6396), .A(n6411), .ZN(
        n6397) );
  INV_X1 U7989 ( .A(n6397), .ZN(n9636) );
  NAND2_X1 U7990 ( .A1(n6482), .A2(n9636), .ZN(n6401) );
  NAND2_X1 U7991 ( .A1(n6480), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6400) );
  NAND2_X1 U7992 ( .A1(n9280), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6399) );
  NAND2_X1 U7993 ( .A1(n9279), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6398) );
  NAND4_X1 U7994 ( .A1(n6401), .A2(n6400), .A3(n6399), .A4(n6398), .ZN(n9430)
         );
  NAND2_X1 U7995 ( .A1(n9430), .A2(n6436), .ZN(n6402) );
  NAND2_X1 U7996 ( .A1(n6403), .A2(n6402), .ZN(n6404) );
  XNOR2_X1 U7997 ( .A(n6404), .B(n6418), .ZN(n6423) );
  AND2_X1 U7998 ( .A1(n9430), .A2(n4424), .ZN(n6405) );
  AOI21_X1 U7999 ( .B1(n9771), .B2(n6436), .A(n6405), .ZN(n6424) );
  XNOR2_X1 U8000 ( .A(n6423), .B(n6424), .ZN(n9147) );
  NOR2_X1 U8001 ( .A1(n6407), .A2(n6406), .ZN(n9148) );
  NOR2_X2 U8002 ( .A1(n9064), .A2(n6408), .ZN(n6676) );
  OR2_X1 U8003 ( .A1(n6003), .A2(n8148), .ZN(n6409) );
  NAND2_X1 U8004 ( .A1(n9766), .A2(n6430), .ZN(n6417) );
  INV_X1 U8005 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6988) );
  AOI21_X1 U8006 ( .B1(n6988), .B2(n6411), .A(n6481), .ZN(n9625) );
  NAND2_X1 U8007 ( .A1(n6482), .A2(n9625), .ZN(n6415) );
  NAND2_X1 U8008 ( .A1(n6480), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6414) );
  NAND2_X1 U8009 ( .A1(n9279), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6413) );
  NAND2_X1 U8010 ( .A1(n9280), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6412) );
  NAND4_X1 U8011 ( .A1(n6415), .A2(n6414), .A3(n6413), .A4(n6412), .ZN(n9429)
         );
  NAND2_X1 U8012 ( .A1(n9429), .A2(n6436), .ZN(n6416) );
  NAND2_X1 U8013 ( .A1(n6417), .A2(n6416), .ZN(n6419) );
  XNOR2_X1 U8014 ( .A(n6419), .B(n6418), .ZN(n6422) );
  AND2_X1 U8015 ( .A1(n9429), .A2(n4424), .ZN(n6420) );
  AOI21_X1 U8016 ( .B1(n9766), .B2(n6436), .A(n6420), .ZN(n6421) );
  NAND2_X1 U8017 ( .A1(n6422), .A2(n6421), .ZN(n6491) );
  OAI21_X1 U8018 ( .B1(n6422), .B2(n6421), .A(n6491), .ZN(n6678) );
  INV_X1 U8019 ( .A(n6423), .ZN(n6426) );
  INV_X1 U8020 ( .A(n6424), .ZN(n6425) );
  NOR2_X2 U8021 ( .A1(n6676), .A2(n6427), .ZN(n6681) );
  NAND2_X1 U8022 ( .A1(n8217), .A2(n9176), .ZN(n6429) );
  OR2_X1 U8023 ( .A1(n6003), .A2(n8219), .ZN(n6428) );
  NAND2_X1 U8024 ( .A1(n9759), .A2(n6430), .ZN(n6438) );
  INV_X1 U8025 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6432) );
  INV_X1 U8026 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n6431) );
  OAI22_X1 U8027 ( .A1(n9284), .A2(n6432), .B1(n6009), .B2(n6431), .ZN(n6435)
         );
  XNOR2_X1 U8028 ( .A(P1_REG3_REG_28__SCAN_IN), .B(n6481), .ZN(n8522) );
  INV_X1 U8029 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n6433) );
  OAI22_X1 U8030 ( .A1(n6006), .A2(n8522), .B1(n6742), .B2(n6433), .ZN(n6434)
         );
  NAND2_X1 U8031 ( .A1(n9605), .A2(n6436), .ZN(n6437) );
  NAND2_X1 U8032 ( .A1(n6438), .A2(n6437), .ZN(n6440) );
  XNOR2_X1 U8033 ( .A(n6440), .B(n6439), .ZN(n6443) );
  AOI22_X1 U8034 ( .A1(n9759), .A2(n6436), .B1(n4424), .B2(n9605), .ZN(n6442)
         );
  XNOR2_X1 U8035 ( .A(n6443), .B(n6442), .ZN(n6469) );
  INV_X1 U8036 ( .A(n6469), .ZN(n6492) );
  NAND2_X1 U8037 ( .A1(n8061), .A2(P1_B_REG_SCAN_IN), .ZN(n6445) );
  INV_X1 U8038 ( .A(n8027), .ZN(n6444) );
  MUX2_X1 U8039 ( .A(n6445), .B(P1_B_REG_SCAN_IN), .S(n6444), .Z(n6447) );
  INV_X1 U8040 ( .A(n8100), .ZN(n6446) );
  AND2_X1 U8041 ( .A1(n6447), .A2(n6446), .ZN(n6734) );
  INV_X1 U8042 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6738) );
  NAND2_X1 U8043 ( .A1(n6734), .A2(n6738), .ZN(n6448) );
  NAND2_X1 U8044 ( .A1(n8100), .A2(n8061), .ZN(n6736) );
  NAND2_X1 U8045 ( .A1(n6448), .A2(n6736), .ZN(n7435) );
  INV_X1 U8046 ( .A(n7435), .ZN(n6461) );
  INV_X1 U8047 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6449) );
  NAND2_X1 U8048 ( .A1(n6734), .A2(n6449), .ZN(n6451) );
  NAND2_X1 U8049 ( .A1(n8100), .A2(n8027), .ZN(n6450) );
  AND2_X1 U8050 ( .A1(n6451), .A2(n6450), .ZN(n9829) );
  NOR2_X1 U8051 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .ZN(
        n6791) );
  NOR4_X1 U8052 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6454) );
  NOR4_X1 U8053 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6453) );
  NOR4_X1 U8054 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6452) );
  NAND4_X1 U8055 ( .A1(n6791), .A2(n6454), .A3(n6453), .A4(n6452), .ZN(n6460)
         );
  NOR4_X1 U8056 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n6458) );
  NOR4_X1 U8057 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n6457) );
  NOR4_X1 U8058 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6456) );
  NOR4_X1 U8059 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n6455) );
  NAND4_X1 U8060 ( .A1(n6458), .A2(n6457), .A3(n6456), .A4(n6455), .ZN(n6459)
         );
  OAI21_X1 U8061 ( .B1(n6460), .B2(n6459), .A(n6734), .ZN(n7104) );
  AND3_X1 U8062 ( .A1(n6461), .A2(n9829), .A3(n7104), .ZN(n6474) );
  INV_X1 U8063 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6462) );
  NAND2_X1 U8064 ( .A1(n6463), .A2(n6462), .ZN(n6464) );
  NAND2_X1 U8065 ( .A1(n6464), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6465) );
  XNOR2_X1 U8066 ( .A(n6465), .B(n6937), .ZN(n7910) );
  AND2_X1 U8067 ( .A1(n6705), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6466) );
  AND2_X1 U8068 ( .A1(n6474), .A2(n9828), .ZN(n6479) );
  INV_X1 U8069 ( .A(n9361), .ZN(n9294) );
  NAND2_X1 U8070 ( .A1(n7854), .A2(n9294), .ZN(n7481) );
  INV_X1 U8071 ( .A(n7481), .ZN(n7552) );
  INV_X1 U8072 ( .A(n9415), .ZN(n7111) );
  NAND2_X1 U8073 ( .A1(n4429), .A2(n9361), .ZN(n9356) );
  INV_X1 U8074 ( .A(n9356), .ZN(n6752) );
  NOR2_X1 U8075 ( .A1(n10059), .A2(n6752), .ZN(n6468) );
  NAND3_X1 U8076 ( .A1(n6492), .A2(n9150), .A3(n6491), .ZN(n6497) );
  NAND2_X1 U8077 ( .A1(n6681), .A2(n6470), .ZN(n6496) );
  OR2_X1 U8078 ( .A1(n7481), .A2(n9321), .ZN(n7483) );
  INV_X1 U8079 ( .A(n7483), .ZN(n6471) );
  NAND2_X1 U8080 ( .A1(n6479), .A2(n6471), .ZN(n6473) );
  INV_X1 U8081 ( .A(n9321), .ZN(n9410) );
  INV_X1 U8082 ( .A(n7107), .ZN(n6472) );
  NAND2_X1 U8083 ( .A1(n6472), .A2(n9828), .ZN(n8523) );
  INV_X1 U8084 ( .A(n6474), .ZN(n6475) );
  NAND2_X1 U8085 ( .A1(n7107), .A2(n6475), .ZN(n6478) );
  OR2_X1 U8086 ( .A1(n9356), .A2(n9415), .ZN(n6476) );
  NAND3_X1 U8087 ( .A1(n6476), .A2(n7910), .A3(n6705), .ZN(n7106) );
  INV_X1 U8088 ( .A(n7106), .ZN(n6477) );
  NAND2_X1 U8089 ( .A1(n6478), .A2(n6477), .ZN(n9089) );
  INV_X1 U8090 ( .A(n9158), .ZN(n9168) );
  NAND2_X1 U8091 ( .A1(n6479), .A2(n9415), .ZN(n9156) );
  INV_X1 U8092 ( .A(n9156), .ZN(n9165) );
  NAND2_X1 U8093 ( .A1(n6480), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6486) );
  AND2_X1 U8094 ( .A1(n6481), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9613) );
  NAND2_X1 U8095 ( .A1(n6482), .A2(n9613), .ZN(n6485) );
  NAND2_X1 U8096 ( .A1(n9279), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6484) );
  NAND2_X1 U8097 ( .A1(n9280), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6483) );
  NAND4_X1 U8098 ( .A1(n6486), .A2(n6485), .A3(n6484), .A4(n6483), .ZN(n9428)
         );
  INV_X1 U8099 ( .A(n6487), .ZN(n7064) );
  OR2_X1 U8100 ( .A1(n9356), .A2(n7064), .ZN(n9128) );
  INV_X1 U8101 ( .A(n9128), .ZN(n9152) );
  NAND2_X1 U8102 ( .A1(n9428), .A2(n9152), .ZN(n6489) );
  NAND2_X1 U8103 ( .A1(n9429), .A2(n9604), .ZN(n6488) );
  NAND2_X1 U8104 ( .A1(n6489), .A2(n6488), .ZN(n8503) );
  AOI22_X1 U8105 ( .A1(n9165), .A2(n8503), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6490) );
  OAI21_X1 U8106 ( .B1(n8522), .B2(n9168), .A(n6490), .ZN(n6494) );
  NOR3_X1 U8107 ( .A1(n6492), .A2(n9174), .A3(n6491), .ZN(n6493) );
  AOI211_X1 U8108 ( .C1(n9759), .C2(n9171), .A(n6494), .B(n6493), .ZN(n6495)
         );
  OAI211_X1 U8109 ( .C1(n6681), .C2(n6497), .A(n6496), .B(n6495), .ZN(P1_U3220) );
  NAND2_X1 U8110 ( .A1(n6700), .A2(n6509), .ZN(n6498) );
  AOI22_X1 U8111 ( .A1(n6499), .A2(n6498), .B1(n8654), .B2(n8378), .ZN(n6508)
         );
  INV_X1 U8112 ( .A(SI_28_), .ZN(n6502) );
  NAND2_X1 U8113 ( .A1(n6503), .A2(n6502), .ZN(n6504) );
  INV_X1 U8114 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8221) );
  INV_X1 U8115 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8539) );
  MUX2_X1 U8116 ( .A(n8221), .B(n8539), .S(n5186), .Z(n8368) );
  XNOR2_X1 U8117 ( .A(n8367), .B(SI_29_), .ZN(n8220) );
  NAND2_X1 U8118 ( .A1(n8220), .A2(n8396), .ZN(n6507) );
  OR2_X1 U8119 ( .A1(n4421), .A2(n8221), .ZN(n6506) );
  NAND2_X1 U8120 ( .A1(n6518), .A2(n8234), .ZN(n8381) );
  NAND2_X1 U8121 ( .A1(n8378), .A2(n6509), .ZN(n6510) );
  AND2_X1 U8122 ( .A1(n5134), .A2(P2_B_REG_SCAN_IN), .ZN(n6512) );
  NOR2_X1 U8123 ( .A1(n10171), .A2(n6512), .ZN(n8747) );
  INV_X1 U8124 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8754) );
  NAND2_X1 U8125 ( .A1(n5155), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6514) );
  NAND2_X1 U8126 ( .A1(n5176), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6513) );
  OAI211_X1 U8127 ( .C1(n8754), .C2(n4529), .A(n6514), .B(n6513), .ZN(n6515)
         );
  INV_X1 U8128 ( .A(n6515), .ZN(n6516) );
  NAND2_X1 U8129 ( .A1(n7521), .A2(n6516), .ZN(n8652) );
  AOI22_X1 U8130 ( .A1(n8654), .A2(n8891), .B1(n8747), .B2(n8652), .ZN(n6517)
         );
  INV_X1 U8131 ( .A(n10205), .ZN(n10216) );
  INV_X1 U8132 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6520) );
  OAI21_X1 U8133 ( .B1(n6693), .B2(n10240), .A(n6522), .ZN(P2_U3456) );
  INV_X1 U8134 ( .A(n6732), .ZN(n6523) );
  OR2_X1 U8135 ( .A1(n6524), .A2(n6523), .ZN(n8732) );
  INV_X2 U8136 ( .A(n8732), .ZN(P2_U3893) );
  INV_X1 U8137 ( .A(n6525), .ZN(n7914) );
  OR2_X1 U8138 ( .A1(n8399), .A2(n7914), .ZN(n6527) );
  INV_X1 U8139 ( .A(n6524), .ZN(n6526) );
  NAND2_X1 U8140 ( .A1(n6526), .A2(n6525), .ZN(n6662) );
  NAND2_X1 U8141 ( .A1(n6527), .A2(n6662), .ZN(n6664) );
  OR2_X1 U8142 ( .A1(n6664), .A2(n5169), .ZN(n6528) );
  NAND2_X1 U8143 ( .A1(n6528), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U8144 ( .A(n8698), .ZN(n7307) );
  INV_X1 U8145 ( .A(n6618), .ZN(n10161) );
  INV_X1 U8146 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6628) );
  OAI21_X1 U8147 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n6628), .A(n6564), .ZN(n6529) );
  NAND2_X1 U8148 ( .A1(n6566), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6530) );
  NAND2_X1 U8149 ( .A1(n6529), .A2(n6530), .ZN(n7174) );
  INV_X1 U8150 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10241) );
  INV_X1 U8151 ( .A(n6530), .ZN(n6531) );
  INV_X1 U8152 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6532) );
  MUX2_X1 U8153 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6532), .S(n6632), .Z(n7190)
         );
  INV_X1 U8154 ( .A(n6632), .ZN(n7185) );
  NAND2_X1 U8155 ( .A1(n7252), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7160) );
  XNOR2_X1 U8156 ( .A(n7164), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n7161) );
  NOR2_X1 U8157 ( .A1(n7159), .A2(n5017), .ZN(n6536) );
  XNOR2_X1 U8158 ( .A(n6536), .B(n8483), .ZN(n8475) );
  INV_X1 U8159 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10246) );
  NOR2_X1 U8160 ( .A1(n8475), .A2(n10246), .ZN(n8474) );
  INV_X1 U8161 ( .A(n6536), .ZN(n6537) );
  INV_X1 U8162 ( .A(n8483), .ZN(n6714) );
  NOR2_X1 U8163 ( .A1(n8474), .A2(n5007), .ZN(n7220) );
  INV_X1 U8164 ( .A(n7220), .ZN(n6539) );
  INV_X1 U8165 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10248) );
  INV_X1 U8166 ( .A(n6642), .ZN(n7216) );
  AOI22_X1 U8167 ( .A1(n6642), .A2(P2_REG1_REG_6__SCAN_IN), .B1(n10248), .B2(
        n7216), .ZN(n7219) );
  INV_X1 U8168 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10250) );
  NAND2_X1 U8169 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n10140), .ZN(n6542) );
  OAI21_X1 U8170 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n10140), .A(n6542), .ZN(
        n10133) );
  INV_X1 U8171 ( .A(n6542), .ZN(n6543) );
  INV_X1 U8172 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10254) );
  INV_X1 U8173 ( .A(n6544), .ZN(n6545) );
  NOR2_X1 U8174 ( .A1(n6625), .A2(n6545), .ZN(n6546) );
  INV_X1 U8175 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10256) );
  AOI22_X1 U8176 ( .A1(n7704), .A2(P2_REG1_REG_10__SCAN_IN), .B1(n10256), .B2(
        n7020), .ZN(n7699) );
  INV_X1 U8177 ( .A(n7698), .ZN(n6547) );
  INV_X1 U8178 ( .A(n7993), .ZN(n7073) );
  OR2_X2 U8179 ( .A1(n6548), .A2(n7073), .ZN(n6549) );
  INV_X1 U8180 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10258) );
  INV_X1 U8181 ( .A(n6550), .ZN(n6551) );
  INV_X1 U8182 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6552) );
  MUX2_X1 U8183 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n6552), .S(n6622), .Z(n8133)
         );
  INV_X1 U8184 ( .A(n6622), .ZN(n8136) );
  NOR2_X1 U8185 ( .A1(n8186), .A2(n6553), .ZN(n6556) );
  INV_X1 U8186 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9841) );
  XNOR2_X2 U8187 ( .A(n6555), .B(n6554), .ZN(n8178) );
  INV_X1 U8188 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8113) );
  AOI22_X1 U8189 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n6618), .B1(n10161), .B2(
        n8113), .ZN(n10145) );
  NOR2_X1 U8190 ( .A1(n8679), .A2(n6557), .ZN(n6558) );
  INV_X1 U8191 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8942) );
  XNOR2_X1 U8192 ( .A(n6557), .B(n8679), .ZN(n8684) );
  NOR2_X1 U8193 ( .A1(n8942), .A2(n8684), .ZN(n8683) );
  NOR2_X1 U8194 ( .A1(n6558), .A2(n8683), .ZN(n8693) );
  INV_X1 U8195 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8936) );
  AOI22_X1 U8196 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8698), .B1(n7307), .B2(
        n8936), .ZN(n8692) );
  NOR2_X1 U8197 ( .A1(n8693), .A2(n8692), .ZN(n8691) );
  INV_X1 U8198 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8933) );
  INV_X1 U8199 ( .A(n6614), .ZN(n8720) );
  INV_X1 U8200 ( .A(n8734), .ZN(n7331) );
  NAND2_X1 U8201 ( .A1(n7331), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6560) );
  OAI21_X1 U8202 ( .B1(n7331), .B2(P2_REG1_REG_18__SCAN_IN), .A(n6560), .ZN(
        n8724) );
  NOR2_X1 U8203 ( .A1(n8725), .A2(n8724), .ZN(n8723) );
  INV_X1 U8204 ( .A(n6560), .ZN(n6561) );
  XNOR2_X1 U8205 ( .A(n7409), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n6612) );
  XNOR2_X1 U8206 ( .A(n6562), .B(n6612), .ZN(n6675) );
  NOR2_X1 U8207 ( .A1(n5110), .A2(P2_U3151), .ZN(n6665) );
  INV_X1 U8208 ( .A(n6665), .ZN(n8160) );
  NOR2_X1 U8209 ( .A1(n6664), .A2(n8160), .ZN(n10123) );
  INV_X1 U8210 ( .A(n10123), .ZN(n6563) );
  INV_X1 U8211 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8673) );
  INV_X1 U8212 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6565) );
  NAND2_X1 U8213 ( .A1(n6566), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6568) );
  INV_X1 U8214 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7385) );
  INV_X1 U8215 ( .A(n6568), .ZN(n6569) );
  INV_X1 U8216 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6570) );
  MUX2_X1 U8217 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n6570), .S(n6632), .Z(n7186)
         );
  AOI21_X1 U8218 ( .B1(n6571), .B2(n6708), .A(n6572), .ZN(n7254) );
  INV_X1 U8219 ( .A(n6572), .ZN(n7155) );
  XNOR2_X1 U8220 ( .A(n7164), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n7156) );
  INV_X1 U8221 ( .A(n6573), .ZN(n6574) );
  INV_X1 U8222 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n8478) );
  INV_X1 U8223 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6575) );
  AOI22_X1 U8224 ( .A1(n6642), .A2(P2_REG2_REG_6__SCAN_IN), .B1(n6575), .B2(
        n7216), .ZN(n7222) );
  INV_X1 U8225 ( .A(n7221), .ZN(n6577) );
  INV_X1 U8226 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7240) );
  NAND2_X1 U8227 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n10140), .ZN(n6580) );
  OAI21_X1 U8228 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n10140), .A(n6580), .ZN(
        n10131) );
  INV_X1 U8229 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7785) );
  NOR2_X1 U8230 ( .A1(n6625), .A2(n6584), .ZN(n6585) );
  INV_X1 U8231 ( .A(n7709), .ZN(n6588) );
  INV_X1 U8232 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6586) );
  MUX2_X1 U8233 ( .A(n6586), .B(P2_REG2_REG_10__SCAN_IN), .S(n7020), .Z(n7708)
         );
  NAND2_X1 U8234 ( .A1(n7020), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6589) );
  INV_X1 U8235 ( .A(n6591), .ZN(n6590) );
  NAND2_X1 U8236 ( .A1(n6590), .A2(n7993), .ZN(n6592) );
  NAND2_X1 U8237 ( .A1(n7073), .A2(n6591), .ZN(n6593) );
  INV_X1 U8238 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7989) );
  INV_X1 U8239 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6594) );
  MUX2_X1 U8240 ( .A(n6594), .B(P2_REG2_REG_12__SCAN_IN), .S(n6622), .Z(n8131)
         );
  NAND2_X1 U8241 ( .A1(n8130), .A2(n8131), .ZN(n8129) );
  NAND2_X1 U8242 ( .A1(n8136), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6595) );
  NOR2_X1 U8243 ( .A1(n8186), .A2(n6596), .ZN(n6597) );
  INV_X1 U8244 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8183) );
  INV_X1 U8245 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6598) );
  AOI22_X1 U8246 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n6618), .B1(n10161), .B2(
        n6598), .ZN(n10143) );
  NOR2_X1 U8247 ( .A1(n8679), .A2(n6601), .ZN(n6602) );
  INV_X1 U8248 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n6603) );
  MUX2_X1 U8249 ( .A(n6603), .B(P2_REG2_REG_16__SCAN_IN), .S(n8698), .Z(n6604)
         );
  INV_X1 U8250 ( .A(n6604), .ZN(n8703) );
  INV_X1 U8251 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8882) );
  NOR2_X1 U8252 ( .A1(n6614), .A2(n6606), .ZN(n6607) );
  NAND2_X1 U8253 ( .A1(n7331), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6608) );
  OAI21_X1 U8254 ( .B1(n7331), .B2(P2_REG2_REG_18__SCAN_IN), .A(n6608), .ZN(
        n8739) );
  INV_X1 U8255 ( .A(n6608), .ZN(n6609) );
  XNOR2_X1 U8256 ( .A(n7409), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n6613) );
  XNOR2_X1 U8257 ( .A(n6610), .B(n6613), .ZN(n6673) );
  AND2_X1 U8258 ( .A1(n10123), .A2(n6611), .ZN(n8741) );
  MUX2_X1 U8259 ( .A(n6613), .B(n6612), .S(n8460), .Z(n6661) );
  MUX2_X1 U8260 ( .A(n8882), .B(n8933), .S(n8460), .Z(n6615) );
  NAND2_X1 U8261 ( .A1(n6615), .A2(n6614), .ZN(n6655) );
  XNOR2_X1 U8262 ( .A(n6615), .B(n8720), .ZN(n8713) );
  MUX2_X1 U8263 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8460), .Z(n6616) );
  OR2_X1 U8264 ( .A1(n6616), .A2(n7307), .ZN(n6654) );
  XNOR2_X1 U8265 ( .A(n6616), .B(n8698), .ZN(n8696) );
  MUX2_X1 U8266 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8460), .Z(n6617) );
  OR2_X1 U8267 ( .A1(n6617), .A2(n6599), .ZN(n6653) );
  XNOR2_X1 U8268 ( .A(n6617), .B(n8679), .ZN(n8677) );
  MUX2_X1 U8269 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8460), .Z(n6619) );
  OR2_X1 U8270 ( .A1(n6619), .A2(n10161), .ZN(n6652) );
  XNOR2_X1 U8271 ( .A(n6619), .B(n6618), .ZN(n10151) );
  MUX2_X1 U8272 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8460), .Z(n6621) );
  INV_X1 U8273 ( .A(n6621), .ZN(n6620) );
  NAND2_X1 U8274 ( .A1(n8186), .A2(n6620), .ZN(n6651) );
  XNOR2_X1 U8275 ( .A(n6621), .B(n8186), .ZN(n8181) );
  MUX2_X1 U8276 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8460), .Z(n6623) );
  OR2_X1 U8277 ( .A1(n6623), .A2(n8136), .ZN(n6650) );
  XNOR2_X1 U8278 ( .A(n6623), .B(n6622), .ZN(n8141) );
  MUX2_X1 U8279 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8460), .Z(n6649) );
  XNOR2_X1 U8280 ( .A(n6649), .B(n7993), .ZN(n7986) );
  MUX2_X1 U8281 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8460), .Z(n6624) );
  OR2_X1 U8282 ( .A1(n6624), .A2(n7020), .ZN(n6648) );
  XNOR2_X1 U8283 ( .A(n6624), .B(n7704), .ZN(n7702) );
  MUX2_X1 U8284 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8460), .Z(n6626) );
  OR2_X1 U8285 ( .A1(n6626), .A2(n6582), .ZN(n6647) );
  XNOR2_X1 U8286 ( .A(n6626), .B(n6625), .ZN(n7528) );
  MUX2_X1 U8287 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8460), .Z(n6645) );
  OR2_X1 U8288 ( .A1(n6645), .A2(n10140), .ZN(n6646) );
  MUX2_X1 U8289 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8460), .Z(n6640) );
  INV_X1 U8290 ( .A(n6640), .ZN(n6641) );
  MUX2_X1 U8291 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8460), .Z(n6638) );
  INV_X1 U8292 ( .A(n6638), .ZN(n6639) );
  INV_X1 U8293 ( .A(n7164), .ZN(n6637) );
  MUX2_X1 U8294 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8460), .Z(n6635) );
  INV_X1 U8295 ( .A(n6635), .ZN(n6636) );
  MUX2_X1 U8296 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8460), .Z(n6633) );
  INV_X1 U8297 ( .A(n6633), .ZN(n6634) );
  MUX2_X1 U8298 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8460), .Z(n6630) );
  INV_X1 U8299 ( .A(n6630), .ZN(n6631) );
  MUX2_X1 U8300 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n8460), .Z(n6627) );
  INV_X1 U8301 ( .A(n6627), .ZN(n6629) );
  XNOR2_X1 U8302 ( .A(n6627), .B(n6564), .ZN(n7182) );
  MUX2_X1 U8303 ( .A(n6565), .B(n6628), .S(n8460), .Z(n10121) );
  NAND2_X1 U8304 ( .A1(n10121), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7181) );
  NAND2_X1 U8305 ( .A1(n7182), .A2(n7181), .ZN(n7180) );
  OAI21_X1 U8306 ( .B1(n6564), .B2(n6629), .A(n7180), .ZN(n7197) );
  XNOR2_X1 U8307 ( .A(n6630), .B(n6632), .ZN(n7196) );
  NAND2_X1 U8308 ( .A1(n7197), .A2(n7196), .ZN(n7195) );
  OAI21_X1 U8309 ( .B1(n6632), .B2(n6631), .A(n7195), .ZN(n7250) );
  XOR2_X1 U8310 ( .A(n6633), .B(n6708), .Z(n7251) );
  NOR2_X1 U8311 ( .A1(n7250), .A2(n7251), .ZN(n7249) );
  AOI21_X1 U8312 ( .B1(n6708), .B2(n6634), .A(n7249), .ZN(n7152) );
  XOR2_X1 U8313 ( .A(n7164), .B(n6635), .Z(n7151) );
  NAND2_X1 U8314 ( .A1(n7152), .A2(n7151), .ZN(n7150) );
  OAI21_X1 U8315 ( .B1(n6637), .B2(n6636), .A(n7150), .ZN(n8486) );
  XNOR2_X1 U8316 ( .A(n6638), .B(n8483), .ZN(n8485) );
  NAND2_X1 U8317 ( .A1(n8486), .A2(n8485), .ZN(n8484) );
  OAI21_X1 U8318 ( .B1(n8483), .B2(n6639), .A(n8484), .ZN(n7214) );
  XNOR2_X1 U8319 ( .A(n6640), .B(n7216), .ZN(n7215) );
  NOR2_X1 U8320 ( .A1(n7214), .A2(n7215), .ZN(n7213) );
  AOI21_X1 U8321 ( .B1(n6642), .B2(n6641), .A(n7213), .ZN(n7235) );
  MUX2_X1 U8322 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8460), .Z(n6643) );
  XNOR2_X1 U8323 ( .A(n6643), .B(n7237), .ZN(n7236) );
  OAI22_X1 U8324 ( .A1(n7235), .A2(n7236), .B1(n6643), .B2(n7237), .ZN(n10128)
         );
  XNOR2_X1 U8325 ( .A(n6645), .B(n6644), .ZN(n10127) );
  NAND2_X1 U8326 ( .A1(n10128), .A2(n10127), .ZN(n10126) );
  NAND2_X1 U8327 ( .A1(n6646), .A2(n10126), .ZN(n7527) );
  NAND2_X1 U8328 ( .A1(n7528), .A2(n7527), .ZN(n7526) );
  NAND2_X1 U8329 ( .A1(n6647), .A2(n7526), .ZN(n7701) );
  NAND2_X1 U8330 ( .A1(n7702), .A2(n7701), .ZN(n7700) );
  NAND2_X1 U8331 ( .A1(n6648), .A2(n7700), .ZN(n7985) );
  NAND2_X1 U8332 ( .A1(n7986), .A2(n7985), .ZN(n7984) );
  OAI21_X1 U8333 ( .B1(n6649), .B2(n7073), .A(n7984), .ZN(n8142) );
  NAND2_X1 U8334 ( .A1(n8141), .A2(n8142), .ZN(n8140) );
  NAND2_X1 U8335 ( .A1(n6650), .A2(n8140), .ZN(n8180) );
  NAND2_X1 U8336 ( .A1(n8181), .A2(n8180), .ZN(n8179) );
  NAND2_X1 U8337 ( .A1(n6651), .A2(n8179), .ZN(n10150) );
  NAND2_X1 U8338 ( .A1(n10151), .A2(n10150), .ZN(n10149) );
  NAND2_X1 U8339 ( .A1(n6652), .A2(n10149), .ZN(n8676) );
  NAND2_X1 U8340 ( .A1(n8677), .A2(n8676), .ZN(n8675) );
  NAND2_X1 U8341 ( .A1(n6653), .A2(n8675), .ZN(n8695) );
  NAND2_X1 U8342 ( .A1(n8696), .A2(n8695), .ZN(n8694) );
  NAND2_X1 U8343 ( .A1(n6654), .A2(n8694), .ZN(n8712) );
  NAND2_X1 U8344 ( .A1(n8713), .A2(n8712), .ZN(n8714) );
  NAND2_X1 U8345 ( .A1(n6655), .A2(n8714), .ZN(n6659) );
  INV_X1 U8346 ( .A(n6659), .ZN(n6657) );
  INV_X1 U8347 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8869) );
  INV_X1 U8348 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8931) );
  MUX2_X1 U8349 ( .A(n8869), .B(n8931), .S(n8460), .Z(n6658) );
  INV_X1 U8350 ( .A(n6658), .ZN(n6656) );
  NAND2_X1 U8351 ( .A1(n6657), .A2(n6656), .ZN(n8728) );
  AND2_X1 U8352 ( .A1(n6659), .A2(n6658), .ZN(n8727) );
  AOI21_X1 U8353 ( .B1(n8734), .B2(n8728), .A(n8727), .ZN(n6660) );
  XOR2_X1 U8354 ( .A(n6661), .B(n6660), .Z(n6671) );
  NAND2_X1 U8355 ( .A1(P2_U3893), .A2(n5110), .ZN(n8730) );
  INV_X1 U8356 ( .A(n6662), .ZN(n6666) );
  NOR2_X2 U8357 ( .A1(P2_U3150), .A2(n6666), .ZN(n10141) );
  NOR2_X1 U8358 ( .A1(n8460), .A2(P2_U3151), .ZN(n8127) );
  NAND2_X1 U8359 ( .A1(n8127), .A2(n5110), .ZN(n6663) );
  OR2_X1 U8360 ( .A1(n6664), .A2(n6663), .ZN(n6668) );
  NAND2_X1 U8361 ( .A1(n6666), .A2(n6665), .ZN(n6667) );
  NAND2_X1 U8362 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8570) );
  OAI21_X1 U8363 ( .B1(n10162), .B2(n7409), .A(n8570), .ZN(n6669) );
  AOI21_X1 U8364 ( .B1(P2_ADDR_REG_19__SCAN_IN), .B2(n10141), .A(n6669), .ZN(
        n6670) );
  OAI21_X1 U8365 ( .B1(n6671), .B2(n8730), .A(n6670), .ZN(n6672) );
  AOI21_X1 U8366 ( .B1(n6673), .B2(n8741), .A(n6672), .ZN(n6674) );
  OAI21_X1 U8367 ( .B1(n6675), .B2(n10147), .A(n6674), .ZN(P2_U3201) );
  INV_X1 U8368 ( .A(n6677), .ZN(n6680) );
  INV_X1 U8369 ( .A(n6678), .ZN(n6679) );
  AOI21_X1 U8370 ( .B1(n9151), .B2(n6680), .A(n6679), .ZN(n6682) );
  OAI21_X1 U8371 ( .B1(n6682), .B2(n6681), .A(n9150), .ZN(n6689) );
  INV_X1 U8372 ( .A(n9766), .ZN(n9628) );
  NAND2_X1 U8373 ( .A1(n9430), .A2(n9604), .ZN(n6684) );
  NAND2_X1 U8374 ( .A1(n9605), .A2(n9152), .ZN(n6683) );
  AND2_X1 U8375 ( .A1(n6684), .A2(n6683), .ZN(n9623) );
  OAI22_X1 U8376 ( .A1(n9156), .A2(n9623), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6988), .ZN(n6685) );
  AOI21_X1 U8377 ( .B1(n9625), .B2(n9158), .A(n6685), .ZN(n6686) );
  OAI21_X1 U8378 ( .B1(n9628), .B2(n9161), .A(n6686), .ZN(n6687) );
  NAND2_X1 U8379 ( .A1(n6689), .A2(n6688), .ZN(P1_U3214) );
  INV_X1 U8380 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6821) );
  OAI21_X1 U8381 ( .B1(n6693), .B2(n6692), .A(n6691), .ZN(P2_U3488) );
  INV_X1 U8382 ( .A(n6694), .ZN(n6697) );
  NAND2_X1 U8383 ( .A1(n10261), .A2(n10234), .ZN(n8944) );
  OAI22_X1 U8384 ( .A1(n6701), .A2(n8944), .B1(n6700), .B2(n8925), .ZN(n6695)
         );
  INV_X1 U8385 ( .A(n6695), .ZN(n6696) );
  NAND2_X1 U8386 ( .A1(n6697), .A2(n6696), .ZN(P2_U3487) );
  OR2_X1 U8387 ( .A1(n6698), .A2(n10240), .ZN(n6699) );
  NAND2_X1 U8388 ( .A1(n6699), .A2(n5004), .ZN(n6704) );
  NAND2_X1 U8389 ( .A1(n10238), .A2(n10234), .ZN(n9017) );
  OAI22_X1 U8390 ( .A1(n6701), .A2(n9017), .B1(n6700), .B2(n8989), .ZN(n6702)
         );
  INV_X1 U8391 ( .A(n6702), .ZN(n6703) );
  NAND2_X1 U8392 ( .A1(n6704), .A2(n6703), .ZN(P2_U3455) );
  NOR2_X1 U8393 ( .A1(n6705), .A2(P1_U3086), .ZN(n6706) );
  NOR2_X1 U8394 ( .A1(n8392), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9022) );
  INV_X2 U8395 ( .A(n9022), .ZN(n8549) );
  AND2_X1 U8396 ( .A1(n8392), .A2(P2_U3151), .ZN(n8159) );
  INV_X2 U8397 ( .A(n8159), .ZN(n9024) );
  OAI222_X1 U8398 ( .A1(n8549), .A2(n5121), .B1(n9024), .B2(n6722), .C1(
        P2_U3151), .C2(n6707), .ZN(P2_U3294) );
  OAI222_X1 U8399 ( .A1(n8549), .A2(n6784), .B1(n9024), .B2(n6710), .C1(
        P2_U3151), .C2(n7185), .ZN(P2_U3293) );
  OAI222_X1 U8400 ( .A1(n8549), .A2(n6709), .B1(n9024), .B2(n6712), .C1(
        P2_U3151), .C2(n4846), .ZN(P2_U3292) );
  AND2_X1 U8401 ( .A1(n8392), .A2(P1_U3086), .ZN(n9832) );
  NAND2_X1 U8402 ( .A1(n5186), .A2(P1_U3086), .ZN(n8472) );
  OAI222_X1 U8403 ( .A1(n4428), .A2(n6711), .B1(n8472), .B2(n6710), .C1(
        P1_U3086), .C2(n7054), .ZN(P1_U3353) );
  OAI222_X1 U8404 ( .A1(n4428), .A2(n6713), .B1(n8472), .B2(n6712), .C1(
        P1_U3086), .C2(n9453), .ZN(P1_U3352) );
  OAI222_X1 U8405 ( .A1(n8549), .A2(n6715), .B1(n9024), .B2(n6716), .C1(
        P2_U3151), .C2(n6714), .ZN(P2_U3290) );
  OAI222_X1 U8406 ( .A1(n4428), .A2(n6717), .B1(n8472), .B2(n6716), .C1(
        P1_U3086), .C2(n7085), .ZN(P1_U3350) );
  OAI222_X1 U8407 ( .A1(n8549), .A2(n6718), .B1(n9024), .B2(n8490), .C1(
        P2_U3151), .C2(n7164), .ZN(P2_U3291) );
  INV_X1 U8408 ( .A(n7093), .ZN(n7050) );
  OAI222_X1 U8409 ( .A1(n4428), .A2(n6719), .B1(n8472), .B2(n6720), .C1(
        P1_U3086), .C2(n7050), .ZN(P1_U3349) );
  OAI222_X1 U8410 ( .A1(n8549), .A2(n6721), .B1(n9024), .B2(n6720), .C1(
        P2_U3151), .C2(n7216), .ZN(P2_U3289) );
  INV_X1 U8411 ( .A(n8472), .ZN(n7909) );
  INV_X1 U8412 ( .A(n7909), .ZN(n9834) );
  OAI222_X1 U8413 ( .A1(n4428), .A2(n5120), .B1(n9834), .B2(n6722), .C1(
        P1_U3086), .C2(n7036), .ZN(P1_U3354) );
  INV_X1 U8414 ( .A(n7205), .ZN(n7103) );
  OAI222_X1 U8415 ( .A1(n4428), .A2(n6964), .B1(n8472), .B2(n6723), .C1(
        P1_U3086), .C2(n7103), .ZN(P1_U3348) );
  OAI222_X1 U8416 ( .A1(n8549), .A2(n6809), .B1(n9024), .B2(n6723), .C1(
        P2_U3151), .C2(n7237), .ZN(P2_U3288) );
  INV_X1 U8417 ( .A(n6724), .ZN(n6725) );
  NAND2_X1 U8418 ( .A1(n6726), .A2(n6725), .ZN(n6748) );
  INV_X1 U8419 ( .A(n6727), .ZN(n6728) );
  AOI22_X1 U8420 ( .A1(n6748), .A2(n6729), .B1(n6732), .B2(n6728), .ZN(
        P2_U3377) );
  INV_X1 U8421 ( .A(n6730), .ZN(n6731) );
  AOI22_X1 U8422 ( .A1(n6748), .A2(n6733), .B1(n6732), .B2(n6731), .ZN(
        P2_U3376) );
  INV_X1 U8423 ( .A(n6734), .ZN(n6735) );
  AND2_X1 U8424 ( .A1(n9828), .A2(n6735), .ZN(n9998) );
  NAND2_X1 U8425 ( .A1(n9998), .A2(n6736), .ZN(n6737) );
  OAI21_X1 U8426 ( .B1(n9998), .B2(n6738), .A(n6737), .ZN(P1_U3440) );
  AND2_X1 U8427 ( .A1(n6748), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8428 ( .A1(n6748), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8429 ( .A1(n6748), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8430 ( .A1(n6748), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8431 ( .A1(n6748), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8432 ( .A1(n6748), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8433 ( .A1(n6748), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8434 ( .A1(n6748), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8435 ( .A1(n6748), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8436 ( .A1(n6748), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8437 ( .A1(n6748), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8438 ( .A1(n6748), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8439 ( .A1(n6748), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8440 ( .A1(n6748), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8441 ( .A1(n6748), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8442 ( .A1(n6748), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8443 ( .A1(n6748), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8444 ( .A1(n6748), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8445 ( .A1(n6748), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8446 ( .A1(n6748), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8447 ( .A1(n6748), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8448 ( .A1(n6748), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8449 ( .A1(n6748), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  INV_X1 U8450 ( .A(n7274), .ZN(n7269) );
  OAI222_X1 U8451 ( .A1(n4428), .A2(n6939), .B1(n8472), .B2(n6739), .C1(
        P1_U3086), .C2(n7269), .ZN(P1_U3347) );
  OAI222_X1 U8452 ( .A1(n8549), .A2(n6740), .B1(n9024), .B2(n6739), .C1(
        P2_U3151), .C2(n10140), .ZN(P2_U3287) );
  INV_X1 U8453 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6747) );
  INV_X1 U8454 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6745) );
  INV_X1 U8455 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9593) );
  OR2_X1 U8456 ( .A1(n6009), .A2(n9593), .ZN(n6744) );
  INV_X1 U8457 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6741) );
  OR2_X1 U8458 ( .A1(n6742), .A2(n6741), .ZN(n6743) );
  OAI211_X1 U8459 ( .C1(n9284), .C2(n6745), .A(n6744), .B(n6743), .ZN(n9289)
         );
  NAND2_X1 U8460 ( .A1(n9289), .A2(P1_U3973), .ZN(n6746) );
  OAI21_X1 U8461 ( .B1(P1_U3973), .B2(n6747), .A(n6746), .ZN(P1_U3585) );
  INV_X1 U8462 ( .A(n6748), .ZN(n6749) );
  INV_X1 U8463 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n6914) );
  NOR2_X1 U8464 ( .A1(n6749), .A2(n6914), .ZN(P2_U3236) );
  INV_X1 U8465 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n6875) );
  NOR2_X1 U8466 ( .A1(n6749), .A2(n6875), .ZN(P2_U3248) );
  INV_X1 U8467 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n6818) );
  NOR2_X1 U8468 ( .A1(n6749), .A2(n6818), .ZN(P2_U3249) );
  INV_X1 U8469 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n6860) );
  NOR2_X1 U8470 ( .A1(n6749), .A2(n6860), .ZN(P2_U3261) );
  INV_X1 U8471 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n6862) );
  NOR2_X1 U8472 ( .A1(n6749), .A2(n6862), .ZN(P2_U3237) );
  INV_X1 U8473 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n6924) );
  NOR2_X1 U8474 ( .A1(n6749), .A2(n6924), .ZN(P2_U3242) );
  INV_X1 U8475 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n6932) );
  NOR2_X1 U8476 ( .A1(n6749), .A2(n6932), .ZN(P2_U3259) );
  NAND2_X1 U8477 ( .A1(n7910), .A2(n6750), .ZN(n6751) );
  NAND2_X1 U8478 ( .A1(n6751), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7023) );
  INV_X1 U8479 ( .A(n7023), .ZN(n6755) );
  NAND2_X1 U8480 ( .A1(n6752), .A2(n7910), .ZN(n6754) );
  NAND2_X1 U8481 ( .A1(n6754), .A2(n6753), .ZN(n7024) );
  NAND2_X1 U8482 ( .A1(n6755), .A2(n7024), .ZN(n9589) );
  INV_X1 U8483 ( .A(n9589), .ZN(n9878) );
  NOR2_X1 U8484 ( .A1(n9878), .A2(P1_U3973), .ZN(P1_U3085) );
  MUX2_X1 U8485 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n7444), .S(P1_U3973), .Z(
        n7013) );
  NAND4_X1 U8486 ( .A1(P2_REG2_REG_30__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), 
        .A3(P1_REG1_REG_29__SCAN_IN), .A4(P1_REG0_REG_21__SCAN_IN), .ZN(n6759)
         );
  NAND4_X1 U8487 ( .A1(n6866), .A2(n6887), .A3(n6937), .A4(
        P1_IR_REG_6__SCAN_IN), .ZN(n6758) );
  NAND4_X1 U8488 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(P1_REG2_REG_11__SCAN_IN), 
        .A3(P1_REG0_REG_7__SCAN_IN), .A4(P1_STATE_REG_SCAN_IN), .ZN(n6757) );
  NAND4_X1 U8489 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_1__SCAN_IN), 
        .A3(P1_WR_REG_SCAN_IN), .A4(P1_ADDR_REG_4__SCAN_IN), .ZN(n6756) );
  OR4_X1 U8490 ( .A1(n6759), .A2(n6758), .A3(n6757), .A4(n6756), .ZN(n6762) );
  INV_X1 U8491 ( .A(SI_12_), .ZN(n6949) );
  NAND4_X1 U8492 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(P2_DATAO_REG_8__SCAN_IN), 
        .A3(P1_D_REG_29__SCAN_IN), .A4(n6949), .ZN(n6761) );
  INV_X1 U8493 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6830) );
  NAND4_X1 U8494 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), 
        .A3(P1_ADDR_REG_17__SCAN_IN), .A4(n6830), .ZN(n6760) );
  NOR4_X1 U8495 ( .A1(n6762), .A2(n6761), .A3(n6760), .A4(P2_D_REG_6__SCAN_IN), 
        .ZN(n6793) );
  INV_X1 U8496 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6845) );
  INV_X1 U8497 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6848) );
  NAND4_X1 U8498 ( .A1(SI_26_), .A2(P1_REG2_REG_26__SCAN_IN), .A3(n6845), .A4(
        n6848), .ZN(n6766) );
  INV_X1 U8499 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8850) );
  NAND4_X1 U8500 ( .A1(SI_11_), .A2(n8850), .A3(n7022), .A4(n5940), .ZN(n6765)
         );
  INV_X1 U8501 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8536) );
  NAND4_X1 U8502 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P1_REG2_REG_6__SCAN_IN), 
        .A3(n6877), .A4(n8536), .ZN(n6764) );
  NAND4_X1 U8503 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_REG2_REG_24__SCAN_IN), .A4(P1_REG2_REG_22__SCAN_IN), .ZN(n6763) );
  NOR4_X1 U8504 ( .A1(n6766), .A2(n6765), .A3(n6764), .A4(n6763), .ZN(n6792)
         );
  INV_X1 U8505 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7265) );
  NAND4_X1 U8506 ( .A1(P1_REG1_REG_6__SCAN_IN), .A2(P2_REG1_REG_31__SCAN_IN), 
        .A3(n7265), .A4(n6964), .ZN(n6769) );
  INV_X1 U8507 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9554) );
  NAND4_X1 U8508 ( .A1(P2_REG2_REG_20__SCAN_IN), .A2(P1_DATAO_REG_26__SCAN_IN), 
        .A3(P1_REG0_REG_30__SCAN_IN), .A4(n9554), .ZN(n6768) );
  NOR2_X1 U8509 ( .A1(n6769), .A2(n6768), .ZN(n6773) );
  NOR4_X1 U8510 ( .A1(SI_29_), .A2(P1_DATAO_REG_19__SCAN_IN), .A3(SI_7_), .A4(
        P1_REG0_REG_27__SCAN_IN), .ZN(n6772) );
  NOR4_X1 U8511 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), 
        .A3(P1_IR_REG_24__SCAN_IN), .A4(P1_IR_REG_27__SCAN_IN), .ZN(n6771) );
  INV_X1 U8512 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9283) );
  NOR4_X1 U8513 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_DATAO_REG_31__SCAN_IN), 
        .A3(n7332), .A4(n9283), .ZN(n6770) );
  NAND4_X1 U8514 ( .A1(n6773), .A2(n6772), .A3(n6771), .A4(n6770), .ZN(n6781)
         );
  INV_X1 U8515 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n6833) );
  NAND4_X1 U8516 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P1_REG0_REG_19__SCAN_IN), 
        .A3(n6829), .A4(n6833), .ZN(n6777) );
  INV_X1 U8517 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6911) );
  NAND4_X1 U8518 ( .A1(P2_REG1_REG_22__SCAN_IN), .A2(P2_DATAO_REG_26__SCAN_IN), 
        .A3(P2_REG0_REG_10__SCAN_IN), .A4(n6911), .ZN(n6776) );
  INV_X1 U8519 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n7372) );
  NAND4_X1 U8520 ( .A1(SI_13_), .A2(P1_REG0_REG_14__SCAN_IN), .A3(
        P1_ADDR_REG_18__SCAN_IN), .A4(n7372), .ZN(n6775) );
  NAND2_X1 U8521 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P2_U3151), .ZN(n6774) );
  NOR4_X1 U8522 ( .A1(n6777), .A2(n6776), .A3(n6775), .A4(n6774), .ZN(n6779)
         );
  INV_X1 U8523 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10007) );
  NOR2_X1 U8524 ( .A1(n5614), .A2(n10007), .ZN(n6778) );
  INV_X1 U8525 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10071) );
  NAND4_X1 U8526 ( .A1(n6779), .A2(n6778), .A3(n5154), .A4(n10071), .ZN(n6780)
         );
  NOR3_X1 U8527 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(n6781), .A3(n6780), .ZN(n6783) );
  NAND4_X1 U8528 ( .A1(n4562), .A2(n6783), .A3(n6782), .A4(n5064), .ZN(n6789)
         );
  INV_X1 U8529 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10166) );
  INV_X1 U8530 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n6923) );
  NAND4_X1 U8531 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P1_REG3_REG_25__SCAN_IN), 
        .A3(n10166), .A4(n6923), .ZN(n6788) );
  NAND4_X1 U8532 ( .A1(n6808), .A2(n6784), .A3(n6821), .A4(
        P2_REG2_REG_17__SCAN_IN), .ZN(n6787) );
  NAND4_X1 U8533 ( .A1(n6785), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P2_IR_REG_11__SCAN_IN), .A4(P1_IR_REG_16__SCAN_IN), .ZN(n6786) );
  NOR4_X1 U8534 ( .A1(n6789), .A2(n6788), .A3(n6787), .A4(n6786), .ZN(n6790)
         );
  AND4_X1 U8535 ( .A1(n6793), .A2(n6792), .A3(n6791), .A4(n6790), .ZN(n6803)
         );
  INV_X1 U8536 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7201) );
  NAND4_X1 U8537 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(P2_REG3_REG_14__SCAN_IN), 
        .A3(P1_REG2_REG_4__SCAN_IN), .A4(n7201), .ZN(n6797) );
  INV_X1 U8538 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8197) );
  INV_X1 U8539 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8976) );
  NAND4_X1 U8540 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(P2_REG2_REG_1__SCAN_IN), 
        .A3(n8197), .A4(n8976), .ZN(n6796) );
  NAND4_X1 U8541 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_REG1_REG_12__SCAN_IN), 
        .A3(P1_REG3_REG_22__SCAN_IN), .A4(P2_ADDR_REG_18__SCAN_IN), .ZN(n6795)
         );
  NAND4_X1 U8542 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .A3(n6988), .A4(n5953), .ZN(n6794) );
  NOR4_X1 U8543 ( .A1(n6797), .A2(n6796), .A3(n6795), .A4(n6794), .ZN(n6801)
         );
  NOR4_X1 U8544 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(P2_REG2_REG_23__SCAN_IN), 
        .A3(P1_REG2_REG_31__SCAN_IN), .A4(n7072), .ZN(n6798) );
  NAND3_X1 U8545 ( .A1(P2_REG2_REG_25__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), 
        .A3(n6798), .ZN(n6799) );
  NOR3_X1 U8546 ( .A1(P2_REG1_REG_24__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .A3(n6799), .ZN(n6800) );
  NAND4_X1 U8547 ( .A1(n6803), .A2(n6802), .A3(n6801), .A4(n6800), .ZN(n7011)
         );
  AOI22_X1 U8548 ( .A1(n10007), .A2(keyinput88), .B1(n5614), .B2(keyinput103), 
        .ZN(n6804) );
  OAI221_X1 U8549 ( .B1(n10007), .B2(keyinput88), .C1(n5614), .C2(keyinput103), 
        .A(n6804), .ZN(n6815) );
  INV_X1 U8550 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7315) );
  INV_X1 U8551 ( .A(keyinput119), .ZN(n6806) );
  AOI22_X1 U8552 ( .A1(n7315), .A2(keyinput122), .B1(P1_WR_REG_SCAN_IN), .B2(
        n6806), .ZN(n6805) );
  OAI221_X1 U8553 ( .B1(n7315), .B2(keyinput122), .C1(n6806), .C2(
        P1_WR_REG_SCAN_IN), .A(n6805), .ZN(n6814) );
  AOI22_X1 U8554 ( .A1(n6809), .A2(keyinput11), .B1(n6808), .B2(keyinput53), 
        .ZN(n6807) );
  OAI221_X1 U8555 ( .B1(n6809), .B2(keyinput11), .C1(n6808), .C2(keyinput53), 
        .A(n6807), .ZN(n6813) );
  XNOR2_X1 U8556 ( .A(P2_IR_REG_11__SCAN_IN), .B(keyinput72), .ZN(n6811) );
  XNOR2_X1 U8557 ( .A(P2_IR_REG_7__SCAN_IN), .B(keyinput111), .ZN(n6810) );
  NAND2_X1 U8558 ( .A1(n6811), .A2(n6810), .ZN(n6812) );
  NOR4_X1 U8559 ( .A1(n6815), .A2(n6814), .A3(n6813), .A4(n6812), .ZN(n6857)
         );
  INV_X1 U8560 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n9996) );
  INV_X1 U8561 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n7848) );
  AOI22_X1 U8562 ( .A1(n9996), .A2(keyinput97), .B1(keyinput61), .B2(n7848), 
        .ZN(n6816) );
  OAI221_X1 U8563 ( .B1(n9996), .B2(keyinput97), .C1(n7848), .C2(keyinput61), 
        .A(n6816), .ZN(n6827) );
  INV_X1 U8564 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6819) );
  AOI22_X1 U8565 ( .A1(n6819), .A2(keyinput75), .B1(n6818), .B2(keyinput48), 
        .ZN(n6817) );
  OAI221_X1 U8566 ( .B1(n6819), .B2(keyinput75), .C1(n6818), .C2(keyinput48), 
        .A(n6817), .ZN(n6826) );
  AOI22_X1 U8567 ( .A1(n6821), .A2(keyinput57), .B1(n8754), .B2(keyinput6), 
        .ZN(n6820) );
  OAI221_X1 U8568 ( .B1(n6821), .B2(keyinput57), .C1(n8754), .C2(keyinput6), 
        .A(n6820), .ZN(n6825) );
  XNOR2_X1 U8569 ( .A(P1_REG0_REG_21__SCAN_IN), .B(keyinput55), .ZN(n6823) );
  XNOR2_X1 U8570 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput33), .ZN(n6822) );
  NAND2_X1 U8571 ( .A1(n6823), .A2(n6822), .ZN(n6824) );
  NOR4_X1 U8572 ( .A1(n6827), .A2(n6826), .A3(n6825), .A4(n6824), .ZN(n6856)
         );
  AOI22_X1 U8573 ( .A1(n6830), .A2(keyinput77), .B1(n6829), .B2(keyinput102), 
        .ZN(n6828) );
  OAI221_X1 U8574 ( .B1(n6830), .B2(keyinput77), .C1(n6829), .C2(keyinput102), 
        .A(n6828), .ZN(n6840) );
  INV_X1 U8575 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n6832) );
  AOI22_X1 U8576 ( .A1(n6833), .A2(keyinput10), .B1(n6832), .B2(keyinput93), 
        .ZN(n6831) );
  OAI221_X1 U8577 ( .B1(n6833), .B2(keyinput10), .C1(n6832), .C2(keyinput93), 
        .A(n6831), .ZN(n6839) );
  XNOR2_X1 U8578 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput47), .ZN(n6837) );
  XNOR2_X1 U8579 ( .A(P2_IR_REG_15__SCAN_IN), .B(keyinput44), .ZN(n6836) );
  XNOR2_X1 U8580 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(keyinput71), .ZN(n6835) );
  XNOR2_X1 U8581 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput23), .ZN(n6834) );
  NAND4_X1 U8582 ( .A1(n6837), .A2(n6836), .A3(n6835), .A4(n6834), .ZN(n6838)
         );
  NOR3_X1 U8583 ( .A1(n6840), .A2(n6839), .A3(n6838), .ZN(n6855) );
  AOI22_X1 U8584 ( .A1(n6842), .A2(keyinput2), .B1(keyinput25), .B2(n7022), 
        .ZN(n6841) );
  OAI221_X1 U8585 ( .B1(n6842), .B2(keyinput2), .C1(n7022), .C2(keyinput25), 
        .A(n6841), .ZN(n6853) );
  AOI22_X1 U8586 ( .A1(n5940), .A2(keyinput52), .B1(n8850), .B2(keyinput76), 
        .ZN(n6843) );
  OAI221_X1 U8587 ( .B1(n5940), .B2(keyinput52), .C1(n8850), .C2(keyinput76), 
        .A(n6843), .ZN(n6852) );
  AOI22_X1 U8588 ( .A1(n6846), .A2(keyinput120), .B1(n6845), .B2(keyinput118), 
        .ZN(n6844) );
  OAI221_X1 U8589 ( .B1(n6846), .B2(keyinput120), .C1(n6845), .C2(keyinput118), 
        .A(n6844), .ZN(n6851) );
  AOI22_X1 U8590 ( .A1(n6849), .A2(keyinput79), .B1(keyinput0), .B2(n6848), 
        .ZN(n6847) );
  OAI221_X1 U8591 ( .B1(n6849), .B2(keyinput79), .C1(n6848), .C2(keyinput0), 
        .A(n6847), .ZN(n6850) );
  NOR4_X1 U8592 ( .A1(n6853), .A2(n6852), .A3(n6851), .A4(n6850), .ZN(n6854)
         );
  NAND4_X1 U8593 ( .A1(n6857), .A2(n6856), .A3(n6855), .A4(n6854), .ZN(n7009)
         );
  INV_X1 U8594 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n6859) );
  AOI22_X1 U8595 ( .A1(n6860), .A2(keyinput126), .B1(keyinput51), .B2(n6859), 
        .ZN(n6858) );
  OAI221_X1 U8596 ( .B1(n6860), .B2(keyinput126), .C1(n6859), .C2(keyinput51), 
        .A(n6858), .ZN(n6872) );
  INV_X1 U8597 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6863) );
  AOI22_X1 U8598 ( .A1(n6863), .A2(keyinput89), .B1(n6862), .B2(keyinput54), 
        .ZN(n6861) );
  OAI221_X1 U8599 ( .B1(n6863), .B2(keyinput89), .C1(n6862), .C2(keyinput54), 
        .A(n6861), .ZN(n6871) );
  INV_X1 U8600 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n6865) );
  AOI22_X1 U8601 ( .A1(n6866), .A2(keyinput92), .B1(keyinput85), .B2(n6865), 
        .ZN(n6864) );
  OAI221_X1 U8602 ( .B1(n6866), .B2(keyinput92), .C1(n6865), .C2(keyinput85), 
        .A(n6864), .ZN(n6870) );
  XNOR2_X1 U8603 ( .A(P2_IR_REG_12__SCAN_IN), .B(keyinput7), .ZN(n6868) );
  XNOR2_X1 U8604 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput32), .ZN(n6867) );
  NAND2_X1 U8605 ( .A1(n6868), .A2(n6867), .ZN(n6869) );
  NOR4_X1 U8606 ( .A1(n6872), .A2(n6871), .A3(n6870), .A4(n6869), .ZN(n6909)
         );
  INV_X1 U8607 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6874) );
  AOI22_X1 U8608 ( .A1(n6875), .A2(keyinput105), .B1(keyinput121), .B2(n6874), 
        .ZN(n6873) );
  OAI221_X1 U8609 ( .B1(n6875), .B2(keyinput105), .C1(n6874), .C2(keyinput121), 
        .A(n6873), .ZN(n6884) );
  AOI22_X1 U8610 ( .A1(n8536), .A2(keyinput26), .B1(n6877), .B2(keyinput24), 
        .ZN(n6876) );
  OAI221_X1 U8611 ( .B1(n8536), .B2(keyinput26), .C1(n6877), .C2(keyinput24), 
        .A(n6876), .ZN(n6883) );
  AOI22_X1 U8612 ( .A1(n5034), .A2(keyinput104), .B1(keyinput78), .B2(n6879), 
        .ZN(n6878) );
  OAI221_X1 U8613 ( .B1(n5034), .B2(keyinput104), .C1(n6879), .C2(keyinput78), 
        .A(n6878), .ZN(n6882) );
  INV_X1 U8614 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8911) );
  INV_X1 U8615 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7830) );
  AOI22_X1 U8616 ( .A1(n8911), .A2(keyinput125), .B1(keyinput42), .B2(n7830), 
        .ZN(n6880) );
  OAI221_X1 U8617 ( .B1(n8911), .B2(keyinput125), .C1(n7830), .C2(keyinput42), 
        .A(n6880), .ZN(n6881) );
  NOR4_X1 U8618 ( .A1(n6884), .A2(n6883), .A3(n6882), .A4(n6881), .ZN(n6908)
         );
  AOI22_X1 U8619 ( .A1(n7072), .A2(keyinput28), .B1(n7297), .B2(keyinput74), 
        .ZN(n6885) );
  OAI221_X1 U8620 ( .B1(n7072), .B2(keyinput28), .C1(n7297), .C2(keyinput74), 
        .A(n6885), .ZN(n6893) );
  AOI22_X1 U8621 ( .A1(n9593), .A2(keyinput22), .B1(n6887), .B2(keyinput117), 
        .ZN(n6886) );
  OAI221_X1 U8622 ( .B1(n9593), .B2(keyinput22), .C1(n6887), .C2(keyinput117), 
        .A(n6886), .ZN(n6892) );
  INV_X1 U8623 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n9995) );
  AOI22_X1 U8624 ( .A1(n8799), .A2(keyinput5), .B1(keyinput45), .B2(n9995), 
        .ZN(n6888) );
  OAI221_X1 U8625 ( .B1(n8799), .B2(keyinput5), .C1(n9995), .C2(keyinput45), 
        .A(n6888), .ZN(n6891) );
  INV_X1 U8626 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n7523) );
  AOI22_X1 U8627 ( .A1(n5598), .A2(keyinput13), .B1(keyinput115), .B2(n7523), 
        .ZN(n6889) );
  OAI221_X1 U8628 ( .B1(n5598), .B2(keyinput13), .C1(n7523), .C2(keyinput115), 
        .A(n6889), .ZN(n6890) );
  NOR4_X1 U8629 ( .A1(n6893), .A2(n6892), .A3(n6891), .A4(n6890), .ZN(n6907)
         );
  AOI22_X1 U8630 ( .A1(n7332), .A2(keyinput46), .B1(keyinput21), .B2(n9283), 
        .ZN(n6894) );
  OAI221_X1 U8631 ( .B1(n7332), .B2(keyinput46), .C1(n9283), .C2(keyinput21), 
        .A(n6894), .ZN(n6905) );
  INV_X1 U8632 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6897) );
  INV_X1 U8633 ( .A(SI_7_), .ZN(n6896) );
  AOI22_X1 U8634 ( .A1(n6897), .A2(keyinput56), .B1(keyinput87), .B2(n6896), 
        .ZN(n6895) );
  OAI221_X1 U8635 ( .B1(n6897), .B2(keyinput56), .C1(n6896), .C2(keyinput87), 
        .A(n6895), .ZN(n6904) );
  INV_X1 U8636 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9471) );
  AOI22_X1 U8637 ( .A1(n7410), .A2(keyinput108), .B1(keyinput107), .B2(n9471), 
        .ZN(n6898) );
  OAI221_X1 U8638 ( .B1(n7410), .B2(keyinput108), .C1(n9471), .C2(keyinput107), 
        .A(n6898), .ZN(n6903) );
  INV_X1 U8639 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n6901) );
  INV_X1 U8640 ( .A(SI_29_), .ZN(n6900) );
  AOI22_X1 U8641 ( .A1(n6901), .A2(keyinput14), .B1(n6900), .B2(keyinput19), 
        .ZN(n6899) );
  OAI221_X1 U8642 ( .B1(n6901), .B2(keyinput14), .C1(n6900), .C2(keyinput19), 
        .A(n6899), .ZN(n6902) );
  NOR4_X1 U8643 ( .A1(n6905), .A2(n6904), .A3(n6903), .A4(n6902), .ZN(n6906)
         );
  NAND4_X1 U8644 ( .A1(n6909), .A2(n6908), .A3(n6907), .A4(n6906), .ZN(n7008)
         );
  AOI22_X1 U8645 ( .A1(n6911), .A2(keyinput98), .B1(keyinput90), .B2(n6207), 
        .ZN(n6910) );
  OAI221_X1 U8646 ( .B1(n6911), .B2(keyinput98), .C1(n6207), .C2(keyinput90), 
        .A(n6910), .ZN(n6921) );
  INV_X1 U8647 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10225) );
  AOI22_X1 U8648 ( .A1(n8098), .A2(keyinput64), .B1(keyinput20), .B2(n10225), 
        .ZN(n6912) );
  OAI221_X1 U8649 ( .B1(n8098), .B2(keyinput64), .C1(n10225), .C2(keyinput20), 
        .A(n6912), .ZN(n6920) );
  INV_X1 U8650 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8916) );
  AOI22_X1 U8651 ( .A1(n6914), .A2(keyinput58), .B1(keyinput8), .B2(n8916), 
        .ZN(n6913) );
  OAI221_X1 U8652 ( .B1(n6914), .B2(keyinput58), .C1(n8916), .C2(keyinput8), 
        .A(n6913), .ZN(n6919) );
  INV_X1 U8653 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n6915) );
  XOR2_X1 U8654 ( .A(n6915), .B(keyinput73), .Z(n6917) );
  XNOR2_X1 U8655 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput34), .ZN(n6916) );
  NAND2_X1 U8656 ( .A1(n6917), .A2(n6916), .ZN(n6918) );
  NOR4_X1 U8657 ( .A1(n6921), .A2(n6920), .A3(n6919), .A4(n6918), .ZN(n6960)
         );
  AOI22_X1 U8658 ( .A1(n6924), .A2(keyinput3), .B1(keyinput31), .B2(n6923), 
        .ZN(n6922) );
  OAI221_X1 U8659 ( .B1(n6924), .B2(keyinput3), .C1(n6923), .C2(keyinput31), 
        .A(n6922), .ZN(n6929) );
  INV_X1 U8660 ( .A(SI_13_), .ZN(n6926) );
  AOI22_X1 U8661 ( .A1(n7372), .A2(keyinput84), .B1(n6926), .B2(keyinput81), 
        .ZN(n6925) );
  OAI221_X1 U8662 ( .B1(n7372), .B2(keyinput84), .C1(n6926), .C2(keyinput81), 
        .A(n6925), .ZN(n6928) );
  XOR2_X1 U8663 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput39), .Z(n6927) );
  OR3_X1 U8664 ( .A1(n6929), .A2(n6928), .A3(n6927), .ZN(n6935) );
  AOI22_X1 U8665 ( .A1(n6931), .A2(keyinput15), .B1(n10166), .B2(keyinput35), 
        .ZN(n6930) );
  OAI221_X1 U8666 ( .B1(n6931), .B2(keyinput15), .C1(n10166), .C2(keyinput35), 
        .A(n6930), .ZN(n6934) );
  XNOR2_X1 U8667 ( .A(n6932), .B(keyinput95), .ZN(n6933) );
  NOR3_X1 U8668 ( .A1(n6935), .A2(n6934), .A3(n6933), .ZN(n6959) );
  INV_X1 U8669 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10047) );
  AOI22_X1 U8670 ( .A1(n6937), .A2(keyinput12), .B1(keyinput17), .B2(n10047), 
        .ZN(n6936) );
  OAI221_X1 U8671 ( .B1(n6937), .B2(keyinput12), .C1(n10047), .C2(keyinput17), 
        .A(n6936), .ZN(n6946) );
  INV_X1 U8672 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7313) );
  AOI22_X1 U8673 ( .A1(n6939), .A2(keyinput112), .B1(n7313), .B2(keyinput29), 
        .ZN(n6938) );
  OAI221_X1 U8674 ( .B1(n6939), .B2(keyinput112), .C1(n7313), .C2(keyinput29), 
        .A(n6938), .ZN(n6945) );
  INV_X1 U8675 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10267) );
  XOR2_X1 U8676 ( .A(n10267), .B(keyinput116), .Z(n6943) );
  XOR2_X1 U8677 ( .A(n5154), .B(keyinput101), .Z(n6942) );
  XNOR2_X1 U8678 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput36), .ZN(n6941) );
  XNOR2_X1 U8679 ( .A(P2_IR_REG_19__SCAN_IN), .B(keyinput82), .ZN(n6940) );
  NAND4_X1 U8680 ( .A1(n6943), .A2(n6942), .A3(n6941), .A4(n6940), .ZN(n6944)
         );
  NOR3_X1 U8681 ( .A1(n6946), .A2(n6945), .A3(n6944), .ZN(n6958) );
  INV_X1 U8682 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7802) );
  AOI22_X1 U8683 ( .A1(P1_U3086), .A2(keyinput66), .B1(keyinput91), .B2(n7802), 
        .ZN(n6947) );
  OAI221_X1 U8684 ( .B1(P1_U3086), .B2(keyinput66), .C1(n7802), .C2(keyinput91), .A(n6947), .ZN(n6956) );
  INV_X1 U8685 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n9993) );
  AOI22_X1 U8686 ( .A1(n9993), .A2(keyinput9), .B1(n6949), .B2(keyinput68), 
        .ZN(n6948) );
  OAI221_X1 U8687 ( .B1(n9993), .B2(keyinput9), .C1(n6949), .C2(keyinput68), 
        .A(n6948), .ZN(n6955) );
  XNOR2_X1 U8688 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput27), .ZN(n6953) );
  XNOR2_X1 U8689 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput1), .ZN(n6952) );
  XNOR2_X1 U8690 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput127), .ZN(n6951) );
  XNOR2_X1 U8691 ( .A(P2_REG3_REG_25__SCAN_IN), .B(keyinput59), .ZN(n6950) );
  NAND4_X1 U8692 ( .A1(n6953), .A2(n6952), .A3(n6951), .A4(n6950), .ZN(n6954)
         );
  NOR3_X1 U8693 ( .A1(n6956), .A2(n6955), .A3(n6954), .ZN(n6957) );
  NAND4_X1 U8694 ( .A1(n6960), .A2(n6959), .A3(n6958), .A4(n6957), .ZN(n7007)
         );
  INV_X1 U8695 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6962) );
  AOI22_X1 U8696 ( .A1(n6962), .A2(keyinput109), .B1(keyinput38), .B2(n10071), 
        .ZN(n6961) );
  OAI221_X1 U8697 ( .B1(n6962), .B2(keyinput109), .C1(n10071), .C2(keyinput38), 
        .A(n6961), .ZN(n6971) );
  AOI22_X1 U8698 ( .A1(n8882), .A2(keyinput60), .B1(n6964), .B2(keyinput49), 
        .ZN(n6963) );
  OAI221_X1 U8699 ( .B1(n8882), .B2(keyinput60), .C1(n6964), .C2(keyinput49), 
        .A(n6963), .ZN(n6970) );
  INV_X1 U8700 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8903) );
  AOI22_X1 U8701 ( .A1(n8903), .A2(keyinput94), .B1(n7265), .B2(keyinput70), 
        .ZN(n6965) );
  OAI221_X1 U8702 ( .B1(n8903), .B2(keyinput94), .C1(n7265), .C2(keyinput70), 
        .A(n6965), .ZN(n6969) );
  XNOR2_X1 U8703 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput114), .ZN(n6967) );
  XNOR2_X1 U8704 ( .A(keyinput99), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n6966) );
  NAND2_X1 U8705 ( .A1(n6967), .A2(n6966), .ZN(n6968) );
  NOR4_X1 U8706 ( .A1(n6971), .A2(n6970), .A3(n6969), .A4(n6968), .ZN(n7005)
         );
  INV_X1 U8707 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n6974) );
  INV_X1 U8708 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n6973) );
  AOI22_X1 U8709 ( .A1(n6974), .A2(keyinput65), .B1(keyinput80), .B2(n6973), 
        .ZN(n6972) );
  OAI221_X1 U8710 ( .B1(n6974), .B2(keyinput65), .C1(n6973), .C2(keyinput80), 
        .A(n6972), .ZN(n6981) );
  AOI22_X1 U8711 ( .A1(P2_U3151), .A2(keyinput100), .B1(keyinput41), .B2(n9554), .ZN(n6975) );
  OAI221_X1 U8712 ( .B1(P2_U3151), .B2(keyinput100), .C1(n9554), .C2(
        keyinput41), .A(n6975), .ZN(n6980) );
  AOI22_X1 U8713 ( .A1(n8083), .A2(keyinput106), .B1(n8197), .B2(keyinput96), 
        .ZN(n6976) );
  OAI221_X1 U8714 ( .B1(n8083), .B2(keyinput106), .C1(n8197), .C2(keyinput96), 
        .A(n6976), .ZN(n6979) );
  AOI22_X1 U8715 ( .A1(n8976), .A2(keyinput62), .B1(keyinput69), .B2(n7385), 
        .ZN(n6977) );
  OAI221_X1 U8716 ( .B1(n8976), .B2(keyinput62), .C1(n7385), .C2(keyinput69), 
        .A(n6977), .ZN(n6978) );
  NOR4_X1 U8717 ( .A1(n6981), .A2(n6980), .A3(n6979), .A4(n6978), .ZN(n7004)
         );
  AOI22_X1 U8718 ( .A1(n6983), .A2(keyinput86), .B1(n8931), .B2(keyinput124), 
        .ZN(n6982) );
  OAI221_X1 U8719 ( .B1(n6983), .B2(keyinput86), .C1(n8931), .C2(keyinput124), 
        .A(n6982), .ZN(n6992) );
  INV_X1 U8720 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7026) );
  AOI22_X1 U8721 ( .A1(n8942), .A2(keyinput30), .B1(keyinput123), .B2(n7026), 
        .ZN(n6984) );
  OAI221_X1 U8722 ( .B1(n8942), .B2(keyinput30), .C1(n7026), .C2(keyinput123), 
        .A(n6984), .ZN(n6991) );
  INV_X1 U8723 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n6986) );
  AOI22_X1 U8724 ( .A1(n7201), .A2(keyinput37), .B1(n6986), .B2(keyinput40), 
        .ZN(n6985) );
  OAI221_X1 U8725 ( .B1(n7201), .B2(keyinput37), .C1(n6986), .C2(keyinput40), 
        .A(n6985), .ZN(n6990) );
  INV_X1 U8726 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n9997) );
  AOI22_X1 U8727 ( .A1(n6988), .A2(keyinput83), .B1(n9997), .B2(keyinput67), 
        .ZN(n6987) );
  OAI221_X1 U8728 ( .B1(n6988), .B2(keyinput83), .C1(n9997), .C2(keyinput67), 
        .A(n6987), .ZN(n6989) );
  NOR4_X1 U8729 ( .A1(n6992), .A2(n6991), .A3(n6990), .A4(n6989), .ZN(n7003)
         );
  INV_X1 U8730 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10270) );
  INV_X1 U8731 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n9994) );
  AOI22_X1 U8732 ( .A1(n10270), .A2(keyinput63), .B1(n9994), .B2(keyinput18), 
        .ZN(n6993) );
  OAI221_X1 U8733 ( .B1(n10270), .B2(keyinput63), .C1(n9994), .C2(keyinput18), 
        .A(n6993), .ZN(n7001) );
  INV_X1 U8734 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7837) );
  AOI22_X1 U8735 ( .A1(n7837), .A2(keyinput4), .B1(n5953), .B2(keyinput43), 
        .ZN(n6994) );
  OAI221_X1 U8736 ( .B1(n7837), .B2(keyinput4), .C1(n5953), .C2(keyinput43), 
        .A(n6994), .ZN(n7000) );
  AOI22_X1 U8737 ( .A1(n6552), .A2(keyinput110), .B1(keyinput113), .B2(n9132), 
        .ZN(n6995) );
  OAI221_X1 U8738 ( .B1(n6552), .B2(keyinput110), .C1(n9132), .C2(keyinput113), 
        .A(n6995), .ZN(n6999) );
  INV_X1 U8739 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9559) );
  XOR2_X1 U8740 ( .A(n9559), .B(keyinput50), .Z(n6997) );
  XNOR2_X1 U8741 ( .A(P2_IR_REG_18__SCAN_IN), .B(keyinput16), .ZN(n6996) );
  NAND2_X1 U8742 ( .A1(n6997), .A2(n6996), .ZN(n6998) );
  NOR4_X1 U8743 ( .A1(n7001), .A2(n7000), .A3(n6999), .A4(n6998), .ZN(n7002)
         );
  NAND4_X1 U8744 ( .A1(n7005), .A2(n7004), .A3(n7003), .A4(n7002), .ZN(n7006)
         );
  NOR4_X1 U8745 ( .A1(n7009), .A2(n7008), .A3(n7007), .A4(n7006), .ZN(n7010)
         );
  XOR2_X1 U8746 ( .A(n7011), .B(n7010), .Z(n7012) );
  XNOR2_X1 U8747 ( .A(n7013), .B(n7012), .ZN(P1_U3556) );
  INV_X1 U8748 ( .A(n7014), .ZN(n7016) );
  OAI222_X1 U8749 ( .A1(n9024), .A2(n7016), .B1(n6582), .B2(P2_U3151), .C1(
        n7015), .C2(n8549), .ZN(P2_U3286) );
  INV_X1 U8750 ( .A(n7337), .ZN(n7279) );
  OAI222_X1 U8751 ( .A1(n4428), .A2(n7017), .B1(n8472), .B2(n7016), .C1(n7279), 
        .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U8752 ( .A(n7018), .ZN(n7021) );
  OAI222_X1 U8753 ( .A1(n9024), .A2(n7021), .B1(n7020), .B2(P2_U3151), .C1(
        n7019), .C2(n8549), .ZN(P2_U3285) );
  INV_X1 U8754 ( .A(n7565), .ZN(n7346) );
  OAI222_X1 U8755 ( .A1(n4428), .A2(n7022), .B1(n8472), .B2(n7021), .C1(n7346), 
        .C2(P1_U3086), .ZN(P1_U3345) );
  OR2_X1 U8756 ( .A1(n7024), .A2(n7023), .ZN(n9877) );
  OR2_X1 U8757 ( .A1(n9877), .A2(n7064), .ZN(n9578) );
  AOI22_X1 U8758 ( .A1(n9884), .A2(n5926), .B1(P1_REG2_REG_1__SCAN_IN), .B2(
        n7036), .ZN(n9881) );
  NAND2_X1 U8759 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9882) );
  NOR2_X1 U8760 ( .A1(n9881), .A2(n9882), .ZN(n9880) );
  AOI21_X1 U8761 ( .B1(P1_REG2_REG_1__SCAN_IN), .B2(n9884), .A(n9880), .ZN(
        n7057) );
  AOI22_X1 U8762 ( .A1(n7035), .A2(n5963), .B1(P1_REG2_REG_2__SCAN_IN), .B2(
        n7054), .ZN(n7056) );
  NOR2_X1 U8763 ( .A1(n7057), .A2(n7056), .ZN(n7055) );
  NAND2_X1 U8764 ( .A1(n7033), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7025) );
  OAI21_X1 U8765 ( .B1(n7033), .B2(P1_REG2_REG_3__SCAN_IN), .A(n7025), .ZN(
        n9457) );
  NOR2_X1 U8766 ( .A1(n9458), .A2(n9457), .ZN(n9456) );
  AOI21_X1 U8767 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(n7033), .A(n9456), .ZN(
        n9468) );
  AOI22_X1 U8768 ( .A1(n9473), .A2(n7026), .B1(P1_REG2_REG_4__SCAN_IN), .B2(
        n8491), .ZN(n9467) );
  NAND2_X1 U8769 ( .A1(n7031), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n7027) );
  OAI21_X1 U8770 ( .B1(n7031), .B2(P1_REG2_REG_5__SCAN_IN), .A(n7027), .ZN(
        n7077) );
  XNOR2_X1 U8771 ( .A(n7093), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n7029) );
  NOR2_X1 U8772 ( .A1(n7029), .A2(n7030), .ZN(n7088) );
  OR2_X1 U8773 ( .A1(n6487), .A2(n4426), .ZN(n7065) );
  OR2_X1 U8774 ( .A1(n9877), .A2(n7065), .ZN(n9879) );
  AOI211_X1 U8775 ( .C1(n7030), .C2(n7029), .A(n7088), .B(n9879), .ZN(n7046)
         );
  NAND2_X1 U8776 ( .A1(n7031), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n7039) );
  INV_X1 U8777 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7032) );
  MUX2_X1 U8778 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n7032), .S(n7031), .Z(n7080)
         );
  INV_X1 U8779 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10103) );
  MUX2_X1 U8780 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10103), .S(n9473), .Z(n9475)
         );
  NAND2_X1 U8781 ( .A1(n7033), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7038) );
  MUX2_X1 U8782 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n7034), .S(n7033), .Z(n9461)
         );
  AOI22_X1 U8783 ( .A1(n7035), .A2(P1_REG1_REG_2__SCAN_IN), .B1(n5967), .B2(
        n7054), .ZN(n7052) );
  INV_X1 U8784 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10099) );
  MUX2_X1 U8785 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n10099), .S(n9884), .Z(n9889)
         );
  NAND3_X1 U8786 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .A3(n9889), .ZN(n9887) );
  OAI21_X1 U8787 ( .B1(n10099), .B2(n7036), .A(n9887), .ZN(n7051) );
  NAND2_X1 U8788 ( .A1(n7052), .A2(n7051), .ZN(n7037) );
  OAI21_X1 U8789 ( .B1(n5967), .B2(n7054), .A(n7037), .ZN(n9462) );
  NAND2_X1 U8790 ( .A1(n9461), .A2(n9462), .ZN(n9460) );
  NAND2_X1 U8791 ( .A1(n7038), .A2(n9460), .ZN(n9476) );
  NAND2_X1 U8792 ( .A1(n9475), .A2(n9476), .ZN(n9474) );
  OAI21_X1 U8793 ( .B1(n8491), .B2(n10103), .A(n9474), .ZN(n7081) );
  NAND2_X1 U8794 ( .A1(n7080), .A2(n7081), .ZN(n7079) );
  NAND2_X1 U8795 ( .A1(n7039), .A2(n7079), .ZN(n7041) );
  INV_X1 U8796 ( .A(n7041), .ZN(n7044) );
  INV_X1 U8797 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10106) );
  MUX2_X1 U8798 ( .A(n10106), .B(P1_REG1_REG_6__SCAN_IN), .S(n7093), .Z(n7043)
         );
  MUX2_X1 U8799 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10106), .S(n7093), .Z(n7040)
         );
  NAND2_X1 U8800 ( .A1(n7041), .A2(n7040), .ZN(n7096) );
  INV_X1 U8801 ( .A(n7096), .ZN(n7042) );
  INV_X1 U8802 ( .A(n4426), .ZN(n8544) );
  OR2_X1 U8803 ( .A1(n9877), .A2(n8544), .ZN(n9579) );
  AOI211_X1 U8804 ( .C1(n7044), .C2(n7043), .A(n7042), .B(n9579), .ZN(n7045)
         );
  NOR2_X1 U8805 ( .A1(n7046), .A2(n7045), .ZN(n7049) );
  AND2_X1 U8806 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7047) );
  AOI21_X1 U8807 ( .B1(n9878), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n7047), .ZN(
        n7048) );
  OAI211_X1 U8808 ( .C1(n7050), .C2(n9578), .A(n7049), .B(n7048), .ZN(P1_U3249) );
  INV_X1 U8809 ( .A(n9579), .ZN(n9888) );
  XOR2_X1 U8810 ( .A(n7052), .B(n7051), .Z(n7060) );
  AOI22_X1 U8811 ( .A1(n9878), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n7053) );
  OAI21_X1 U8812 ( .B1(n7054), .B2(n9578), .A(n7053), .ZN(n7059) );
  AOI211_X1 U8813 ( .C1(n7057), .C2(n7056), .A(n7055), .B(n9879), .ZN(n7058)
         );
  AOI211_X1 U8814 ( .C1(n9888), .C2(n7060), .A(n7059), .B(n7058), .ZN(n7070)
         );
  OAI21_X1 U8815 ( .B1(n7063), .B2(n7062), .A(n7061), .ZN(n7135) );
  NAND3_X1 U8816 ( .A1(n7135), .A2(n7064), .A3(n4426), .ZN(n7069) );
  INV_X1 U8817 ( .A(n7065), .ZN(n9411) );
  INV_X1 U8818 ( .A(n9882), .ZN(n7067) );
  NOR2_X1 U8819 ( .A1(n4426), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n7066) );
  NOR2_X1 U8820 ( .A1(n7066), .A2(n6487), .ZN(n9870) );
  NOR2_X1 U8821 ( .A1(n9870), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n9869) );
  AOI21_X1 U8822 ( .B1(n9411), .B2(n7067), .A(n9869), .ZN(n7068) );
  NAND3_X1 U8823 ( .A1(n7069), .A2(P1_U3973), .A3(n7068), .ZN(n9478) );
  NAND2_X1 U8824 ( .A1(n7070), .A2(n9478), .ZN(P1_U3245) );
  INV_X1 U8825 ( .A(n7071), .ZN(n7074) );
  INV_X1 U8826 ( .A(n7666), .ZN(n7660) );
  OAI222_X1 U8827 ( .A1(n4428), .A2(n7072), .B1(n9834), .B2(n7074), .C1(
        P1_U3086), .C2(n7660), .ZN(P1_U3344) );
  OAI222_X1 U8828 ( .A1(n8549), .A2(n7075), .B1(n9024), .B2(n7074), .C1(
        P2_U3151), .C2(n7073), .ZN(P2_U3284) );
  AOI211_X1 U8829 ( .C1(n7078), .C2(n7077), .A(n7076), .B(n9879), .ZN(n7087)
         );
  OAI211_X1 U8830 ( .C1(n7081), .C2(n7080), .A(n9888), .B(n7079), .ZN(n7084)
         );
  NOR2_X1 U8831 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7372), .ZN(n7082) );
  AOI21_X1 U8832 ( .B1(n9878), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n7082), .ZN(
        n7083) );
  OAI211_X1 U8833 ( .C1(n9578), .C2(n7085), .A(n7084), .B(n7083), .ZN(n7086)
         );
  OR2_X1 U8834 ( .A1(n7087), .A2(n7086), .ZN(P1_U3248) );
  INV_X1 U8835 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7089) );
  MUX2_X1 U8836 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n7089), .S(n7205), .Z(n7090)
         );
  INV_X1 U8837 ( .A(n7090), .ZN(n7091) );
  NOR2_X1 U8838 ( .A1(n7092), .A2(n7091), .ZN(n7204) );
  AOI211_X1 U8839 ( .C1(n7092), .C2(n7091), .A(n7204), .B(n9879), .ZN(n7099)
         );
  NAND2_X1 U8840 ( .A1(n7093), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7095) );
  INV_X1 U8841 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10108) );
  MUX2_X1 U8842 ( .A(n10108), .B(P1_REG1_REG_7__SCAN_IN), .S(n7205), .Z(n7094)
         );
  AOI21_X1 U8843 ( .B1(n7096), .B2(n7095), .A(n7094), .ZN(n7200) );
  AND3_X1 U8844 ( .A1(n7096), .A2(n7095), .A3(n7094), .ZN(n7097) );
  NOR3_X1 U8845 ( .A1(n9579), .A2(n7200), .A3(n7097), .ZN(n7098) );
  NOR2_X1 U8846 ( .A1(n7099), .A2(n7098), .ZN(n7102) );
  NOR2_X1 U8847 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7545), .ZN(n7100) );
  AOI21_X1 U8848 ( .B1(n9878), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n7100), .ZN(
        n7101) );
  OAI211_X1 U8849 ( .C1(n7103), .C2(n9578), .A(n7102), .B(n7101), .ZN(P1_U3250) );
  NAND2_X1 U8850 ( .A1(n7104), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7105) );
  OR2_X1 U8851 ( .A1(n7106), .A2(n7105), .ZN(n7434) );
  NAND2_X1 U8852 ( .A1(n7107), .A2(n7435), .ZN(n7108) );
  NOR2_X1 U8853 ( .A1(n7434), .A2(n7108), .ZN(n7118) );
  INV_X1 U8854 ( .A(n9829), .ZN(n7109) );
  AND2_X2 U8855 ( .A1(n7118), .A2(n7109), .ZN(n10098) );
  INV_X1 U8856 ( .A(n7550), .ZN(n9986) );
  NAND2_X1 U8857 ( .A1(n4429), .A2(n9584), .ZN(n7110) );
  NAND2_X1 U8858 ( .A1(n9361), .A2(n9410), .ZN(n9326) );
  NAND2_X1 U8859 ( .A1(n7110), .A2(n9326), .ZN(n9980) );
  OR2_X1 U8860 ( .A1(n7112), .A2(n7477), .ZN(n7551) );
  NAND2_X1 U8861 ( .A1(n7112), .A2(n7111), .ZN(n7113) );
  NAND3_X1 U8862 ( .A1(n7551), .A2(n7481), .A3(n7113), .ZN(n10048) );
  OAI21_X1 U8863 ( .B1(n7114), .B2(n7550), .A(n9974), .ZN(n9295) );
  INV_X1 U8864 ( .A(n9295), .ZN(n7115) );
  OAI21_X1 U8865 ( .B1(n9980), .B2(n10095), .A(n7115), .ZN(n7116) );
  NAND2_X1 U8866 ( .A1(n7440), .A2(n9152), .ZN(n7553) );
  OAI211_X1 U8867 ( .C1(n7481), .C2(n9986), .A(n7116), .B(n7553), .ZN(n7119)
         );
  NAND2_X1 U8868 ( .A1(n7119), .A2(n10098), .ZN(n7117) );
  OAI21_X1 U8869 ( .B1(n10098), .B2(n5941), .A(n7117), .ZN(P1_U3453) );
  AND2_X2 U8870 ( .A1(n7118), .A2(n9829), .ZN(n10120) );
  NAND2_X1 U8871 ( .A1(n7119), .A2(n10120), .ZN(n7120) );
  OAI21_X1 U8872 ( .B1(n10120), .B2(n5953), .A(n7120), .ZN(P1_U3522) );
  OAI21_X1 U8873 ( .B1(n7123), .B2(n7122), .A(n7121), .ZN(n7124) );
  NAND2_X1 U8874 ( .A1(n7124), .A2(n9150), .ZN(n7128) );
  INV_X1 U8875 ( .A(n7114), .ZN(n7125) );
  INV_X1 U8876 ( .A(n9604), .ZN(n9114) );
  OAI22_X1 U8877 ( .A1(n7125), .A2(n9114), .B1(n7443), .B2(n9128), .ZN(n9978)
         );
  INV_X1 U8878 ( .A(n9089), .ZN(n7126) );
  NAND2_X1 U8879 ( .A1(n7126), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7145) );
  AOI22_X1 U8880 ( .A1(n9978), .A2(n9165), .B1(n7145), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n7127) );
  OAI211_X1 U8881 ( .C1(n7439), .C2(n9161), .A(n7128), .B(n7127), .ZN(P1_U3222) );
  INV_X1 U8882 ( .A(P1_U3973), .ZN(n9452) );
  NAND2_X1 U8883 ( .A1(n9452), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7129) );
  OAI21_X1 U8884 ( .B1(n9129), .B2(n9452), .A(n7129), .ZN(P1_U3577) );
  INV_X1 U8885 ( .A(n7130), .ZN(n7136) );
  OAI222_X1 U8886 ( .A1(n9024), .A2(n7136), .B1(n8136), .B2(P2_U3151), .C1(
        n7131), .C2(n8549), .ZN(P2_U3283) );
  INV_X1 U8887 ( .A(n7145), .ZN(n7132) );
  OAI22_X1 U8888 ( .A1(n7132), .A2(n7554), .B1(n9156), .B2(n7553), .ZN(n7133)
         );
  AOI21_X1 U8889 ( .B1(n7550), .B2(n9171), .A(n7133), .ZN(n7134) );
  OAI21_X1 U8890 ( .B1(n9174), .B2(n7135), .A(n7134), .ZN(P1_U3232) );
  INV_X1 U8891 ( .A(n7921), .ZN(n7661) );
  OAI222_X1 U8892 ( .A1(n4428), .A2(n7137), .B1(n9834), .B2(n7136), .C1(n7661), 
        .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U8893 ( .A(n7138), .ZN(n7148) );
  AOI22_X1 U8894 ( .A1(n8186), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n9022), .ZN(n7139) );
  OAI21_X1 U8895 ( .B1(n7148), .B2(n9024), .A(n7139), .ZN(P2_U3282) );
  INV_X1 U8896 ( .A(n7442), .ZN(n7460) );
  XNOR2_X1 U8897 ( .A(n7141), .B(n7140), .ZN(n7142) );
  NAND2_X1 U8898 ( .A1(n7142), .A2(n9150), .ZN(n7147) );
  NAND2_X1 U8899 ( .A1(n7440), .A2(n9604), .ZN(n7144) );
  NAND2_X1 U8900 ( .A1(n7463), .A2(n9152), .ZN(n7143) );
  NAND2_X1 U8901 ( .A1(n7144), .A2(n7143), .ZN(n7594) );
  AOI22_X1 U8902 ( .A1(n9165), .A2(n7594), .B1(n7145), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n7146) );
  OAI211_X1 U8903 ( .C1(n7460), .C2(n9161), .A(n7147), .B(n7146), .ZN(P1_U3237) );
  INV_X1 U8904 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n7149) );
  INV_X1 U8905 ( .A(n9484), .ZN(n9492) );
  OAI222_X1 U8906 ( .A1(n4428), .A2(n7149), .B1(n9834), .B2(n7148), .C1(
        P1_U3086), .C2(n9492), .ZN(P1_U3342) );
  INV_X1 U8907 ( .A(n10141), .ZN(n8682) );
  INV_X1 U8908 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7170) );
  INV_X1 U8909 ( .A(n8730), .ZN(n10152) );
  OAI211_X1 U8910 ( .C1(n7152), .C2(n7151), .A(n7150), .B(n10152), .ZN(n7169)
         );
  INV_X1 U8911 ( .A(n7153), .ZN(n7158) );
  NAND3_X1 U8912 ( .A1(n7154), .A2(n7156), .A3(n7155), .ZN(n7157) );
  INV_X1 U8913 ( .A(n8741), .ZN(n10156) );
  AOI21_X1 U8914 ( .B1(n7158), .B2(n7157), .A(n10156), .ZN(n7167) );
  INV_X1 U8915 ( .A(n7159), .ZN(n7163) );
  NAND3_X1 U8916 ( .A1(n7253), .A2(n7161), .A3(n4848), .ZN(n7162) );
  AOI21_X1 U8917 ( .B1(n7163), .B2(n7162), .A(n10147), .ZN(n7166) );
  NAND2_X1 U8918 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3151), .ZN(n7324) );
  OAI21_X1 U8919 ( .B1(n10162), .B2(n7164), .A(n7324), .ZN(n7165) );
  NOR3_X1 U8920 ( .A1(n7167), .A2(n7166), .A3(n7165), .ZN(n7168) );
  OAI211_X1 U8921 ( .C1(n8682), .C2(n7170), .A(n7169), .B(n7168), .ZN(P2_U3186) );
  INV_X1 U8922 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7171) );
  OAI22_X1 U8923 ( .A1(n10162), .A2(n6707), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7171), .ZN(n7179) );
  AOI21_X1 U8924 ( .B1(n7385), .B2(n7173), .A(n7172), .ZN(n7177) );
  AOI21_X1 U8925 ( .B1(n10241), .B2(n7174), .A(n7175), .ZN(n7176) );
  OAI22_X1 U8926 ( .A1(n10156), .A2(n7177), .B1(n7176), .B2(n10147), .ZN(n7178) );
  AOI211_X1 U8927 ( .C1(n10141), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n7179), .B(
        n7178), .ZN(n7184) );
  OAI211_X1 U8928 ( .C1(n7182), .C2(n7181), .A(n7180), .B(n10152), .ZN(n7183)
         );
  NAND2_X1 U8929 ( .A1(n7184), .A2(n7183), .ZN(P2_U3183) );
  OAI22_X1 U8930 ( .A1(n10162), .A2(n7185), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10166), .ZN(n7194) );
  AOI21_X1 U8931 ( .B1(n7187), .B2(n7186), .A(n4525), .ZN(n7192) );
  AOI21_X1 U8932 ( .B1(n7188), .B2(n7190), .A(n7189), .ZN(n7191) );
  OAI22_X1 U8933 ( .A1(n10156), .A2(n7192), .B1(n7191), .B2(n10147), .ZN(n7193) );
  AOI211_X1 U8934 ( .C1(n10141), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n7194), .B(
        n7193), .ZN(n7199) );
  OAI211_X1 U8935 ( .C1(n7197), .C2(n7196), .A(n7195), .B(n10152), .ZN(n7198)
         );
  NAND2_X1 U8936 ( .A1(n7199), .A2(n7198), .ZN(P2_U3184) );
  INV_X1 U8937 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10110) );
  MUX2_X1 U8938 ( .A(n10110), .B(P1_REG1_REG_8__SCAN_IN), .S(n7274), .Z(n7266)
         );
  AOI21_X1 U8939 ( .B1(n7205), .B2(P1_REG1_REG_7__SCAN_IN), .A(n7200), .ZN(
        n7267) );
  XOR2_X1 U8940 ( .A(n7266), .B(n7267), .Z(n7211) );
  NOR2_X1 U8941 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7201), .ZN(n7202) );
  AOI21_X1 U8942 ( .B1(n9878), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n7202), .ZN(
        n7203) );
  OAI21_X1 U8943 ( .B1(n7269), .B2(n9578), .A(n7203), .ZN(n7210) );
  INV_X1 U8944 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7206) );
  AOI22_X1 U8945 ( .A1(n7274), .A2(n7206), .B1(P1_REG2_REG_8__SCAN_IN), .B2(
        n7269), .ZN(n7207) );
  AOI211_X1 U8946 ( .C1(n7208), .C2(n7207), .A(n7273), .B(n9879), .ZN(n7209)
         );
  AOI211_X1 U8947 ( .C1(n7211), .C2(n9888), .A(n7210), .B(n7209), .ZN(n7212)
         );
  INV_X1 U8948 ( .A(n7212), .ZN(P1_U3251) );
  AOI21_X1 U8949 ( .B1(n7215), .B2(n7214), .A(n7213), .ZN(n7229) );
  NAND2_X1 U8950 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3151), .ZN(n7414) );
  OAI21_X1 U8951 ( .B1(n10162), .B2(n7216), .A(n7414), .ZN(n7227) );
  INV_X1 U8952 ( .A(n7217), .ZN(n7218) );
  AOI21_X1 U8953 ( .B1(n7220), .B2(n7219), .A(n7218), .ZN(n7225) );
  AOI21_X1 U8954 ( .B1(n7223), .B2(n7222), .A(n7221), .ZN(n7224) );
  OAI22_X1 U8955 ( .A1(n7225), .A2(n10147), .B1(n7224), .B2(n10156), .ZN(n7226) );
  AOI211_X1 U8956 ( .C1(n10141), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n7227), .B(
        n7226), .ZN(n7228) );
  OAI21_X1 U8957 ( .B1(n7229), .B2(n8730), .A(n7228), .ZN(P2_U3188) );
  XOR2_X1 U8958 ( .A(n7231), .B(n7230), .Z(n7234) );
  OAI22_X1 U8959 ( .A1(n7467), .A2(n9128), .B1(n7443), .B2(n9114), .ZN(n9958)
         );
  AOI22_X1 U8960 ( .A1(n9171), .A2(n9960), .B1(n9165), .B2(n9958), .ZN(n7233)
         );
  MUX2_X1 U8961 ( .A(n9168), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n7232) );
  OAI211_X1 U8962 ( .C1(n7234), .C2(n9174), .A(n7233), .B(n7232), .ZN(P1_U3218) );
  XOR2_X1 U8963 ( .A(n7236), .B(n7235), .Z(n7248) );
  NAND2_X1 U8964 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7508) );
  OAI21_X1 U8965 ( .B1(n10162), .B2(n7237), .A(n7508), .ZN(n7246) );
  AOI21_X1 U8966 ( .B1(n7240), .B2(n7239), .A(n7238), .ZN(n7244) );
  AOI21_X1 U8967 ( .B1(n10250), .B2(n7242), .A(n7241), .ZN(n7243) );
  OAI22_X1 U8968 ( .A1(n10156), .A2(n7244), .B1(n7243), .B2(n10147), .ZN(n7245) );
  AOI211_X1 U8969 ( .C1(n10141), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n7246), .B(
        n7245), .ZN(n7247) );
  OAI21_X1 U8970 ( .B1(n7248), .B2(n8730), .A(n7247), .ZN(P2_U3189) );
  AOI21_X1 U8971 ( .B1(n7251), .B2(n7250), .A(n7249), .ZN(n7261) );
  INV_X1 U8972 ( .A(n10147), .ZN(n7257) );
  OAI21_X1 U8973 ( .B1(n7252), .B2(P2_REG1_REG_3__SCAN_IN), .A(n7253), .ZN(
        n7256) );
  OAI21_X1 U8974 ( .B1(n7254), .B2(P2_REG2_REG_3__SCAN_IN), .A(n7154), .ZN(
        n7255) );
  AOI22_X1 U8975 ( .A1(n7257), .A2(n7256), .B1(n8741), .B2(n7255), .ZN(n7258)
         );
  NAND2_X1 U8976 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7391) );
  OAI211_X1 U8977 ( .C1(n10162), .C2(n4846), .A(n7258), .B(n7391), .ZN(n7259)
         );
  AOI21_X1 U8978 ( .B1(n10141), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n7259), .ZN(
        n7260) );
  OAI21_X1 U8979 ( .B1(n7261), .B2(n8730), .A(n7260), .ZN(P2_U3185) );
  INV_X1 U8980 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7263) );
  INV_X1 U8981 ( .A(n7262), .ZN(n7264) );
  OAI222_X1 U8982 ( .A1(n4428), .A2(n7263), .B1(n9834), .B2(n7264), .C1(
        P1_U3086), .C2(n9505), .ZN(P1_U3341) );
  OAI222_X1 U8983 ( .A1(n8549), .A2(n7265), .B1(n9024), .B2(n7264), .C1(
        P2_U3151), .C2(n10161), .ZN(P2_U3281) );
  INV_X1 U8984 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10112) );
  AOI22_X1 U8985 ( .A1(n7337), .A2(n10112), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n7279), .ZN(n7271) );
  OR2_X1 U8986 ( .A1(n7267), .A2(n7266), .ZN(n7268) );
  OAI21_X1 U8987 ( .B1(n10110), .B2(n7269), .A(n7268), .ZN(n7270) );
  NOR2_X1 U8988 ( .A1(n7271), .A2(n7270), .ZN(n7338) );
  AOI21_X1 U8989 ( .B1(n7271), .B2(n7270), .A(n7338), .ZN(n7283) );
  NOR2_X1 U8990 ( .A1(n7337), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7272) );
  AOI21_X1 U8991 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n7337), .A(n7272), .ZN(
        n7276) );
  OAI21_X1 U8992 ( .B1(n7276), .B2(n7275), .A(n7333), .ZN(n7277) );
  INV_X1 U8993 ( .A(n9879), .ZN(n9582) );
  NAND2_X1 U8994 ( .A1(n7277), .A2(n9582), .ZN(n7282) );
  NOR2_X1 U8995 ( .A1(n7278), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8013) );
  NOR2_X1 U8996 ( .A1(n9578), .A2(n7279), .ZN(n7280) );
  AOI211_X1 U8997 ( .C1(n9878), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n8013), .B(
        n7280), .ZN(n7281) );
  OAI211_X1 U8998 ( .C1(n7283), .C2(n9579), .A(n7282), .B(n7281), .ZN(P1_U3252) );
  AOI21_X1 U8999 ( .B1(n7285), .B2(n7284), .A(n9174), .ZN(n7287) );
  NAND2_X1 U9000 ( .A1(n7287), .A2(n7286), .ZN(n7293) );
  NAND2_X1 U9001 ( .A1(n9450), .A2(n9152), .ZN(n7289) );
  NAND2_X1 U9002 ( .A1(n7463), .A2(n9604), .ZN(n7288) );
  AND2_X1 U9003 ( .A1(n7289), .A2(n7288), .ZN(n7611) );
  INV_X1 U9004 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n7290) );
  OAI22_X1 U9005 ( .A1(n9156), .A2(n7611), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7290), .ZN(n7291) );
  AOI21_X1 U9006 ( .B1(n7618), .B2(n9158), .A(n7291), .ZN(n7292) );
  OAI211_X1 U9007 ( .C1(n10021), .C2(n9161), .A(n7293), .B(n7292), .ZN(
        P1_U3230) );
  INV_X1 U9008 ( .A(n7294), .ZN(n7296) );
  OAI222_X1 U9009 ( .A1(n8549), .A2(n7295), .B1(n9024), .B2(n7296), .C1(
        P2_U3151), .C2(n8720), .ZN(P2_U3278) );
  INV_X1 U9010 ( .A(n9561), .ZN(n9547) );
  OAI222_X1 U9011 ( .A1(n4428), .A2(n7297), .B1(n9834), .B2(n7296), .C1(
        P1_U3086), .C2(n9547), .ZN(P1_U3338) );
  OAI21_X1 U9012 ( .B1(n7299), .B2(n8412), .A(n7298), .ZN(n7873) );
  XNOR2_X1 U9013 ( .A(n7301), .B(n7300), .ZN(n7302) );
  OAI222_X1 U9014 ( .A1(n10171), .A2(n7402), .B1(n5626), .B2(n7303), .C1(n5628), .C2(n7302), .ZN(n7870) );
  AOI21_X1 U9015 ( .B1(n10234), .B2(n7873), .A(n7870), .ZN(n7367) );
  AOI22_X1 U9016 ( .A1(n8937), .A2(n7395), .B1(n6692), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n7304) );
  OAI21_X1 U9017 ( .B1(n7367), .B2(n6692), .A(n7304), .ZN(P2_U3462) );
  INV_X1 U9018 ( .A(n7305), .ZN(n7317) );
  INV_X1 U9019 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7306) );
  OAI222_X1 U9020 ( .A1(n9024), .A2(n7317), .B1(n7307), .B2(P2_U3151), .C1(
        n7306), .C2(n8549), .ZN(P2_U3279) );
  INV_X1 U9021 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7311) );
  NAND2_X1 U9022 ( .A1(n8671), .A2(n7309), .ZN(n8253) );
  NAND2_X1 U9023 ( .A1(n8250), .A2(n8253), .ZN(n8409) );
  OAI21_X1 U9024 ( .B1(n8894), .B2(n10234), .A(n8409), .ZN(n7308) );
  NAND2_X1 U9025 ( .A1(n5135), .A2(n8889), .ZN(n7579) );
  OAI211_X1 U9026 ( .C1(n10226), .C2(n7309), .A(n7308), .B(n7579), .ZN(n8945)
         );
  NAND2_X1 U9027 ( .A1(n8945), .A2(n10238), .ZN(n7310) );
  OAI21_X1 U9028 ( .B1(n7311), .B2(n10238), .A(n7310), .ZN(P2_U3390) );
  INV_X1 U9029 ( .A(n7312), .ZN(n7314) );
  OAI222_X1 U9030 ( .A1(n8549), .A2(n7313), .B1(n9024), .B2(n7314), .C1(
        P2_U3151), .C2(n6599), .ZN(P2_U3280) );
  OAI222_X1 U9031 ( .A1(n4428), .A2(n7315), .B1(n9834), .B2(n7314), .C1(
        P1_U3086), .C2(n4609), .ZN(P1_U3340) );
  INV_X1 U9032 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7316) );
  OAI222_X1 U9033 ( .A1(P1_U3086), .A2(n9537), .B1(n9834), .B2(n7317), .C1(
        n7316), .C2(n4428), .ZN(P1_U3339) );
  INV_X1 U9034 ( .A(n7318), .ZN(n7330) );
  AOI22_X1 U9035 ( .A1(n9575), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9832), .ZN(n7319) );
  OAI21_X1 U9036 ( .B1(n7330), .B2(n9834), .A(n7319), .ZN(P1_U3337) );
  INV_X1 U9037 ( .A(n7320), .ZN(n7321) );
  AOI21_X1 U9038 ( .B1(n7323), .B2(n7322), .A(n7321), .ZN(n7329) );
  INV_X1 U9039 ( .A(n8648), .ZN(n8592) );
  OAI21_X1 U9040 ( .B1(n10170), .B2(n8635), .A(n7324), .ZN(n7325) );
  AOI21_X1 U9041 ( .B1(n8632), .B2(n8667), .A(n7325), .ZN(n7326) );
  OAI21_X1 U9042 ( .B1(n10189), .B2(n8592), .A(n7326), .ZN(n7327) );
  AOI21_X1 U9043 ( .B1(n7726), .B2(n8641), .A(n7327), .ZN(n7328) );
  OAI21_X1 U9044 ( .B1(n7329), .B2(n8650), .A(n7328), .ZN(P2_U3170) );
  OAI222_X1 U9045 ( .A1(n8549), .A2(n7332), .B1(n7331), .B2(P2_U3151), .C1(
        n9024), .C2(n7330), .ZN(P2_U3277) );
  OAI21_X1 U9046 ( .B1(n7337), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7333), .ZN(
        n7336) );
  NAND2_X1 U9047 ( .A1(n7565), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7334) );
  OAI21_X1 U9048 ( .B1(n7565), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7334), .ZN(
        n7335) );
  NOR2_X1 U9049 ( .A1(n7335), .A2(n7336), .ZN(n7564) );
  AOI211_X1 U9050 ( .C1(n7336), .C2(n7335), .A(n7564), .B(n9879), .ZN(n7348)
         );
  NOR2_X1 U9051 ( .A1(n7337), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7339) );
  NOR2_X1 U9052 ( .A1(n7339), .A2(n7338), .ZN(n7342) );
  INV_X1 U9053 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7340) );
  MUX2_X1 U9054 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n7340), .S(n7565), .Z(n7341)
         );
  NAND2_X1 U9055 ( .A1(n7341), .A2(n7342), .ZN(n7559) );
  OAI211_X1 U9056 ( .C1(n7342), .C2(n7341), .A(n9888), .B(n7559), .ZN(n7345)
         );
  AND2_X1 U9057 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7343) );
  AOI21_X1 U9058 ( .B1(n9878), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n7343), .ZN(
        n7344) );
  OAI211_X1 U9059 ( .C1(n9578), .C2(n7346), .A(n7345), .B(n7344), .ZN(n7347)
         );
  OR2_X1 U9060 ( .A1(n7348), .A2(n7347), .ZN(P1_U3253) );
  INV_X1 U9061 ( .A(n8409), .ZN(n7578) );
  INV_X1 U9062 ( .A(n8641), .ZN(n8558) );
  NAND2_X1 U9063 ( .A1(n8558), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7361) );
  NAND2_X1 U9064 ( .A1(n7361), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7350) );
  AOI22_X1 U9065 ( .A1(n8632), .A2(n5135), .B1(n8648), .B2(n7582), .ZN(n7349)
         );
  OAI211_X1 U9066 ( .C1(n7578), .C2(n8650), .A(n7350), .B(n7349), .ZN(P2_U3172) );
  XOR2_X1 U9067 ( .A(n7351), .B(n7352), .Z(n7356) );
  AOI22_X1 U9068 ( .A1(n8640), .A2(n8671), .B1(n8632), .B2(n8670), .ZN(n7353)
         );
  OAI21_X1 U9069 ( .B1(n8592), .B2(n5136), .A(n7353), .ZN(n7354) );
  AOI21_X1 U9070 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n7361), .A(n7354), .ZN(
        n7355) );
  OAI21_X1 U9071 ( .B1(n7356), .B2(n8650), .A(n7355), .ZN(P2_U3162) );
  XOR2_X1 U9072 ( .A(n7358), .B(n7357), .Z(n7363) );
  AOI22_X1 U9073 ( .A1(n8640), .A2(n5135), .B1(n8632), .B2(n8669), .ZN(n7359)
         );
  OAI21_X1 U9074 ( .B1(n10182), .B2(n8592), .A(n7359), .ZN(n7360) );
  AOI21_X1 U9075 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n7361), .A(n7360), .ZN(
        n7362) );
  OAI21_X1 U9076 ( .B1(n7363), .B2(n8650), .A(n7362), .ZN(P2_U3177) );
  INV_X1 U9077 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7364) );
  OAI22_X1 U9078 ( .A1(n8989), .A2(n7869), .B1(n7364), .B2(n10238), .ZN(n7365)
         );
  INV_X1 U9079 ( .A(n7365), .ZN(n7366) );
  OAI21_X1 U9080 ( .B1(n7367), .B2(n10240), .A(n7366), .ZN(P2_U3399) );
  NAND2_X1 U9081 ( .A1(n7369), .A2(n7368), .ZN(n7371) );
  XNOR2_X1 U9082 ( .A(n7371), .B(n7370), .ZN(n7376) );
  AOI22_X1 U9083 ( .A1(n9604), .A2(n9451), .B1(n9449), .B2(n9152), .ZN(n9943)
         );
  OAI22_X1 U9084 ( .A1(n9943), .A2(n9156), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7372), .ZN(n7374) );
  INV_X1 U9085 ( .A(n9948), .ZN(n10028) );
  NOR2_X1 U9086 ( .A1(n9161), .A2(n10028), .ZN(n7373) );
  AOI211_X1 U9087 ( .C1(n9158), .C2(n9946), .A(n7374), .B(n7373), .ZN(n7375)
         );
  OAI21_X1 U9088 ( .B1(n7376), .B2(n9174), .A(n7375), .ZN(P1_U3227) );
  XNOR2_X1 U9089 ( .A(n7377), .B(n8408), .ZN(n7382) );
  INV_X1 U9090 ( .A(n7378), .ZN(n7379) );
  AOI21_X1 U9091 ( .B1(n8250), .B2(n8408), .A(n7379), .ZN(n10178) );
  AOI22_X1 U9092 ( .A1(n8891), .A2(n8671), .B1(n8670), .B2(n8889), .ZN(n7380)
         );
  OAI21_X1 U9093 ( .B1(n10178), .B2(n7777), .A(n7380), .ZN(n7381) );
  AOI21_X1 U9094 ( .B1(n8894), .B2(n7382), .A(n7381), .ZN(n10177) );
  INV_X1 U9095 ( .A(n10178), .ZN(n7383) );
  AOI22_X1 U9096 ( .A1(n7383), .A2(n7626), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8897), .ZN(n7384) );
  AOI21_X1 U9097 ( .B1(n10177), .B2(n7384), .A(n10176), .ZN(n7387) );
  OAI22_X1 U9098 ( .A1(n8839), .A2(n5136), .B1(n8895), .B2(n7385), .ZN(n7386)
         );
  OR2_X1 U9099 ( .A1(n7387), .A2(n7386), .ZN(P2_U3232) );
  OAI211_X1 U9100 ( .C1(n7390), .C2(n7389), .A(n7388), .B(n8616), .ZN(n7397)
         );
  NAND2_X1 U9101 ( .A1(n8640), .A2(n8670), .ZN(n7392) );
  OAI211_X1 U9102 ( .C1(n7402), .C2(n8645), .A(n7392), .B(n7391), .ZN(n7394)
         );
  NOR2_X1 U9103 ( .A1(n8558), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7393) );
  AOI211_X1 U9104 ( .C1(n7395), .C2(n8648), .A(n7394), .B(n7393), .ZN(n7396)
         );
  NAND2_X1 U9105 ( .A1(n7397), .A2(n7396), .ZN(P2_U3158) );
  XOR2_X1 U9106 ( .A(n7399), .B(n7398), .Z(n7407) );
  NAND2_X1 U9107 ( .A1(n8632), .A2(n8666), .ZN(n7401) );
  AND2_X1 U9108 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8482) );
  INV_X1 U9109 ( .A(n8482), .ZN(n7400) );
  OAI211_X1 U9110 ( .C1(n7402), .C2(n8635), .A(n7401), .B(n7400), .ZN(n7405)
         );
  INV_X1 U9111 ( .A(n7759), .ZN(n7403) );
  NOR2_X1 U9112 ( .A1(n8558), .A2(n7403), .ZN(n7404) );
  AOI211_X1 U9113 ( .C1(n7760), .C2(n8648), .A(n7405), .B(n7404), .ZN(n7406)
         );
  OAI21_X1 U9114 ( .B1(n7407), .B2(n8650), .A(n7406), .ZN(P2_U3167) );
  INV_X1 U9115 ( .A(n7408), .ZN(n8471) );
  OAI222_X1 U9116 ( .A1(n8549), .A2(n7410), .B1(n9024), .B2(n8471), .C1(
        P2_U3151), .C2(n7409), .ZN(P2_U3276) );
  AOI21_X1 U9117 ( .B1(n7412), .B2(n7411), .A(n8650), .ZN(n7413) );
  OR2_X1 U9118 ( .A1(n7412), .A2(n7411), .ZN(n7504) );
  NAND2_X1 U9119 ( .A1(n7413), .A2(n7504), .ZN(n7420) );
  NAND2_X1 U9120 ( .A1(n8640), .A2(n8667), .ZN(n7415) );
  OAI211_X1 U9121 ( .C1(n7416), .C2(n8645), .A(n7415), .B(n7414), .ZN(n7418)
         );
  NOR2_X1 U9122 ( .A1(n8592), .A2(n10198), .ZN(n7417) );
  AOI211_X1 U9123 ( .C1(n7745), .C2(n8641), .A(n7418), .B(n7417), .ZN(n7419)
         );
  NAND2_X1 U9124 ( .A1(n7420), .A2(n7419), .ZN(P2_U3179) );
  XNOR2_X1 U9125 ( .A(n7422), .B(n7421), .ZN(n7423) );
  XNOR2_X1 U9126 ( .A(n7424), .B(n7423), .ZN(n7431) );
  INV_X1 U9127 ( .A(n10035), .ZN(n7605) );
  NAND2_X1 U9128 ( .A1(n9450), .A2(n9604), .ZN(n7426) );
  NAND2_X1 U9129 ( .A1(n9448), .A2(n9152), .ZN(n7425) );
  NAND2_X1 U9130 ( .A1(n7426), .A2(n7425), .ZN(n7600) );
  AOI22_X1 U9131 ( .A1(n9165), .A2(n7600), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3086), .ZN(n7427) );
  OAI21_X1 U9132 ( .B1(n7428), .B2(n9168), .A(n7427), .ZN(n7429) );
  AOI21_X1 U9133 ( .B1(n7605), .B2(n9171), .A(n7429), .ZN(n7430) );
  OAI21_X1 U9134 ( .B1(n7431), .B2(n9174), .A(n7430), .ZN(P1_U3239) );
  INV_X1 U9135 ( .A(n7432), .ZN(n7539) );
  OAI222_X1 U9136 ( .A1(n9024), .A2(n7539), .B1(n5754), .B2(P2_U3151), .C1(
        n7433), .C2(n8549), .ZN(P2_U3275) );
  INV_X1 U9137 ( .A(n7434), .ZN(n7437) );
  NOR2_X1 U9138 ( .A1(n9829), .A2(n7435), .ZN(n7436) );
  NAND2_X1 U9139 ( .A1(n7437), .A2(n7436), .ZN(n7438) );
  INV_X2 U9140 ( .A(n9744), .ZN(n9992) );
  INV_X1 U9141 ( .A(n9976), .ZN(n9973) );
  NOR2_X1 U9142 ( .A1(n7114), .A2(n9986), .ZN(n9972) );
  NAND2_X1 U9143 ( .A1(n9973), .A2(n9972), .ZN(n9971) );
  NAND2_X1 U9144 ( .A1(n7456), .A2(n9982), .ZN(n7441) );
  NAND2_X1 U9145 ( .A1(n9971), .A2(n7441), .ZN(n7593) );
  NAND2_X1 U9146 ( .A1(n7445), .A2(n9364), .ZN(n7459) );
  INV_X1 U9147 ( .A(n7459), .ZN(n9297) );
  NAND2_X1 U9148 ( .A1(n7463), .A2(n10015), .ZN(n9366) );
  INV_X1 U9149 ( .A(n7463), .ZN(n7464) );
  NAND2_X1 U9150 ( .A1(n7464), .A2(n9960), .ZN(n7446) );
  NAND2_X1 U9151 ( .A1(n7467), .A2(n7617), .ZN(n9185) );
  INV_X1 U9152 ( .A(n9450), .ZN(n7470) );
  NAND2_X1 U9153 ( .A1(n7470), .A2(n9948), .ZN(n9184) );
  INV_X1 U9154 ( .A(n9184), .ZN(n9192) );
  NAND2_X1 U9155 ( .A1(n9450), .A2(n10028), .ZN(n9365) );
  INV_X1 U9156 ( .A(n9449), .ZN(n7473) );
  NAND2_X1 U9157 ( .A1(n7473), .A2(n7605), .ZN(n9194) );
  NAND2_X1 U9158 ( .A1(n7599), .A2(n9194), .ZN(n7496) );
  INV_X1 U9159 ( .A(n9446), .ZN(n7448) );
  NOR2_X1 U9160 ( .A1(n10058), .A2(n7448), .ZN(n7476) );
  INV_X1 U9161 ( .A(n7476), .ZN(n9204) );
  INV_X1 U9162 ( .A(n9447), .ZN(n7475) );
  OR2_X1 U9163 ( .A1(n7866), .A2(n7475), .ZN(n9198) );
  NAND2_X1 U9164 ( .A1(n9204), .A2(n9198), .ZN(n9190) );
  NAND2_X1 U9165 ( .A1(n7866), .A2(n7475), .ZN(n9180) );
  INV_X1 U9166 ( .A(n10042), .ZN(n9934) );
  AND2_X1 U9167 ( .A1(n9934), .A2(n7447), .ZN(n7474) );
  INV_X1 U9168 ( .A(n7474), .ZN(n9195) );
  AND2_X1 U9169 ( .A1(n9180), .A2(n9195), .ZN(n9188) );
  AND2_X1 U9170 ( .A1(n10058), .A2(n7448), .ZN(n9182) );
  INV_X1 U9171 ( .A(n9182), .ZN(n9200) );
  AND2_X1 U9172 ( .A1(n10042), .A2(n9448), .ZN(n9197) );
  NAND2_X1 U9173 ( .A1(n10035), .A2(n9449), .ZN(n9186) );
  NAND2_X1 U9174 ( .A1(n9371), .A2(n9369), .ZN(n7451) );
  INV_X1 U9175 ( .A(n9445), .ZN(n8069) );
  OR2_X1 U9176 ( .A1(n7480), .A2(n8069), .ZN(n9208) );
  NAND2_X1 U9177 ( .A1(n7480), .A2(n8069), .ZN(n9206) );
  NAND2_X1 U9178 ( .A1(n9208), .A2(n9206), .ZN(n7643) );
  XNOR2_X1 U9179 ( .A(n7451), .B(n7643), .ZN(n7455) );
  NAND2_X1 U9180 ( .A1(n9446), .A2(n9604), .ZN(n7453) );
  NAND2_X1 U9181 ( .A1(n9444), .A2(n9152), .ZN(n7452) );
  AND2_X1 U9182 ( .A1(n7453), .A2(n7452), .ZN(n7967) );
  INV_X1 U9183 ( .A(n7967), .ZN(n7454) );
  AOI21_X1 U9184 ( .B1(n7455), .B2(n9980), .A(n7454), .ZN(n10067) );
  INV_X1 U9185 ( .A(n7440), .ZN(n7456) );
  NAND2_X1 U9186 ( .A1(n7456), .A2(n7439), .ZN(n7457) );
  NAND2_X1 U9187 ( .A1(n7458), .A2(n7457), .ZN(n7587) );
  NAND2_X1 U9188 ( .A1(n7587), .A2(n7459), .ZN(n7462) );
  NAND2_X1 U9189 ( .A1(n7443), .A2(n7460), .ZN(n7461) );
  NAND2_X1 U9190 ( .A1(n7462), .A2(n7461), .ZN(n9962) );
  NAND2_X1 U9191 ( .A1(n9962), .A2(n9963), .ZN(n7466) );
  NAND2_X1 U9192 ( .A1(n7464), .A2(n10015), .ZN(n7465) );
  NAND2_X1 U9193 ( .A1(n7466), .A2(n7465), .ZN(n7614) );
  NAND2_X1 U9194 ( .A1(n9185), .A2(n9367), .ZN(n7615) );
  NAND2_X1 U9195 ( .A1(n7614), .A2(n7615), .ZN(n7469) );
  NAND2_X1 U9196 ( .A1(n7467), .A2(n10021), .ZN(n7468) );
  NAND2_X1 U9197 ( .A1(n7469), .A2(n7468), .ZN(n9949) );
  NAND2_X1 U9198 ( .A1(n9949), .A2(n9950), .ZN(n7472) );
  NAND2_X1 U9199 ( .A1(n7470), .A2(n10028), .ZN(n7471) );
  NAND2_X1 U9200 ( .A1(n9186), .A2(n9194), .ZN(n9299) );
  NOR2_X1 U9201 ( .A1(n9197), .A2(n7474), .ZN(n9928) );
  NAND2_X1 U9202 ( .A1(n9198), .A2(n9180), .ZN(n7676) );
  INV_X1 U9203 ( .A(n7866), .ZN(n10052) );
  NOR2_X1 U9204 ( .A1(n7476), .A2(n9182), .ZN(n7497) );
  XNOR2_X1 U9205 ( .A(n7641), .B(n7643), .ZN(n10070) );
  OR2_X1 U9206 ( .A1(n7477), .A2(n6284), .ZN(n7478) );
  OR2_X1 U9207 ( .A1(n9992), .A2(n7478), .ZN(n9988) );
  OR2_X1 U9208 ( .A1(n9992), .A2(n10048), .ZN(n7479) );
  NAND2_X1 U9209 ( .A1(n9988), .A2(n7479), .ZN(n9968) );
  NAND2_X1 U9210 ( .A1(n10070), .A2(n9968), .ZN(n7488) );
  NAND2_X1 U9211 ( .A1(n9965), .A2(n10015), .ZN(n9964) );
  INV_X1 U9212 ( .A(n9921), .ZN(n7482) );
  OR2_X1 U9213 ( .A1(n7481), .A2(n9410), .ZN(n9737) );
  INV_X1 U9214 ( .A(n9737), .ZN(n9985) );
  OAI211_X1 U9215 ( .C1(n10068), .C2(n7491), .A(n7482), .B(n9985), .ZN(n10066)
         );
  INV_X1 U9216 ( .A(n10066), .ZN(n7486) );
  OR2_X1 U9217 ( .A1(n9992), .A2(n9584), .ZN(n9987) );
  INV_X1 U9218 ( .A(n9744), .ZN(n9947) );
  INV_X1 U9219 ( .A(n8523), .ZN(n9983) );
  AOI22_X1 U9220 ( .A1(n9947), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7970), .B2(
        n9983), .ZN(n7484) );
  OAI21_X1 U9221 ( .B1(n10068), .B2(n9741), .A(n7484), .ZN(n7485) );
  AOI21_X1 U9222 ( .B1(n7486), .B2(n9967), .A(n7485), .ZN(n7487) );
  OAI211_X1 U9223 ( .C1(n9992), .C2(n10067), .A(n7488), .B(n7487), .ZN(
        P1_U3283) );
  XOR2_X1 U9224 ( .A(n7489), .B(n7497), .Z(n10062) );
  INV_X1 U9225 ( .A(n7682), .ZN(n7490) );
  INV_X1 U9226 ( .A(n10058), .ZN(n7494) );
  OAI21_X1 U9227 ( .B1(n7490), .B2(n7494), .A(n9985), .ZN(n7492) );
  NAND2_X1 U9228 ( .A1(n9445), .A2(n9152), .ZN(n8011) );
  OAI21_X1 U9229 ( .B1(n7492), .B2(n7491), .A(n8011), .ZN(n10057) );
  AOI22_X1 U9230 ( .A1(n9992), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n8014), .B2(
        n9983), .ZN(n7493) );
  OAI21_X1 U9231 ( .B1(n7494), .B2(n9741), .A(n7493), .ZN(n7495) );
  AOI21_X1 U9232 ( .B1(n10057), .B2(n9967), .A(n7495), .ZN(n7501) );
  AND2_X1 U9233 ( .A1(n7496), .A2(n9186), .ZN(n9926) );
  NAND2_X1 U9234 ( .A1(n9926), .A2(n4427), .ZN(n9925) );
  NAND2_X1 U9235 ( .A1(n9925), .A2(n9188), .ZN(n7675) );
  NAND2_X1 U9236 ( .A1(n7675), .A2(n9198), .ZN(n7498) );
  XNOR2_X1 U9237 ( .A(n7498), .B(n7497), .ZN(n7499) );
  INV_X1 U9238 ( .A(n9980), .ZN(n9913) );
  NAND2_X1 U9239 ( .A1(n9447), .A2(n9604), .ZN(n8010) );
  OAI21_X1 U9240 ( .B1(n7499), .B2(n9913), .A(n8010), .ZN(n10063) );
  NAND2_X1 U9241 ( .A1(n10063), .A2(n9744), .ZN(n7500) );
  OAI211_X1 U9242 ( .C1(n10062), .C2(n9746), .A(n7501), .B(n7500), .ZN(
        P1_U3284) );
  AND2_X1 U9243 ( .A1(n7504), .A2(n7502), .ZN(n7507) );
  NAND2_X1 U9244 ( .A1(n7504), .A2(n7503), .ZN(n7505) );
  OAI21_X1 U9245 ( .B1(n7507), .B2(n7506), .A(n7505), .ZN(n7515) );
  INV_X1 U9246 ( .A(n7508), .ZN(n7509) );
  AOI21_X1 U9247 ( .B1(n8640), .B2(n8666), .A(n7509), .ZN(n7513) );
  NAND2_X1 U9248 ( .A1(n8641), .A2(n7636), .ZN(n7512) );
  NAND2_X1 U9249 ( .A1(n8648), .A2(n7637), .ZN(n7511) );
  NAND2_X1 U9250 ( .A1(n8632), .A2(n8664), .ZN(n7510) );
  NAND4_X1 U9251 ( .A1(n7513), .A2(n7512), .A3(n7511), .A4(n7510), .ZN(n7514)
         );
  AOI21_X1 U9252 ( .B1(n7515), .B2(n8616), .A(n7514), .ZN(n7516) );
  INV_X1 U9253 ( .A(n7516), .ZN(P2_U3153) );
  NAND2_X1 U9254 ( .A1(n5178), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n7519) );
  NAND2_X1 U9255 ( .A1(n5155), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7518) );
  NAND2_X1 U9256 ( .A1(n5177), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n7517) );
  AND3_X1 U9257 ( .A1(n7519), .A2(n7518), .A3(n7517), .ZN(n7520) );
  NAND2_X1 U9258 ( .A1(n7521), .A2(n7520), .ZN(n8748) );
  NAND2_X1 U9259 ( .A1(n8748), .A2(P2_U3893), .ZN(n7522) );
  OAI21_X1 U9260 ( .B1(P2_U3893), .B2(n7523), .A(n7522), .ZN(P2_U3522) );
  AOI21_X1 U9261 ( .B1(n10254), .B2(n7525), .A(n7524), .ZN(n7537) );
  OAI21_X1 U9262 ( .B1(n7528), .B2(n7527), .A(n7526), .ZN(n7535) );
  AND2_X1 U9263 ( .A1(n10141), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7534) );
  AND2_X1 U9264 ( .A1(n7530), .A2(n7785), .ZN(n7531) );
  OAI21_X1 U9265 ( .B1(n7529), .B2(n7531), .A(n8741), .ZN(n7532) );
  NAND2_X1 U9266 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7770) );
  OAI211_X1 U9267 ( .C1(n10162), .C2(n6582), .A(n7532), .B(n7770), .ZN(n7533)
         );
  AOI211_X1 U9268 ( .C1(n10152), .C2(n7535), .A(n7534), .B(n7533), .ZN(n7536)
         );
  OAI21_X1 U9269 ( .B1(n7537), .B2(n10147), .A(n7536), .ZN(P2_U3191) );
  OAI222_X1 U9270 ( .A1(n9321), .A2(P1_U3086), .B1(n9834), .B2(n7539), .C1(
        n7538), .C2(n4428), .ZN(P1_U3335) );
  NOR2_X1 U9271 ( .A1(n4514), .A2(n7540), .ZN(n7541) );
  XNOR2_X1 U9272 ( .A(n7542), .B(n7541), .ZN(n7549) );
  NAND2_X1 U9273 ( .A1(n9449), .A2(n9604), .ZN(n7544) );
  NAND2_X1 U9274 ( .A1(n9447), .A2(n9152), .ZN(n7543) );
  AND2_X1 U9275 ( .A1(n7544), .A2(n7543), .ZN(n9927) );
  OAI22_X1 U9276 ( .A1(n9156), .A2(n9927), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7545), .ZN(n7547) );
  NOR2_X1 U9277 ( .A1(n9161), .A2(n10042), .ZN(n7546) );
  AOI211_X1 U9278 ( .C1(n9158), .C2(n9933), .A(n7547), .B(n7546), .ZN(n7548)
         );
  OAI21_X1 U9279 ( .B1(n7549), .B2(n9174), .A(n7548), .ZN(P1_U3213) );
  NOR2_X1 U9280 ( .A1(n9987), .A2(n9737), .ZN(n9715) );
  OAI21_X1 U9281 ( .B1(n9715), .B2(n9981), .A(n7550), .ZN(n7558) );
  INV_X1 U9282 ( .A(n7551), .ZN(n9412) );
  NOR3_X1 U9283 ( .A1(n9295), .A2(n9412), .A3(n7552), .ZN(n7556) );
  OAI21_X1 U9284 ( .B1(n8523), .B2(n7554), .A(n7553), .ZN(n7555) );
  OAI21_X1 U9285 ( .B1(n7556), .B2(n7555), .A(n9744), .ZN(n7557) );
  OAI211_X1 U9286 ( .C1(n5940), .C2(n9744), .A(n7558), .B(n7557), .ZN(P1_U3293) );
  NAND2_X1 U9287 ( .A1(n7565), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7560) );
  NAND2_X1 U9288 ( .A1(n7560), .A2(n7559), .ZN(n7563) );
  INV_X1 U9289 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7561) );
  MUX2_X1 U9290 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n7561), .S(n7666), .Z(n7562)
         );
  NAND2_X1 U9291 ( .A1(n7562), .A2(n7563), .ZN(n7659) );
  OAI211_X1 U9292 ( .C1(n7563), .C2(n7562), .A(n9888), .B(n7659), .ZN(n7575)
         );
  NAND2_X1 U9293 ( .A1(n7666), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7566) );
  OAI21_X1 U9294 ( .B1(n7666), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7566), .ZN(
        n7567) );
  AOI211_X1 U9295 ( .C1(n7568), .C2(n7567), .A(n7665), .B(n9879), .ZN(n7573)
         );
  INV_X1 U9296 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7569) );
  NOR2_X1 U9297 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7569), .ZN(n7570) );
  AOI21_X1 U9298 ( .B1(n9878), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n7570), .ZN(
        n7571) );
  OAI21_X1 U9299 ( .B1(n7660), .B2(n9578), .A(n7571), .ZN(n7572) );
  NOR2_X1 U9300 ( .A1(n7573), .A2(n7572), .ZN(n7574) );
  NAND2_X1 U9301 ( .A1(n7575), .A2(n7574), .ZN(P1_U3254) );
  INV_X1 U9302 ( .A(n7576), .ZN(n7577) );
  NOR3_X1 U9303 ( .A1(n7578), .A2(n7577), .A3(n10233), .ZN(n7581) );
  INV_X1 U9304 ( .A(n7579), .ZN(n7580) );
  OAI21_X1 U9305 ( .B1(n7581), .B2(n7580), .A(n10174), .ZN(n7584) );
  AOI22_X1 U9306 ( .A1(n8898), .A2(n7582), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n8897), .ZN(n7583) );
  OAI211_X1 U9307 ( .C1(n6565), .C2(n10174), .A(n7584), .B(n7583), .ZN(
        P2_U3233) );
  INV_X1 U9308 ( .A(n7585), .ZN(n8552) );
  OAI222_X1 U9309 ( .A1(n4428), .A2(n7586), .B1(n8472), .B2(n8552), .C1(n9294), 
        .C2(P1_U3086), .ZN(P1_U3334) );
  XNOR2_X1 U9310 ( .A(n7459), .B(n7587), .ZN(n10010) );
  INV_X1 U9311 ( .A(n9965), .ZN(n7589) );
  AOI21_X1 U9312 ( .B1(n9984), .B2(n7442), .A(n9737), .ZN(n7588) );
  NAND2_X1 U9313 ( .A1(n7589), .A2(n7588), .ZN(n10009) );
  NAND2_X1 U9314 ( .A1(n9981), .A2(n7442), .ZN(n7591) );
  AOI22_X1 U9315 ( .A1(n9947), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9983), .ZN(n7590) );
  OAI211_X1 U9316 ( .C1(n10009), .C2(n9987), .A(n7591), .B(n7590), .ZN(n7597)
         );
  OAI21_X1 U9317 ( .B1(n9297), .B2(n7593), .A(n7592), .ZN(n7595) );
  AOI21_X1 U9318 ( .B1(n7595), .B2(n9980), .A(n7594), .ZN(n10013) );
  NOR2_X1 U9319 ( .A1(n10013), .A2(n9947), .ZN(n7596) );
  AOI211_X1 U9320 ( .C1(n9968), .C2(n10010), .A(n7597), .B(n7596), .ZN(n7598)
         );
  INV_X1 U9321 ( .A(n7598), .ZN(P1_U3291) );
  XNOR2_X1 U9322 ( .A(n7599), .B(n9299), .ZN(n7601) );
  AOI21_X1 U9323 ( .B1(n7601), .B2(n9980), .A(n7600), .ZN(n10039) );
  XNOR2_X1 U9324 ( .A(n7602), .B(n9299), .ZN(n10037) );
  OAI21_X1 U9325 ( .B1(n9952), .B2(n10035), .A(n9985), .ZN(n7603) );
  OR2_X1 U9326 ( .A1(n7603), .A2(n9937), .ZN(n10034) );
  AOI22_X1 U9327 ( .A1(n9992), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7604), .B2(
        n9983), .ZN(n7607) );
  NAND2_X1 U9328 ( .A1(n9981), .A2(n7605), .ZN(n7606) );
  OAI211_X1 U9329 ( .C1(n10034), .C2(n9987), .A(n7607), .B(n7606), .ZN(n7608)
         );
  AOI21_X1 U9330 ( .B1(n10037), .B2(n9968), .A(n7608), .ZN(n7609) );
  OAI21_X1 U9331 ( .B1(n10039), .B2(n9947), .A(n7609), .ZN(P1_U3287) );
  INV_X1 U9332 ( .A(n7615), .ZN(n9298) );
  XNOR2_X1 U9333 ( .A(n7610), .B(n9298), .ZN(n7613) );
  INV_X1 U9334 ( .A(n7611), .ZN(n7612) );
  AOI21_X1 U9335 ( .B1(n7613), .B2(n9980), .A(n7612), .ZN(n10025) );
  XNOR2_X1 U9336 ( .A(n7615), .B(n7614), .ZN(n10023) );
  AOI21_X1 U9337 ( .B1(n9964), .B2(n7617), .A(n9737), .ZN(n7616) );
  NAND2_X1 U9338 ( .A1(n7616), .A2(n9951), .ZN(n10020) );
  NAND2_X1 U9339 ( .A1(n9981), .A2(n7617), .ZN(n7620) );
  AOI22_X1 U9340 ( .A1(n9947), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7618), .B2(
        n9983), .ZN(n7619) );
  OAI211_X1 U9341 ( .C1(n10020), .C2(n9987), .A(n7620), .B(n7619), .ZN(n7621)
         );
  AOI21_X1 U9342 ( .B1(n10023), .B2(n9968), .A(n7621), .ZN(n7622) );
  OAI21_X1 U9343 ( .B1(n10025), .B2(n9947), .A(n7622), .ZN(P1_U3289) );
  NAND2_X1 U9344 ( .A1(n7742), .A2(n8277), .ZN(n7623) );
  NAND2_X1 U9345 ( .A1(n7623), .A2(n8416), .ZN(n7625) );
  NAND2_X1 U9346 ( .A1(n7625), .A2(n7624), .ZN(n10206) );
  NAND2_X1 U9347 ( .A1(n10174), .A2(n7626), .ZN(n8760) );
  OR2_X1 U9348 ( .A1(n10206), .A2(n7777), .ZN(n7634) );
  NAND2_X1 U9349 ( .A1(n7627), .A2(n8285), .ZN(n7628) );
  NAND2_X1 U9350 ( .A1(n7733), .A2(n7628), .ZN(n7632) );
  NAND2_X1 U9351 ( .A1(n8666), .A2(n8891), .ZN(n7630) );
  NAND2_X1 U9352 ( .A1(n8664), .A2(n8889), .ZN(n7629) );
  NAND2_X1 U9353 ( .A1(n7630), .A2(n7629), .ZN(n7631) );
  AOI21_X1 U9354 ( .B1(n7632), .B2(n8894), .A(n7631), .ZN(n7633) );
  NAND2_X1 U9355 ( .A1(n7634), .A2(n7633), .ZN(n10208) );
  MUX2_X1 U9356 ( .A(n10208), .B(P2_REG2_REG_7__SCAN_IN), .S(n10176), .Z(n7635) );
  INV_X1 U9357 ( .A(n7635), .ZN(n7639) );
  AOI22_X1 U9358 ( .A1(n8898), .A2(n7637), .B1(n8897), .B2(n7636), .ZN(n7638)
         );
  OAI211_X1 U9359 ( .C1(n10206), .C2(n8760), .A(n7639), .B(n7638), .ZN(
        P2_U3226) );
  INV_X1 U9360 ( .A(n9444), .ZN(n7642) );
  NAND2_X1 U9361 ( .A1(n9920), .A2(n7642), .ZN(n9210) );
  OAI22_X2 U9362 ( .A1(n9911), .A2(n9910), .B1(n9920), .B2(n9444), .ZN(n7877)
         );
  INV_X1 U9363 ( .A(n9443), .ZN(n8068) );
  NAND2_X1 U9364 ( .A1(n7947), .A2(n8068), .ZN(n9211) );
  NAND2_X1 U9365 ( .A1(n9894), .A2(n9211), .ZN(n7876) );
  XNOR2_X1 U9366 ( .A(n7877), .B(n7876), .ZN(n10084) );
  INV_X1 U9367 ( .A(n10084), .ZN(n7658) );
  INV_X1 U9368 ( .A(n7643), .ZN(n9302) );
  INV_X1 U9369 ( .A(n9910), .ZN(n9915) );
  NAND2_X1 U9370 ( .A1(n7645), .A2(n9209), .ZN(n7644) );
  INV_X1 U9371 ( .A(n7876), .ZN(n9304) );
  NAND2_X1 U9372 ( .A1(n7644), .A2(n9304), .ZN(n9895) );
  NAND3_X1 U9373 ( .A1(n7645), .A2(n9209), .A3(n7876), .ZN(n7646) );
  NAND3_X1 U9374 ( .A1(n9895), .A2(n9980), .A3(n7646), .ZN(n7650) );
  NAND2_X1 U9375 ( .A1(n9444), .A2(n9604), .ZN(n7648) );
  NAND2_X1 U9376 ( .A1(n9442), .A2(n9152), .ZN(n7647) );
  NAND2_X1 U9377 ( .A1(n7648), .A2(n7647), .ZN(n7942) );
  INV_X1 U9378 ( .A(n7942), .ZN(n7649) );
  NAND2_X1 U9379 ( .A1(n7650), .A2(n7649), .ZN(n10083) );
  INV_X1 U9380 ( .A(n9920), .ZN(n10073) );
  NAND2_X1 U9381 ( .A1(n9921), .A2(n10073), .ZN(n7651) );
  INV_X1 U9382 ( .A(n7651), .ZN(n7652) );
  INV_X1 U9383 ( .A(n7947), .ZN(n10081) );
  OAI211_X1 U9384 ( .C1(n7652), .C2(n10081), .A(n9985), .B(n9904), .ZN(n10080)
         );
  OAI22_X1 U9385 ( .A1(n9744), .A2(n7653), .B1(n7945), .B2(n8523), .ZN(n7654)
         );
  AOI21_X1 U9386 ( .B1(n7947), .B2(n9981), .A(n7654), .ZN(n7655) );
  OAI21_X1 U9387 ( .B1(n10080), .B2(n9987), .A(n7655), .ZN(n7656) );
  AOI21_X1 U9388 ( .B1(n10083), .B2(n9744), .A(n7656), .ZN(n7657) );
  OAI21_X1 U9389 ( .B1(n7658), .B2(n9746), .A(n7657), .ZN(P1_U3281) );
  OAI21_X1 U9390 ( .B1(n7561), .B2(n7660), .A(n7659), .ZN(n7663) );
  AOI22_X1 U9391 ( .A1(n7921), .A2(n6170), .B1(P1_REG1_REG_12__SCAN_IN), .B2(
        n7661), .ZN(n7662) );
  NOR2_X1 U9392 ( .A1(n7663), .A2(n7662), .ZN(n7923) );
  AOI21_X1 U9393 ( .B1(n7663), .B2(n7662), .A(n7923), .ZN(n7673) );
  NOR2_X1 U9394 ( .A1(n7921), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7664) );
  AOI21_X1 U9395 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7921), .A(n7664), .ZN(
        n7668) );
  OAI21_X1 U9396 ( .B1(n7668), .B2(n7667), .A(n7917), .ZN(n7669) );
  NAND2_X1 U9397 ( .A1(n7669), .A2(n9582), .ZN(n7672) );
  INV_X1 U9398 ( .A(n9578), .ZN(n9885) );
  NAND2_X1 U9399 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7944) );
  OAI21_X1 U9400 ( .B1(n9589), .B2(n7830), .A(n7944), .ZN(n7670) );
  AOI21_X1 U9401 ( .B1(n9885), .B2(n7921), .A(n7670), .ZN(n7671) );
  OAI211_X1 U9402 ( .C1(n7673), .C2(n9579), .A(n7672), .B(n7671), .ZN(P1_U3255) );
  XOR2_X1 U9403 ( .A(n7674), .B(n7676), .Z(n10049) );
  INV_X1 U9404 ( .A(n7675), .ZN(n7678) );
  AOI21_X1 U9405 ( .B1(n9925), .B2(n9195), .A(n4933), .ZN(n7677) );
  AOI211_X1 U9406 ( .C1(n7678), .C2(n9198), .A(n9913), .B(n7677), .ZN(n7681)
         );
  NAND2_X1 U9407 ( .A1(n9448), .A2(n9604), .ZN(n7680) );
  NAND2_X1 U9408 ( .A1(n9446), .A2(n9152), .ZN(n7679) );
  NAND2_X1 U9409 ( .A1(n7680), .A2(n7679), .ZN(n7862) );
  NOR2_X1 U9410 ( .A1(n7681), .A2(n7862), .ZN(n10051) );
  INV_X1 U9411 ( .A(n10051), .ZN(n7687) );
  AOI21_X1 U9412 ( .B1(n9936), .B2(n7866), .A(n9737), .ZN(n7683) );
  NAND2_X1 U9413 ( .A1(n7683), .A2(n7682), .ZN(n10050) );
  AOI22_X1 U9414 ( .A1(n9992), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7861), .B2(
        n9983), .ZN(n7685) );
  NAND2_X1 U9415 ( .A1(n9981), .A2(n7866), .ZN(n7684) );
  OAI211_X1 U9416 ( .C1(n10050), .C2(n9987), .A(n7685), .B(n7684), .ZN(n7686)
         );
  AOI21_X1 U9417 ( .B1(n7687), .B2(n9744), .A(n7686), .ZN(n7688) );
  OAI21_X1 U9418 ( .B1(n9746), .B2(n10049), .A(n7688), .ZN(P1_U3285) );
  XNOR2_X1 U9419 ( .A(n7765), .B(n7764), .ZN(n7766) );
  XNOR2_X1 U9420 ( .A(n7766), .B(n7689), .ZN(n7697) );
  NAND2_X1 U9421 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n10138) );
  INV_X1 U9422 ( .A(n10138), .ZN(n7690) );
  AOI21_X1 U9423 ( .B1(n8640), .B2(n8665), .A(n7690), .ZN(n7693) );
  NAND2_X1 U9424 ( .A1(n8641), .A2(n7737), .ZN(n7692) );
  NAND2_X1 U9425 ( .A1(n8632), .A2(n8663), .ZN(n7691) );
  NAND3_X1 U9426 ( .A1(n7693), .A2(n7692), .A3(n7691), .ZN(n7694) );
  AOI21_X1 U9427 ( .B1(n7695), .B2(n8648), .A(n7694), .ZN(n7696) );
  OAI21_X1 U9428 ( .B1(n7697), .B2(n8650), .A(n7696), .ZN(P2_U3161) );
  AOI21_X1 U9429 ( .B1(n4517), .B2(n7699), .A(n7698), .ZN(n7715) );
  OAI21_X1 U9430 ( .B1(n7702), .B2(n7701), .A(n7700), .ZN(n7713) );
  INV_X1 U9431 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7822) );
  INV_X1 U9432 ( .A(n10162), .ZN(n8699) );
  INV_X1 U9433 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7703) );
  NOR2_X1 U9434 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7703), .ZN(n7794) );
  AOI21_X1 U9435 ( .B1(n8699), .B2(n7704), .A(n7794), .ZN(n7705) );
  OAI21_X1 U9436 ( .B1(n8682), .B2(n7822), .A(n7705), .ZN(n7712) );
  AOI21_X1 U9437 ( .B1(n7709), .B2(n7708), .A(n7707), .ZN(n7710) );
  NOR2_X1 U9438 ( .A1(n7710), .A2(n10156), .ZN(n7711) );
  AOI211_X1 U9439 ( .C1(n10152), .C2(n7713), .A(n7712), .B(n7711), .ZN(n7714)
         );
  OAI21_X1 U9440 ( .B1(n7715), .B2(n10147), .A(n7714), .ZN(P2_U3192) );
  NAND2_X1 U9441 ( .A1(n8272), .A2(n8265), .ZN(n8410) );
  XNOR2_X1 U9442 ( .A(n7716), .B(n8410), .ZN(n10187) );
  INV_X1 U9443 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7725) );
  INV_X1 U9444 ( .A(n7717), .ZN(n7721) );
  OAI21_X1 U9445 ( .B1(n7718), .B2(n8410), .A(n8894), .ZN(n7719) );
  AOI21_X1 U9446 ( .B1(n7721), .B2(n7720), .A(n7719), .ZN(n7724) );
  OAI22_X1 U9447 ( .A1(n10170), .A2(n5626), .B1(n7722), .B2(n10171), .ZN(n7723) );
  NOR2_X1 U9448 ( .A1(n7724), .A2(n7723), .ZN(n10188) );
  MUX2_X1 U9449 ( .A(n7725), .B(n10188), .S(n8895), .Z(n7729) );
  AOI22_X1 U9450 ( .A1(n8898), .A2(n7727), .B1(n8897), .B2(n7726), .ZN(n7728)
         );
  OAI211_X1 U9451 ( .C1(n8901), .C2(n10187), .A(n7729), .B(n7728), .ZN(
        P2_U3229) );
  XNOR2_X1 U9452 ( .A(n7730), .B(n8415), .ZN(n10213) );
  INV_X1 U9453 ( .A(n10213), .ZN(n7741) );
  NAND2_X1 U9454 ( .A1(n7731), .A2(n8894), .ZN(n7736) );
  AOI21_X1 U9455 ( .B1(n7733), .B2(n7732), .A(n8415), .ZN(n7735) );
  AOI22_X1 U9456 ( .A1(n8889), .A2(n8663), .B1(n8665), .B2(n8891), .ZN(n7734)
         );
  OAI21_X1 U9457 ( .B1(n7736), .B2(n7735), .A(n7734), .ZN(n10211) );
  AOI22_X1 U9458 ( .A1(n10176), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n8897), .B2(
        n7737), .ZN(n7738) );
  OAI21_X1 U9459 ( .B1(n10210), .B2(n8839), .A(n7738), .ZN(n7739) );
  AOI21_X1 U9460 ( .B1(n10211), .B2(n8895), .A(n7739), .ZN(n7740) );
  OAI21_X1 U9461 ( .B1(n7741), .B2(n8901), .A(n7740), .ZN(P2_U3225) );
  INV_X1 U9462 ( .A(n7742), .ZN(n7743) );
  AOI21_X1 U9463 ( .B1(n8414), .B2(n7744), .A(n7743), .ZN(n10200) );
  AOI22_X1 U9464 ( .A1(n8898), .A2(n7746), .B1(n8897), .B2(n7745), .ZN(n7753)
         );
  XNOR2_X1 U9465 ( .A(n7747), .B(n4820), .ZN(n7748) );
  NAND2_X1 U9466 ( .A1(n7748), .A2(n8894), .ZN(n7750) );
  AOI22_X1 U9467 ( .A1(n8891), .A2(n8667), .B1(n8665), .B2(n8889), .ZN(n7749)
         );
  NAND2_X1 U9468 ( .A1(n7750), .A2(n7749), .ZN(n10201) );
  INV_X1 U9469 ( .A(n10201), .ZN(n7751) );
  MUX2_X1 U9470 ( .A(n6575), .B(n7751), .S(n8895), .Z(n7752) );
  OAI211_X1 U9471 ( .C1(n10200), .C2(n8901), .A(n7753), .B(n7752), .ZN(
        P2_U3227) );
  NAND2_X1 U9472 ( .A1(n7755), .A2(n7754), .ZN(n8411) );
  XNOR2_X1 U9473 ( .A(n7756), .B(n8411), .ZN(n10196) );
  INV_X1 U9474 ( .A(n10196), .ZN(n7763) );
  XNOR2_X1 U9475 ( .A(n7757), .B(n8411), .ZN(n7758) );
  AOI222_X1 U9476 ( .A1(n8894), .A2(n7758), .B1(n8666), .B2(n8889), .C1(n8668), 
        .C2(n8891), .ZN(n10193) );
  MUX2_X1 U9477 ( .A(n8478), .B(n10193), .S(n8895), .Z(n7762) );
  AOI22_X1 U9478 ( .A1(n8898), .A2(n7760), .B1(n8897), .B2(n7759), .ZN(n7761)
         );
  OAI211_X1 U9479 ( .C1(n7763), .C2(n8901), .A(n7762), .B(n7761), .ZN(P2_U3228) );
  OAI22_X1 U9480 ( .A1(n7766), .A2(n8664), .B1(n7765), .B2(n7764), .ZN(n7769)
         );
  XNOR2_X1 U9481 ( .A(n7767), .B(n8663), .ZN(n7768) );
  XNOR2_X1 U9482 ( .A(n7769), .B(n7768), .ZN(n7775) );
  NAND2_X1 U9483 ( .A1(n8640), .A2(n8664), .ZN(n7771) );
  OAI211_X1 U9484 ( .C1(n8620), .C2(n8645), .A(n7771), .B(n7770), .ZN(n7773)
         );
  NOR2_X1 U9485 ( .A1(n8592), .A2(n7782), .ZN(n7772) );
  AOI211_X1 U9486 ( .C1(n7783), .C2(n8641), .A(n7773), .B(n7772), .ZN(n7774)
         );
  OAI21_X1 U9487 ( .B1(n7775), .B2(n8650), .A(n7774), .ZN(P2_U3171) );
  INV_X1 U9488 ( .A(n8283), .ZN(n8420) );
  XNOR2_X1 U9489 ( .A(n7776), .B(n8420), .ZN(n10217) );
  XNOR2_X1 U9490 ( .A(n7778), .B(n8283), .ZN(n7780) );
  AOI22_X1 U9491 ( .A1(n8662), .A2(n8889), .B1(n8891), .B2(n8664), .ZN(n7779)
         );
  OAI21_X1 U9492 ( .B1(n7780), .B2(n5628), .A(n7779), .ZN(n7781) );
  AOI21_X1 U9493 ( .B1(n10217), .B2(n4842), .A(n7781), .ZN(n10219) );
  INV_X1 U9494 ( .A(n8760), .ZN(n7788) );
  NOR2_X1 U9495 ( .A1(n8839), .A2(n7782), .ZN(n7787) );
  INV_X1 U9496 ( .A(n7783), .ZN(n7784) );
  OAI22_X1 U9497 ( .A1(n10174), .A2(n7785), .B1(n7784), .B2(n10165), .ZN(n7786) );
  AOI211_X1 U9498 ( .C1(n10217), .C2(n7788), .A(n7787), .B(n7786), .ZN(n7789)
         );
  OAI21_X1 U9499 ( .B1(n10219), .B2(n10176), .A(n7789), .ZN(P2_U3224) );
  NAND2_X1 U9500 ( .A1(n7791), .A2(n7790), .ZN(n7792) );
  XOR2_X1 U9501 ( .A(n7793), .B(n7792), .Z(n7801) );
  NAND2_X1 U9502 ( .A1(n8640), .A2(n8663), .ZN(n7796) );
  INV_X1 U9503 ( .A(n7794), .ZN(n7795) );
  OAI211_X1 U9504 ( .C1(n7951), .C2(n8645), .A(n7796), .B(n7795), .ZN(n7799)
         );
  INV_X1 U9505 ( .A(n7797), .ZN(n10222) );
  NOR2_X1 U9506 ( .A1(n8592), .A2(n10222), .ZN(n7798) );
  AOI211_X1 U9507 ( .C1(n7904), .C2(n8641), .A(n7799), .B(n7798), .ZN(n7800)
         );
  OAI21_X1 U9508 ( .B1(n7801), .B2(n8650), .A(n7800), .ZN(P2_U3157) );
  INV_X1 U9509 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n7849) );
  NOR2_X1 U9510 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7846) );
  NOR2_X1 U9511 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7842) );
  NOR2_X1 U9512 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7839) );
  NOR2_X1 U9513 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7836) );
  NOR2_X1 U9514 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7832) );
  NOR2_X1 U9515 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7829) );
  NOR2_X1 U9516 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7825) );
  NOR2_X1 U9517 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7821) );
  NOR2_X1 U9518 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7817) );
  NOR2_X1 U9519 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7815) );
  NOR2_X1 U9520 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7813) );
  NOR2_X1 U9521 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7811) );
  NOR2_X1 U9522 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7809) );
  NAND2_X1 U9523 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7807) );
  XOR2_X1 U9524 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10301) );
  NAND2_X1 U9525 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7805) );
  XOR2_X1 U9526 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10299) );
  INV_X1 U9527 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10266) );
  OAI21_X1 U9528 ( .B1(n10267), .B2(n10266), .A(n7802), .ZN(n10262) );
  INV_X1 U9529 ( .A(n10262), .ZN(n7803) );
  INV_X1 U9530 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10265) );
  NAND3_X1 U9531 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10263) );
  OAI21_X1 U9532 ( .B1(n7803), .B2(n10265), .A(n10263), .ZN(n10298) );
  NAND2_X1 U9533 ( .A1(n10299), .A2(n10298), .ZN(n7804) );
  NAND2_X1 U9534 ( .A1(n7805), .A2(n7804), .ZN(n10300) );
  NAND2_X1 U9535 ( .A1(n10301), .A2(n10300), .ZN(n7806) );
  NAND2_X1 U9536 ( .A1(n7807), .A2(n7806), .ZN(n10303) );
  XOR2_X1 U9537 ( .A(n9471), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n10302) );
  NOR2_X1 U9538 ( .A1(n10303), .A2(n10302), .ZN(n7808) );
  NOR2_X1 U9539 ( .A1(n7809), .A2(n7808), .ZN(n10291) );
  XNOR2_X1 U9540 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10290) );
  NOR2_X1 U9541 ( .A1(n10291), .A2(n10290), .ZN(n7810) );
  NOR2_X1 U9542 ( .A1(n7811), .A2(n7810), .ZN(n10289) );
  XNOR2_X1 U9543 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n10288) );
  NOR2_X1 U9544 ( .A1(n10289), .A2(n10288), .ZN(n7812) );
  NOR2_X1 U9545 ( .A1(n7813), .A2(n7812), .ZN(n10295) );
  XNOR2_X1 U9546 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10294) );
  NOR2_X1 U9547 ( .A1(n10295), .A2(n10294), .ZN(n7814) );
  NOR2_X1 U9548 ( .A1(n7815), .A2(n7814), .ZN(n10297) );
  XNOR2_X1 U9549 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10296) );
  NOR2_X1 U9550 ( .A1(n10297), .A2(n10296), .ZN(n7816) );
  NOR2_X1 U9551 ( .A1(n7817), .A2(n7816), .ZN(n10293) );
  INV_X1 U9552 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n7819) );
  INV_X1 U9553 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7818) );
  AOI22_X1 U9554 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7819), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n7818), .ZN(n10292) );
  NOR2_X1 U9555 ( .A1(n10293), .A2(n10292), .ZN(n7820) );
  NOR2_X1 U9556 ( .A1(n7821), .A2(n7820), .ZN(n10287) );
  INV_X1 U9557 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7823) );
  AOI22_X1 U9558 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n7823), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n7822), .ZN(n10286) );
  NOR2_X1 U9559 ( .A1(n10287), .A2(n10286), .ZN(n7824) );
  NOR2_X1 U9560 ( .A1(n7825), .A2(n7824), .ZN(n10285) );
  INV_X1 U9561 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7827) );
  INV_X1 U9562 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7826) );
  AOI22_X1 U9563 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n7827), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n7826), .ZN(n10284) );
  NOR2_X1 U9564 ( .A1(n10285), .A2(n10284), .ZN(n7828) );
  NOR2_X1 U9565 ( .A1(n7829), .A2(n7828), .ZN(n10283) );
  XOR2_X1 U9566 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n7830), .Z(n10282) );
  NOR2_X1 U9567 ( .A1(n10283), .A2(n10282), .ZN(n7831) );
  NOR2_X1 U9568 ( .A1(n7832), .A2(n7831), .ZN(n10281) );
  INV_X1 U9569 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7834) );
  INV_X1 U9570 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7833) );
  AOI22_X1 U9571 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(n7834), .B1(
        P1_ADDR_REG_13__SCAN_IN), .B2(n7833), .ZN(n10280) );
  NOR2_X1 U9572 ( .A1(n10281), .A2(n10280), .ZN(n7835) );
  NOR2_X1 U9573 ( .A1(n7836), .A2(n7835), .ZN(n10279) );
  XOR2_X1 U9574 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(n7837), .Z(n10278) );
  NOR2_X1 U9575 ( .A1(n10279), .A2(n10278), .ZN(n7838) );
  NOR2_X1 U9576 ( .A1(n7839), .A2(n7838), .ZN(n10277) );
  INV_X1 U9577 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7840) );
  INV_X1 U9578 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8681) );
  AOI22_X1 U9579 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n7840), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n8681), .ZN(n10276) );
  NOR2_X1 U9580 ( .A1(n10277), .A2(n10276), .ZN(n7841) );
  NOR2_X1 U9581 ( .A1(n7842), .A2(n7841), .ZN(n10275) );
  INV_X1 U9582 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7844) );
  INV_X1 U9583 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7843) );
  AOI22_X1 U9584 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n7844), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n7843), .ZN(n10274) );
  NOR2_X1 U9585 ( .A1(n10275), .A2(n10274), .ZN(n7845) );
  NOR2_X1 U9586 ( .A1(n7846), .A2(n7845), .ZN(n10273) );
  AOI22_X1 U9587 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n7848), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(n7849), .ZN(n10272) );
  NOR2_X1 U9588 ( .A1(n10273), .A2(n10272), .ZN(n7847) );
  AOI21_X1 U9589 ( .B1(n7849), .B2(n7848), .A(n7847), .ZN(n10269) );
  NOR2_X1 U9590 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10269), .ZN(n7850) );
  NAND2_X1 U9591 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10269), .ZN(n10268) );
  OAI21_X1 U9592 ( .B1(n10270), .B2(n7850), .A(n10268), .ZN(n7852) );
  XNOR2_X1 U9593 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7851) );
  XNOR2_X1 U9594 ( .A(n7852), .B(n7851), .ZN(ADD_1068_U4) );
  INV_X1 U9595 ( .A(n7853), .ZN(n7856) );
  OAI222_X1 U9596 ( .A1(n4428), .A2(n7855), .B1(n8472), .B2(n7856), .C1(
        P1_U3086), .C2(n7854), .ZN(P1_U3333) );
  OAI222_X1 U9597 ( .A1(n8549), .A2(n7857), .B1(n9024), .B2(n7856), .C1(
        P2_U3151), .C2(n8248), .ZN(P2_U3273) );
  XNOR2_X1 U9598 ( .A(n7858), .B(n8005), .ZN(n7859) );
  NOR2_X1 U9599 ( .A1(n7859), .A2(n7860), .ZN(n8004) );
  AOI21_X1 U9600 ( .B1(n7860), .B2(n7859), .A(n8004), .ZN(n7868) );
  INV_X1 U9601 ( .A(n7861), .ZN(n7864) );
  AOI22_X1 U9602 ( .A1(n9165), .A2(n7862), .B1(P1_REG3_REG_8__SCAN_IN), .B2(
        P1_U3086), .ZN(n7863) );
  OAI21_X1 U9603 ( .B1(n7864), .B2(n9168), .A(n7863), .ZN(n7865) );
  AOI21_X1 U9604 ( .B1(n7866), .B2(n9171), .A(n7865), .ZN(n7867) );
  OAI21_X1 U9605 ( .B1(n7868), .B2(n9174), .A(n7867), .ZN(P1_U3221) );
  OAI22_X1 U9606 ( .A1(n8839), .A2(n7869), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n10165), .ZN(n7872) );
  MUX2_X1 U9607 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n7870), .S(n8895), .Z(n7871)
         );
  AOI211_X1 U9608 ( .C1(n5715), .C2(n7873), .A(n7872), .B(n7871), .ZN(n7874)
         );
  INV_X1 U9609 ( .A(n7874), .ZN(P2_U3230) );
  OR2_X1 U9610 ( .A1(n8045), .A2(n8044), .ZN(n9224) );
  NAND2_X1 U9611 ( .A1(n8045), .A2(n8044), .ZN(n9219) );
  AOI21_X2 U9612 ( .B1(n7877), .B2(n7876), .A(n7875), .ZN(n9903) );
  INV_X1 U9613 ( .A(n9442), .ZN(n7878) );
  NAND2_X1 U9614 ( .A1(n9905), .A2(n7878), .ZN(n9213) );
  OAI22_X2 U9615 ( .A1(n9903), .A2(n9902), .B1(n9905), .B2(n9442), .ZN(n8043)
         );
  XOR2_X1 U9616 ( .A(n9306), .B(n8043), .Z(n10096) );
  INV_X1 U9617 ( .A(n10096), .ZN(n7891) );
  INV_X1 U9618 ( .A(n9894), .ZN(n9212) );
  INV_X1 U9619 ( .A(n9213), .ZN(n9220) );
  NAND2_X1 U9620 ( .A1(n7880), .A2(n9306), .ZN(n8038) );
  OAI211_X1 U9621 ( .C1(n7880), .C2(n9306), .A(n8038), .B(n9980), .ZN(n7883)
         );
  NAND2_X1 U9622 ( .A1(n9440), .A2(n9152), .ZN(n7882) );
  NAND2_X1 U9623 ( .A1(n9442), .A2(n9604), .ZN(n7881) );
  AND2_X1 U9624 ( .A1(n7882), .A2(n7881), .ZN(n9033) );
  NAND2_X1 U9625 ( .A1(n7883), .A2(n9033), .ZN(n10094) );
  INV_X1 U9626 ( .A(n9906), .ZN(n7885) );
  INV_X1 U9627 ( .A(n8051), .ZN(n7884) );
  OAI211_X1 U9628 ( .C1(n10092), .C2(n7885), .A(n7884), .B(n9985), .ZN(n10090)
         );
  OAI22_X1 U9629 ( .A1(n9744), .A2(n7886), .B1(n9031), .B2(n8523), .ZN(n7887)
         );
  AOI21_X1 U9630 ( .B1(n8045), .B2(n9981), .A(n7887), .ZN(n7888) );
  OAI21_X1 U9631 ( .B1(n10090), .B2(n9987), .A(n7888), .ZN(n7889) );
  AOI21_X1 U9632 ( .B1(n10094), .B2(n9744), .A(n7889), .ZN(n7890) );
  OAI21_X1 U9633 ( .B1(n7891), .B2(n9746), .A(n7890), .ZN(P1_U3279) );
  XNOR2_X1 U9634 ( .A(n7893), .B(n7892), .ZN(n7894) );
  OAI222_X1 U9635 ( .A1(n10171), .A2(n8621), .B1(n5626), .B2(n8620), .C1(n7894), .C2(n5628), .ZN(n10228) );
  INV_X1 U9636 ( .A(n10228), .ZN(n7900) );
  OAI21_X1 U9637 ( .B1(n7896), .B2(n8419), .A(n7895), .ZN(n10230) );
  INV_X1 U9638 ( .A(n8624), .ZN(n10227) );
  AOI22_X1 U9639 ( .A1(n10176), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n8897), .B2(
        n8625), .ZN(n7897) );
  OAI21_X1 U9640 ( .B1(n10227), .B2(n8839), .A(n7897), .ZN(n7898) );
  AOI21_X1 U9641 ( .B1(n10230), .B2(n5715), .A(n7898), .ZN(n7899) );
  OAI21_X1 U9642 ( .B1(n7900), .B2(n10176), .A(n7899), .ZN(P2_U3222) );
  XNOR2_X1 U9643 ( .A(n7901), .B(n8418), .ZN(n7902) );
  AOI222_X1 U9644 ( .A1(n8894), .A2(n7902), .B1(n8661), .B2(n8889), .C1(n8663), 
        .C2(n8891), .ZN(n10221) );
  XNOR2_X1 U9645 ( .A(n7903), .B(n8418), .ZN(n10224) );
  NOR2_X1 U9646 ( .A1(n10222), .A2(n8839), .ZN(n7907) );
  INV_X1 U9647 ( .A(n7904), .ZN(n7905) );
  OAI22_X1 U9648 ( .A1(n10174), .A2(n6586), .B1(n7905), .B2(n10165), .ZN(n7906) );
  AOI211_X1 U9649 ( .C1(n10224), .C2(n5715), .A(n7907), .B(n7906), .ZN(n7908)
         );
  OAI21_X1 U9650 ( .B1(n10221), .B2(n10176), .A(n7908), .ZN(P2_U3223) );
  NAND2_X1 U9651 ( .A1(n7913), .A2(n7909), .ZN(n7911) );
  OR2_X1 U9652 ( .A1(n7910), .A2(P1_U3086), .ZN(n9414) );
  OAI211_X1 U9653 ( .C1(n7912), .C2(n4428), .A(n7911), .B(n9414), .ZN(P1_U3332) );
  NAND2_X1 U9654 ( .A1(n7913), .A2(n8159), .ZN(n7915) );
  NAND2_X1 U9655 ( .A1(n7914), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8466) );
  OAI211_X1 U9656 ( .C1(n7916), .C2(n8549), .A(n7915), .B(n8466), .ZN(P2_U3272) );
  OAI21_X1 U9657 ( .B1(n7921), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7917), .ZN(
        n7920) );
  INV_X1 U9658 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7918) );
  AOI22_X1 U9659 ( .A1(n9484), .A2(n7918), .B1(P1_REG2_REG_13__SCAN_IN), .B2(
        n9492), .ZN(n7919) );
  NOR2_X1 U9660 ( .A1(n7919), .A2(n7920), .ZN(n9483) );
  AOI211_X1 U9661 ( .C1(n7920), .C2(n7919), .A(n9483), .B(n9879), .ZN(n7931)
         );
  NOR2_X1 U9662 ( .A1(n7921), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7922) );
  NOR2_X1 U9663 ( .A1(n7923), .A2(n7922), .ZN(n7926) );
  INV_X1 U9664 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7924) );
  MUX2_X1 U9665 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n7924), .S(n9484), .Z(n7925)
         );
  NAND2_X1 U9666 ( .A1(n7925), .A2(n7926), .ZN(n9491) );
  OAI211_X1 U9667 ( .C1(n7926), .C2(n7925), .A(n9888), .B(n9491), .ZN(n7929)
         );
  NOR2_X1 U9668 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8020), .ZN(n7927) );
  AOI21_X1 U9669 ( .B1(n9878), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n7927), .ZN(
        n7928) );
  OAI211_X1 U9670 ( .C1(n9578), .C2(n9492), .A(n7929), .B(n7928), .ZN(n7930)
         );
  OR2_X1 U9671 ( .A1(n7931), .A2(n7930), .ZN(P1_U3256) );
  XNOR2_X1 U9672 ( .A(n7932), .B(n8621), .ZN(n7933) );
  XNOR2_X1 U9673 ( .A(n7934), .B(n7933), .ZN(n7939) );
  NAND2_X1 U9674 ( .A1(n5372), .A2(n8632), .ZN(n7935) );
  NAND2_X1 U9675 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3151), .ZN(n8135) );
  OAI211_X1 U9676 ( .C1(n7951), .C2(n8635), .A(n7935), .B(n8135), .ZN(n7936)
         );
  AOI21_X1 U9677 ( .B1(n7958), .B2(n8641), .A(n7936), .ZN(n7938) );
  NAND2_X1 U9678 ( .A1(n10232), .A2(n8648), .ZN(n7937) );
  OAI211_X1 U9679 ( .C1(n7939), .C2(n8650), .A(n7938), .B(n7937), .ZN(P2_U3164) );
  XOR2_X1 U9680 ( .A(n7940), .B(n7941), .Z(n7949) );
  NAND2_X1 U9681 ( .A1(n9165), .A2(n7942), .ZN(n7943) );
  OAI211_X1 U9682 ( .C1(n9168), .C2(n7945), .A(n7944), .B(n7943), .ZN(n7946)
         );
  AOI21_X1 U9683 ( .B1(n7947), .B2(n9171), .A(n7946), .ZN(n7948) );
  OAI21_X1 U9684 ( .B1(n7949), .B2(n9174), .A(n7948), .ZN(P1_U3224) );
  XNOR2_X1 U9685 ( .A(n7950), .B(n8308), .ZN(n7954) );
  OAI22_X1 U9686 ( .A1(n7952), .A2(n10171), .B1(n7951), .B2(n5626), .ZN(n7953)
         );
  AOI21_X1 U9687 ( .B1(n7954), .B2(n8894), .A(n7953), .ZN(n10236) );
  OAI21_X1 U9688 ( .B1(n7956), .B2(n8308), .A(n7955), .ZN(n7957) );
  INV_X1 U9689 ( .A(n7957), .ZN(n10235) );
  INV_X1 U9690 ( .A(n10232), .ZN(n7960) );
  AOI22_X1 U9691 ( .A1(n10176), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n8897), .B2(
        n7958), .ZN(n7959) );
  OAI21_X1 U9692 ( .B1(n7960), .B2(n8839), .A(n7959), .ZN(n7961) );
  AOI21_X1 U9693 ( .B1(n10235), .B2(n5715), .A(n7961), .ZN(n7962) );
  OAI21_X1 U9694 ( .B1(n10176), .B2(n10236), .A(n7962), .ZN(P2_U3221) );
  XNOR2_X1 U9695 ( .A(n7963), .B(n8063), .ZN(n7965) );
  NOR2_X1 U9696 ( .A1(n7965), .A2(n7964), .ZN(n8062) );
  AOI21_X1 U9697 ( .B1(n7965), .B2(n7964), .A(n8062), .ZN(n7972) );
  OAI22_X1 U9698 ( .A1(n9156), .A2(n7967), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7966), .ZN(n7969) );
  NOR2_X1 U9699 ( .A1(n10068), .A2(n9161), .ZN(n7968) );
  AOI211_X1 U9700 ( .C1(n9158), .C2(n7970), .A(n7969), .B(n7968), .ZN(n7971)
         );
  OAI21_X1 U9701 ( .B1(n7972), .B2(n9174), .A(n7971), .ZN(P1_U3217) );
  INV_X1 U9702 ( .A(n7973), .ZN(n8313) );
  OR2_X1 U9703 ( .A1(n8314), .A2(n8313), .ZN(n8423) );
  INV_X1 U9704 ( .A(n8423), .ZN(n8312) );
  XNOR2_X1 U9705 ( .A(n7974), .B(n8312), .ZN(n9837) );
  XNOR2_X1 U9706 ( .A(n7975), .B(n8312), .ZN(n7976) );
  OAI222_X1 U9707 ( .A1(n5626), .A2(n8621), .B1(n10171), .B2(n8123), .C1(n5628), .C2(n7976), .ZN(n9839) );
  INV_X1 U9708 ( .A(n8032), .ZN(n7977) );
  OAI22_X1 U9709 ( .A1(n4894), .A2(n10167), .B1(n7977), .B2(n10165), .ZN(n7978) );
  OAI21_X1 U9710 ( .B1(n9839), .B2(n7978), .A(n10174), .ZN(n7980) );
  NAND2_X1 U9711 ( .A1(n10176), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7979) );
  OAI211_X1 U9712 ( .C1(n9837), .C2(n8901), .A(n7980), .B(n7979), .ZN(P2_U3220) );
  INV_X1 U9713 ( .A(n7981), .ZN(n8026) );
  OAI222_X1 U9714 ( .A1(n9024), .A2(n8026), .B1(P2_U3151), .B2(n7983), .C1(
        n7982), .C2(n8549), .ZN(P2_U3271) );
  OAI21_X1 U9715 ( .B1(n7986), .B2(n7985), .A(n7984), .ZN(n8002) );
  NAND2_X1 U9716 ( .A1(n10141), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n7996) );
  INV_X1 U9717 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7987) );
  OR2_X1 U9718 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7987), .ZN(n8619) );
  NAND2_X1 U9719 ( .A1(n7990), .A2(n7989), .ZN(n7991) );
  NAND2_X1 U9720 ( .A1(n7988), .A2(n7991), .ZN(n7992) );
  NAND2_X1 U9721 ( .A1(n8741), .A2(n7992), .ZN(n7995) );
  NAND2_X1 U9722 ( .A1(n8699), .A2(n7993), .ZN(n7994) );
  NAND4_X1 U9723 ( .A1(n7996), .A2(n8619), .A3(n7995), .A4(n7994), .ZN(n8001)
         );
  AOI21_X1 U9724 ( .B1(n7998), .B2(n10258), .A(n7997), .ZN(n7999) );
  NOR2_X1 U9725 ( .A1(n7999), .A2(n10147), .ZN(n8000) );
  AOI211_X1 U9726 ( .C1(n10152), .C2(n8002), .A(n8001), .B(n8000), .ZN(n8003)
         );
  INV_X1 U9727 ( .A(n8003), .ZN(P2_U3193) );
  AOI21_X1 U9728 ( .B1(n8005), .B2(n7858), .A(n8004), .ZN(n8009) );
  XNOR2_X1 U9729 ( .A(n8007), .B(n8006), .ZN(n8008) );
  XNOR2_X1 U9730 ( .A(n8009), .B(n8008), .ZN(n8017) );
  AOI21_X1 U9731 ( .B1(n8011), .B2(n8010), .A(n9156), .ZN(n8012) );
  AOI211_X1 U9732 ( .C1(n9158), .C2(n8014), .A(n8013), .B(n8012), .ZN(n8016)
         );
  NAND2_X1 U9733 ( .A1(n10058), .A2(n9171), .ZN(n8015) );
  OAI211_X1 U9734 ( .C1(n8017), .C2(n9174), .A(n8016), .B(n8015), .ZN(P1_U3231) );
  XOR2_X1 U9735 ( .A(n8018), .B(n8019), .Z(n8024) );
  AOI22_X1 U9736 ( .A1(n9152), .A2(n9441), .B1(n9443), .B2(n9604), .ZN(n9898)
         );
  OAI22_X1 U9737 ( .A1(n9898), .A2(n9156), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8020), .ZN(n8021) );
  AOI21_X1 U9738 ( .B1(n9901), .B2(n9158), .A(n8021), .ZN(n8023) );
  NAND2_X1 U9739 ( .A1(n9905), .A2(n9171), .ZN(n8022) );
  OAI211_X1 U9740 ( .C1(n8024), .C2(n9174), .A(n8023), .B(n8022), .ZN(P1_U3234) );
  OAI222_X1 U9741 ( .A1(n8027), .A2(P1_U3086), .B1(n8472), .B2(n8026), .C1(
        n8025), .C2(n4428), .ZN(P1_U3331) );
  NAND2_X1 U9742 ( .A1(n8029), .A2(n8028), .ZN(n8031) );
  XOR2_X1 U9743 ( .A(n8031), .B(n8030), .Z(n8037) );
  NOR2_X1 U9744 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5034), .ZN(n8185) );
  AOI21_X1 U9745 ( .B1(n8660), .B2(n8640), .A(n8185), .ZN(n8034) );
  NAND2_X1 U9746 ( .A1(n8641), .A2(n8032), .ZN(n8033) );
  OAI211_X1 U9747 ( .C1(n8123), .C2(n8645), .A(n8034), .B(n8033), .ZN(n8035)
         );
  AOI21_X1 U9748 ( .B1(n9840), .B2(n8648), .A(n8035), .ZN(n8036) );
  OAI21_X1 U9749 ( .B1(n8037), .B2(n8650), .A(n8036), .ZN(P2_U3174) );
  NAND2_X1 U9750 ( .A1(n8038), .A2(n9224), .ZN(n8040) );
  INV_X1 U9751 ( .A(n8040), .ZN(n8041) );
  OR2_X1 U9752 ( .A1(n9172), .A2(n8039), .ZN(n9379) );
  NAND2_X1 U9753 ( .A1(n9172), .A2(n8039), .ZN(n9225) );
  NAND2_X1 U9754 ( .A1(n9379), .A2(n9225), .ZN(n8048) );
  INV_X1 U9755 ( .A(n8048), .ZN(n9307) );
  OAI21_X1 U9756 ( .B1(n8041), .B2(n9307), .A(n8084), .ZN(n8042) );
  OAI22_X1 U9757 ( .A1(n8169), .A2(n9128), .B1(n8044), .B2(n9114), .ZN(n9166)
         );
  AOI21_X1 U9758 ( .B1(n8042), .B2(n9980), .A(n9166), .ZN(n9858) );
  AOI21_X1 U9759 ( .B1(n10092), .B2(n8044), .A(n8043), .ZN(n8047) );
  XNOR2_X1 U9760 ( .A(n8088), .B(n8048), .ZN(n9861) );
  NAND2_X1 U9761 ( .A1(n9861), .A2(n9968), .ZN(n8055) );
  INV_X1 U9762 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8050) );
  INV_X1 U9763 ( .A(n8049), .ZN(n9169) );
  OAI22_X1 U9764 ( .A1(n9744), .A2(n8050), .B1(n9169), .B2(n8523), .ZN(n8053)
         );
  OAI211_X1 U9765 ( .C1(n9859), .C2(n8051), .A(n4661), .B(n9985), .ZN(n9857)
         );
  NOR2_X1 U9766 ( .A1(n9857), .A2(n9987), .ZN(n8052) );
  AOI211_X1 U9767 ( .C1(n9981), .C2(n9172), .A(n8053), .B(n8052), .ZN(n8054)
         );
  OAI211_X1 U9768 ( .C1(n9992), .C2(n9858), .A(n8055), .B(n8054), .ZN(P1_U3278) );
  INV_X1 U9769 ( .A(n8056), .ZN(n8060) );
  OAI222_X1 U9770 ( .A1(n9024), .A2(n8060), .B1(P2_U3151), .B2(n8058), .C1(
        n8057), .C2(n8549), .ZN(P2_U3270) );
  OAI222_X1 U9771 ( .A1(n8061), .A2(P1_U3086), .B1(n8472), .B2(n8060), .C1(
        n8059), .C2(n4428), .ZN(P1_U3330) );
  AOI21_X1 U9772 ( .B1(n8063), .B2(n7963), .A(n8062), .ZN(n8067) );
  XNOR2_X1 U9773 ( .A(n8065), .B(n8064), .ZN(n8066) );
  XNOR2_X1 U9774 ( .A(n8067), .B(n8066), .ZN(n8074) );
  OAI22_X1 U9775 ( .A1(n8069), .A2(n9114), .B1(n8068), .B2(n9128), .ZN(n9916)
         );
  AOI22_X1 U9776 ( .A1(n9916), .A2(n9165), .B1(P1_REG3_REG_11__SCAN_IN), .B2(
        P1_U3086), .ZN(n8070) );
  OAI21_X1 U9777 ( .B1(n8071), .B2(n9168), .A(n8070), .ZN(n8072) );
  AOI21_X1 U9778 ( .B1(n9920), .B2(n9171), .A(n8072), .ZN(n8073) );
  OAI21_X1 U9779 ( .B1(n8074), .B2(n9174), .A(n8073), .ZN(P1_U3236) );
  XOR2_X1 U9780 ( .A(n8075), .B(n8076), .Z(n8081) );
  AOI22_X1 U9781 ( .A1(n5372), .A2(n8640), .B1(P2_REG3_REG_14__SCAN_IN), .B2(
        P2_U3151), .ZN(n8078) );
  NAND2_X1 U9782 ( .A1(n8641), .A2(n8103), .ZN(n8077) );
  OAI211_X1 U9783 ( .C1(n8200), .C2(n8645), .A(n8078), .B(n8077), .ZN(n8079)
         );
  AOI21_X1 U9784 ( .B1(n8114), .B2(n8648), .A(n8079), .ZN(n8080) );
  OAI21_X1 U9785 ( .B1(n8081), .B2(n8650), .A(n8080), .ZN(P2_U3155) );
  INV_X1 U9786 ( .A(n8082), .ZN(n8099) );
  OAI222_X1 U9787 ( .A1(n9024), .A2(n8099), .B1(P2_U3151), .B2(n5632), .C1(
        n8083), .C2(n8549), .ZN(P2_U3269) );
  NAND2_X1 U9788 ( .A1(n9083), .A2(n8169), .ZN(n9383) );
  OAI21_X1 U9789 ( .B1(n9308), .B2(n8085), .A(n8165), .ZN(n8087) );
  AOI22_X1 U9790 ( .A1(n9438), .A2(n9152), .B1(n9604), .B2(n9440), .ZN(n9080)
         );
  INV_X1 U9791 ( .A(n9080), .ZN(n8086) );
  AOI21_X1 U9792 ( .B1(n8087), .B2(n9980), .A(n8086), .ZN(n9852) );
  NOR2_X1 U9793 ( .A1(n8088), .A2(n9859), .ZN(n8090) );
  AND2_X1 U9794 ( .A1(n8091), .A2(n9308), .ZN(n9849) );
  OR3_X1 U9795 ( .A1(n9850), .A2(n9746), .A3(n9849), .ZN(n8097) );
  INV_X1 U9796 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9523) );
  OAI22_X1 U9797 ( .A1(n9744), .A2(n9523), .B1(n9078), .B2(n8523), .ZN(n8095)
         );
  INV_X1 U9798 ( .A(n9083), .ZN(n9853) );
  INV_X1 U9799 ( .A(n8170), .ZN(n8092) );
  OAI211_X1 U9800 ( .C1(n9853), .C2(n8093), .A(n8092), .B(n9985), .ZN(n9851)
         );
  NOR2_X1 U9801 ( .A1(n9851), .A2(n9987), .ZN(n8094) );
  AOI211_X1 U9802 ( .C1(n9981), .C2(n9083), .A(n8095), .B(n8094), .ZN(n8096)
         );
  OAI211_X1 U9803 ( .C1(n9992), .C2(n9852), .A(n8097), .B(n8096), .ZN(P1_U3277) );
  OAI222_X1 U9804 ( .A1(n8100), .A2(P1_U3086), .B1(n8472), .B2(n8099), .C1(
        n8098), .C2(n4428), .ZN(P1_U3329) );
  NAND2_X1 U9805 ( .A1(n8320), .A2(n8317), .ZN(n8425) );
  XOR2_X1 U9806 ( .A(n8101), .B(n8425), .Z(n8102) );
  AOI222_X1 U9807 ( .A1(n8894), .A2(n8102), .B1(n5372), .B2(n8891), .C1(n8892), 
        .C2(n8889), .ZN(n8112) );
  AOI22_X1 U9808 ( .A1(n8114), .A2(n8104), .B1(n8897), .B2(n8103), .ZN(n8105)
         );
  AOI21_X1 U9809 ( .B1(n8112), .B2(n8105), .A(n10176), .ZN(n8108) );
  XNOR2_X1 U9810 ( .A(n8106), .B(n8425), .ZN(n8117) );
  OAI22_X1 U9811 ( .A1(n8117), .A2(n8901), .B1(n6598), .B2(n8895), .ZN(n8107)
         );
  OR2_X1 U9812 ( .A1(n8108), .A2(n8107), .ZN(P2_U3219) );
  INV_X1 U9813 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8109) );
  MUX2_X1 U9814 ( .A(n8109), .B(n8112), .S(n10238), .Z(n8111) );
  NAND2_X1 U9815 ( .A1(n8114), .A2(n9009), .ZN(n8110) );
  OAI211_X1 U9816 ( .C1(n8117), .C2(n9017), .A(n8111), .B(n8110), .ZN(P2_U3432) );
  MUX2_X1 U9817 ( .A(n8113), .B(n8112), .S(n10261), .Z(n8116) );
  NAND2_X1 U9818 ( .A1(n8114), .A2(n8937), .ZN(n8115) );
  OAI211_X1 U9819 ( .C1(n8944), .C2(n8117), .A(n8116), .B(n8115), .ZN(P2_U3473) );
  XNOR2_X1 U9820 ( .A(n8941), .B(n8892), .ZN(n8426) );
  XOR2_X1 U9821 ( .A(n8426), .B(n8118), .Z(n9018) );
  INV_X1 U9822 ( .A(n8155), .ZN(n8119) );
  OAI22_X1 U9823 ( .A1(n10174), .A2(n8673), .B1(n8119), .B2(n10165), .ZN(n8120) );
  AOI21_X1 U9824 ( .B1(n8941), .B2(n8898), .A(n8120), .ZN(n8125) );
  XNOR2_X1 U9825 ( .A(n8121), .B(n8426), .ZN(n8122) );
  OAI222_X1 U9826 ( .A1(n10171), .A2(n8227), .B1(n5626), .B2(n8123), .C1(n8122), .C2(n5628), .ZN(n8940) );
  NAND2_X1 U9827 ( .A1(n8940), .A2(n8895), .ZN(n8124) );
  OAI211_X1 U9828 ( .C1(n9018), .C2(n8901), .A(n8125), .B(n8124), .ZN(P2_U3218) );
  INV_X1 U9829 ( .A(n8126), .ZN(n8147) );
  AOI21_X1 U9830 ( .B1(n9022), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n8127), .ZN(
        n8128) );
  OAI21_X1 U9831 ( .B1(n8147), .B2(n9024), .A(n8128), .ZN(P2_U3268) );
  INV_X1 U9832 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n8146) );
  OAI21_X1 U9833 ( .B1(n8131), .B2(n8130), .A(n8129), .ZN(n8139) );
  AOI21_X1 U9834 ( .B1(n4449), .B2(n8133), .A(n8132), .ZN(n8134) );
  NOR2_X1 U9835 ( .A1(n10147), .A2(n8134), .ZN(n8138) );
  OAI21_X1 U9836 ( .B1(n10162), .B2(n8136), .A(n8135), .ZN(n8137) );
  AOI211_X1 U9837 ( .C1(n8741), .C2(n8139), .A(n8138), .B(n8137), .ZN(n8145)
         );
  OAI21_X1 U9838 ( .B1(n8142), .B2(n8141), .A(n8140), .ZN(n8143) );
  NAND2_X1 U9839 ( .A1(n8143), .A2(n10152), .ZN(n8144) );
  OAI211_X1 U9840 ( .C1(n8682), .C2(n8146), .A(n8145), .B(n8144), .ZN(P2_U3194) );
  OAI222_X1 U9841 ( .A1(n4428), .A2(n8148), .B1(n9834), .B2(n8147), .C1(n4426), 
        .C2(P1_U3086), .ZN(P1_U3328) );
  INV_X1 U9842 ( .A(n8941), .ZN(n8158) );
  AOI21_X1 U9843 ( .B1(n8150), .B2(n8149), .A(n8650), .ZN(n8152) );
  NAND2_X1 U9844 ( .A1(n8152), .A2(n8151), .ZN(n8157) );
  AND2_X1 U9845 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8678) );
  AOI21_X1 U9846 ( .B1(n8659), .B2(n8640), .A(n8678), .ZN(n8153) );
  OAI21_X1 U9847 ( .B1(n8227), .B2(n8645), .A(n8153), .ZN(n8154) );
  AOI21_X1 U9848 ( .B1(n8155), .B2(n8641), .A(n8154), .ZN(n8156) );
  OAI211_X1 U9849 ( .C1(n8158), .C2(n8592), .A(n8157), .B(n8156), .ZN(P2_U3181) );
  NAND2_X1 U9850 ( .A1(n8217), .A2(n8159), .ZN(n8161) );
  OAI211_X1 U9851 ( .C1(n8549), .C2(n8162), .A(n8161), .B(n8160), .ZN(P2_U3267) );
  NAND2_X1 U9852 ( .A1(n8165), .A2(n9383), .ZN(n8163) );
  OR2_X1 U9853 ( .A1(n9097), .A2(n8204), .ZN(n9243) );
  NAND2_X1 U9854 ( .A1(n9097), .A2(n8204), .ZN(n9231) );
  NAND2_X1 U9855 ( .A1(n9243), .A2(n9231), .ZN(n9310) );
  AOI21_X1 U9856 ( .B1(n8163), .B2(n9310), .A(n9913), .ZN(n8168) );
  INV_X1 U9857 ( .A(n9383), .ZN(n9228) );
  NOR2_X1 U9858 ( .A1(n9310), .A2(n9228), .ZN(n8164) );
  NAND2_X1 U9859 ( .A1(n9437), .A2(n9152), .ZN(n8167) );
  OR2_X1 U9860 ( .A1(n8169), .A2(n9114), .ZN(n8166) );
  NAND2_X1 U9861 ( .A1(n8167), .A2(n8166), .ZN(n9090) );
  AOI21_X1 U9862 ( .B1(n8168), .B2(n8495), .A(n9090), .ZN(n9845) );
  INV_X1 U9863 ( .A(n8169), .ZN(n9439) );
  XNOR2_X1 U9864 ( .A(n8206), .B(n9310), .ZN(n9848) );
  NAND2_X1 U9865 ( .A1(n9848), .A2(n9968), .ZN(n8176) );
  OAI211_X1 U9866 ( .C1(n9846), .C2(n8170), .A(n9985), .B(n8209), .ZN(n9844)
         );
  INV_X1 U9867 ( .A(n9844), .ZN(n8174) );
  AOI22_X1 U9868 ( .A1(n9947), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n8171), .B2(
        n9983), .ZN(n8172) );
  OAI21_X1 U9869 ( .B1(n9846), .B2(n9741), .A(n8172), .ZN(n8173) );
  AOI21_X1 U9870 ( .B1(n8174), .B2(n9967), .A(n8173), .ZN(n8175) );
  OAI211_X1 U9871 ( .C1(n9992), .C2(n9845), .A(n8176), .B(n8175), .ZN(P1_U3276) );
  AOI21_X1 U9872 ( .B1(n9841), .B2(n8178), .A(n8177), .ZN(n8193) );
  OAI21_X1 U9873 ( .B1(n8181), .B2(n8180), .A(n8179), .ZN(n8191) );
  AOI21_X1 U9874 ( .B1(n8184), .B2(n8183), .A(n8182), .ZN(n8189) );
  AOI21_X1 U9875 ( .B1(n8699), .B2(n8186), .A(n8185), .ZN(n8188) );
  NAND2_X1 U9876 ( .A1(n10141), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n8187) );
  OAI211_X1 U9877 ( .C1(n10156), .C2(n8189), .A(n8188), .B(n8187), .ZN(n8190)
         );
  AOI21_X1 U9878 ( .B1(n10152), .B2(n8191), .A(n8190), .ZN(n8192) );
  OAI21_X1 U9879 ( .B1(n8193), .B2(n10147), .A(n8192), .ZN(P2_U3195) );
  XNOR2_X1 U9880 ( .A(n8194), .B(n8227), .ZN(n8195) );
  XNOR2_X1 U9881 ( .A(n8196), .B(n8195), .ZN(n8203) );
  NOR2_X1 U9882 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8197), .ZN(n8697) );
  AOI21_X1 U9883 ( .B1(n8890), .B2(n8632), .A(n8697), .ZN(n8199) );
  NAND2_X1 U9884 ( .A1(n8641), .A2(n8896), .ZN(n8198) );
  OAI211_X1 U9885 ( .C1(n8200), .C2(n8635), .A(n8199), .B(n8198), .ZN(n8201)
         );
  AOI21_X1 U9886 ( .B1(n9010), .B2(n8648), .A(n8201), .ZN(n8202) );
  OAI21_X1 U9887 ( .B1(n8203), .B2(n8650), .A(n8202), .ZN(P2_U3166) );
  NAND2_X1 U9888 ( .A1(n8205), .A2(n9438), .ZN(n8208) );
  OR2_X1 U9889 ( .A1(n8206), .A2(n9846), .ZN(n8207) );
  NAND2_X1 U9890 ( .A1(n8208), .A2(n8207), .ZN(n8505) );
  INV_X1 U9891 ( .A(n9437), .ZN(n8507) );
  OR2_X1 U9892 ( .A1(n9810), .A2(n8507), .ZN(n9389) );
  NAND2_X1 U9893 ( .A1(n9810), .A2(n8507), .ZN(n9244) );
  NAND2_X1 U9894 ( .A1(n9389), .A2(n9244), .ZN(n9293) );
  XNOR2_X1 U9895 ( .A(n8505), .B(n9293), .ZN(n9813) );
  AOI211_X1 U9896 ( .C1(n9810), .C2(n8209), .A(n9737), .B(n9734), .ZN(n9809)
         );
  INV_X1 U9897 ( .A(n9810), .ZN(n8506) );
  INV_X1 U9898 ( .A(n9143), .ZN(n8210) );
  AOI22_X1 U9899 ( .A1(n9947), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n8210), .B2(
        n9983), .ZN(n8211) );
  OAI21_X1 U9900 ( .B1(n8506), .B2(n9741), .A(n8211), .ZN(n8215) );
  NAND2_X1 U9901 ( .A1(n8495), .A2(n9243), .ZN(n8212) );
  XNOR2_X1 U9902 ( .A(n8212), .B(n9293), .ZN(n8213) );
  OAI22_X1 U9903 ( .A1(n9115), .A2(n9128), .B1(n8204), .B2(n9114), .ZN(n9140)
         );
  AOI21_X1 U9904 ( .B1(n8213), .B2(n9980), .A(n9140), .ZN(n9812) );
  NOR2_X1 U9905 ( .A1(n9812), .A2(n9947), .ZN(n8214) );
  AOI211_X1 U9906 ( .C1(n9809), .C2(n9967), .A(n8215), .B(n8214), .ZN(n8216)
         );
  OAI21_X1 U9907 ( .B1(n9813), .B2(n9746), .A(n8216), .ZN(P1_U3275) );
  INV_X1 U9908 ( .A(n8217), .ZN(n8218) );
  OAI222_X1 U9909 ( .A1(n4428), .A2(n8219), .B1(P1_U3086), .B2(n6487), .C1(
        n8218), .C2(n9834), .ZN(P1_U3327) );
  INV_X1 U9910 ( .A(n8220), .ZN(n8232) );
  OAI222_X1 U9911 ( .A1(n9024), .A2(n8232), .B1(n8222), .B2(P2_U3151), .C1(
        n8221), .C2(n8549), .ZN(P2_U3266) );
  XNOR2_X1 U9912 ( .A(n8223), .B(n8866), .ZN(n8224) );
  XNOR2_X1 U9913 ( .A(n8225), .B(n8224), .ZN(n8231) );
  NAND2_X1 U9914 ( .A1(n8879), .A2(n8632), .ZN(n8226) );
  NAND2_X1 U9915 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8719) );
  OAI211_X1 U9916 ( .C1(n8227), .C2(n8635), .A(n8226), .B(n8719), .ZN(n8228)
         );
  AOI21_X1 U9917 ( .B1(n8883), .B2(n8641), .A(n8228), .ZN(n8230) );
  NAND2_X1 U9918 ( .A1(n9003), .A2(n8648), .ZN(n8229) );
  OAI211_X1 U9919 ( .C1(n8231), .C2(n8650), .A(n8230), .B(n8229), .ZN(P2_U3168) );
  OAI222_X1 U9920 ( .A1(n4428), .A2(n8539), .B1(n9834), .B2(n8232), .C1(n5930), 
        .C2(P1_U3086), .ZN(P1_U3326) );
  OAI21_X1 U9921 ( .B1(n8233), .B2(n8399), .A(n8445), .ZN(n8235) );
  NAND2_X1 U9922 ( .A1(n8235), .A2(n4438), .ZN(n8364) );
  MUX2_X1 U9923 ( .A(n8654), .B(n8378), .S(n8399), .Z(n8385) );
  INV_X1 U9924 ( .A(n8385), .ZN(n8365) );
  NAND2_X1 U9925 ( .A1(n8350), .A2(n8383), .ZN(n8241) );
  OAI21_X1 U9926 ( .B1(n8236), .B2(n8383), .A(n8357), .ZN(n8238) );
  NAND2_X1 U9927 ( .A1(n8238), .A2(n8237), .ZN(n8240) );
  NAND2_X1 U9928 ( .A1(n8352), .A2(n8399), .ZN(n8239) );
  OAI211_X1 U9929 ( .C1(n8352), .C2(n8241), .A(n8240), .B(n8239), .ZN(n8243)
         );
  INV_X1 U9930 ( .A(n8243), .ZN(n8247) );
  MUX2_X1 U9931 ( .A(n8655), .B(n8765), .S(n8399), .Z(n8242) );
  OAI21_X1 U9932 ( .B1(n8244), .B2(n8243), .A(n8242), .ZN(n8245) );
  OAI21_X1 U9933 ( .B1(n8247), .B2(n8246), .A(n8245), .ZN(n8363) );
  NAND2_X1 U9934 ( .A1(n8253), .A2(n8248), .ZN(n8249) );
  MUX2_X1 U9935 ( .A(n8250), .B(n8249), .S(n5753), .Z(n8257) );
  INV_X1 U9936 ( .A(n8251), .ZN(n8252) );
  INV_X1 U9937 ( .A(n8253), .ZN(n8254) );
  NOR2_X1 U9938 ( .A1(n8408), .A2(n8254), .ZN(n8256) );
  AOI21_X1 U9939 ( .B1(n8257), .B2(n8256), .A(n8255), .ZN(n8263) );
  NAND2_X1 U9940 ( .A1(n8264), .A2(n8258), .ZN(n8261) );
  NAND2_X1 U9941 ( .A1(n8274), .A2(n8259), .ZN(n8260) );
  MUX2_X1 U9942 ( .A(n8261), .B(n8260), .S(n8383), .Z(n8262) );
  NAND2_X1 U9943 ( .A1(n8275), .A2(n8264), .ZN(n8266) );
  NAND3_X1 U9944 ( .A1(n8266), .A2(n8276), .A3(n8265), .ZN(n8270) );
  NOR2_X1 U9945 ( .A1(n8271), .A2(n8267), .ZN(n8269) );
  INV_X1 U9946 ( .A(n8279), .ZN(n8268) );
  AOI21_X1 U9947 ( .B1(n8270), .B2(n8269), .A(n8268), .ZN(n8280) );
  NAND2_X1 U9948 ( .A1(n4818), .A2(n8272), .ZN(n8273) );
  AOI21_X1 U9949 ( .B1(n8275), .B2(n8274), .A(n8273), .ZN(n8278) );
  INV_X1 U9950 ( .A(n8292), .ZN(n8282) );
  MUX2_X1 U9951 ( .A(n8282), .B(n8281), .S(n8383), .Z(n8284) );
  NAND2_X1 U9952 ( .A1(n8287), .A2(n8286), .ZN(n8290) );
  NAND2_X1 U9953 ( .A1(n8303), .A2(n8288), .ZN(n8289) );
  AOI21_X1 U9954 ( .B1(n8296), .B2(n8290), .A(n8289), .ZN(n8298) );
  NAND2_X1 U9955 ( .A1(n8292), .A2(n8291), .ZN(n8295) );
  NAND2_X1 U9956 ( .A1(n8301), .A2(n8293), .ZN(n8294) );
  AOI21_X1 U9957 ( .B1(n8296), .B2(n8295), .A(n8294), .ZN(n8297) );
  MUX2_X1 U9958 ( .A(n8298), .B(n8297), .S(n8383), .Z(n8299) );
  NAND2_X1 U9959 ( .A1(n8300), .A2(n8299), .ZN(n8305) );
  NAND3_X1 U9960 ( .A1(n8305), .A2(n8301), .A3(n8306), .ZN(n8302) );
  NAND3_X1 U9961 ( .A1(n8305), .A2(n8304), .A3(n8303), .ZN(n8307) );
  INV_X1 U9962 ( .A(n8308), .ZN(n8422) );
  MUX2_X1 U9963 ( .A(n8310), .B(n8309), .S(n8383), .Z(n8311) );
  MUX2_X1 U9964 ( .A(n8314), .B(n8313), .S(n8383), .Z(n8315) );
  NOR2_X1 U9965 ( .A1(n8425), .A2(n8315), .ZN(n8316) );
  NAND3_X1 U9966 ( .A1(n8321), .A2(n8317), .A3(n8426), .ZN(n8319) );
  NAND3_X1 U9967 ( .A1(n8321), .A2(n8320), .A3(n8426), .ZN(n8323) );
  INV_X1 U9968 ( .A(n8874), .ZN(n8324) );
  MUX2_X1 U9969 ( .A(n8873), .B(n8324), .S(n8383), .Z(n8325) );
  NOR2_X1 U9970 ( .A1(n8878), .A2(n8325), .ZN(n8326) );
  NAND2_X1 U9971 ( .A1(n8329), .A2(n8327), .ZN(n8430) );
  NAND2_X1 U9972 ( .A1(n8430), .A2(n8399), .ZN(n8328) );
  NAND2_X1 U9973 ( .A1(n8407), .A2(n8428), .ZN(n8330) );
  OAI211_X1 U9974 ( .C1(n8333), .C2(n8330), .A(n8329), .B(n8334), .ZN(n8331)
         );
  NAND3_X1 U9975 ( .A1(n8333), .A2(n8407), .A3(n8332), .ZN(n8336) );
  NAND3_X1 U9976 ( .A1(n8336), .A2(n8335), .A3(n8334), .ZN(n8338) );
  NAND2_X1 U9977 ( .A1(n8338), .A2(n8337), .ZN(n8339) );
  MUX2_X1 U9978 ( .A(n8341), .B(n8340), .S(n8383), .Z(n8342) );
  INV_X1 U9979 ( .A(n8342), .ZN(n8343) );
  NOR2_X1 U9980 ( .A1(n8806), .A2(n8343), .ZN(n8344) );
  AND2_X1 U9981 ( .A1(n8404), .A2(n8345), .ZN(n8347) );
  MUX2_X1 U9982 ( .A(n8347), .B(n8346), .S(n8383), .Z(n8348) );
  NAND2_X1 U9983 ( .A1(n8349), .A2(n8348), .ZN(n8356) );
  NAND3_X1 U9984 ( .A1(n8356), .A2(n4826), .A3(n8401), .ZN(n8354) );
  INV_X1 U9985 ( .A(n8402), .ZN(n8355) );
  NAND3_X1 U9986 ( .A1(n8350), .A2(n8355), .A3(n8399), .ZN(n8351) );
  NOR2_X1 U9987 ( .A1(n8352), .A2(n8351), .ZN(n8353) );
  NAND3_X1 U9988 ( .A1(n8354), .A2(n8353), .A3(n8434), .ZN(n8362) );
  OAI211_X1 U9989 ( .C1(n8356), .C2(n8406), .A(n8355), .B(n8404), .ZN(n8360)
         );
  AND4_X1 U9990 ( .A1(n8358), .A2(n8357), .A3(n8383), .A4(n8401), .ZN(n8359)
         );
  NAND3_X1 U9991 ( .A1(n8360), .A2(n8359), .A3(n8434), .ZN(n8361) );
  NAND2_X1 U9992 ( .A1(n8369), .A2(n8368), .ZN(n8370) );
  INV_X1 U9993 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8469) );
  MUX2_X1 U9994 ( .A(n8536), .B(n8469), .S(n8392), .Z(n8373) );
  INV_X1 U9995 ( .A(SI_30_), .ZN(n8372) );
  NAND2_X1 U9996 ( .A1(n8373), .A2(n8372), .ZN(n8390) );
  INV_X1 U9997 ( .A(n8373), .ZN(n8374) );
  NAND2_X1 U9998 ( .A1(n8374), .A2(SI_30_), .ZN(n8375) );
  AND2_X1 U9999 ( .A1(n8390), .A2(n8375), .ZN(n8388) );
  NAND2_X1 U10000 ( .A1(n8535), .A2(n8396), .ZN(n8377) );
  OR2_X1 U10001 ( .A1(n4422), .A2(n8469), .ZN(n8376) );
  NAND2_X1 U10002 ( .A1(n8952), .A2(n8652), .ZN(n8454) );
  OAI211_X1 U10003 ( .C1(n8382), .C2(n8378), .A(n8445), .B(n8454), .ZN(n8379)
         );
  INV_X1 U10004 ( .A(n8652), .ZN(n8380) );
  NAND2_X1 U10005 ( .A1(n8751), .A2(n8380), .ZN(n8400) );
  AND2_X1 U10006 ( .A1(n8400), .A2(n8381), .ZN(n8451) );
  NAND2_X1 U10007 ( .A1(n8389), .A2(n8388), .ZN(n8391) );
  MUX2_X1 U10008 ( .A(n7523), .B(n6747), .S(n8392), .Z(n8393) );
  XNOR2_X1 U10009 ( .A(n8393), .B(SI_31_), .ZN(n8394) );
  NAND2_X1 U10010 ( .A1(n9177), .A2(n8396), .ZN(n8398) );
  OR2_X1 U10011 ( .A1(n4421), .A2(n6747), .ZN(n8397) );
  INV_X1 U10012 ( .A(n8748), .ZN(n8455) );
  NAND2_X1 U10013 ( .A1(n8399), .A2(n5754), .ZN(n8453) );
  INV_X1 U10014 ( .A(n8454), .ZN(n8456) );
  INV_X1 U10015 ( .A(n8400), .ZN(n8440) );
  INV_X1 U10016 ( .A(n8401), .ZN(n8403) );
  INV_X1 U10017 ( .A(n8404), .ZN(n8405) );
  NOR2_X1 U10018 ( .A1(n8406), .A2(n8405), .ZN(n8795) );
  INV_X1 U10019 ( .A(n8816), .ZN(n8819) );
  INV_X1 U10020 ( .A(n8844), .ZN(n8846) );
  INV_X1 U10021 ( .A(n8407), .ZN(n8431) );
  INV_X1 U10022 ( .A(n8886), .ZN(n8887) );
  NOR3_X1 U10023 ( .A1(n8410), .A2(n8409), .A3(n8408), .ZN(n8413) );
  NAND4_X1 U10024 ( .A1(n8413), .A2(n4543), .A3(n8412), .A4(n8411), .ZN(n8417)
         );
  NOR4_X1 U10025 ( .A1(n8417), .A2(n8416), .A3(n8415), .A4(n8414), .ZN(n8421)
         );
  NAND4_X1 U10026 ( .A1(n8421), .A2(n8420), .A3(n8419), .A4(n4835), .ZN(n8424)
         );
  NOR4_X1 U10027 ( .A1(n8425), .A2(n8424), .A3(n8423), .A4(n8422), .ZN(n8427)
         );
  NAND4_X1 U10028 ( .A1(n8428), .A2(n8887), .A3(n8427), .A4(n8426), .ZN(n8429)
         );
  NOR4_X1 U10029 ( .A1(n8846), .A2(n8431), .A3(n8430), .A4(n8429), .ZN(n8432)
         );
  NAND4_X1 U10030 ( .A1(n8795), .A2(n8819), .A3(n8833), .A4(n8432), .ZN(n8433)
         );
  NOR4_X1 U10031 ( .A1(n8771), .A2(n8780), .A3(n8433), .A4(n8806), .ZN(n8435)
         );
  NAND4_X1 U10032 ( .A1(n8437), .A2(n8436), .A3(n8435), .A4(n8434), .ZN(n8438)
         );
  NOR4_X1 U10033 ( .A1(n8456), .A2(n8440), .A3(n8439), .A4(n8438), .ZN(n8443)
         );
  INV_X1 U10034 ( .A(n8441), .ZN(n8442) );
  AOI211_X1 U10035 ( .C1(n8443), .C2(n8442), .A(n5753), .B(n5754), .ZN(n8444)
         );
  NAND2_X1 U10036 ( .A1(n8446), .A2(n8445), .ZN(n8452) );
  INV_X1 U10037 ( .A(n8447), .ZN(n8450) );
  NAND2_X1 U10038 ( .A1(n8452), .A2(n5020), .ZN(n8459) );
  NOR3_X1 U10039 ( .A1(n8454), .A2(n8453), .A3(n8748), .ZN(n8457) );
  OAI22_X1 U10040 ( .A1(n8457), .A2(n8946), .B1(n8456), .B2(n8455), .ZN(n8458)
         );
  NAND3_X1 U10041 ( .A1(n8462), .A2(n8461), .A3(n8460), .ZN(n8463) );
  OAI211_X1 U10042 ( .C1(n8464), .C2(n8466), .A(n8463), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8465) );
  OAI21_X1 U10043 ( .B1(n8467), .B2(n8466), .A(n8465), .ZN(P2_U3296) );
  INV_X1 U10044 ( .A(n8535), .ZN(n8470) );
  OAI222_X1 U10045 ( .A1(n4428), .A2(n8536), .B1(n8472), .B2(n8470), .C1(n8468), .C2(P1_U3086), .ZN(P1_U3325) );
  OAI222_X1 U10046 ( .A1(n9024), .A2(n8470), .B1(n5102), .B2(P2_U3151), .C1(
        n8469), .C2(n8549), .ZN(P2_U3265) );
  OAI222_X1 U10047 ( .A1(n4428), .A2(n8473), .B1(n8472), .B2(n8471), .C1(
        P1_U3086), .C2(n6284), .ZN(P1_U3336) );
  INV_X1 U10048 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n8489) );
  AOI21_X1 U10049 ( .B1(n10246), .B2(n8475), .A(n8474), .ZN(n8480) );
  AOI21_X1 U10050 ( .B1(n8478), .B2(n8477), .A(n8476), .ZN(n8479) );
  OAI22_X1 U10051 ( .A1(n8480), .A2(n10147), .B1(n8479), .B2(n10156), .ZN(
        n8481) );
  AOI211_X1 U10052 ( .C1(n8483), .C2(n8699), .A(n8482), .B(n8481), .ZN(n8488)
         );
  OAI211_X1 U10053 ( .C1(n8486), .C2(n8485), .A(n8484), .B(n10152), .ZN(n8487)
         );
  OAI211_X1 U10054 ( .C1(n8682), .C2(n8489), .A(n8488), .B(n8487), .ZN(
        P2_U3187) );
  OAI222_X1 U10055 ( .A1(n8492), .A2(n4428), .B1(P1_U3086), .B2(n8491), .C1(
        n9834), .C2(n8490), .ZN(P1_U3351) );
  NAND2_X1 U10056 ( .A1(n9759), .A2(n9606), .ZN(n9598) );
  OR2_X1 U10057 ( .A1(n9785), .A2(n9129), .ZN(n9259) );
  NAND2_X1 U10058 ( .A1(n9785), .A2(n9129), .ZN(n9258) );
  NAND2_X1 U10059 ( .A1(n9259), .A2(n9258), .ZN(n9314) );
  INV_X1 U10060 ( .A(n9314), .ZN(n9680) );
  OR2_X1 U10061 ( .A1(n9790), .A2(n9256), .ZN(n9678) );
  NAND2_X1 U10062 ( .A1(n9680), .A2(n9678), .ZN(n8498) );
  OR2_X1 U10063 ( .A1(n9794), .A2(n9116), .ZN(n9238) );
  INV_X1 U10064 ( .A(n9435), .ZN(n8496) );
  OR2_X1 U10065 ( .A1(n9800), .A2(n8496), .ZN(n9706) );
  NAND2_X1 U10066 ( .A1(n9238), .A2(n9706), .ZN(n9347) );
  INV_X1 U10067 ( .A(n9243), .ZN(n8493) );
  NOR2_X1 U10068 ( .A1(n9293), .A2(n8493), .ZN(n8494) );
  OR2_X1 U10069 ( .A1(n9806), .A2(n9115), .ZN(n9390) );
  NAND2_X1 U10070 ( .A1(n9806), .A2(n9115), .ZN(n9392) );
  INV_X1 U10071 ( .A(n9392), .ZN(n9246) );
  AND2_X1 U10072 ( .A1(n9800), .A2(n8496), .ZN(n9235) );
  NAND2_X1 U10073 ( .A1(n9238), .A2(n9235), .ZN(n8497) );
  NAND2_X1 U10074 ( .A1(n9794), .A2(n9116), .ZN(n9237) );
  AND2_X1 U10075 ( .A1(n8497), .A2(n9237), .ZN(n9338) );
  XNOR2_X1 U10076 ( .A(n9790), .B(n9256), .ZN(n9694) );
  INV_X1 U10077 ( .A(n9432), .ZN(n8499) );
  OR2_X1 U10078 ( .A1(n9780), .A2(n8499), .ZN(n9333) );
  NAND2_X1 U10079 ( .A1(n9780), .A2(n8499), .ZN(n9340) );
  NAND2_X1 U10080 ( .A1(n9333), .A2(n9340), .ZN(n9666) );
  INV_X1 U10081 ( .A(n9333), .ZN(n8500) );
  NAND2_X1 U10082 ( .A1(n9776), .A2(n9104), .ZN(n9341) );
  NAND2_X1 U10083 ( .A1(n9336), .A2(n9341), .ZN(n9643) );
  XNOR2_X1 U10084 ( .A(n9771), .B(n9430), .ZN(n9632) );
  INV_X1 U10085 ( .A(n9430), .ZN(n9261) );
  INV_X1 U10086 ( .A(n9429), .ZN(n8501) );
  NAND2_X1 U10087 ( .A1(n9766), .A2(n8501), .ZN(n9267) );
  NAND2_X1 U10088 ( .A1(n8502), .A2(n9317), .ZN(n9599) );
  OAI21_X1 U10089 ( .B1(n9317), .B2(n8502), .A(n9599), .ZN(n8504) );
  AOI21_X1 U10090 ( .B1(n8504), .B2(n9980), .A(n8503), .ZN(n9762) );
  NAND2_X1 U10091 ( .A1(n9742), .A2(n9115), .ZN(n8508) );
  NAND2_X1 U10092 ( .A1(n9705), .A2(n9116), .ZN(n8509) );
  NAND2_X1 U10093 ( .A1(n9700), .A2(n8509), .ZN(n8511) );
  NAND2_X1 U10094 ( .A1(n9794), .A2(n9434), .ZN(n8510) );
  NAND2_X1 U10095 ( .A1(n8511), .A2(n8510), .ZN(n9687) );
  NOR2_X1 U10096 ( .A1(n9691), .A2(n9256), .ZN(n8513) );
  NAND2_X1 U10097 ( .A1(n9691), .A2(n9256), .ZN(n8512) );
  NOR2_X1 U10098 ( .A1(n9771), .A2(n9430), .ZN(n8516) );
  NAND2_X1 U10099 ( .A1(n9771), .A2(n9430), .ZN(n8515) );
  INV_X1 U10100 ( .A(n9317), .ZN(n8518) );
  NAND2_X1 U10101 ( .A1(n8519), .A2(n9317), .ZN(n8520) );
  INV_X1 U10102 ( .A(n9780), .ZN(n9663) );
  OAI211_X1 U10103 ( .C1(n9607), .C2(n4454), .A(n9985), .B(n9611), .ZN(n9760)
         );
  NAND2_X1 U10104 ( .A1(n9947), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n8521) );
  OAI21_X1 U10105 ( .B1(n8523), .B2(n8522), .A(n8521), .ZN(n8524) );
  AOI21_X1 U10106 ( .B1(n9759), .B2(n9981), .A(n8524), .ZN(n8525) );
  OAI21_X1 U10107 ( .B1(n9760), .B2(n9987), .A(n8525), .ZN(n8526) );
  AOI21_X1 U10108 ( .B1(n9758), .B2(n9968), .A(n8526), .ZN(n8527) );
  OAI21_X1 U10109 ( .B1(n9992), .B2(n9762), .A(n8527), .ZN(P1_U3265) );
  AOI21_X1 U10110 ( .B1(n8529), .B2(n8528), .A(n4452), .ZN(n8534) );
  AOI22_X1 U10111 ( .A1(n8807), .A2(n8632), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8531) );
  NAND2_X1 U10112 ( .A1(n8641), .A2(n8837), .ZN(n8530) );
  OAI211_X1 U10113 ( .C1(n8865), .C2(n8635), .A(n8531), .B(n8530), .ZN(n8532)
         );
  AOI21_X1 U10114 ( .B1(n8836), .B2(n8648), .A(n8532), .ZN(n8533) );
  OAI21_X1 U10115 ( .B1(n8534), .B2(n8650), .A(n8533), .ZN(P2_U3173) );
  NAND2_X1 U10116 ( .A1(n8535), .A2(n9176), .ZN(n8538) );
  OR2_X1 U10117 ( .A1(n6003), .A2(n8536), .ZN(n8537) );
  NAND2_X1 U10118 ( .A1(n8220), .A2(n9176), .ZN(n8541) );
  OR2_X1 U10119 ( .A1(n6003), .A2(n8539), .ZN(n8540) );
  INV_X1 U10120 ( .A(n5012), .ZN(n8543) );
  INV_X1 U10121 ( .A(n9591), .ZN(n8542) );
  OAI211_X1 U10122 ( .C1(n9751), .C2(n8543), .A(n8542), .B(n9985), .ZN(n9750)
         );
  AND2_X1 U10123 ( .A1(n8544), .A2(P1_B_REG_SCAN_IN), .ZN(n8545) );
  NOR2_X1 U10124 ( .A1(n9128), .A2(n8545), .ZN(n9602) );
  NAND2_X1 U10125 ( .A1(n9602), .A2(n9289), .ZN(n9749) );
  NOR2_X1 U10126 ( .A1(n9947), .A2(n9749), .ZN(n9594) );
  AND2_X1 U10127 ( .A1(n9992), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8546) );
  NOR2_X1 U10128 ( .A1(n9594), .A2(n8546), .ZN(n8548) );
  NAND2_X1 U10129 ( .A1(n9354), .A2(n9981), .ZN(n8547) );
  OAI211_X1 U10130 ( .C1(n9750), .C2(n9987), .A(n8548), .B(n8547), .ZN(
        P1_U3264) );
  OAI222_X1 U10131 ( .A1(n9024), .A2(n8552), .B1(n5750), .B2(P2_U3151), .C1(
        n8550), .C2(n8549), .ZN(P2_U3274) );
  OAI211_X1 U10132 ( .C1(n8555), .C2(n8554), .A(n8553), .B(n8616), .ZN(n8561)
         );
  INV_X1 U10133 ( .A(n8556), .ZN(n8763) );
  AOI22_X1 U10134 ( .A1(n4713), .A2(n8640), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8557) );
  OAI21_X1 U10135 ( .B1(n8763), .B2(n8558), .A(n8557), .ZN(n8559) );
  AOI21_X1 U10136 ( .B1(n8632), .B2(n8654), .A(n8559), .ZN(n8560) );
  OAI211_X1 U10137 ( .C1(n5749), .C2(n8592), .A(n8561), .B(n8560), .ZN(
        P2_U3154) );
  XNOR2_X1 U10138 ( .A(n8597), .B(n8596), .ZN(n8598) );
  XNOR2_X1 U10139 ( .A(n8598), .B(n8785), .ZN(n8566) );
  AOI22_X1 U10140 ( .A1(n8657), .A2(n8640), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8563) );
  NAND2_X1 U10141 ( .A1(n8641), .A2(n8800), .ZN(n8562) );
  OAI211_X1 U10142 ( .C1(n8797), .C2(n8645), .A(n8563), .B(n8562), .ZN(n8564)
         );
  AOI21_X1 U10143 ( .B1(n8801), .B2(n8648), .A(n8564), .ZN(n8565) );
  OAI21_X1 U10144 ( .B1(n8566), .B2(n8650), .A(n8565), .ZN(P2_U3156) );
  XNOR2_X1 U10145 ( .A(n8567), .B(n8865), .ZN(n8568) );
  XNOR2_X1 U10146 ( .A(n8569), .B(n8568), .ZN(n8575) );
  NAND2_X1 U10147 ( .A1(n8879), .A2(n8640), .ZN(n8571) );
  OAI211_X1 U10148 ( .C1(n8822), .C2(n8645), .A(n8571), .B(n8570), .ZN(n8572)
         );
  AOI21_X1 U10149 ( .B1(n8851), .B2(n8641), .A(n8572), .ZN(n8574) );
  NAND2_X1 U10150 ( .A1(n8993), .A2(n8648), .ZN(n8573) );
  OAI211_X1 U10151 ( .C1(n8575), .C2(n8650), .A(n8574), .B(n8573), .ZN(
        P2_U3159) );
  INV_X1 U10152 ( .A(n8826), .ZN(n8982) );
  INV_X1 U10153 ( .A(n8576), .ZN(n8578) );
  NOR3_X1 U10154 ( .A1(n4452), .A2(n8578), .A3(n8577), .ZN(n8581) );
  OAI21_X1 U10155 ( .B1(n8581), .B2(n4488), .A(n8616), .ZN(n8585) );
  AOI22_X1 U10156 ( .A1(n8657), .A2(n8632), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8582) );
  OAI21_X1 U10157 ( .B1(n8822), .B2(n8635), .A(n8582), .ZN(n8583) );
  AOI21_X1 U10158 ( .B1(n8825), .B2(n8641), .A(n8583), .ZN(n8584) );
  OAI211_X1 U10159 ( .C1(n8982), .C2(n8592), .A(n8585), .B(n8584), .ZN(
        P2_U3163) );
  XNOR2_X1 U10160 ( .A(n8587), .B(n8586), .ZN(n8594) );
  INV_X1 U10161 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8588) );
  OAI22_X1 U10162 ( .A1(n8797), .A2(n8635), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8588), .ZN(n8589) );
  AOI21_X1 U10163 ( .B1(n4713), .B2(n8632), .A(n8589), .ZN(n8591) );
  NAND2_X1 U10164 ( .A1(n8641), .A2(n8776), .ZN(n8590) );
  OAI211_X1 U10165 ( .C1(n8960), .C2(n8592), .A(n8591), .B(n8590), .ZN(n8593)
         );
  AOI21_X1 U10166 ( .B1(n8594), .B2(n8616), .A(n8593), .ZN(n8595) );
  INV_X1 U10167 ( .A(n8595), .ZN(P2_U3165) );
  OAI22_X1 U10168 ( .A1(n8598), .A2(n8808), .B1(n8597), .B2(n8596), .ZN(n8601)
         );
  XNOR2_X1 U10169 ( .A(n8599), .B(n8797), .ZN(n8600) );
  XNOR2_X1 U10170 ( .A(n8601), .B(n8600), .ZN(n8606) );
  AOI22_X1 U10171 ( .A1(n8783), .A2(n8632), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8603) );
  NAND2_X1 U10172 ( .A1(n8641), .A2(n8790), .ZN(n8602) );
  OAI211_X1 U10173 ( .C1(n8785), .C2(n8635), .A(n8603), .B(n8602), .ZN(n8604)
         );
  AOI21_X1 U10174 ( .B1(n8966), .B2(n8648), .A(n8604), .ZN(n8605) );
  OAI21_X1 U10175 ( .B1(n8606), .B2(n8650), .A(n8605), .ZN(P2_U3169) );
  XNOR2_X1 U10176 ( .A(n8608), .B(n8821), .ZN(n8609) );
  XNOR2_X1 U10177 ( .A(n8607), .B(n8609), .ZN(n8614) );
  AOI22_X1 U10178 ( .A1(n8807), .A2(n8640), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8611) );
  NAND2_X1 U10179 ( .A1(n8641), .A2(n8811), .ZN(n8610) );
  OAI211_X1 U10180 ( .C1(n8785), .C2(n8645), .A(n8611), .B(n8610), .ZN(n8612)
         );
  AOI21_X1 U10181 ( .B1(n8977), .B2(n8648), .A(n8612), .ZN(n8613) );
  OAI21_X1 U10182 ( .B1(n8614), .B2(n8650), .A(n8613), .ZN(P2_U3175) );
  OAI211_X1 U10183 ( .C1(n8615), .C2(n8618), .A(n8617), .B(n8616), .ZN(n8629)
         );
  OAI21_X1 U10184 ( .B1(n8620), .B2(n8635), .A(n8619), .ZN(n8623) );
  NOR2_X1 U10185 ( .A1(n8621), .A2(n8645), .ZN(n8622) );
  NOR2_X1 U10186 ( .A1(n8623), .A2(n8622), .ZN(n8628) );
  NAND2_X1 U10187 ( .A1(n8624), .A2(n8648), .ZN(n8627) );
  NAND2_X1 U10188 ( .A1(n8641), .A2(n8625), .ZN(n8626) );
  NAND4_X1 U10189 ( .A1(n8629), .A2(n8628), .A3(n8627), .A4(n8626), .ZN(
        P2_U3176) );
  XOR2_X1 U10190 ( .A(n8631), .B(n8630), .Z(n8638) );
  AOI22_X1 U10191 ( .A1(n8658), .A2(n8632), .B1(P2_REG3_REG_18__SCAN_IN), .B2(
        P2_U3151), .ZN(n8634) );
  NAND2_X1 U10192 ( .A1(n8641), .A2(n8867), .ZN(n8633) );
  OAI211_X1 U10193 ( .C1(n8866), .C2(n8635), .A(n8634), .B(n8633), .ZN(n8636)
         );
  AOI21_X1 U10194 ( .B1(n8930), .B2(n8648), .A(n8636), .ZN(n8637) );
  OAI21_X1 U10195 ( .B1(n8638), .B2(n8650), .A(n8637), .ZN(P2_U3178) );
  XNOR2_X1 U10196 ( .A(n8639), .B(n4713), .ZN(n8651) );
  AOI22_X1 U10197 ( .A1(n8783), .A2(n8640), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8644) );
  NAND2_X1 U10198 ( .A1(n8642), .A2(n8641), .ZN(n8643) );
  OAI211_X1 U10199 ( .C1(n8646), .C2(n8645), .A(n8644), .B(n8643), .ZN(n8647)
         );
  AOI21_X1 U10200 ( .B1(n8955), .B2(n8648), .A(n8647), .ZN(n8649) );
  OAI21_X1 U10201 ( .B1(n8651), .B2(n8650), .A(n8649), .ZN(P2_U3180) );
  MUX2_X1 U10202 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8652), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10203 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8653), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10204 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8654), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U10205 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8655), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10206 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n4713), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10207 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8783), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10208 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8656), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10209 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8808), .S(P2_U3893), .Z(
        P2_U3514) );
  MUX2_X1 U10210 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8657), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10211 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8807), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10212 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8848), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10213 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8658), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10214 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8879), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10215 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8890), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10216 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8880), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U10217 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8892), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10218 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8659), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U10219 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n5372), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U10220 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8660), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U10221 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8661), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U10222 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8662), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U10223 ( .A(n8663), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8732), .Z(
        P2_U3500) );
  MUX2_X1 U10224 ( .A(n8664), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8732), .Z(
        P2_U3499) );
  MUX2_X1 U10225 ( .A(n8665), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8732), .Z(
        P2_U3498) );
  MUX2_X1 U10226 ( .A(n8666), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8732), .Z(
        P2_U3497) );
  MUX2_X1 U10227 ( .A(n8667), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8732), .Z(
        P2_U3496) );
  MUX2_X1 U10228 ( .A(n8668), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8732), .Z(
        P2_U3495) );
  MUX2_X1 U10229 ( .A(n8669), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8732), .Z(
        P2_U3494) );
  MUX2_X1 U10230 ( .A(n8670), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8732), .Z(
        P2_U3493) );
  MUX2_X1 U10231 ( .A(n5135), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8732), .Z(
        P2_U3492) );
  MUX2_X1 U10232 ( .A(n8671), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8732), .Z(
        P2_U3491) );
  AOI21_X1 U10233 ( .B1(n8674), .B2(n8673), .A(n8672), .ZN(n8690) );
  OAI21_X1 U10234 ( .B1(n8677), .B2(n8676), .A(n8675), .ZN(n8688) );
  AOI21_X1 U10235 ( .B1(n8699), .B2(n8679), .A(n8678), .ZN(n8680) );
  OAI21_X1 U10236 ( .B1(n8682), .B2(n8681), .A(n8680), .ZN(n8687) );
  AOI21_X1 U10237 ( .B1(n8942), .B2(n8684), .A(n8683), .ZN(n8685) );
  NOR2_X1 U10238 ( .A1(n8685), .A2(n10147), .ZN(n8686) );
  AOI211_X1 U10239 ( .C1(n10152), .C2(n8688), .A(n8687), .B(n8686), .ZN(n8689)
         );
  OAI21_X1 U10240 ( .B1(n8690), .B2(n10156), .A(n8689), .ZN(P2_U3197) );
  AOI21_X1 U10241 ( .B1(n8693), .B2(n8692), .A(n8691), .ZN(n8709) );
  OAI21_X1 U10242 ( .B1(n8696), .B2(n8695), .A(n8694), .ZN(n8707) );
  AOI21_X1 U10243 ( .B1(n8699), .B2(n8698), .A(n8697), .ZN(n8701) );
  NAND2_X1 U10244 ( .A1(n10141), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n8700) );
  NAND2_X1 U10245 ( .A1(n8701), .A2(n8700), .ZN(n8706) );
  AOI21_X1 U10246 ( .B1(n4465), .B2(n8703), .A(n8702), .ZN(n8704) );
  NOR2_X1 U10247 ( .A1(n8704), .A2(n10156), .ZN(n8705) );
  AOI211_X1 U10248 ( .C1(n10152), .C2(n8707), .A(n8706), .B(n8705), .ZN(n8708)
         );
  OAI21_X1 U10249 ( .B1(n8709), .B2(n10147), .A(n8708), .ZN(P2_U3198) );
  AOI21_X1 U10250 ( .B1(n8933), .B2(n8711), .A(n8710), .ZN(n8722) );
  OR2_X1 U10251 ( .A1(n8713), .A2(n8712), .ZN(n8715) );
  AOI21_X1 U10252 ( .B1(n8715), .B2(n8714), .A(n8730), .ZN(n8721) );
  AND2_X1 U10253 ( .A1(n8716), .A2(n8882), .ZN(n8717) );
  AOI21_X1 U10254 ( .B1(n8725), .B2(n8724), .A(n8723), .ZN(n8746) );
  INV_X1 U10255 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8726) );
  NOR2_X1 U10256 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8726), .ZN(n8738) );
  INV_X1 U10257 ( .A(n8727), .ZN(n8729) );
  AND2_X1 U10258 ( .A1(n8729), .A2(n8728), .ZN(n8731) );
  NOR2_X1 U10259 ( .A1(n8731), .A2(n8730), .ZN(n8736) );
  INV_X1 U10260 ( .A(n8731), .ZN(n8733) );
  OAI21_X1 U10261 ( .B1(n8733), .B2(n8732), .A(n10162), .ZN(n8735) );
  MUX2_X1 U10262 ( .A(n8736), .B(n8735), .S(n8734), .Z(n8737) );
  AOI211_X1 U10263 ( .C1(n10141), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n8738), .B(
        n8737), .ZN(n8745) );
  AND2_X1 U10264 ( .A1(n8740), .A2(n8739), .ZN(n8742) );
  OAI21_X1 U10265 ( .B1(n8743), .B2(n8742), .A(n8741), .ZN(n8744) );
  OAI211_X1 U10266 ( .C1(n8746), .C2(n10147), .A(n8745), .B(n8744), .ZN(
        P2_U3200) );
  AND2_X1 U10267 ( .A1(n8748), .A2(n8747), .ZN(n8947) );
  NOR3_X1 U10268 ( .A1(n8749), .A2(P2_REG3_REG_28__SCAN_IN), .A3(n10165), .ZN(
        n8757) );
  AOI21_X1 U10269 ( .B1(n8947), .B2(n8895), .A(n8757), .ZN(n8752) );
  NAND2_X1 U10270 ( .A1(n10176), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8750) );
  OAI211_X1 U10271 ( .C1(n8448), .C2(n8839), .A(n8752), .B(n8750), .ZN(
        P2_U3202) );
  NAND2_X1 U10272 ( .A1(n8751), .A2(n8898), .ZN(n8753) );
  OAI211_X1 U10273 ( .C1(n8895), .C2(n8754), .A(n8753), .B(n8752), .ZN(
        P2_U3203) );
  NAND2_X1 U10274 ( .A1(n8755), .A2(n8895), .ZN(n8759) );
  NOR2_X1 U10275 ( .A1(n8233), .A2(n8839), .ZN(n8756) );
  AOI211_X1 U10276 ( .C1(n10176), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8757), .B(
        n8756), .ZN(n8758) );
  OAI211_X1 U10277 ( .C1(n8761), .C2(n8760), .A(n8759), .B(n8758), .ZN(
        P2_U3204) );
  INV_X1 U10278 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8762) );
  OAI22_X1 U10279 ( .A1(n8763), .A2(n10165), .B1(n8895), .B2(n8762), .ZN(n8764) );
  AOI21_X1 U10280 ( .B1(n8765), .B2(n8898), .A(n8764), .ZN(n8768) );
  NAND3_X1 U10281 ( .A1(n8766), .A2(n5715), .A3(n5733), .ZN(n8767) );
  OAI211_X1 U10282 ( .C1(n8769), .C2(n10176), .A(n8768), .B(n8767), .ZN(
        P2_U3206) );
  XOR2_X1 U10283 ( .A(n8770), .B(n8771), .Z(n8961) );
  XOR2_X1 U10284 ( .A(n8772), .B(n8771), .Z(n8773) );
  OAI222_X1 U10285 ( .A1(n5626), .A2(n8797), .B1(n10171), .B2(n8774), .C1(
        n5628), .C2(n8773), .ZN(n8959) );
  NOR2_X1 U10286 ( .A1(n8960), .A2(n10167), .ZN(n8775) );
  OAI21_X1 U10287 ( .B1(n8959), .B2(n8775), .A(n10174), .ZN(n8778) );
  AOI22_X1 U10288 ( .A1(n8897), .A2(n8776), .B1(n10176), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n8777) );
  OAI211_X1 U10289 ( .C1(n8961), .C2(n8901), .A(n8778), .B(n8777), .ZN(
        P2_U3208) );
  XNOR2_X1 U10290 ( .A(n8779), .B(n8780), .ZN(n8969) );
  INV_X1 U10291 ( .A(n8966), .ZN(n8788) );
  INV_X1 U10292 ( .A(n8780), .ZN(n8781) );
  XNOR2_X1 U10293 ( .A(n8782), .B(n8781), .ZN(n8787) );
  NAND2_X1 U10294 ( .A1(n8783), .A2(n8889), .ZN(n8784) );
  OAI21_X1 U10295 ( .B1(n8785), .B2(n5626), .A(n8784), .ZN(n8786) );
  AOI21_X1 U10296 ( .B1(n8787), .B2(n8894), .A(n8786), .ZN(n8965) );
  OAI21_X1 U10297 ( .B1(n8788), .B2(n10167), .A(n8965), .ZN(n8789) );
  NAND2_X1 U10298 ( .A1(n8789), .A2(n8895), .ZN(n8792) );
  AOI22_X1 U10299 ( .A1(n10176), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8897), 
        .B2(n8790), .ZN(n8791) );
  OAI211_X1 U10300 ( .C1(n8969), .C2(n8901), .A(n8792), .B(n8791), .ZN(
        P2_U3209) );
  XNOR2_X1 U10301 ( .A(n8793), .B(n8795), .ZN(n8972) );
  XNOR2_X1 U10302 ( .A(n8794), .B(n8795), .ZN(n8796) );
  OAI222_X1 U10303 ( .A1(n5626), .A2(n8821), .B1(n10171), .B2(n8797), .C1(
        n5628), .C2(n8796), .ZN(n8970) );
  INV_X1 U10304 ( .A(n8970), .ZN(n8798) );
  MUX2_X1 U10305 ( .A(n8799), .B(n8798), .S(n8895), .Z(n8803) );
  AOI22_X1 U10306 ( .A1(n8801), .A2(n8898), .B1(n8897), .B2(n8800), .ZN(n8802)
         );
  OAI211_X1 U10307 ( .C1(n8972), .C2(n8901), .A(n8803), .B(n8802), .ZN(
        P2_U3210) );
  XOR2_X1 U10308 ( .A(n8804), .B(n8806), .Z(n8980) );
  INV_X1 U10309 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8810) );
  XNOR2_X1 U10310 ( .A(n8805), .B(n8806), .ZN(n8809) );
  AOI222_X1 U10311 ( .A1(n8894), .A2(n8809), .B1(n8808), .B2(n8889), .C1(n8807), .C2(n8891), .ZN(n8975) );
  MUX2_X1 U10312 ( .A(n8810), .B(n8975), .S(n8895), .Z(n8813) );
  AOI22_X1 U10313 ( .A1(n8977), .A2(n8898), .B1(n8897), .B2(n8811), .ZN(n8812)
         );
  OAI211_X1 U10314 ( .C1(n8980), .C2(n8901), .A(n8813), .B(n8812), .ZN(
        P2_U3211) );
  NAND2_X1 U10315 ( .A1(n8815), .A2(n8814), .ZN(n8817) );
  XNOR2_X1 U10316 ( .A(n8817), .B(n8816), .ZN(n8983) );
  INV_X1 U10317 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8824) );
  XNOR2_X1 U10318 ( .A(n8818), .B(n8819), .ZN(n8820) );
  OAI222_X1 U10319 ( .A1(n5626), .A2(n8822), .B1(n10171), .B2(n8821), .C1(
        n5628), .C2(n8820), .ZN(n8981) );
  INV_X1 U10320 ( .A(n8981), .ZN(n8823) );
  MUX2_X1 U10321 ( .A(n8824), .B(n8823), .S(n8895), .Z(n8828) );
  AOI22_X1 U10322 ( .A1(n8826), .A2(n8898), .B1(n8897), .B2(n8825), .ZN(n8827)
         );
  OAI211_X1 U10323 ( .C1(n8983), .C2(n8901), .A(n8828), .B(n8827), .ZN(
        P2_U3212) );
  XNOR2_X1 U10324 ( .A(n8829), .B(n8833), .ZN(n8922) );
  INV_X1 U10325 ( .A(n8922), .ZN(n8842) );
  INV_X1 U10326 ( .A(n8830), .ZN(n8831) );
  AOI21_X1 U10327 ( .B1(n8833), .B2(n8832), .A(n8831), .ZN(n8834) );
  OAI222_X1 U10328 ( .A1(n10171), .A2(n8835), .B1(n5626), .B2(n8865), .C1(
        n5628), .C2(n8834), .ZN(n8921) );
  INV_X1 U10329 ( .A(n8836), .ZN(n8990) );
  AOI22_X1 U10330 ( .A1(n10176), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8897), 
        .B2(n8837), .ZN(n8838) );
  OAI21_X1 U10331 ( .B1(n8990), .B2(n8839), .A(n8838), .ZN(n8840) );
  AOI21_X1 U10332 ( .B1(n8921), .B2(n8895), .A(n8840), .ZN(n8841) );
  OAI21_X1 U10333 ( .B1(n8842), .B2(n8901), .A(n8841), .ZN(P2_U3213) );
  OAI21_X1 U10334 ( .B1(n8845), .B2(n8844), .A(n8843), .ZN(n8996) );
  XNOR2_X1 U10335 ( .A(n8847), .B(n8846), .ZN(n8849) );
  AOI222_X1 U10336 ( .A1(n8894), .A2(n8849), .B1(n8848), .B2(n8889), .C1(n8879), .C2(n8891), .ZN(n8991) );
  MUX2_X1 U10337 ( .A(n8850), .B(n8991), .S(n8895), .Z(n8853) );
  AOI22_X1 U10338 ( .A1(n8993), .A2(n8898), .B1(n8897), .B2(n8851), .ZN(n8852)
         );
  OAI211_X1 U10339 ( .C1(n8901), .C2(n8996), .A(n8853), .B(n8852), .ZN(
        P2_U3214) );
  OR2_X1 U10340 ( .A1(n8854), .A2(n8855), .ZN(n8857) );
  INV_X1 U10341 ( .A(n8862), .ZN(n8861) );
  AND2_X1 U10342 ( .A1(n8859), .A2(n8858), .ZN(n8860) );
  OAI21_X1 U10343 ( .B1(n5015), .B2(n8861), .A(n8860), .ZN(n9000) );
  XNOR2_X1 U10344 ( .A(n8863), .B(n8862), .ZN(n8864) );
  OAI222_X1 U10345 ( .A1(n5626), .A2(n8866), .B1(n10171), .B2(n8865), .C1(
        n8864), .C2(n5628), .ZN(n8929) );
  NAND2_X1 U10346 ( .A1(n8929), .A2(n8895), .ZN(n8872) );
  INV_X1 U10347 ( .A(n8867), .ZN(n8868) );
  OAI22_X1 U10348 ( .A1(n10174), .A2(n8869), .B1(n8868), .B2(n10165), .ZN(
        n8870) );
  AOI21_X1 U10349 ( .B1(n8930), .B2(n8898), .A(n8870), .ZN(n8871) );
  OAI211_X1 U10350 ( .C1(n9000), .C2(n8901), .A(n8872), .B(n8871), .ZN(
        P2_U3215) );
  OR2_X1 U10351 ( .A1(n8854), .A2(n8873), .ZN(n8875) );
  NAND2_X1 U10352 ( .A1(n8875), .A2(n8874), .ZN(n8876) );
  XOR2_X1 U10353 ( .A(n8878), .B(n8876), .Z(n9006) );
  XOR2_X1 U10354 ( .A(n8877), .B(n8878), .Z(n8881) );
  AOI222_X1 U10355 ( .A1(n8894), .A2(n8881), .B1(n8880), .B2(n8891), .C1(n8879), .C2(n8889), .ZN(n9001) );
  MUX2_X1 U10356 ( .A(n8882), .B(n9001), .S(n8895), .Z(n8885) );
  AOI22_X1 U10357 ( .A1(n9003), .A2(n8898), .B1(n8897), .B2(n8883), .ZN(n8884)
         );
  OAI211_X1 U10358 ( .C1(n9006), .C2(n8901), .A(n8885), .B(n8884), .ZN(
        P2_U3216) );
  XNOR2_X1 U10359 ( .A(n8854), .B(n8886), .ZN(n9013) );
  XNOR2_X1 U10360 ( .A(n8888), .B(n8887), .ZN(n8893) );
  AOI222_X1 U10361 ( .A1(n8894), .A2(n8893), .B1(n8892), .B2(n8891), .C1(n8890), .C2(n8889), .ZN(n9007) );
  MUX2_X1 U10362 ( .A(n6603), .B(n9007), .S(n8895), .Z(n8900) );
  AOI22_X1 U10363 ( .A1(n9010), .A2(n8898), .B1(n8897), .B2(n8896), .ZN(n8899)
         );
  OAI211_X1 U10364 ( .C1(n9013), .C2(n8901), .A(n8900), .B(n8899), .ZN(
        P2_U3217) );
  NAND2_X1 U10365 ( .A1(n8946), .A2(n8937), .ZN(n8902) );
  NAND2_X1 U10366 ( .A1(n8947), .A2(n10261), .ZN(n8904) );
  OAI211_X1 U10367 ( .C1(n10261), .C2(n8903), .A(n8902), .B(n8904), .ZN(
        P2_U3490) );
  NAND2_X1 U10368 ( .A1(n6692), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8905) );
  OAI211_X1 U10369 ( .C1(n8952), .C2(n8925), .A(n8905), .B(n8904), .ZN(
        P2_U3489) );
  INV_X1 U10370 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8906) );
  MUX2_X1 U10371 ( .A(n8906), .B(n8953), .S(n10261), .Z(n8908) );
  NAND2_X1 U10372 ( .A1(n8955), .A2(n8937), .ZN(n8907) );
  OAI211_X1 U10373 ( .C1(n8944), .C2(n8958), .A(n8908), .B(n8907), .ZN(
        P2_U3485) );
  MUX2_X1 U10374 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8959), .S(n10261), .Z(
        n8910) );
  OAI22_X1 U10375 ( .A1(n8961), .A2(n8944), .B1(n8960), .B2(n8925), .ZN(n8909)
         );
  OR2_X1 U10376 ( .A1(n8910), .A2(n8909), .ZN(P2_U3484) );
  MUX2_X1 U10377 ( .A(n8911), .B(n8965), .S(n10261), .Z(n8913) );
  NAND2_X1 U10378 ( .A1(n8966), .A2(n8937), .ZN(n8912) );
  OAI211_X1 U10379 ( .C1(n8944), .C2(n8969), .A(n8913), .B(n8912), .ZN(
        P2_U3483) );
  MUX2_X1 U10380 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8970), .S(n10261), .Z(
        n8915) );
  OAI22_X1 U10381 ( .A1(n8972), .A2(n8944), .B1(n8971), .B2(n8925), .ZN(n8914)
         );
  OR2_X1 U10382 ( .A1(n8915), .A2(n8914), .ZN(P2_U3482) );
  MUX2_X1 U10383 ( .A(n8916), .B(n8975), .S(n10261), .Z(n8918) );
  NAND2_X1 U10384 ( .A1(n8977), .A2(n8937), .ZN(n8917) );
  OAI211_X1 U10385 ( .C1(n8980), .C2(n8944), .A(n8918), .B(n8917), .ZN(
        P2_U3481) );
  MUX2_X1 U10386 ( .A(n8981), .B(P2_REG1_REG_21__SCAN_IN), .S(n6692), .Z(n8920) );
  OAI22_X1 U10387 ( .A1(n8983), .A2(n8944), .B1(n8982), .B2(n8925), .ZN(n8919)
         );
  OR2_X1 U10388 ( .A1(n8920), .A2(n8919), .ZN(P2_U3480) );
  INV_X1 U10389 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8923) );
  AOI21_X1 U10390 ( .B1(n10234), .B2(n8922), .A(n8921), .ZN(n8986) );
  MUX2_X1 U10391 ( .A(n8923), .B(n8986), .S(n10261), .Z(n8924) );
  OAI21_X1 U10392 ( .B1(n8990), .B2(n8925), .A(n8924), .ZN(P2_U3479) );
  INV_X1 U10393 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8926) );
  MUX2_X1 U10394 ( .A(n8926), .B(n8991), .S(n10261), .Z(n8928) );
  NAND2_X1 U10395 ( .A1(n8993), .A2(n8937), .ZN(n8927) );
  OAI211_X1 U10396 ( .C1(n8996), .C2(n8944), .A(n8928), .B(n8927), .ZN(
        P2_U3478) );
  AOI21_X1 U10397 ( .B1(n10233), .B2(n8930), .A(n8929), .ZN(n8997) );
  MUX2_X1 U10398 ( .A(n8931), .B(n8997), .S(n10261), .Z(n8932) );
  OAI21_X1 U10399 ( .B1(n8944), .B2(n9000), .A(n8932), .ZN(P2_U3477) );
  MUX2_X1 U10400 ( .A(n8933), .B(n9001), .S(n10261), .Z(n8935) );
  NAND2_X1 U10401 ( .A1(n9003), .A2(n8937), .ZN(n8934) );
  OAI211_X1 U10402 ( .C1(n9006), .C2(n8944), .A(n8935), .B(n8934), .ZN(
        P2_U3476) );
  MUX2_X1 U10403 ( .A(n8936), .B(n9007), .S(n10261), .Z(n8939) );
  NAND2_X1 U10404 ( .A1(n9010), .A2(n8937), .ZN(n8938) );
  OAI211_X1 U10405 ( .C1(n8944), .C2(n9013), .A(n8939), .B(n8938), .ZN(
        P2_U3475) );
  AOI21_X1 U10406 ( .B1(n10233), .B2(n8941), .A(n8940), .ZN(n9014) );
  MUX2_X1 U10407 ( .A(n8942), .B(n9014), .S(n10261), .Z(n8943) );
  OAI21_X1 U10408 ( .B1(n9018), .B2(n8944), .A(n8943), .ZN(P2_U3474) );
  MUX2_X1 U10409 ( .A(n8945), .B(P2_REG1_REG_0__SCAN_IN), .S(n6692), .Z(
        P2_U3459) );
  INV_X1 U10410 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8949) );
  NAND2_X1 U10411 ( .A1(n8946), .A2(n9009), .ZN(n8948) );
  NAND2_X1 U10412 ( .A1(n8947), .A2(n10238), .ZN(n8950) );
  OAI211_X1 U10413 ( .C1(n8949), .C2(n10238), .A(n8948), .B(n8950), .ZN(
        P2_U3458) );
  NAND2_X1 U10414 ( .A1(n10240), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8951) );
  OAI211_X1 U10415 ( .C1(n8952), .C2(n8989), .A(n8951), .B(n8950), .ZN(
        P2_U3457) );
  INV_X1 U10416 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8954) );
  MUX2_X1 U10417 ( .A(n8954), .B(n8953), .S(n10238), .Z(n8957) );
  NAND2_X1 U10418 ( .A1(n8955), .A2(n9009), .ZN(n8956) );
  OAI211_X1 U10419 ( .C1(n8958), .C2(n9017), .A(n8957), .B(n8956), .ZN(
        P2_U3453) );
  MUX2_X1 U10420 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8959), .S(n10238), .Z(
        n8963) );
  OAI22_X1 U10421 ( .A1(n8961), .A2(n9017), .B1(n8960), .B2(n8989), .ZN(n8962)
         );
  OR2_X1 U10422 ( .A1(n8963), .A2(n8962), .ZN(P2_U3452) );
  INV_X1 U10423 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8964) );
  MUX2_X1 U10424 ( .A(n8965), .B(n8964), .S(n10240), .Z(n8968) );
  NAND2_X1 U10425 ( .A1(n8966), .A2(n9009), .ZN(n8967) );
  OAI211_X1 U10426 ( .C1(n8969), .C2(n9017), .A(n8968), .B(n8967), .ZN(
        P2_U3451) );
  MUX2_X1 U10427 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8970), .S(n10238), .Z(
        n8974) );
  OAI22_X1 U10428 ( .A1(n8972), .A2(n9017), .B1(n8971), .B2(n8989), .ZN(n8973)
         );
  OR2_X1 U10429 ( .A1(n8974), .A2(n8973), .ZN(P2_U3450) );
  MUX2_X1 U10430 ( .A(n8976), .B(n8975), .S(n10238), .Z(n8979) );
  NAND2_X1 U10431 ( .A1(n8977), .A2(n9009), .ZN(n8978) );
  OAI211_X1 U10432 ( .C1(n8980), .C2(n9017), .A(n8979), .B(n8978), .ZN(
        P2_U3449) );
  MUX2_X1 U10433 ( .A(n8981), .B(P2_REG0_REG_21__SCAN_IN), .S(n10240), .Z(
        n8985) );
  OAI22_X1 U10434 ( .A1(n8983), .A2(n9017), .B1(n8982), .B2(n8989), .ZN(n8984)
         );
  OR2_X1 U10435 ( .A1(n8985), .A2(n8984), .ZN(P2_U3448) );
  INV_X1 U10436 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8987) );
  MUX2_X1 U10437 ( .A(n8987), .B(n8986), .S(n10238), .Z(n8988) );
  OAI21_X1 U10438 ( .B1(n8990), .B2(n8989), .A(n8988), .ZN(P2_U3447) );
  INV_X1 U10439 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8992) );
  MUX2_X1 U10440 ( .A(n8992), .B(n8991), .S(n10238), .Z(n8995) );
  NAND2_X1 U10441 ( .A1(n8993), .A2(n9009), .ZN(n8994) );
  OAI211_X1 U10442 ( .C1(n8996), .C2(n9017), .A(n8995), .B(n8994), .ZN(
        P2_U3446) );
  INV_X1 U10443 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8998) );
  MUX2_X1 U10444 ( .A(n8998), .B(n8997), .S(n10238), .Z(n8999) );
  OAI21_X1 U10445 ( .B1(n9000), .B2(n9017), .A(n8999), .ZN(P2_U3444) );
  INV_X1 U10446 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9002) );
  MUX2_X1 U10447 ( .A(n9002), .B(n9001), .S(n10238), .Z(n9005) );
  NAND2_X1 U10448 ( .A1(n9003), .A2(n9009), .ZN(n9004) );
  OAI211_X1 U10449 ( .C1(n9006), .C2(n9017), .A(n9005), .B(n9004), .ZN(
        P2_U3441) );
  INV_X1 U10450 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9008) );
  MUX2_X1 U10451 ( .A(n9008), .B(n9007), .S(n10238), .Z(n9012) );
  NAND2_X1 U10452 ( .A1(n9010), .A2(n9009), .ZN(n9011) );
  OAI211_X1 U10453 ( .C1(n9013), .C2(n9017), .A(n9012), .B(n9011), .ZN(
        P2_U3438) );
  INV_X1 U10454 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9015) );
  MUX2_X1 U10455 ( .A(n9015), .B(n9014), .S(n10238), .Z(n9016) );
  OAI21_X1 U10456 ( .B1(n9018), .B2(n9017), .A(n9016), .ZN(P2_U3435) );
  INV_X1 U10457 ( .A(n9177), .ZN(n9835) );
  NOR4_X1 U10458 ( .A1(n9019), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n9020), .ZN(n9021) );
  AOI21_X1 U10459 ( .B1(n9022), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9021), .ZN(
        n9023) );
  OAI21_X1 U10460 ( .B1(n9835), .B2(n9024), .A(n9023), .ZN(P2_U3264) );
  INV_X1 U10461 ( .A(n9025), .ZN(n9026) );
  MUX2_X1 U10462 ( .A(n9026), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  OAI21_X1 U10463 ( .B1(n9029), .B2(n9028), .A(n9027), .ZN(n9030) );
  NAND2_X1 U10464 ( .A1(n9030), .A2(n9150), .ZN(n9037) );
  INV_X1 U10465 ( .A(n9031), .ZN(n9035) );
  OAI22_X1 U10466 ( .A1(n9156), .A2(n9033), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9032), .ZN(n9034) );
  AOI21_X1 U10467 ( .B1(n9035), .B2(n9158), .A(n9034), .ZN(n9036) );
  OAI211_X1 U10468 ( .C1(n10092), .C2(n9161), .A(n9037), .B(n9036), .ZN(
        P1_U3215) );
  INV_X1 U10469 ( .A(n9038), .ZN(n9042) );
  NOR3_X1 U10470 ( .A1(n9039), .A2(n9125), .A3(n9040), .ZN(n9041) );
  OAI21_X1 U10471 ( .B1(n9042), .B2(n9041), .A(n9150), .ZN(n9049) );
  NAND2_X1 U10472 ( .A1(n9432), .A2(n9152), .ZN(n9044) );
  OR2_X1 U10473 ( .A1(n9256), .A2(n9114), .ZN(n9043) );
  NAND2_X1 U10474 ( .A1(n9044), .A2(n9043), .ZN(n9682) );
  INV_X1 U10475 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9045) );
  OAI22_X1 U10476 ( .A1(n9046), .A2(n9168), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9045), .ZN(n9047) );
  AOI21_X1 U10477 ( .B1(n9682), .B2(n9165), .A(n9047), .ZN(n9048) );
  OAI211_X1 U10478 ( .C1(n9677), .C2(n9161), .A(n9049), .B(n9048), .ZN(
        P1_U3216) );
  XOR2_X1 U10479 ( .A(n9051), .B(n9050), .Z(n9055) );
  AOI22_X1 U10480 ( .A1(n9435), .A2(n9152), .B1(n9604), .B2(n9437), .ZN(n9732)
         );
  AOI22_X1 U10481 ( .A1(n9158), .A2(n9738), .B1(P1_REG3_REG_19__SCAN_IN), .B2(
        P1_U3086), .ZN(n9052) );
  OAI21_X1 U10482 ( .B1(n9732), .B2(n9156), .A(n9052), .ZN(n9053) );
  AOI21_X1 U10483 ( .B1(n9806), .B2(n9171), .A(n9053), .ZN(n9054) );
  OAI21_X1 U10484 ( .B1(n9055), .B2(n9174), .A(n9054), .ZN(P1_U3219) );
  XOR2_X1 U10485 ( .A(n9057), .B(n9056), .Z(n9063) );
  OR2_X1 U10486 ( .A1(n9256), .A2(n9128), .ZN(n9059) );
  NAND2_X1 U10487 ( .A1(n9435), .A2(n9604), .ZN(n9058) );
  AND2_X1 U10488 ( .A1(n9059), .A2(n9058), .ZN(n9710) );
  AOI22_X1 U10489 ( .A1(n9158), .A2(n9703), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n9060) );
  OAI21_X1 U10490 ( .B1(n9710), .B2(n9156), .A(n9060), .ZN(n9061) );
  AOI21_X1 U10491 ( .B1(n9794), .B2(n9171), .A(n9061), .ZN(n9062) );
  OAI21_X1 U10492 ( .B1(n9063), .B2(n9174), .A(n9062), .ZN(P1_U3223) );
  AOI21_X1 U10493 ( .B1(n9066), .B2(n9065), .A(n9064), .ZN(n9071) );
  AND2_X1 U10494 ( .A1(n9430), .A2(n9152), .ZN(n9067) );
  AOI21_X1 U10495 ( .B1(n9432), .B2(n9604), .A(n9067), .ZN(n9646) );
  AOI22_X1 U10496 ( .A1(n9158), .A2(n9652), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n9068) );
  OAI21_X1 U10497 ( .B1(n9646), .B2(n9156), .A(n9068), .ZN(n9069) );
  AOI21_X1 U10498 ( .B1(n9776), .B2(n9171), .A(n9069), .ZN(n9070) );
  OAI21_X1 U10499 ( .B1(n9071), .B2(n9174), .A(n9070), .ZN(P1_U3225) );
  XNOR2_X1 U10500 ( .A(n9072), .B(n9073), .ZN(n9164) );
  NOR2_X1 U10501 ( .A1(n9164), .A2(n9163), .ZN(n9162) );
  AOI21_X1 U10502 ( .B1(n9073), .B2(n9072), .A(n9162), .ZN(n9077) );
  XNOR2_X1 U10503 ( .A(n9075), .B(n9074), .ZN(n9076) );
  XNOR2_X1 U10504 ( .A(n9077), .B(n9076), .ZN(n9085) );
  NOR2_X1 U10505 ( .A1(n9168), .A2(n9078), .ZN(n9082) );
  INV_X1 U10506 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9079) );
  OAI22_X1 U10507 ( .A1(n9080), .A2(n9156), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9079), .ZN(n9081) );
  AOI211_X1 U10508 ( .C1(n9083), .C2(n9171), .A(n9082), .B(n9081), .ZN(n9084)
         );
  OAI21_X1 U10509 ( .B1(n9085), .B2(n9174), .A(n9084), .ZN(P1_U3226) );
  XOR2_X1 U10510 ( .A(n9087), .B(n9086), .Z(n9099) );
  INV_X1 U10511 ( .A(n9091), .ZN(n9088) );
  AOI21_X1 U10512 ( .B1(n9089), .B2(n9088), .A(P1_U3086), .ZN(n9095) );
  NAND2_X1 U10513 ( .A1(n9090), .A2(n9165), .ZN(n9093) );
  NAND3_X1 U10514 ( .A1(n9158), .A2(n9091), .A3(n9094), .ZN(n9092) );
  OAI211_X1 U10515 ( .C1(n9095), .C2(n9094), .A(n9093), .B(n9092), .ZN(n9096)
         );
  AOI21_X1 U10516 ( .B1(n9097), .B2(n9171), .A(n9096), .ZN(n9098) );
  OAI21_X1 U10517 ( .B1(n9099), .B2(n9174), .A(n9098), .ZN(P1_U3228) );
  AND3_X1 U10518 ( .A1(n9038), .A2(n9101), .A3(n9100), .ZN(n9102) );
  OAI21_X1 U10519 ( .B1(n9103), .B2(n9102), .A(n9150), .ZN(n9109) );
  OAI22_X1 U10520 ( .A1(n9129), .A2(n9114), .B1(n9104), .B2(n9128), .ZN(n9667)
         );
  INV_X1 U10521 ( .A(n9661), .ZN(n9106) );
  INV_X1 U10522 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9105) );
  OAI22_X1 U10523 ( .A1(n9106), .A2(n9168), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9105), .ZN(n9107) );
  AOI21_X1 U10524 ( .B1(n9667), .B2(n9165), .A(n9107), .ZN(n9108) );
  OAI211_X1 U10525 ( .C1(n9663), .C2(n9161), .A(n9109), .B(n9108), .ZN(
        P1_U3229) );
  XNOR2_X1 U10526 ( .A(n9111), .B(n9110), .ZN(n9112) );
  XNOR2_X1 U10527 ( .A(n9113), .B(n9112), .ZN(n9121) );
  INV_X1 U10528 ( .A(n9721), .ZN(n9118) );
  OAI22_X1 U10529 ( .A1(n9116), .A2(n9128), .B1(n9115), .B2(n9114), .ZN(n9725)
         );
  AOI22_X1 U10530 ( .A1(n9725), .A2(n9165), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n9117) );
  OAI21_X1 U10531 ( .B1(n9118), .B2(n9168), .A(n9117), .ZN(n9119) );
  AOI21_X1 U10532 ( .B1(n9800), .B2(n9171), .A(n9119), .ZN(n9120) );
  OAI21_X1 U10533 ( .B1(n9121), .B2(n9174), .A(n9120), .ZN(P1_U3233) );
  INV_X1 U10534 ( .A(n9039), .ZN(n9126) );
  OAI21_X1 U10535 ( .B1(n9123), .B2(n9125), .A(n9122), .ZN(n9124) );
  OAI21_X1 U10536 ( .B1(n9126), .B2(n9125), .A(n9124), .ZN(n9127) );
  NAND2_X1 U10537 ( .A1(n9127), .A2(n9150), .ZN(n9136) );
  OR2_X1 U10538 ( .A1(n9129), .A2(n9128), .ZN(n9131) );
  NAND2_X1 U10539 ( .A1(n9434), .A2(n9604), .ZN(n9130) );
  NAND2_X1 U10540 ( .A1(n9131), .A2(n9130), .ZN(n9695) );
  OAI22_X1 U10541 ( .A1(n9168), .A2(n9133), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9132), .ZN(n9134) );
  AOI21_X1 U10542 ( .B1(n9695), .B2(n9165), .A(n9134), .ZN(n9135) );
  OAI211_X1 U10543 ( .C1(n9691), .C2(n9161), .A(n9136), .B(n9135), .ZN(
        P1_U3235) );
  OAI21_X1 U10544 ( .B1(n9139), .B2(n9138), .A(n9137), .ZN(n9145) );
  NAND2_X1 U10545 ( .A1(n9810), .A2(n9171), .ZN(n9142) );
  AOI22_X1 U10546 ( .A1(n9140), .A2(n9165), .B1(P1_REG3_REG_18__SCAN_IN), .B2(
        P1_U3086), .ZN(n9141) );
  OAI211_X1 U10547 ( .C1(n9168), .C2(n9143), .A(n9142), .B(n9141), .ZN(n9144)
         );
  AOI21_X1 U10548 ( .B1(n9145), .B2(n9150), .A(n9144), .ZN(n9146) );
  INV_X1 U10549 ( .A(n9146), .ZN(P1_U3238) );
  INV_X1 U10550 ( .A(n9771), .ZN(n9639) );
  OAI21_X1 U10551 ( .B1(n9064), .B2(n9148), .A(n9147), .ZN(n9149) );
  NAND3_X1 U10552 ( .A1(n9151), .A2(n9150), .A3(n9149), .ZN(n9160) );
  NAND2_X1 U10553 ( .A1(n9429), .A2(n9152), .ZN(n9154) );
  NAND2_X1 U10554 ( .A1(n9431), .A2(n9604), .ZN(n9153) );
  AND2_X1 U10555 ( .A1(n9154), .A2(n9153), .ZN(n9633) );
  INV_X1 U10556 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9155) );
  OAI22_X1 U10557 ( .A1(n9156), .A2(n9633), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9155), .ZN(n9157) );
  AOI21_X1 U10558 ( .B1(n9636), .B2(n9158), .A(n9157), .ZN(n9159) );
  OAI211_X1 U10559 ( .C1(n9639), .C2(n9161), .A(n9160), .B(n9159), .ZN(
        P1_U3240) );
  AOI21_X1 U10560 ( .B1(n9164), .B2(n9163), .A(n9162), .ZN(n9175) );
  AOI22_X1 U10561 ( .A1(n9166), .A2(n9165), .B1(P1_REG3_REG_15__SCAN_IN), .B2(
        P1_U3086), .ZN(n9167) );
  OAI21_X1 U10562 ( .B1(n9169), .B2(n9168), .A(n9167), .ZN(n9170) );
  AOI21_X1 U10563 ( .B1(n9172), .B2(n9171), .A(n9170), .ZN(n9173) );
  OAI21_X1 U10564 ( .B1(n9175), .B2(n9174), .A(n9173), .ZN(P1_U3241) );
  NAND2_X1 U10565 ( .A1(n9177), .A2(n9176), .ZN(n9179) );
  OR2_X1 U10566 ( .A1(n6003), .A2(n7523), .ZN(n9178) );
  INV_X1 U10567 ( .A(n9596), .ZN(n9748) );
  INV_X1 U10568 ( .A(n9379), .ZN(n9217) );
  INV_X1 U10569 ( .A(n9380), .ZN(n9216) );
  INV_X1 U10570 ( .A(n9180), .ZN(n9181) );
  NOR2_X1 U10571 ( .A1(n9182), .A2(n9181), .ZN(n9189) );
  MUX2_X1 U10572 ( .A(n9183), .B(n9942), .S(n9287), .Z(n9193) );
  NAND3_X1 U10573 ( .A1(n9193), .A2(n9185), .A3(n9184), .ZN(n9187) );
  AND2_X1 U10574 ( .A1(n9186), .A2(n9365), .ZN(n9191) );
  INV_X1 U10575 ( .A(n9190), .ZN(n9199) );
  OAI21_X1 U10576 ( .B1(n9193), .B2(n9192), .A(n9191), .ZN(n9196) );
  AND2_X1 U10577 ( .A1(n9210), .A2(n9206), .ZN(n9372) );
  NAND3_X1 U10578 ( .A1(n9205), .A2(n9372), .A3(n9200), .ZN(n9203) );
  INV_X1 U10579 ( .A(n9372), .ZN(n9201) );
  OR2_X1 U10580 ( .A1(n9201), .A2(n9208), .ZN(n9202) );
  AND3_X1 U10581 ( .A1(n9894), .A2(n9209), .A3(n9202), .ZN(n9375) );
  INV_X1 U10582 ( .A(n9211), .ZN(n9374) );
  NAND2_X1 U10583 ( .A1(n9205), .A2(n9204), .ZN(n9207) );
  NAND2_X1 U10584 ( .A1(n9224), .A2(n9222), .ZN(n9377) );
  INV_X1 U10585 ( .A(n9377), .ZN(n9214) );
  OAI211_X1 U10586 ( .C1(n9377), .C2(n9213), .A(n9225), .B(n9219), .ZN(n9382)
         );
  AOI211_X1 U10587 ( .C1(n9218), .C2(n9214), .A(n9228), .B(n9382), .ZN(n9215)
         );
  AOI211_X1 U10588 ( .C1(n9217), .C2(n9383), .A(n9216), .B(n9215), .ZN(n9230)
         );
  INV_X1 U10589 ( .A(n9219), .ZN(n9221) );
  AOI211_X1 U10590 ( .C1(n9223), .C2(n9222), .A(n9221), .B(n9220), .ZN(n9227)
         );
  NAND2_X1 U10591 ( .A1(n9379), .A2(n9224), .ZN(n9226) );
  OAI21_X1 U10592 ( .B1(n9227), .B2(n9226), .A(n9225), .ZN(n9229) );
  NAND2_X1 U10593 ( .A1(n9244), .A2(n9231), .ZN(n9385) );
  NOR2_X1 U10594 ( .A1(n9249), .A2(n9385), .ZN(n9253) );
  INV_X1 U10595 ( .A(n9347), .ZN(n9232) );
  NAND4_X1 U10596 ( .A1(n9232), .A2(n9285), .A3(n9390), .A4(n9389), .ZN(n9252)
         );
  NAND3_X1 U10597 ( .A1(n9347), .A2(n9285), .A3(n9237), .ZN(n9242) );
  INV_X1 U10598 ( .A(n9237), .ZN(n9233) );
  NOR2_X1 U10599 ( .A1(n9233), .A2(n9235), .ZN(n9248) );
  INV_X1 U10600 ( .A(n9248), .ZN(n9234) );
  NAND3_X1 U10601 ( .A1(n9234), .A2(n9287), .A3(n9238), .ZN(n9241) );
  INV_X1 U10602 ( .A(n9235), .ZN(n9236) );
  NAND4_X1 U10603 ( .A1(n9237), .A2(n9285), .A3(n9236), .A4(n9392), .ZN(n9240)
         );
  NAND4_X1 U10604 ( .A1(n9238), .A2(n9287), .A3(n9706), .A4(n9390), .ZN(n9239)
         );
  NAND4_X1 U10605 ( .A1(n9242), .A2(n9241), .A3(n9240), .A4(n9239), .ZN(n9251)
         );
  NAND2_X1 U10606 ( .A1(n9389), .A2(n9243), .ZN(n9388) );
  INV_X1 U10607 ( .A(n9244), .ZN(n9245) );
  NOR3_X1 U10608 ( .A1(n9246), .A2(n9245), .A3(n9285), .ZN(n9247) );
  INV_X1 U10609 ( .A(n9694), .ZN(n9254) );
  NAND2_X1 U10610 ( .A1(n9259), .A2(n9678), .ZN(n9255) );
  INV_X1 U10611 ( .A(n9256), .ZN(n9433) );
  OR2_X1 U10612 ( .A1(n9691), .A2(n9433), .ZN(n9257) );
  NAND2_X1 U10613 ( .A1(n9258), .A2(n9257), .ZN(n9337) );
  MUX2_X1 U10614 ( .A(n9333), .B(n9340), .S(n9285), .Z(n9260) );
  OR2_X1 U10615 ( .A1(n9771), .A2(n9261), .ZN(n9330) );
  NAND2_X1 U10616 ( .A1(n9330), .A2(n9336), .ZN(n9264) );
  AOI21_X1 U10617 ( .B1(n9263), .B2(n9341), .A(n9264), .ZN(n9262) );
  NOR2_X1 U10618 ( .A1(n9262), .A2(n9394), .ZN(n9266) );
  MUX2_X1 U10619 ( .A(n9266), .B(n9265), .S(n9285), .Z(n9269) );
  NAND2_X1 U10620 ( .A1(n9598), .A2(n9267), .ZN(n9345) );
  AOI21_X1 U10621 ( .B1(n9269), .B2(n9331), .A(n9345), .ZN(n9268) );
  NOR2_X1 U10622 ( .A1(n9268), .A2(n9287), .ZN(n9273) );
  NAND2_X1 U10623 ( .A1(n9273), .A2(n9328), .ZN(n9275) );
  INV_X1 U10624 ( .A(n9328), .ZN(n9272) );
  INV_X1 U10625 ( .A(n9269), .ZN(n9270) );
  AOI21_X1 U10626 ( .B1(n9270), .B2(n9331), .A(n9345), .ZN(n9271) );
  NOR3_X1 U10627 ( .A1(n9273), .A2(n9272), .A3(n9271), .ZN(n9274) );
  AOI21_X1 U10628 ( .B1(n9285), .B2(n9275), .A(n9274), .ZN(n9278) );
  INV_X1 U10629 ( .A(n9428), .ZN(n9276) );
  NAND2_X1 U10630 ( .A1(n9754), .A2(n9276), .ZN(n9402) );
  MUX2_X1 U10631 ( .A(n9402), .B(n9329), .S(n9285), .Z(n9277) );
  NAND2_X1 U10632 ( .A1(n9279), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9282) );
  NAND2_X1 U10633 ( .A1(n9280), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n9281) );
  OAI211_X1 U10634 ( .C1(n9284), .C2(n9283), .A(n9282), .B(n9281), .ZN(n9603)
         );
  INV_X1 U10635 ( .A(n9603), .ZN(n9318) );
  NOR2_X1 U10636 ( .A1(n9751), .A2(n9318), .ZN(n9286) );
  NOR2_X1 U10637 ( .A1(n9354), .A2(n9318), .ZN(n9292) );
  AOI22_X1 U10638 ( .A1(n9288), .A2(n9286), .B1(n9292), .B2(n9285), .ZN(n9291)
         );
  INV_X1 U10639 ( .A(n9289), .ZN(n9290) );
  AND2_X1 U10640 ( .A1(n9596), .A2(n9290), .ZN(n9324) );
  NAND2_X1 U10641 ( .A1(n9289), .A2(n9603), .ZN(n9355) );
  AOI21_X1 U10642 ( .B1(n9325), .B2(n4429), .A(n9294), .ZN(n9427) );
  INV_X1 U10643 ( .A(n9292), .ZN(n9405) );
  XNOR2_X1 U10644 ( .A(n9705), .B(n9434), .ZN(n9708) );
  XNOR2_X1 U10645 ( .A(n9800), .B(n9435), .ZN(n9717) );
  INV_X1 U10646 ( .A(n9293), .ZN(n9312) );
  AND2_X1 U10647 ( .A1(n9295), .A2(n9294), .ZN(n9296) );
  NAND4_X1 U10648 ( .A1(n9298), .A2(n9297), .A3(n9296), .A4(n9973), .ZN(n9300)
         );
  NOR4_X1 U10649 ( .A1(n9300), .A2(n9299), .A3(n9950), .A4(n9963), .ZN(n9301)
         );
  AND4_X1 U10650 ( .A1(n5002), .A2(n9302), .A3(n4512), .A4(n9301), .ZN(n9303)
         );
  AND4_X1 U10651 ( .A1(n9902), .A2(n9304), .A3(n9910), .A4(n9303), .ZN(n9305)
         );
  NAND4_X1 U10652 ( .A1(n9308), .A2(n9307), .A3(n9306), .A4(n9305), .ZN(n9309)
         );
  NOR2_X1 U10653 ( .A1(n9310), .A2(n9309), .ZN(n9311) );
  NAND4_X1 U10654 ( .A1(n9717), .A2(n9731), .A3(n9312), .A4(n9311), .ZN(n9313)
         );
  NOR4_X1 U10655 ( .A1(n9314), .A2(n9694), .A3(n9708), .A4(n9313), .ZN(n9315)
         );
  AND4_X1 U10656 ( .A1(n9621), .A2(n4593), .A3(n4753), .A4(n9315), .ZN(n9316)
         );
  AND3_X1 U10657 ( .A1(n9317), .A2(n9316), .A3(n9632), .ZN(n9319) );
  NAND2_X1 U10658 ( .A1(n9354), .A2(n9318), .ZN(n9401) );
  AND4_X1 U10659 ( .A1(n9609), .A2(n9405), .A3(n9319), .A4(n9401), .ZN(n9320)
         );
  AND2_X1 U10660 ( .A1(n9320), .A2(n9408), .ZN(n9359) );
  INV_X1 U10661 ( .A(n9359), .ZN(n9323) );
  NOR3_X1 U10662 ( .A1(n9414), .A2(n6284), .A3(n9321), .ZN(n9322) );
  OAI21_X1 U10663 ( .B1(n9323), .B2(n9324), .A(n9322), .ZN(n9426) );
  INV_X1 U10664 ( .A(n9324), .ZN(n9407) );
  OAI21_X1 U10665 ( .B1(n6284), .B2(n9407), .A(n9325), .ZN(n9424) );
  NOR2_X1 U10666 ( .A1(n9408), .A2(n6284), .ZN(n9327) );
  NOR4_X1 U10667 ( .A1(n9327), .A2(n4429), .A3(n9414), .A4(n9326), .ZN(n9423)
         );
  NAND2_X1 U10668 ( .A1(n9329), .A2(n9328), .ZN(n9404) );
  NAND2_X1 U10669 ( .A1(n9331), .A2(n9330), .ZN(n9397) );
  NAND2_X1 U10670 ( .A1(n9333), .A2(n9332), .ZN(n9334) );
  NAND2_X1 U10671 ( .A1(n9334), .A2(n9340), .ZN(n9335) );
  AND2_X1 U10672 ( .A1(n9336), .A2(n9335), .ZN(n9346) );
  INV_X1 U10673 ( .A(n9337), .ZN(n9339) );
  NAND3_X1 U10674 ( .A1(n9340), .A2(n9339), .A3(n9338), .ZN(n9342) );
  AOI21_X1 U10675 ( .B1(n9346), .B2(n9342), .A(n4734), .ZN(n9343) );
  NOR2_X1 U10676 ( .A1(n9397), .A2(n9343), .ZN(n9344) );
  OR2_X1 U10677 ( .A1(n9345), .A2(n9344), .ZN(n9400) );
  INV_X1 U10678 ( .A(n9346), .ZN(n9348) );
  NOR2_X1 U10679 ( .A1(n9348), .A2(n9347), .ZN(n9396) );
  INV_X1 U10680 ( .A(n9724), .ZN(n9707) );
  AOI21_X1 U10681 ( .B1(n9396), .B2(n9707), .A(n9394), .ZN(n9349) );
  NOR2_X1 U10682 ( .A1(n9349), .A2(n9397), .ZN(n9350) );
  NOR2_X1 U10683 ( .A1(n9400), .A2(n9350), .ZN(n9352) );
  NAND2_X1 U10684 ( .A1(n9354), .A2(n9355), .ZN(n9351) );
  OAI211_X1 U10685 ( .C1(n9404), .C2(n9352), .A(n9402), .B(n9351), .ZN(n9353)
         );
  OAI21_X1 U10686 ( .B1(n9355), .B2(n9354), .A(n9353), .ZN(n9357) );
  AOI21_X1 U10687 ( .B1(n9357), .B2(n9408), .A(n9356), .ZN(n9360) );
  INV_X1 U10688 ( .A(n9414), .ZN(n9416) );
  AND4_X1 U10689 ( .A1(n9407), .A2(n9416), .A3(n9410), .A4(n6284), .ZN(n9358)
         );
  OAI21_X1 U10690 ( .B1(n9360), .B2(n9359), .A(n9358), .ZN(n9421) );
  NAND2_X1 U10691 ( .A1(n7114), .A2(n9986), .ZN(n9363) );
  NAND2_X1 U10692 ( .A1(n7440), .A2(n7439), .ZN(n9362) );
  AND4_X1 U10693 ( .A1(n9364), .A2(n9363), .A3(n9362), .A4(n9361), .ZN(n9368)
         );
  AND4_X1 U10694 ( .A1(n9368), .A2(n9367), .A3(n9366), .A4(n9365), .ZN(n9370)
         );
  OAI21_X1 U10695 ( .B1(n9371), .B2(n9370), .A(n9369), .ZN(n9373) );
  NAND2_X1 U10696 ( .A1(n9373), .A2(n9372), .ZN(n9376) );
  AOI21_X1 U10697 ( .B1(n9376), .B2(n9375), .A(n9374), .ZN(n9378) );
  NOR2_X1 U10698 ( .A1(n9378), .A2(n9377), .ZN(n9381) );
  OAI211_X1 U10699 ( .C1(n9382), .C2(n9381), .A(n9380), .B(n9379), .ZN(n9384)
         );
  AND2_X1 U10700 ( .A1(n9384), .A2(n9383), .ZN(n9387) );
  INV_X1 U10701 ( .A(n9385), .ZN(n9386) );
  OAI21_X1 U10702 ( .B1(n9388), .B2(n9387), .A(n9386), .ZN(n9391) );
  NAND3_X1 U10703 ( .A1(n9391), .A2(n9390), .A3(n9389), .ZN(n9393) );
  NAND2_X1 U10704 ( .A1(n9393), .A2(n9392), .ZN(n9395) );
  AOI21_X1 U10705 ( .B1(n9396), .B2(n9395), .A(n9394), .ZN(n9398) );
  NOR2_X1 U10706 ( .A1(n9398), .A2(n9397), .ZN(n9399) );
  NOR2_X1 U10707 ( .A1(n9400), .A2(n9399), .ZN(n9403) );
  OAI211_X1 U10708 ( .C1(n9404), .C2(n9403), .A(n9402), .B(n9401), .ZN(n9406)
         );
  NAND3_X1 U10709 ( .A1(n9407), .A2(n9406), .A3(n9405), .ZN(n9409) );
  NAND2_X1 U10710 ( .A1(n9409), .A2(n9408), .ZN(n9417) );
  OR4_X1 U10711 ( .A1(n9417), .A2(n9410), .A3(n9414), .A4(n6284), .ZN(n9420)
         );
  NAND3_X1 U10712 ( .A1(n9412), .A2(n9828), .A3(n9411), .ZN(n9413) );
  OAI211_X1 U10713 ( .C1(n4429), .C2(n9414), .A(n9413), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9419) );
  NAND3_X1 U10714 ( .A1(n9417), .A2(n9416), .A3(n9415), .ZN(n9418) );
  NAND4_X1 U10715 ( .A1(n9421), .A2(n9420), .A3(n9419), .A4(n9418), .ZN(n9422)
         );
  AOI21_X1 U10716 ( .B1(n9424), .B2(n9423), .A(n9422), .ZN(n9425) );
  OAI21_X1 U10717 ( .B1(n9427), .B2(n9426), .A(n9425), .ZN(P1_U3242) );
  MUX2_X1 U10718 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9603), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10719 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9428), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10720 ( .A(n9605), .B(P1_DATAO_REG_28__SCAN_IN), .S(n9452), .Z(
        P1_U3582) );
  MUX2_X1 U10721 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9429), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10722 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9430), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10723 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9431), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10724 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9432), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10725 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9433), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10726 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9434), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10727 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9435), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10728 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9436), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10729 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9437), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10730 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9438), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10731 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9439), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10732 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9440), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10733 ( .A(n9441), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9452), .Z(
        P1_U3568) );
  MUX2_X1 U10734 ( .A(n9442), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9452), .Z(
        P1_U3567) );
  MUX2_X1 U10735 ( .A(n9443), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9452), .Z(
        P1_U3566) );
  MUX2_X1 U10736 ( .A(n9444), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9452), .Z(
        P1_U3565) );
  MUX2_X1 U10737 ( .A(n9445), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9452), .Z(
        P1_U3564) );
  MUX2_X1 U10738 ( .A(n9446), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9452), .Z(
        P1_U3563) );
  MUX2_X1 U10739 ( .A(n9447), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9452), .Z(
        P1_U3562) );
  MUX2_X1 U10740 ( .A(n9448), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9452), .Z(
        P1_U3561) );
  MUX2_X1 U10741 ( .A(n9449), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9452), .Z(
        P1_U3560) );
  MUX2_X1 U10742 ( .A(n9450), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9452), .Z(
        P1_U3559) );
  MUX2_X1 U10743 ( .A(n9451), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9452), .Z(
        P1_U3558) );
  MUX2_X1 U10744 ( .A(n7463), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9452), .Z(
        P1_U3557) );
  MUX2_X1 U10745 ( .A(n7440), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9452), .Z(
        P1_U3555) );
  MUX2_X1 U10746 ( .A(n7114), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9452), .Z(
        P1_U3554) );
  AND2_X1 U10747 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9455) );
  NOR2_X1 U10748 ( .A1(n9578), .A2(n9453), .ZN(n9454) );
  AOI211_X1 U10749 ( .C1(n9878), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n9455), .B(
        n9454), .ZN(n9465) );
  AOI211_X1 U10750 ( .C1(n9458), .C2(n9457), .A(n9456), .B(n9879), .ZN(n9459)
         );
  INV_X1 U10751 ( .A(n9459), .ZN(n9464) );
  OAI211_X1 U10752 ( .C1(n9462), .C2(n9461), .A(n9888), .B(n9460), .ZN(n9463)
         );
  NAND3_X1 U10753 ( .A1(n9465), .A2(n9464), .A3(n9463), .ZN(P1_U3246) );
  AOI211_X1 U10754 ( .C1(n9468), .C2(n9467), .A(n9466), .B(n9879), .ZN(n9469)
         );
  INV_X1 U10755 ( .A(n9469), .ZN(n9480) );
  NAND2_X1 U10756 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n9470) );
  OAI21_X1 U10757 ( .B1(n9589), .B2(n9471), .A(n9470), .ZN(n9472) );
  AOI21_X1 U10758 ( .B1(n9885), .B2(n9473), .A(n9472), .ZN(n9479) );
  OAI211_X1 U10759 ( .C1(n9476), .C2(n9475), .A(n9888), .B(n9474), .ZN(n9477)
         );
  NAND4_X1 U10760 ( .A1(n9480), .A2(n9479), .A3(n9478), .A4(n9477), .ZN(
        P1_U3247) );
  AND2_X1 U10761 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9482) );
  NOR2_X1 U10762 ( .A1(n9578), .A2(n9505), .ZN(n9481) );
  AOI211_X1 U10763 ( .C1(n9878), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n9482), .B(
        n9481), .ZN(n9497) );
  AOI21_X1 U10764 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n9484), .A(n9483), .ZN(
        n9487) );
  NAND2_X1 U10765 ( .A1(n9499), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9485) );
  OAI21_X1 U10766 ( .B1(n9499), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9485), .ZN(
        n9486) );
  NOR2_X1 U10767 ( .A1(n9487), .A2(n9486), .ZN(n9498) );
  AOI211_X1 U10768 ( .C1(n9487), .C2(n9486), .A(n9498), .B(n9879), .ZN(n9488)
         );
  INV_X1 U10769 ( .A(n9488), .ZN(n9496) );
  NOR2_X1 U10770 ( .A1(n9505), .A2(n9489), .ZN(n9490) );
  AOI21_X1 U10771 ( .B1(n9489), .B2(n9505), .A(n9490), .ZN(n9494) );
  OAI21_X1 U10772 ( .B1(n9492), .B2(n7924), .A(n9491), .ZN(n9493) );
  NAND2_X1 U10773 ( .A1(n9494), .A2(n9493), .ZN(n9504) );
  OAI211_X1 U10774 ( .C1(n9494), .C2(n9493), .A(n9888), .B(n9504), .ZN(n9495)
         );
  NAND3_X1 U10775 ( .A1(n9497), .A2(n9496), .A3(n9495), .ZN(P1_U3257) );
  AOI211_X1 U10776 ( .C1(n9500), .C2(n8050), .A(n9521), .B(n9879), .ZN(n9501)
         );
  INV_X1 U10777 ( .A(n9501), .ZN(n9511) );
  NOR2_X1 U10778 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9502), .ZN(n9503) );
  AOI21_X1 U10779 ( .B1(n9878), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n9503), .ZN(
        n9510) );
  OAI21_X1 U10780 ( .B1(n9489), .B2(n9505), .A(n9504), .ZN(n9512) );
  INV_X1 U10781 ( .A(n9512), .ZN(n9506) );
  XNOR2_X1 U10782 ( .A(n9513), .B(n9506), .ZN(n9507) );
  NAND2_X1 U10783 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n9507), .ZN(n9514) );
  OAI211_X1 U10784 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n9507), .A(n9888), .B(
        n9514), .ZN(n9509) );
  NAND2_X1 U10785 ( .A1(n9885), .A2(n9513), .ZN(n9508) );
  NAND4_X1 U10786 ( .A1(n9511), .A2(n9510), .A3(n9509), .A4(n9508), .ZN(
        P1_U3258) );
  INV_X1 U10787 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9856) );
  MUX2_X1 U10788 ( .A(n9856), .B(P1_REG1_REG_16__SCAN_IN), .S(n9537), .Z(n9517) );
  NAND2_X1 U10789 ( .A1(n9513), .A2(n9512), .ZN(n9515) );
  AND2_X1 U10790 ( .A1(n9515), .A2(n9514), .ZN(n9516) );
  NAND2_X1 U10791 ( .A1(n9516), .A2(n9517), .ZN(n9543) );
  OAI21_X1 U10792 ( .B1(n9517), .B2(n9516), .A(n9543), .ZN(n9529) );
  AND2_X1 U10793 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9518) );
  AOI21_X1 U10794 ( .B1(n9878), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n9518), .ZN(
        n9519) );
  OAI21_X1 U10795 ( .B1(n9537), .B2(n9578), .A(n9519), .ZN(n9528) );
  NOR2_X1 U10796 ( .A1(n9520), .A2(n4609), .ZN(n9522) );
  XNOR2_X1 U10797 ( .A(n9537), .B(n9523), .ZN(n9525) );
  INV_X1 U10798 ( .A(n9534), .ZN(n9524) );
  AOI211_X1 U10799 ( .C1(n9526), .C2(n9525), .A(n9879), .B(n9524), .ZN(n9527)
         );
  AOI211_X1 U10800 ( .C1(n9888), .C2(n9529), .A(n9528), .B(n9527), .ZN(n9530)
         );
  INV_X1 U10801 ( .A(n9530), .ZN(P1_U3259) );
  OR2_X1 U10802 ( .A1(n9561), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9552) );
  NAND2_X1 U10803 ( .A1(n9561), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9531) );
  AND2_X1 U10804 ( .A1(n9552), .A2(n9531), .ZN(n9536) );
  NAND2_X1 U10805 ( .A1(n9532), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9533) );
  OAI21_X1 U10806 ( .B1(n9536), .B2(n9535), .A(n9553), .ZN(n9550) );
  NAND2_X1 U10807 ( .A1(n9537), .A2(n9856), .ZN(n9541) );
  OR2_X1 U10808 ( .A1(n9561), .A2(n9538), .ZN(n9540) );
  NAND2_X1 U10809 ( .A1(n9561), .A2(n9538), .ZN(n9539) );
  AND2_X1 U10810 ( .A1(n9540), .A2(n9539), .ZN(n9542) );
  AOI21_X1 U10811 ( .B1(n9543), .B2(n9541), .A(n9542), .ZN(n9564) );
  INV_X1 U10812 ( .A(n9564), .ZN(n9545) );
  NAND3_X1 U10813 ( .A1(n9543), .A2(n9542), .A3(n9541), .ZN(n9544) );
  AOI21_X1 U10814 ( .B1(n9545), .B2(n9544), .A(n9579), .ZN(n9549) );
  AOI22_X1 U10815 ( .A1(n9878), .A2(P1_ADDR_REG_17__SCAN_IN), .B1(
        P1_REG3_REG_17__SCAN_IN), .B2(P1_U3086), .ZN(n9546) );
  OAI21_X1 U10816 ( .B1(n9547), .B2(n9578), .A(n9546), .ZN(n9548) );
  AOI211_X1 U10817 ( .C1(n9550), .C2(n9582), .A(n9549), .B(n9548), .ZN(n9551)
         );
  INV_X1 U10818 ( .A(n9551), .ZN(P1_U3260) );
  OR2_X1 U10819 ( .A1(n9575), .A2(n9554), .ZN(n9556) );
  NAND2_X1 U10820 ( .A1(n9575), .A2(n9554), .ZN(n9555) );
  NAND2_X1 U10821 ( .A1(n9556), .A2(n9555), .ZN(n9557) );
  OAI211_X1 U10822 ( .C1(n9558), .C2(n9557), .A(n9571), .B(n9582), .ZN(n9570)
         );
  NOR2_X1 U10823 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9559), .ZN(n9560) );
  AOI21_X1 U10824 ( .B1(n9878), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n9560), .ZN(
        n9569) );
  NOR2_X1 U10825 ( .A1(n9561), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9563) );
  XNOR2_X1 U10826 ( .A(n9575), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9562) );
  NOR3_X1 U10827 ( .A1(n9564), .A2(n9563), .A3(n9562), .ZN(n9574) );
  INV_X1 U10828 ( .A(n9574), .ZN(n9566) );
  OAI21_X1 U10829 ( .B1(n9564), .B2(n9563), .A(n9562), .ZN(n9565) );
  NAND3_X1 U10830 ( .A1(n9566), .A2(n9888), .A3(n9565), .ZN(n9568) );
  NAND2_X1 U10831 ( .A1(n9885), .A2(n9575), .ZN(n9567) );
  NAND4_X1 U10832 ( .A1(n9570), .A2(n9569), .A3(n9568), .A4(n9567), .ZN(
        P1_U3261) );
  INV_X1 U10833 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9572) );
  XNOR2_X1 U10834 ( .A(n9573), .B(n9572), .ZN(n9577) );
  AOI21_X1 U10835 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n9575), .A(n9574), .ZN(
        n9576) );
  XNOR2_X1 U10836 ( .A(n9576), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9580) );
  AOI22_X1 U10837 ( .A1(n9577), .A2(n9582), .B1(n9888), .B2(n9580), .ZN(n9586)
         );
  INV_X1 U10838 ( .A(n9577), .ZN(n9583) );
  OAI21_X1 U10839 ( .B1(n9580), .B2(n9579), .A(n9578), .ZN(n9581) );
  AOI21_X1 U10840 ( .B1(n9583), .B2(n9582), .A(n9581), .ZN(n9585) );
  MUX2_X1 U10841 ( .A(n9586), .B(n9585), .S(n9584), .Z(n9588) );
  NAND2_X1 U10842 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n9587) );
  OAI211_X1 U10843 ( .C1(n9590), .C2(n9589), .A(n9588), .B(n9587), .ZN(
        P1_U3262) );
  XNOR2_X1 U10844 ( .A(n9591), .B(n9596), .ZN(n9592) );
  NAND2_X1 U10845 ( .A1(n9592), .A2(n9985), .ZN(n9747) );
  NOR2_X1 U10846 ( .A1(n9744), .A2(n9593), .ZN(n9595) );
  AOI211_X1 U10847 ( .C1(n9596), .C2(n9981), .A(n9595), .B(n9594), .ZN(n9597)
         );
  OAI21_X1 U10848 ( .B1(n9747), .B2(n9987), .A(n9597), .ZN(P1_U3263) );
  NAND2_X1 U10849 ( .A1(n9599), .A2(n9598), .ZN(n9600) );
  XNOR2_X1 U10850 ( .A(n9610), .B(n9609), .ZN(n9752) );
  NAND2_X1 U10851 ( .A1(n9752), .A2(n9968), .ZN(n9618) );
  AOI21_X1 U10852 ( .B1(n9754), .B2(n9611), .A(n9737), .ZN(n9612) );
  NAND2_X1 U10853 ( .A1(n9754), .A2(n9981), .ZN(n9615) );
  AOI22_X1 U10854 ( .A1(n9992), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9983), .B2(
        n9613), .ZN(n9614) );
  NAND2_X1 U10855 ( .A1(n9615), .A2(n9614), .ZN(n9616) );
  AOI21_X1 U10856 ( .B1(n9753), .B2(n9967), .A(n9616), .ZN(n9617) );
  OAI211_X1 U10857 ( .C1(n9756), .C2(n9947), .A(n9618), .B(n9617), .ZN(
        P1_U3356) );
  XNOR2_X1 U10858 ( .A(n9620), .B(n9619), .ZN(n9768) );
  XNOR2_X1 U10859 ( .A(n9622), .B(n9621), .ZN(n9624) );
  OAI21_X1 U10860 ( .B1(n9624), .B2(n9913), .A(n9623), .ZN(n9764) );
  AOI211_X1 U10861 ( .C1(n9766), .C2(n9634), .A(n9737), .B(n4454), .ZN(n9765)
         );
  NAND2_X1 U10862 ( .A1(n9765), .A2(n9967), .ZN(n9627) );
  AOI22_X1 U10863 ( .A1(n9992), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9625), .B2(
        n9983), .ZN(n9626) );
  OAI211_X1 U10864 ( .C1(n9628), .C2(n9741), .A(n9627), .B(n9626), .ZN(n9629)
         );
  AOI21_X1 U10865 ( .B1(n9764), .B2(n9744), .A(n9629), .ZN(n9630) );
  OAI21_X1 U10866 ( .B1(n9768), .B2(n9746), .A(n9630), .ZN(P1_U3266) );
  XNOR2_X1 U10867 ( .A(n9631), .B(n9632), .ZN(n9773) );
  INV_X1 U10868 ( .A(n9634), .ZN(n9635) );
  AOI211_X1 U10869 ( .C1(n9771), .C2(n9649), .A(n9737), .B(n9635), .ZN(n9770)
         );
  NAND2_X1 U10870 ( .A1(n9770), .A2(n9967), .ZN(n9638) );
  AOI22_X1 U10871 ( .A1(n9992), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9636), .B2(
        n9983), .ZN(n9637) );
  OAI211_X1 U10872 ( .C1(n9639), .C2(n9741), .A(n9638), .B(n9637), .ZN(n9640)
         );
  AOI21_X1 U10873 ( .B1(n9769), .B2(n9744), .A(n9640), .ZN(n9641) );
  OAI21_X1 U10874 ( .B1(n9773), .B2(n9746), .A(n9641), .ZN(P1_U3267) );
  XNOR2_X1 U10875 ( .A(n9642), .B(n9643), .ZN(n9778) );
  INV_X1 U10876 ( .A(n9644), .ZN(n9645) );
  OAI21_X1 U10877 ( .B1(n9645), .B2(n4753), .A(n9980), .ZN(n9648) );
  OAI21_X1 U10878 ( .B1(n9648), .B2(n9647), .A(n9646), .ZN(n9774) );
  INV_X1 U10879 ( .A(n9659), .ZN(n9651) );
  INV_X1 U10880 ( .A(n9649), .ZN(n9650) );
  AOI211_X1 U10881 ( .C1(n9776), .C2(n9651), .A(n9737), .B(n9650), .ZN(n9775)
         );
  NAND2_X1 U10882 ( .A1(n9775), .A2(n9967), .ZN(n9654) );
  AOI22_X1 U10883 ( .A1(n9992), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9652), .B2(
        n9983), .ZN(n9653) );
  OAI211_X1 U10884 ( .C1(n9655), .C2(n9741), .A(n9654), .B(n9653), .ZN(n9656)
         );
  AOI21_X1 U10885 ( .B1(n9774), .B2(n9744), .A(n9656), .ZN(n9657) );
  OAI21_X1 U10886 ( .B1(n9778), .B2(n9746), .A(n9657), .ZN(P1_U3268) );
  XNOR2_X1 U10887 ( .A(n9658), .B(n4593), .ZN(n9783) );
  INV_X1 U10888 ( .A(n9673), .ZN(n9660) );
  AOI211_X1 U10889 ( .C1(n9780), .C2(n9660), .A(n9737), .B(n9659), .ZN(n9779)
         );
  AOI22_X1 U10890 ( .A1(n9661), .A2(n9983), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9947), .ZN(n9662) );
  OAI21_X1 U10891 ( .B1(n9663), .B2(n9741), .A(n9662), .ZN(n9670) );
  AOI211_X1 U10892 ( .C1(n9666), .C2(n9665), .A(n9913), .B(n9664), .ZN(n9668)
         );
  NOR2_X1 U10893 ( .A1(n9668), .A2(n9667), .ZN(n9782) );
  NOR2_X1 U10894 ( .A1(n9782), .A2(n9947), .ZN(n9669) );
  AOI211_X1 U10895 ( .C1(n9779), .C2(n9967), .A(n9670), .B(n9669), .ZN(n9671)
         );
  OAI21_X1 U10896 ( .B1(n9783), .B2(n9746), .A(n9671), .ZN(P1_U3269) );
  XNOR2_X1 U10897 ( .A(n9672), .B(n9680), .ZN(n9788) );
  INV_X1 U10898 ( .A(n9688), .ZN(n9674) );
  AOI211_X1 U10899 ( .C1(n9785), .C2(n9674), .A(n9737), .B(n9673), .ZN(n9784)
         );
  AOI22_X1 U10900 ( .A1(n9675), .A2(n9983), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9947), .ZN(n9676) );
  OAI21_X1 U10901 ( .B1(n9677), .B2(n9741), .A(n9676), .ZN(n9685) );
  INV_X1 U10902 ( .A(n9678), .ZN(n9679) );
  NOR2_X1 U10903 ( .A1(n9692), .A2(n9679), .ZN(n9681) );
  XNOR2_X1 U10904 ( .A(n9681), .B(n9680), .ZN(n9683) );
  AOI21_X1 U10905 ( .B1(n9683), .B2(n9980), .A(n9682), .ZN(n9787) );
  NOR2_X1 U10906 ( .A1(n9787), .A2(n9947), .ZN(n9684) );
  AOI211_X1 U10907 ( .C1(n9784), .C2(n9967), .A(n9685), .B(n9684), .ZN(n9686)
         );
  OAI21_X1 U10908 ( .B1(n9788), .B2(n9746), .A(n9686), .ZN(P1_U3270) );
  XNOR2_X1 U10909 ( .A(n9687), .B(n9694), .ZN(n9793) );
  AOI211_X1 U10910 ( .C1(n9790), .C2(n9701), .A(n9737), .B(n9688), .ZN(n9789)
         );
  AOI22_X1 U10911 ( .A1(n9689), .A2(n9983), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9947), .ZN(n9690) );
  OAI21_X1 U10912 ( .B1(n9691), .B2(n9741), .A(n9690), .ZN(n9698) );
  AOI211_X1 U10913 ( .C1(n9694), .C2(n9693), .A(n9913), .B(n9692), .ZN(n9696)
         );
  NOR2_X1 U10914 ( .A1(n9696), .A2(n9695), .ZN(n9792) );
  NOR2_X1 U10915 ( .A1(n9792), .A2(n9992), .ZN(n9697) );
  AOI211_X1 U10916 ( .C1(n9789), .C2(n9967), .A(n9698), .B(n9697), .ZN(n9699)
         );
  OAI21_X1 U10917 ( .B1(n9793), .B2(n9746), .A(n9699), .ZN(P1_U3271) );
  XNOR2_X1 U10918 ( .A(n9700), .B(n9708), .ZN(n9798) );
  INV_X1 U10919 ( .A(n9701), .ZN(n9702) );
  AOI21_X1 U10920 ( .B1(n9794), .B2(n9719), .A(n9702), .ZN(n9795) );
  AOI22_X1 U10921 ( .A1(n9947), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9703), .B2(
        n9983), .ZN(n9704) );
  OAI21_X1 U10922 ( .B1(n9705), .B2(n9741), .A(n9704), .ZN(n9714) );
  INV_X1 U10923 ( .A(n9717), .ZN(n9723) );
  OAI21_X1 U10924 ( .B1(n9707), .B2(n9723), .A(n9706), .ZN(n9709) );
  XNOR2_X1 U10925 ( .A(n9709), .B(n9708), .ZN(n9712) );
  INV_X1 U10926 ( .A(n9710), .ZN(n9711) );
  AOI21_X1 U10927 ( .B1(n9712), .B2(n9980), .A(n9711), .ZN(n9797) );
  NOR2_X1 U10928 ( .A1(n9797), .A2(n9992), .ZN(n9713) );
  AOI211_X1 U10929 ( .C1(n9795), .C2(n9715), .A(n9714), .B(n9713), .ZN(n9716)
         );
  OAI21_X1 U10930 ( .B1(n9798), .B2(n9746), .A(n9716), .ZN(P1_U3272) );
  XNOR2_X1 U10931 ( .A(n9718), .B(n9717), .ZN(n9803) );
  INV_X1 U10932 ( .A(n9719), .ZN(n9720) );
  AOI211_X1 U10933 ( .C1(n9800), .C2(n9735), .A(n9737), .B(n9720), .ZN(n9799)
         );
  AOI22_X1 U10934 ( .A1(n9947), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9721), .B2(
        n9983), .ZN(n9722) );
  OAI21_X1 U10935 ( .B1(n4669), .B2(n9741), .A(n9722), .ZN(n9728) );
  XNOR2_X1 U10936 ( .A(n9724), .B(n9723), .ZN(n9726) );
  AOI21_X1 U10937 ( .B1(n9726), .B2(n9980), .A(n9725), .ZN(n9802) );
  NOR2_X1 U10938 ( .A1(n9802), .A2(n9947), .ZN(n9727) );
  AOI211_X1 U10939 ( .C1(n9799), .C2(n9967), .A(n9728), .B(n9727), .ZN(n9729)
         );
  OAI21_X1 U10940 ( .B1(n9803), .B2(n9746), .A(n9729), .ZN(P1_U3273) );
  XOR2_X1 U10941 ( .A(n9731), .B(n4500), .Z(n9808) );
  XOR2_X1 U10942 ( .A(n9731), .B(n9730), .Z(n9733) );
  OAI21_X1 U10943 ( .B1(n9733), .B2(n9913), .A(n9732), .ZN(n9804) );
  INV_X1 U10944 ( .A(n9735), .ZN(n9736) );
  AOI211_X1 U10945 ( .C1(n9806), .C2(n4672), .A(n9737), .B(n9736), .ZN(n9805)
         );
  NAND2_X1 U10946 ( .A1(n9805), .A2(n9967), .ZN(n9740) );
  AOI22_X1 U10947 ( .A1(n9992), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9738), .B2(
        n9983), .ZN(n9739) );
  OAI211_X1 U10948 ( .C1(n9742), .C2(n9741), .A(n9740), .B(n9739), .ZN(n9743)
         );
  AOI21_X1 U10949 ( .B1(n9744), .B2(n9804), .A(n9743), .ZN(n9745) );
  OAI21_X1 U10950 ( .B1(n9808), .B2(n9746), .A(n9745), .ZN(P1_U3274) );
  INV_X1 U10951 ( .A(n10059), .ZN(n10091) );
  OAI211_X1 U10952 ( .C1(n9748), .C2(n10091), .A(n9747), .B(n9749), .ZN(n9814)
         );
  MUX2_X1 U10953 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9814), .S(n10120), .Z(
        P1_U3553) );
  OAI211_X1 U10954 ( .C1(n9751), .C2(n10091), .A(n9750), .B(n9749), .ZN(n9815)
         );
  MUX2_X1 U10955 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9815), .S(n10120), .Z(
        P1_U3552) );
  NAND2_X1 U10956 ( .A1(n9752), .A2(n10095), .ZN(n9757) );
  AOI21_X1 U10957 ( .B1(n10059), .B2(n9754), .A(n9753), .ZN(n9755) );
  MUX2_X1 U10958 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9816), .S(n10120), .Z(
        P1_U3551) );
  NAND2_X1 U10959 ( .A1(n9759), .A2(n10059), .ZN(n9761) );
  MUX2_X1 U10960 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9817), .S(n10120), .Z(
        P1_U3550) );
  INV_X1 U10961 ( .A(n10095), .ZN(n10061) );
  AOI211_X1 U10962 ( .C1(n10059), .C2(n9766), .A(n9765), .B(n9764), .ZN(n9767)
         );
  OAI21_X1 U10963 ( .B1(n9768), .B2(n10061), .A(n9767), .ZN(n9818) );
  MUX2_X1 U10964 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9818), .S(n10120), .Z(
        P1_U3549) );
  OAI21_X1 U10965 ( .B1(n9773), .B2(n10061), .A(n9772), .ZN(n9819) );
  MUX2_X1 U10966 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9819), .S(n10120), .Z(
        P1_U3548) );
  AOI211_X1 U10967 ( .C1(n10059), .C2(n9776), .A(n9775), .B(n9774), .ZN(n9777)
         );
  OAI21_X1 U10968 ( .B1(n9778), .B2(n10061), .A(n9777), .ZN(n9820) );
  MUX2_X1 U10969 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9820), .S(n10120), .Z(
        P1_U3547) );
  AOI21_X1 U10970 ( .B1(n10059), .B2(n9780), .A(n9779), .ZN(n9781) );
  OAI211_X1 U10971 ( .C1(n9783), .C2(n10061), .A(n9782), .B(n9781), .ZN(n9821)
         );
  MUX2_X1 U10972 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9821), .S(n10120), .Z(
        P1_U3546) );
  AOI21_X1 U10973 ( .B1(n10059), .B2(n9785), .A(n9784), .ZN(n9786) );
  OAI211_X1 U10974 ( .C1(n9788), .C2(n10061), .A(n9787), .B(n9786), .ZN(n9822)
         );
  MUX2_X1 U10975 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9822), .S(n10120), .Z(
        P1_U3545) );
  AOI21_X1 U10976 ( .B1(n10059), .B2(n9790), .A(n9789), .ZN(n9791) );
  OAI211_X1 U10977 ( .C1(n9793), .C2(n10061), .A(n9792), .B(n9791), .ZN(n9823)
         );
  MUX2_X1 U10978 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9823), .S(n10120), .Z(
        P1_U3544) );
  AOI22_X1 U10979 ( .A1(n9795), .A2(n9985), .B1(n10059), .B2(n9794), .ZN(n9796) );
  OAI211_X1 U10980 ( .C1(n9798), .C2(n10061), .A(n9797), .B(n9796), .ZN(n9824)
         );
  MUX2_X1 U10981 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9824), .S(n10120), .Z(
        P1_U3543) );
  AOI21_X1 U10982 ( .B1(n10059), .B2(n9800), .A(n9799), .ZN(n9801) );
  OAI211_X1 U10983 ( .C1(n9803), .C2(n10061), .A(n9802), .B(n9801), .ZN(n9825)
         );
  MUX2_X1 U10984 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9825), .S(n10120), .Z(
        P1_U3542) );
  AOI211_X1 U10985 ( .C1(n10059), .C2(n9806), .A(n9805), .B(n9804), .ZN(n9807)
         );
  OAI21_X1 U10986 ( .B1(n9808), .B2(n10061), .A(n9807), .ZN(n9826) );
  MUX2_X1 U10987 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9826), .S(n10120), .Z(
        P1_U3541) );
  AOI21_X1 U10988 ( .B1(n10059), .B2(n9810), .A(n9809), .ZN(n9811) );
  OAI211_X1 U10989 ( .C1(n9813), .C2(n10061), .A(n9812), .B(n9811), .ZN(n9827)
         );
  MUX2_X1 U10990 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9827), .S(n10120), .Z(
        P1_U3540) );
  MUX2_X1 U10991 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9814), .S(n10098), .Z(
        P1_U3521) );
  MUX2_X1 U10992 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9815), .S(n10098), .Z(
        P1_U3520) );
  MUX2_X1 U10993 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9816), .S(n10098), .Z(
        P1_U3519) );
  MUX2_X1 U10994 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9817), .S(n10098), .Z(
        P1_U3518) );
  MUX2_X1 U10995 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9818), .S(n10098), .Z(
        P1_U3517) );
  MUX2_X1 U10996 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9819), .S(n10098), .Z(
        P1_U3516) );
  MUX2_X1 U10997 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9820), .S(n10098), .Z(
        P1_U3515) );
  MUX2_X1 U10998 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9821), .S(n10098), .Z(
        P1_U3514) );
  MUX2_X1 U10999 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9822), .S(n10098), .Z(
        P1_U3513) );
  MUX2_X1 U11000 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9823), .S(n10098), .Z(
        P1_U3512) );
  MUX2_X1 U11001 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9824), .S(n10098), .Z(
        P1_U3511) );
  MUX2_X1 U11002 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9825), .S(n10098), .Z(
        P1_U3510) );
  MUX2_X1 U11003 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9826), .S(n10098), .Z(
        P1_U3509) );
  MUX2_X1 U11004 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9827), .S(n10098), .Z(
        P1_U3507) );
  MUX2_X1 U11005 ( .A(P1_D_REG_0__SCAN_IN), .B(n9829), .S(n9828), .Z(P1_U3439)
         );
  NOR4_X1 U11006 ( .A1(n9830), .A2(P1_IR_REG_30__SCAN_IN), .A3(n5921), .A4(
        P1_U3086), .ZN(n9831) );
  AOI21_X1 U11007 ( .B1(n9832), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9831), .ZN(
        n9833) );
  OAI21_X1 U11008 ( .B1(n9835), .B2(n9834), .A(n9833), .ZN(P1_U3324) );
  MUX2_X1 U11009 ( .A(n9836), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U11010 ( .A(n10234), .ZN(n10199) );
  NOR2_X1 U11011 ( .A1(n9837), .A2(n10199), .ZN(n9838) );
  AOI211_X1 U11012 ( .C1(n10233), .C2(n9840), .A(n9839), .B(n9838), .ZN(n9842)
         );
  AOI22_X1 U11013 ( .A1(n10261), .A2(n9842), .B1(n9841), .B2(n6692), .ZN(
        P2_U3472) );
  INV_X1 U11014 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9843) );
  AOI22_X1 U11015 ( .A1(n10240), .A2(n9843), .B1(n9842), .B2(n10238), .ZN(
        P2_U3429) );
  OAI211_X1 U11016 ( .C1(n9846), .C2(n10091), .A(n9845), .B(n9844), .ZN(n9847)
         );
  AOI21_X1 U11017 ( .B1(n9848), .B2(n10095), .A(n9847), .ZN(n9864) );
  AOI22_X1 U11018 ( .A1(n10120), .A2(n9864), .B1(n9538), .B2(n10118), .ZN(
        P1_U3539) );
  NOR3_X1 U11019 ( .A1(n9850), .A2(n9849), .A3(n10061), .ZN(n9855) );
  OAI211_X1 U11020 ( .C1(n9853), .C2(n10091), .A(n9852), .B(n9851), .ZN(n9854)
         );
  NOR2_X1 U11021 ( .A1(n9855), .A2(n9854), .ZN(n9866) );
  AOI22_X1 U11022 ( .A1(n10120), .A2(n9866), .B1(n9856), .B2(n10118), .ZN(
        P1_U3538) );
  OAI211_X1 U11023 ( .C1(n9859), .C2(n10091), .A(n9858), .B(n9857), .ZN(n9860)
         );
  AOI21_X1 U11024 ( .B1(n9861), .B2(n10095), .A(n9860), .ZN(n9868) );
  INV_X1 U11025 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9862) );
  AOI22_X1 U11026 ( .A1(n10120), .A2(n9868), .B1(n9862), .B2(n10118), .ZN(
        P1_U3537) );
  INV_X1 U11027 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9863) );
  AOI22_X1 U11028 ( .A1(n10098), .A2(n9864), .B1(n9863), .B2(n10097), .ZN(
        P1_U3504) );
  INV_X1 U11029 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9865) );
  AOI22_X1 U11030 ( .A1(n10098), .A2(n9866), .B1(n9865), .B2(n10097), .ZN(
        P1_U3501) );
  INV_X1 U11031 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9867) );
  AOI22_X1 U11032 ( .A1(n10098), .A2(n9868), .B1(n9867), .B2(n10097), .ZN(
        P1_U3498) );
  XNOR2_X1 U11033 ( .A(P1_WR_REG_SCAN_IN), .B(P2_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11034 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U11035 ( .A(n9869), .ZN(n9874) );
  NAND2_X1 U11036 ( .A1(n4426), .A2(n5953), .ZN(n9872) );
  NAND2_X1 U11037 ( .A1(n9870), .A2(n9872), .ZN(n9871) );
  MUX2_X1 U11038 ( .A(n9872), .B(n9871), .S(P1_IR_REG_0__SCAN_IN), .Z(n9873)
         );
  NAND2_X1 U11039 ( .A1(n9874), .A2(n9873), .ZN(n9876) );
  AOI22_X1 U11040 ( .A1(n9878), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9875) );
  OAI21_X1 U11041 ( .B1(n9877), .B2(n9876), .A(n9875), .ZN(P1_U3243) );
  AOI22_X1 U11042 ( .A1(n9878), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9893) );
  AOI211_X1 U11043 ( .C1(n9882), .C2(n9881), .A(n9880), .B(n9879), .ZN(n9883)
         );
  AOI21_X1 U11044 ( .B1(n9885), .B2(n9884), .A(n9883), .ZN(n9892) );
  NOR2_X1 U11045 ( .A1(n9886), .A2(n5953), .ZN(n9890) );
  OAI211_X1 U11046 ( .C1(n9890), .C2(n9889), .A(n9888), .B(n9887), .ZN(n9891)
         );
  NAND3_X1 U11047 ( .A1(n9893), .A2(n9892), .A3(n9891), .ZN(P1_U3244) );
  NAND2_X1 U11048 ( .A1(n9895), .A2(n9894), .ZN(n9897) );
  XNOR2_X1 U11049 ( .A(n9897), .B(n9896), .ZN(n9900) );
  INV_X1 U11050 ( .A(n9898), .ZN(n9899) );
  AOI21_X1 U11051 ( .B1(n9900), .B2(n9980), .A(n9899), .ZN(n10086) );
  AOI222_X1 U11052 ( .A1(n9905), .A2(n9981), .B1(P1_REG2_REG_13__SCAN_IN), 
        .B2(n9992), .C1(n9983), .C2(n9901), .ZN(n9909) );
  XNOR2_X1 U11053 ( .A(n9903), .B(n9902), .ZN(n10088) );
  OAI211_X1 U11054 ( .C1(n4662), .C2(n4627), .A(n9985), .B(n9906), .ZN(n10085)
         );
  INV_X1 U11055 ( .A(n10085), .ZN(n9907) );
  AOI22_X1 U11056 ( .A1(n10088), .A2(n9968), .B1(n9967), .B2(n9907), .ZN(n9908) );
  OAI211_X1 U11057 ( .C1(n9992), .C2(n10086), .A(n9909), .B(n9908), .ZN(
        P1_U3280) );
  XNOR2_X1 U11058 ( .A(n9911), .B(n9910), .ZN(n10077) );
  INV_X1 U11059 ( .A(n10048), .ZN(n9918) );
  INV_X1 U11060 ( .A(n7645), .ZN(n9912) );
  AOI211_X1 U11061 ( .C1(n9915), .C2(n9914), .A(n9913), .B(n9912), .ZN(n9917)
         );
  AOI211_X1 U11062 ( .C1(n10077), .C2(n9918), .A(n9917), .B(n9916), .ZN(n10074) );
  AOI222_X1 U11063 ( .A1(n9920), .A2(n9981), .B1(P1_REG2_REG_11__SCAN_IN), 
        .B2(n9947), .C1(n9983), .C2(n9919), .ZN(n9924) );
  INV_X1 U11064 ( .A(n9988), .ZN(n9939) );
  OAI211_X1 U11065 ( .C1(n9921), .C2(n10073), .A(n9985), .B(n7651), .ZN(n10072) );
  INV_X1 U11066 ( .A(n10072), .ZN(n9922) );
  AOI22_X1 U11067 ( .A1(n10077), .A2(n9939), .B1(n9967), .B2(n9922), .ZN(n9923) );
  OAI211_X1 U11068 ( .C1(n9992), .C2(n10074), .A(n9924), .B(n9923), .ZN(
        P1_U3282) );
  OAI21_X1 U11069 ( .B1(n4427), .B2(n9926), .A(n9925), .ZN(n9932) );
  INV_X1 U11070 ( .A(n9927), .ZN(n9931) );
  XOR2_X1 U11071 ( .A(n9929), .B(n4427), .Z(n9935) );
  NOR2_X1 U11072 ( .A1(n9935), .A2(n10048), .ZN(n9930) );
  AOI211_X1 U11073 ( .C1(n9980), .C2(n9932), .A(n9931), .B(n9930), .ZN(n10043)
         );
  AOI222_X1 U11074 ( .A1(n9934), .A2(n9981), .B1(P1_REG2_REG_7__SCAN_IN), .B2(
        n9992), .C1(n9983), .C2(n9933), .ZN(n9941) );
  INV_X1 U11075 ( .A(n9935), .ZN(n10046) );
  OAI211_X1 U11076 ( .C1(n9937), .C2(n10042), .A(n9985), .B(n9936), .ZN(n10041) );
  INV_X1 U11077 ( .A(n10041), .ZN(n9938) );
  AOI22_X1 U11078 ( .A1(n10046), .A2(n9939), .B1(n9967), .B2(n9938), .ZN(n9940) );
  OAI211_X1 U11079 ( .C1(n9992), .C2(n10043), .A(n9941), .B(n9940), .ZN(
        P1_U3286) );
  XOR2_X1 U11080 ( .A(n9950), .B(n9942), .Z(n9945) );
  INV_X1 U11081 ( .A(n9943), .ZN(n9944) );
  AOI21_X1 U11082 ( .B1(n9945), .B2(n9980), .A(n9944), .ZN(n10029) );
  AOI222_X1 U11083 ( .A1(n9948), .A2(n9981), .B1(P1_REG2_REG_5__SCAN_IN), .B2(
        n9947), .C1(n9983), .C2(n9946), .ZN(n9956) );
  XNOR2_X1 U11084 ( .A(n9949), .B(n9950), .ZN(n10032) );
  INV_X1 U11085 ( .A(n9952), .ZN(n9953) );
  OAI211_X1 U11086 ( .C1(n10028), .C2(n4665), .A(n9953), .B(n9985), .ZN(n10027) );
  INV_X1 U11087 ( .A(n10027), .ZN(n9954) );
  AOI22_X1 U11088 ( .A1(n10032), .A2(n9968), .B1(n9967), .B2(n9954), .ZN(n9955) );
  OAI211_X1 U11089 ( .C1(n9992), .C2(n10029), .A(n9956), .B(n9955), .ZN(
        P1_U3288) );
  XOR2_X1 U11090 ( .A(n9963), .B(n9957), .Z(n9959) );
  AOI21_X1 U11091 ( .B1(n9959), .B2(n9980), .A(n9958), .ZN(n10016) );
  INV_X1 U11092 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9961) );
  AOI222_X1 U11093 ( .A1(n9961), .A2(n9983), .B1(n9992), .B2(
        P1_REG2_REG_3__SCAN_IN), .C1(n9960), .C2(n9981), .ZN(n9970) );
  XNOR2_X1 U11094 ( .A(n9963), .B(n9962), .ZN(n10019) );
  OAI211_X1 U11095 ( .C1(n9965), .C2(n10015), .A(n9964), .B(n9985), .ZN(n10014) );
  INV_X1 U11096 ( .A(n10014), .ZN(n9966) );
  AOI22_X1 U11097 ( .A1(n10019), .A2(n9968), .B1(n9967), .B2(n9966), .ZN(n9969) );
  OAI211_X1 U11098 ( .C1(n9992), .C2(n10016), .A(n9970), .B(n9969), .ZN(
        P1_U3290) );
  OAI21_X1 U11099 ( .B1(n9973), .B2(n9972), .A(n9971), .ZN(n9979) );
  INV_X1 U11100 ( .A(n9974), .ZN(n9975) );
  XNOR2_X1 U11101 ( .A(n9976), .B(n9975), .ZN(n10001) );
  NOR2_X1 U11102 ( .A1(n10001), .A2(n10048), .ZN(n9977) );
  AOI211_X1 U11103 ( .C1(n9980), .C2(n9979), .A(n9978), .B(n9977), .ZN(n10003)
         );
  AOI222_X1 U11104 ( .A1(P1_REG2_REG_1__SCAN_IN), .A2(n9992), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n9983), .C1(n9982), .C2(n9981), .ZN(n9991) );
  OAI211_X1 U11105 ( .C1(n9986), .C2(n7439), .A(n9985), .B(n9984), .ZN(n10002)
         );
  OAI22_X1 U11106 ( .A1(n9988), .A2(n10001), .B1(n9987), .B2(n10002), .ZN(
        n9989) );
  INV_X1 U11107 ( .A(n9989), .ZN(n9990) );
  OAI211_X1 U11108 ( .C1(n9992), .C2(n10003), .A(n9991), .B(n9990), .ZN(
        P1_U3292) );
  AND2_X1 U11109 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9999), .ZN(P1_U3294) );
  AND2_X1 U11110 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9999), .ZN(P1_U3295) );
  NOR2_X1 U11111 ( .A1(n9998), .A2(n9993), .ZN(P1_U3296) );
  AND2_X1 U11112 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9999), .ZN(P1_U3297) );
  AND2_X1 U11113 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9999), .ZN(P1_U3298) );
  NOR2_X1 U11114 ( .A1(n9998), .A2(n9994), .ZN(P1_U3299) );
  AND2_X1 U11115 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9999), .ZN(P1_U3300) );
  AND2_X1 U11116 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9999), .ZN(P1_U3301) );
  AND2_X1 U11117 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9999), .ZN(P1_U3302) );
  AND2_X1 U11118 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9999), .ZN(P1_U3303) );
  NOR2_X1 U11119 ( .A1(n9998), .A2(n9995), .ZN(P1_U3304) );
  AND2_X1 U11120 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9999), .ZN(P1_U3305) );
  AND2_X1 U11121 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9999), .ZN(P1_U3306) );
  AND2_X1 U11122 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9999), .ZN(P1_U3307) );
  AND2_X1 U11123 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9999), .ZN(P1_U3308) );
  NOR2_X1 U11124 ( .A1(n9998), .A2(n9996), .ZN(P1_U3309) );
  AND2_X1 U11125 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9999), .ZN(P1_U3310) );
  AND2_X1 U11126 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9999), .ZN(P1_U3311) );
  AND2_X1 U11127 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9999), .ZN(P1_U3312) );
  AND2_X1 U11128 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9999), .ZN(P1_U3313) );
  AND2_X1 U11129 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9999), .ZN(P1_U3314) );
  AND2_X1 U11130 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9999), .ZN(P1_U3315) );
  AND2_X1 U11131 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9999), .ZN(P1_U3316) );
  AND2_X1 U11132 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9999), .ZN(P1_U3317) );
  AND2_X1 U11133 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9999), .ZN(P1_U3318) );
  AND2_X1 U11134 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9999), .ZN(P1_U3319) );
  AND2_X1 U11135 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9999), .ZN(P1_U3320) );
  NOR2_X1 U11136 ( .A1(n9998), .A2(n9997), .ZN(P1_U3321) );
  AND2_X1 U11137 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9999), .ZN(P1_U3322) );
  AND2_X1 U11138 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9999), .ZN(P1_U3323) );
  INV_X1 U11139 ( .A(n10000), .ZN(n10078) );
  INV_X1 U11140 ( .A(n10001), .ZN(n10006) );
  OAI21_X1 U11141 ( .B1(n7439), .B2(n10091), .A(n10002), .ZN(n10005) );
  INV_X1 U11142 ( .A(n10003), .ZN(n10004) );
  AOI211_X1 U11143 ( .C1(n10078), .C2(n10006), .A(n10005), .B(n10004), .ZN(
        n10100) );
  AOI22_X1 U11144 ( .A1(n10098), .A2(n10100), .B1(n10007), .B2(n10097), .ZN(
        P1_U3456) );
  NAND2_X1 U11145 ( .A1(n10059), .A2(n7442), .ZN(n10008) );
  AND2_X1 U11146 ( .A1(n10009), .A2(n10008), .ZN(n10012) );
  NAND2_X1 U11147 ( .A1(n10010), .A2(n10095), .ZN(n10011) );
  AND3_X1 U11148 ( .A1(n10013), .A2(n10012), .A3(n10011), .ZN(n10101) );
  AOI22_X1 U11149 ( .A1(n10098), .A2(n10101), .B1(n5966), .B2(n10097), .ZN(
        P1_U3459) );
  OAI21_X1 U11150 ( .B1(n10015), .B2(n10091), .A(n10014), .ZN(n10018) );
  INV_X1 U11151 ( .A(n10016), .ZN(n10017) );
  AOI211_X1 U11152 ( .C1(n10019), .C2(n10095), .A(n10018), .B(n10017), .ZN(
        n10102) );
  AOI22_X1 U11153 ( .A1(n10098), .A2(n10102), .B1(n5988), .B2(n10097), .ZN(
        P1_U3462) );
  OAI21_X1 U11154 ( .B1(n10021), .B2(n10091), .A(n10020), .ZN(n10022) );
  AOI21_X1 U11155 ( .B1(n10023), .B2(n10095), .A(n10022), .ZN(n10024) );
  AND2_X1 U11156 ( .A1(n10025), .A2(n10024), .ZN(n10104) );
  INV_X1 U11157 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10026) );
  AOI22_X1 U11158 ( .A1(n10098), .A2(n10104), .B1(n10026), .B2(n10097), .ZN(
        P1_U3465) );
  OAI21_X1 U11159 ( .B1(n10028), .B2(n10091), .A(n10027), .ZN(n10031) );
  INV_X1 U11160 ( .A(n10029), .ZN(n10030) );
  AOI211_X1 U11161 ( .C1(n10095), .C2(n10032), .A(n10031), .B(n10030), .ZN(
        n10105) );
  INV_X1 U11162 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10033) );
  AOI22_X1 U11163 ( .A1(n10098), .A2(n10105), .B1(n10033), .B2(n10097), .ZN(
        P1_U3468) );
  OAI21_X1 U11164 ( .B1(n10035), .B2(n10091), .A(n10034), .ZN(n10036) );
  AOI21_X1 U11165 ( .B1(n10037), .B2(n10095), .A(n10036), .ZN(n10038) );
  AND2_X1 U11166 ( .A1(n10039), .A2(n10038), .ZN(n10107) );
  INV_X1 U11167 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10040) );
  AOI22_X1 U11168 ( .A1(n10098), .A2(n10107), .B1(n10040), .B2(n10097), .ZN(
        P1_U3471) );
  OAI21_X1 U11169 ( .B1(n10042), .B2(n10091), .A(n10041), .ZN(n10045) );
  INV_X1 U11170 ( .A(n10043), .ZN(n10044) );
  AOI211_X1 U11171 ( .C1(n10078), .C2(n10046), .A(n10045), .B(n10044), .ZN(
        n10109) );
  AOI22_X1 U11172 ( .A1(n10098), .A2(n10109), .B1(n10047), .B2(n10097), .ZN(
        P1_U3474) );
  INV_X1 U11173 ( .A(n10049), .ZN(n10055) );
  NOR2_X1 U11174 ( .A1(n10049), .A2(n10048), .ZN(n10054) );
  OAI211_X1 U11175 ( .C1(n10052), .C2(n10091), .A(n10051), .B(n10050), .ZN(
        n10053) );
  AOI211_X1 U11176 ( .C1(n10078), .C2(n10055), .A(n10054), .B(n10053), .ZN(
        n10111) );
  INV_X1 U11177 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10056) );
  AOI22_X1 U11178 ( .A1(n10098), .A2(n10111), .B1(n10056), .B2(n10097), .ZN(
        P1_U3477) );
  AOI21_X1 U11179 ( .B1(n10059), .B2(n10058), .A(n10057), .ZN(n10060) );
  OAI21_X1 U11180 ( .B1(n10062), .B2(n10061), .A(n10060), .ZN(n10064) );
  NOR2_X1 U11181 ( .A1(n10064), .A2(n10063), .ZN(n10113) );
  INV_X1 U11182 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10065) );
  AOI22_X1 U11183 ( .A1(n10098), .A2(n10113), .B1(n10065), .B2(n10097), .ZN(
        P1_U3480) );
  OAI211_X1 U11184 ( .C1(n10068), .C2(n10091), .A(n10067), .B(n10066), .ZN(
        n10069) );
  AOI21_X1 U11185 ( .B1(n10070), .B2(n10095), .A(n10069), .ZN(n10114) );
  AOI22_X1 U11186 ( .A1(n10098), .A2(n10114), .B1(n10071), .B2(n10097), .ZN(
        P1_U3483) );
  OAI21_X1 U11187 ( .B1(n10073), .B2(n10091), .A(n10072), .ZN(n10076) );
  INV_X1 U11188 ( .A(n10074), .ZN(n10075) );
  AOI211_X1 U11189 ( .C1(n10078), .C2(n10077), .A(n10076), .B(n10075), .ZN(
        n10115) );
  INV_X1 U11190 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10079) );
  AOI22_X1 U11191 ( .A1(n10098), .A2(n10115), .B1(n10079), .B2(n10097), .ZN(
        P1_U3486) );
  OAI21_X1 U11192 ( .B1(n10081), .B2(n10091), .A(n10080), .ZN(n10082) );
  AOI211_X1 U11193 ( .C1(n10084), .C2(n10095), .A(n10083), .B(n10082), .ZN(
        n10116) );
  AOI22_X1 U11194 ( .A1(n10098), .A2(n10116), .B1(n6173), .B2(n10097), .ZN(
        P1_U3489) );
  OAI211_X1 U11195 ( .C1(n4627), .C2(n10091), .A(n10086), .B(n10085), .ZN(
        n10087) );
  AOI21_X1 U11196 ( .B1(n10088), .B2(n10095), .A(n10087), .ZN(n10117) );
  INV_X1 U11197 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10089) );
  AOI22_X1 U11198 ( .A1(n10098), .A2(n10117), .B1(n10089), .B2(n10097), .ZN(
        P1_U3492) );
  OAI21_X1 U11199 ( .B1(n10092), .B2(n10091), .A(n10090), .ZN(n10093) );
  AOI211_X1 U11200 ( .C1(n10096), .C2(n10095), .A(n10094), .B(n10093), .ZN(
        n10119) );
  AOI22_X1 U11201 ( .A1(n10098), .A2(n10119), .B1(n6207), .B2(n10097), .ZN(
        P1_U3495) );
  AOI22_X1 U11202 ( .A1(n10120), .A2(n10100), .B1(n10099), .B2(n10118), .ZN(
        P1_U3523) );
  AOI22_X1 U11203 ( .A1(n10120), .A2(n10101), .B1(n5967), .B2(n10118), .ZN(
        P1_U3524) );
  AOI22_X1 U11204 ( .A1(n10120), .A2(n10102), .B1(n7034), .B2(n10118), .ZN(
        P1_U3525) );
  AOI22_X1 U11205 ( .A1(n10120), .A2(n10104), .B1(n10103), .B2(n10118), .ZN(
        P1_U3526) );
  AOI22_X1 U11206 ( .A1(n10120), .A2(n10105), .B1(n7032), .B2(n10118), .ZN(
        P1_U3527) );
  AOI22_X1 U11207 ( .A1(n10120), .A2(n10107), .B1(n10106), .B2(n10118), .ZN(
        P1_U3528) );
  AOI22_X1 U11208 ( .A1(n10120), .A2(n10109), .B1(n10108), .B2(n10118), .ZN(
        P1_U3529) );
  AOI22_X1 U11209 ( .A1(n10120), .A2(n10111), .B1(n10110), .B2(n10118), .ZN(
        P1_U3530) );
  AOI22_X1 U11210 ( .A1(n10120), .A2(n10113), .B1(n10112), .B2(n10118), .ZN(
        P1_U3531) );
  AOI22_X1 U11211 ( .A1(n10120), .A2(n10114), .B1(n7340), .B2(n10118), .ZN(
        P1_U3532) );
  AOI22_X1 U11212 ( .A1(n10120), .A2(n10115), .B1(n7561), .B2(n10118), .ZN(
        P1_U3533) );
  AOI22_X1 U11213 ( .A1(n10120), .A2(n10116), .B1(n6170), .B2(n10118), .ZN(
        P1_U3534) );
  AOI22_X1 U11214 ( .A1(n10120), .A2(n10117), .B1(n7924), .B2(n10118), .ZN(
        P1_U3535) );
  AOI22_X1 U11215 ( .A1(n10120), .A2(n10119), .B1(n9489), .B2(n10118), .ZN(
        P1_U3536) );
  AOI22_X1 U11216 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n10141), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .ZN(n10125) );
  XNOR2_X1 U11217 ( .A(n10121), .B(P2_IR_REG_0__SCAN_IN), .ZN(n10122) );
  OAI21_X1 U11218 ( .B1(n10123), .B2(n10152), .A(n10122), .ZN(n10124) );
  OAI211_X1 U11219 ( .C1(n10162), .C2(n4762), .A(n10125), .B(n10124), .ZN(
        P2_U3182) );
  OAI21_X1 U11220 ( .B1(n10128), .B2(n10127), .A(n10126), .ZN(n10129) );
  AND2_X1 U11221 ( .A1(n10129), .A2(n10152), .ZN(n10137) );
  AOI21_X1 U11222 ( .B1(n4518), .B2(n10131), .A(n10130), .ZN(n10135) );
  AOI21_X1 U11223 ( .B1(n4519), .B2(n10133), .A(n10132), .ZN(n10134) );
  OAI22_X1 U11224 ( .A1(n10156), .A2(n10135), .B1(n10134), .B2(n10147), .ZN(
        n10136) );
  AOI211_X1 U11225 ( .C1(P2_ADDR_REG_8__SCAN_IN), .C2(n10141), .A(n10137), .B(
        n10136), .ZN(n10139) );
  OAI211_X1 U11226 ( .C1(n10162), .C2(n10140), .A(n10139), .B(n10138), .ZN(
        P2_U3190) );
  AOI22_X1 U11227 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n10141), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(P2_U3151), .ZN(n10160) );
  AOI21_X1 U11228 ( .B1(n4511), .B2(n10143), .A(n10142), .ZN(n10157) );
  AOI21_X1 U11229 ( .B1(n10146), .B2(n10145), .A(n10144), .ZN(n10148) );
  OR2_X1 U11230 ( .A1(n10148), .A2(n10147), .ZN(n10155) );
  OAI21_X1 U11231 ( .B1(n10151), .B2(n10150), .A(n10149), .ZN(n10153) );
  NAND2_X1 U11232 ( .A1(n10153), .A2(n10152), .ZN(n10154) );
  OAI211_X1 U11233 ( .C1(n10157), .C2(n10156), .A(n10155), .B(n10154), .ZN(
        n10158) );
  INV_X1 U11234 ( .A(n10158), .ZN(n10159) );
  OAI211_X1 U11235 ( .C1(n10162), .C2(n10161), .A(n10160), .B(n10159), .ZN(
        P2_U3196) );
  OAI21_X1 U11236 ( .B1(n10164), .B2(n4543), .A(n10163), .ZN(n10185) );
  OAI22_X1 U11237 ( .A1(n10182), .A2(n10167), .B1(n10166), .B2(n10165), .ZN(
        n10172) );
  XNOR2_X1 U11238 ( .A(n10168), .B(n4543), .ZN(n10169) );
  OAI222_X1 U11239 ( .A1(n10171), .A2(n10170), .B1(n5626), .B2(n5756), .C1(
        n5628), .C2(n10169), .ZN(n10183) );
  AOI211_X1 U11240 ( .C1(n10173), .C2(n10185), .A(n10172), .B(n10183), .ZN(
        n10175) );
  AOI22_X1 U11241 ( .A1(n10176), .A2(n6570), .B1(n10175), .B2(n10174), .ZN(
        P2_U3231) );
  INV_X1 U11242 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10181) );
  INV_X1 U11243 ( .A(n10177), .ZN(n10180) );
  OAI22_X1 U11244 ( .A1(n10178), .A2(n10205), .B1(n5136), .B2(n10226), .ZN(
        n10179) );
  NOR2_X1 U11245 ( .A1(n10180), .A2(n10179), .ZN(n10242) );
  AOI22_X1 U11246 ( .A1(n10240), .A2(n10181), .B1(n10242), .B2(n10238), .ZN(
        P2_U3393) );
  INV_X1 U11247 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10186) );
  NOR2_X1 U11248 ( .A1(n10182), .A2(n10226), .ZN(n10184) );
  AOI211_X1 U11249 ( .C1(n10234), .C2(n10185), .A(n10184), .B(n10183), .ZN(
        n10243) );
  AOI22_X1 U11250 ( .A1(n10240), .A2(n10186), .B1(n10243), .B2(n10238), .ZN(
        P2_U3396) );
  INV_X1 U11251 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10192) );
  INV_X1 U11252 ( .A(n10187), .ZN(n10191) );
  OAI21_X1 U11253 ( .B1(n10189), .B2(n10226), .A(n10188), .ZN(n10190) );
  AOI21_X1 U11254 ( .B1(n10191), .B2(n10234), .A(n10190), .ZN(n10245) );
  AOI22_X1 U11255 ( .A1(n10240), .A2(n10192), .B1(n10245), .B2(n10238), .ZN(
        P2_U3402) );
  INV_X1 U11256 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10197) );
  OAI21_X1 U11257 ( .B1(n10194), .B2(n10226), .A(n10193), .ZN(n10195) );
  AOI21_X1 U11258 ( .B1(n10234), .B2(n10196), .A(n10195), .ZN(n10247) );
  AOI22_X1 U11259 ( .A1(n10240), .A2(n10197), .B1(n10247), .B2(n10238), .ZN(
        P2_U3405) );
  INV_X1 U11260 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10203) );
  OAI22_X1 U11261 ( .A1(n10200), .A2(n10199), .B1(n10198), .B2(n10226), .ZN(
        n10202) );
  NOR2_X1 U11262 ( .A1(n10202), .A2(n10201), .ZN(n10249) );
  AOI22_X1 U11263 ( .A1(n10240), .A2(n10203), .B1(n10249), .B2(n10238), .ZN(
        P2_U3408) );
  INV_X1 U11264 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10209) );
  OAI22_X1 U11265 ( .A1(n10206), .A2(n10205), .B1(n10204), .B2(n10226), .ZN(
        n10207) );
  NOR2_X1 U11266 ( .A1(n10208), .A2(n10207), .ZN(n10251) );
  AOI22_X1 U11267 ( .A1(n10240), .A2(n10209), .B1(n10251), .B2(n10238), .ZN(
        P2_U3411) );
  INV_X1 U11268 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10214) );
  NOR2_X1 U11269 ( .A1(n10210), .A2(n10226), .ZN(n10212) );
  AOI211_X1 U11270 ( .C1(n10234), .C2(n10213), .A(n10212), .B(n10211), .ZN(
        n10253) );
  AOI22_X1 U11271 ( .A1(n10240), .A2(n10214), .B1(n10253), .B2(n10238), .ZN(
        P2_U3414) );
  INV_X1 U11272 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10220) );
  AOI22_X1 U11273 ( .A1(n10217), .A2(n10216), .B1(n10233), .B2(n10215), .ZN(
        n10218) );
  AND2_X1 U11274 ( .A1(n10219), .A2(n10218), .ZN(n10255) );
  AOI22_X1 U11275 ( .A1(n10240), .A2(n10220), .B1(n10255), .B2(n10238), .ZN(
        P2_U3417) );
  OAI21_X1 U11276 ( .B1(n10222), .B2(n10226), .A(n10221), .ZN(n10223) );
  AOI21_X1 U11277 ( .B1(n10234), .B2(n10224), .A(n10223), .ZN(n10257) );
  AOI22_X1 U11278 ( .A1(n10240), .A2(n10225), .B1(n10257), .B2(n10238), .ZN(
        P2_U3420) );
  INV_X1 U11279 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10231) );
  NOR2_X1 U11280 ( .A1(n10227), .A2(n10226), .ZN(n10229) );
  AOI211_X1 U11281 ( .C1(n10234), .C2(n10230), .A(n10229), .B(n10228), .ZN(
        n10259) );
  AOI22_X1 U11282 ( .A1(n10240), .A2(n10231), .B1(n10259), .B2(n10238), .ZN(
        P2_U3423) );
  INV_X1 U11283 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10239) );
  AOI22_X1 U11284 ( .A1(n10235), .A2(n10234), .B1(n10233), .B2(n10232), .ZN(
        n10237) );
  AND2_X1 U11285 ( .A1(n10237), .A2(n10236), .ZN(n10260) );
  AOI22_X1 U11286 ( .A1(n10240), .A2(n10239), .B1(n10260), .B2(n10238), .ZN(
        P2_U3426) );
  AOI22_X1 U11287 ( .A1(n10261), .A2(n10242), .B1(n10241), .B2(n6692), .ZN(
        P2_U3460) );
  AOI22_X1 U11288 ( .A1(n10261), .A2(n10243), .B1(n6532), .B2(n6692), .ZN(
        P2_U3461) );
  INV_X1 U11289 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10244) );
  AOI22_X1 U11290 ( .A1(n10261), .A2(n10245), .B1(n10244), .B2(n6692), .ZN(
        P2_U3463) );
  AOI22_X1 U11291 ( .A1(n10261), .A2(n10247), .B1(n10246), .B2(n6692), .ZN(
        P2_U3464) );
  AOI22_X1 U11292 ( .A1(n10261), .A2(n10249), .B1(n10248), .B2(n6692), .ZN(
        P2_U3465) );
  AOI22_X1 U11293 ( .A1(n10261), .A2(n10251), .B1(n10250), .B2(n6692), .ZN(
        P2_U3466) );
  INV_X1 U11294 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10252) );
  AOI22_X1 U11295 ( .A1(n10261), .A2(n10253), .B1(n10252), .B2(n6692), .ZN(
        P2_U3467) );
  AOI22_X1 U11296 ( .A1(n10261), .A2(n10255), .B1(n10254), .B2(n6692), .ZN(
        P2_U3468) );
  AOI22_X1 U11297 ( .A1(n10261), .A2(n10257), .B1(n10256), .B2(n6692), .ZN(
        P2_U3469) );
  AOI22_X1 U11298 ( .A1(n10261), .A2(n10259), .B1(n10258), .B2(n6692), .ZN(
        P2_U3470) );
  AOI22_X1 U11299 ( .A1(n10261), .A2(n10260), .B1(n6552), .B2(n6692), .ZN(
        P2_U3471) );
  NAND2_X1 U11300 ( .A1(n10263), .A2(n10262), .ZN(n10264) );
  XOR2_X1 U11301 ( .A(n10265), .B(n10264), .Z(ADD_1068_U5) );
  AOI22_X1 U11302 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .B1(n10267), .B2(n10266), .ZN(ADD_1068_U46) );
  OAI21_X1 U11303 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n10269), .A(n10268), 
        .ZN(n10271) );
  XOR2_X1 U11304 ( .A(n10271), .B(n10270), .Z(ADD_1068_U55) );
  XNOR2_X1 U11305 ( .A(n10273), .B(n10272), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11306 ( .A(n10275), .B(n10274), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11307 ( .A(n10277), .B(n10276), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11308 ( .A(n10279), .B(n10278), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11309 ( .A(n10281), .B(n10280), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11310 ( .A(n10283), .B(n10282), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11311 ( .A(n10285), .B(n10284), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11312 ( .A(n10287), .B(n10286), .ZN(ADD_1068_U63) );
  XNOR2_X1 U11313 ( .A(n10289), .B(n10288), .ZN(ADD_1068_U50) );
  XNOR2_X1 U11314 ( .A(n10291), .B(n10290), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11315 ( .A(n10293), .B(n10292), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11316 ( .A(n10295), .B(n10294), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11317 ( .A(n10297), .B(n10296), .ZN(ADD_1068_U48) );
  XOR2_X1 U11318 ( .A(n10299), .B(n10298), .Z(ADD_1068_U54) );
  XOR2_X1 U11319 ( .A(n10301), .B(n10300), .Z(ADD_1068_U53) );
  XNOR2_X1 U11320 ( .A(n10303), .B(n10302), .ZN(ADD_1068_U52) );
  INV_X1 U4928 ( .A(n5296), .ZN(n8396) );
  CLKBUF_X1 U4942 ( .A(n5987), .Z(n6742) );
  CLKBUF_X1 U4943 ( .A(n9928), .Z(n4427) );
endmodule

