

module b20_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, 
        SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, 
        SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, 
        SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, 
        P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104;

  INV_X4 U5172 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NAND4_X1 U5173 ( .A1(n5781), .A2(n5780), .A3(n5779), .A4(n5778), .ZN(n10168)
         );
  NAND2_X1 U5174 ( .A1(n6711), .A2(n8849), .ZN(n7207) );
  NAND2_X1 U5175 ( .A1(n6234), .A2(n6227), .ZN(n7032) );
  INV_X1 U5176 ( .A(n6951), .ZN(n6953) );
  INV_X2 U5177 ( .A(n9889), .ZN(n5825) );
  NAND2_X1 U5178 ( .A1(n5697), .A2(n5696), .ZN(n10660) );
  AND4_X2 U5179 ( .A1(n6304), .A2(n6303), .A3(n6302), .A4(n6301), .ZN(n6951)
         );
  OR2_X1 U5180 ( .A1(n6352), .A2(n6964), .ZN(n6302) );
  AND2_X1 U5181 ( .A1(n8846), .A2(n8845), .ZN(n8852) );
  INV_X1 U5182 ( .A(n7759), .ZN(n7115) );
  INV_X1 U5183 ( .A(n6803), .ZN(n5987) );
  INV_X2 U5184 ( .A(n7079), .ZN(n9050) );
  INV_X1 U5186 ( .A(n9381), .ZN(n9415) );
  OR2_X1 U5187 ( .A1(n7494), .A2(n7738), .ZN(n8733) );
  NAND2_X1 U5188 ( .A1(n6953), .A2(n10869), .ZN(n8706) );
  INV_X1 U5189 ( .A(n9001), .ZN(n8976) );
  INV_X1 U5190 ( .A(n7115), .ZN(n8961) );
  INV_X1 U5191 ( .A(n7115), .ZN(n8938) );
  INV_X1 U5192 ( .A(n6205), .ZN(n9887) );
  XNOR2_X1 U5193 ( .A(n5184), .B(P2_IR_REG_27__SCAN_IN), .ZN(n6859) );
  NAND2_X1 U5194 ( .A1(n6529), .A2(n6528), .ZN(n9521) );
  OR2_X1 U5195 ( .A1(n6289), .A2(n6269), .ZN(n6291) );
  INV_X2 U5196 ( .A(n9885), .ZN(n6209) );
  CLKBUF_X3 U5197 ( .A(n6352), .Z(n5108) );
  OAI21_X2 U5198 ( .B1(n8852), .B2(n8851), .A(n8854), .ZN(n8853) );
  NAND2_X1 U5199 ( .A1(n9545), .A2(n9551), .ZN(n9480) );
  NAND2_X2 U5201 ( .A1(n5116), .A2(n6261), .ZN(n6442) );
  INV_X2 U5202 ( .A(n6386), .ZN(n6261) );
  NAND2_X2 U5203 ( .A1(n6336), .A2(n6335), .ZN(n7390) );
  INV_X2 U5204 ( .A(n8710), .ZN(n7206) );
  XNOR2_X2 U5205 ( .A(n5841), .B(n5840), .ZN(n6796) );
  XNOR2_X2 U5206 ( .A(n9521), .B(n9503), .ZN(n9519) );
  OR2_X1 U5207 ( .A1(n9607), .A2(n9606), .ZN(n9664) );
  AOI21_X1 U5208 ( .B1(n9385), .B2(n10928), .A(n9384), .ZN(n9603) );
  NAND2_X1 U5209 ( .A1(n5287), .A2(n5288), .ZN(n9379) );
  MUX2_X1 U5210 ( .A(n10475), .B(n10474), .S(n10529), .Z(n10476) );
  AOI21_X1 U5211 ( .B1(n8851), .B2(n9080), .A(n8692), .ZN(n8844) );
  NAND2_X1 U5212 ( .A1(n5199), .A2(n5567), .ZN(n9149) );
  NAND2_X1 U5213 ( .A1(n9573), .A2(n6485), .ZN(n9558) );
  NAND2_X1 U5214 ( .A1(n5519), .A2(n5518), .ZN(n5517) );
  NAND2_X1 U5215 ( .A1(n5202), .A2(n5201), .ZN(n9126) );
  NAND2_X1 U5216 ( .A1(n5203), .A2(n9115), .ZN(n5202) );
  OAI21_X1 U5217 ( .B1(n9864), .B2(n10158), .A(n8143), .ZN(n8152) );
  OR2_X1 U5218 ( .A1(n10491), .A2(n10375), .ZN(n6109) );
  OR2_X1 U5219 ( .A1(n6552), .A2(n6551), .ZN(n9483) );
  AND2_X1 U5220 ( .A1(n10382), .A2(n10400), .ZN(n6085) );
  OAI21_X1 U5221 ( .B1(n7928), .B2(n5590), .A(n5120), .ZN(n5200) );
  NAND2_X1 U5222 ( .A1(n6574), .A2(n6573), .ZN(n9474) );
  NAND2_X1 U5223 ( .A1(n6018), .A2(n6017), .ZN(n10432) );
  XNOR2_X1 U5224 ( .A(n6003), .B(n6002), .ZN(n7534) );
  NAND2_X1 U5225 ( .A1(n5859), .A2(n5858), .ZN(n7773) );
  NAND2_X1 U5226 ( .A1(n6413), .A2(n6412), .ZN(n10997) );
  NOR2_X1 U5227 ( .A1(n11051), .A2(n7459), .ZN(n10458) );
  INV_X1 U5228 ( .A(n7152), .ZN(n7079) );
  NAND2_X1 U5229 ( .A1(n6331), .A2(n5336), .ZN(n9204) );
  NAND2_X1 U5230 ( .A1(n5208), .A2(n6946), .ZN(n5207) );
  AND2_X1 U5231 ( .A1(n6727), .A2(n6810), .ZN(n6946) );
  NAND4_X2 U5232 ( .A1(n6318), .A2(n6317), .A3(n6316), .A4(n6315), .ZN(n10925)
         );
  OAI211_X1 U5233 ( .C1(n6313), .C2(n7338), .A(n6348), .B(n6347), .ZN(n10951)
         );
  NAND4_X1 U5234 ( .A1(n5736), .A2(n5735), .A3(n5734), .A4(n5733), .ZN(n10170)
         );
  CLKBUF_X3 U5235 ( .A(n6478), .Z(n5110) );
  INV_X1 U5236 ( .A(n10884), .ZN(n9848) );
  AND2_X1 U5237 ( .A1(n7207), .A2(n8879), .ZN(n5208) );
  INV_X1 U5238 ( .A(n6338), .ZN(n6300) );
  NAND3_X2 U5239 ( .A1(n7032), .A2(n7458), .A3(n7023), .ZN(n9001) );
  NAND2_X2 U5240 ( .A1(n7029), .A2(n7032), .ZN(n9002) );
  NAND2_X1 U5241 ( .A1(n5604), .A2(n5298), .ZN(n7148) );
  NAND4_X1 U5242 ( .A1(n5724), .A2(n5723), .A3(n5722), .A4(n5721), .ZN(n9906)
         );
  AND3_X1 U5243 ( .A1(n5743), .A2(n5742), .A3(n5741), .ZN(n10884) );
  AND3_X1 U5244 ( .A1(n5758), .A2(n5757), .A3(n5756), .ZN(n10899) );
  INV_X1 U5245 ( .A(n9718), .ZN(n6294) );
  INV_X1 U5246 ( .A(n6293), .ZN(n6292) );
  XNOR2_X1 U5247 ( .A(n6720), .B(n6719), .ZN(n8615) );
  NAND2_X1 U5248 ( .A1(n6803), .A2(n8662), .ZN(n5799) );
  XNOR2_X1 U5249 ( .A(n6288), .B(n9711), .ZN(n6293) );
  NAND2_X1 U5250 ( .A1(n6718), .A2(n6717), .ZN(n8058) );
  NAND2_X1 U5251 ( .A1(n9710), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6288) );
  INV_X2 U5252 ( .A(n6859), .ZN(n9327) );
  XNOR2_X1 U5253 ( .A(n5244), .B(n8369), .ZN(n10598) );
  INV_X1 U5254 ( .A(n6724), .ZN(n6271) );
  MUX2_X1 U5255 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5695), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n5697) );
  AND2_X1 U5256 ( .A1(n6470), .A2(n6469), .ZN(n6487) );
  NAND2_X1 U5257 ( .A1(n5696), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5694) );
  INV_X2 U5258 ( .A(n10592), .ZN(n8657) );
  NAND2_X2 U5259 ( .A1(n8662), .A2(P2_U3151), .ZN(n8618) );
  NAND2_X1 U5260 ( .A1(n6322), .A2(n6321), .ZN(n7339) );
  AND3_X1 U5261 ( .A1(n5563), .A2(n5303), .A3(n5365), .ZN(n5302) );
  AND2_X1 U5262 ( .A1(n5564), .A2(n6734), .ZN(n5563) );
  AND2_X1 U5263 ( .A1(n5132), .A2(n5565), .ZN(n5564) );
  NAND2_X1 U5264 ( .A1(n5369), .A2(n5367), .ZN(n5618) );
  NAND4_X1 U5265 ( .A1(n6511), .A2(n6265), .A3(n6264), .A4(n6263), .ZN(n6266)
         );
  AND3_X1 U5266 ( .A1(n6523), .A2(n6525), .A3(n6262), .ZN(n6511) );
  AND2_X2 U5267 ( .A1(n5182), .A2(n5181), .ZN(n6849) );
  INV_X4 U5268 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U5269 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5680) );
  NOR2_X1 U5270 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5681) );
  NOR2_X1 U5271 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5739) );
  NOR2_X4 U5272 ( .A1(n5783), .A2(n5236), .ZN(n5123) );
  INV_X2 U5273 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n5182) );
  NOR2_X1 U5274 ( .A1(n6442), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n6470) );
  NAND2_X1 U5275 ( .A1(n6724), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5184) );
  XNOR2_X2 U5276 ( .A(n5206), .B(P2_IR_REG_19__SCAN_IN), .ZN(n6711) );
  NAND2_X1 U5277 ( .A1(n6457), .A2(n6456), .ZN(n8010) );
  NAND2_X1 U5278 ( .A1(n6292), .A2(n6294), .ZN(n6352) );
  XNOR2_X2 U5279 ( .A(n10925), .B(n7206), .ZN(n7202) );
  OAI21_X2 U5280 ( .B1(n9558), .B2(n6697), .A(n8784), .ZN(n9545) );
  OAI22_X2 U5281 ( .A1(n9379), .A2(n9387), .B1(n9399), .B2(n9601), .ZN(n9015)
         );
  OAI21_X2 U5282 ( .B1(n8010), .B2(n5172), .A(n6468), .ZN(n9574) );
  NAND2_X4 U5283 ( .A1(n6669), .A2(n6668), .ZN(n6313) );
  XNOR2_X2 U5284 ( .A(n6270), .B(n6287), .ZN(n6668) );
  NAND2_X1 U5285 ( .A1(n6602), .A2(n6601), .ZN(n9435) );
  INV_X1 U5286 ( .A(n6338), .ZN(n5109) );
  OAI222_X1 U5287 ( .A1(n9719), .A2(n10597), .B1(P2_U3151), .B2(n9718), .C1(
        n9717), .C2(n8618), .ZN(P2_U3266) );
  NAND2_X1 U5288 ( .A1(n6292), .A2(n9718), .ZN(n6478) );
  OR2_X1 U5289 ( .A1(n10540), .A2(n9787), .ZN(n10003) );
  OR2_X1 U5290 ( .A1(n5835), .A2(n5642), .ZN(n5647) );
  OR2_X1 U5291 ( .A1(n5834), .A2(n5645), .ZN(n5642) );
  INV_X2 U5292 ( .A(n6377), .ZN(n6416) );
  INV_X1 U5293 ( .A(n8108), .ZN(n6234) );
  INV_X1 U5294 ( .A(n6859), .ZN(n6669) );
  NAND2_X1 U5295 ( .A1(n5282), .A2(n5280), .ZN(n5279) );
  NAND2_X1 U5296 ( .A1(n5284), .A2(n5283), .ZN(n5282) );
  NOR2_X1 U5297 ( .A1(n9974), .A2(n5281), .ZN(n5280) );
  INV_X1 U5298 ( .A(n9968), .ZN(n5283) );
  OR2_X1 U5299 ( .A1(n8941), .A2(n9764), .ZN(n8946) );
  NAND2_X1 U5300 ( .A1(n5158), .A2(n5297), .ZN(n5295) );
  INV_X1 U5301 ( .A(n5838), .ZN(n5645) );
  OR2_X1 U5302 ( .A1(n9596), .A2(n8675), .ZN(n8843) );
  OR2_X1 U5303 ( .A1(n8691), .A2(n8690), .ZN(n8883) );
  NAND2_X1 U5304 ( .A1(n5310), .A2(n5309), .ZN(n7344) );
  OR2_X1 U5305 ( .A1(n10837), .A2(n6337), .ZN(n5309) );
  NAND2_X1 U5306 ( .A1(n10828), .A2(n10829), .ZN(n5310) );
  NOR2_X1 U5307 ( .A1(n9255), .A2(n5176), .ZN(n9256) );
  OR2_X1 U5308 ( .A1(n9601), .A2(n9174), .ZN(n8838) );
  OR2_X1 U5309 ( .A1(n9203), .A2(n10974), .ZN(n8745) );
  INV_X1 U5310 ( .A(n9773), .ZN(n5462) );
  INV_X1 U5311 ( .A(n10446), .ZN(n5518) );
  INV_X1 U5312 ( .A(n10436), .ZN(n5519) );
  AND2_X1 U5313 ( .A1(n5689), .A2(n8359), .ZN(n6215) );
  AND2_X1 U5314 ( .A1(n5420), .A2(n5978), .ZN(n5419) );
  INV_X1 U5315 ( .A(n5998), .ZN(n5420) );
  NAND2_X1 U5316 ( .A1(n5390), .A2(n5388), .ZN(n5677) );
  AOI21_X1 U5317 ( .B1(n5391), .B2(n5125), .A(n5389), .ZN(n5388) );
  NAND2_X1 U5318 ( .A1(n5664), .A2(n5663), .ZN(n5921) );
  INV_X1 U5319 ( .A(n5918), .ZN(n5663) );
  INV_X1 U5320 ( .A(n5919), .ZN(n5664) );
  NAND2_X1 U5321 ( .A1(n5409), .A2(n5649), .ZN(n5408) );
  INV_X1 U5322 ( .A(n5869), .ZN(n5409) );
  INV_X1 U5323 ( .A(n5805), .ZN(n5634) );
  NAND2_X1 U5324 ( .A1(n7712), .A2(n7711), .ZN(n7716) );
  NOR2_X1 U5325 ( .A1(n7954), .A2(n5595), .ZN(n5594) );
  NAND2_X1 U5326 ( .A1(n9149), .A2(n9049), .ZN(n9051) );
  NAND2_X1 U5327 ( .A1(n9048), .A2(n9047), .ZN(n9049) );
  INV_X1 U5328 ( .A(n9046), .ZN(n9048) );
  AND2_X1 U5329 ( .A1(n8688), .A2(n8687), .ZN(n8854) );
  INV_X1 U5330 ( .A(n5108), .ZN(n6671) );
  OR2_X1 U5331 ( .A1(n9256), .A2(n9263), .ZN(n9274) );
  NAND2_X1 U5332 ( .A1(n5160), .A2(n5296), .ZN(n5288) );
  XNOR2_X1 U5333 ( .A(n9601), .B(n9399), .ZN(n9387) );
  INV_X1 U5334 ( .A(n6628), .ZN(n6286) );
  AOI21_X1 U5335 ( .B1(n9536), .B2(n8787), .A(n9519), .ZN(n5354) );
  NAND2_X1 U5336 ( .A1(n9567), .A2(n6700), .ZN(n9552) );
  AND4_X1 U5337 ( .A1(n6440), .A2(n6439), .A3(n6438), .A4(n6437), .ZN(n7962)
         );
  NAND2_X1 U5338 ( .A1(n6557), .A2(n6556), .ZN(n9092) );
  NAND2_X1 U5339 ( .A1(n8122), .A2(n8121), .ZN(n8164) );
  AND2_X1 U5340 ( .A1(n7028), .A2(n7027), .ZN(n7029) );
  AOI21_X1 U5341 ( .B1(n8172), .B2(n5443), .A(n5441), .ZN(n5440) );
  NAND2_X1 U5342 ( .A1(n5442), .A2(n9782), .ZN(n5441) );
  NAND2_X1 U5343 ( .A1(n5445), .A2(n5443), .ZN(n5442) );
  NAND2_X1 U5344 ( .A1(n7242), .A2(n5480), .ZN(n7429) );
  NOR2_X1 U5345 ( .A1(n5481), .A2(n7245), .ZN(n5480) );
  INV_X1 U5346 ( .A(n7241), .ZN(n5481) );
  INV_X1 U5348 ( .A(n5776), .ZN(n9885) );
  NAND2_X1 U5349 ( .A1(n5706), .A2(n5708), .ZN(n5791) );
  NOR2_X1 U5350 ( .A1(n10088), .A2(n5557), .ZN(n5556) );
  INV_X1 U5351 ( .A(n5934), .ZN(n5557) );
  NAND2_X1 U5352 ( .A1(n9884), .A2(n9883), .ZN(n10283) );
  NAND2_X1 U5353 ( .A1(n9897), .A2(n9896), .ZN(n10291) );
  CLKBUF_X2 U5354 ( .A(n5806), .Z(n9893) );
  XNOR2_X1 U5355 ( .A(n6088), .B(n6087), .ZN(n7958) );
  NAND2_X1 U5356 ( .A1(n6070), .A2(n6069), .ZN(n6088) );
  NAND2_X1 U5357 ( .A1(n6604), .A2(n6603), .ZN(n9440) );
  AOI21_X1 U5358 ( .B1(n5582), .B2(n5583), .A(n5581), .ZN(n5580) );
  INV_X1 U5359 ( .A(n5582), .ZN(n5578) );
  INV_X1 U5360 ( .A(n9094), .ZN(n5581) );
  NAND2_X1 U5361 ( .A1(n6540), .A2(n6539), .ZN(n9537) );
  NAND2_X1 U5362 ( .A1(n5279), .A2(n9987), .ZN(n5276) );
  NOR2_X1 U5363 ( .A1(n9986), .A2(n10055), .ZN(n5275) );
  NAND2_X1 U5364 ( .A1(n5279), .A2(n9982), .ZN(n5278) );
  NAND2_X1 U5365 ( .A1(n5264), .A2(n5263), .ZN(n5262) );
  NAND2_X1 U5366 ( .A1(n10031), .A2(n10060), .ZN(n5264) );
  AOI21_X1 U5367 ( .B1(n10032), .B2(n10055), .A(n10428), .ZN(n5263) );
  INV_X1 U5368 ( .A(n10415), .ZN(n5261) );
  NOR2_X1 U5369 ( .A1(n5144), .A2(n5472), .ZN(n5471) );
  NOR2_X1 U5370 ( .A1(n5475), .A2(n5473), .ZN(n5472) );
  INV_X1 U5371 ( .A(n9857), .ZN(n5473) );
  NAND2_X1 U5372 ( .A1(n10046), .A2(n5271), .ZN(n5270) );
  AND2_X1 U5373 ( .A1(n10045), .A2(n5272), .ZN(n5271) );
  INV_X1 U5374 ( .A(n5385), .ZN(n5384) );
  OAI21_X1 U5375 ( .B1(n6135), .B2(n5386), .A(n6160), .ZN(n5385) );
  INV_X1 U5376 ( .A(n6148), .ZN(n5386) );
  AND2_X1 U5377 ( .A1(n9483), .A2(n5136), .ZN(n6566) );
  OR2_X1 U5378 ( .A1(n9002), .A2(n9905), .ZN(n5478) );
  OR2_X1 U5379 ( .A1(n10553), .A2(n10326), .ZN(n10056) );
  NAND2_X1 U5380 ( .A1(n10484), .A2(n10309), .ZN(n5548) );
  OR2_X1 U5381 ( .A1(n10350), .A2(n10325), .ZN(n10049) );
  NOR2_X1 U5382 ( .A1(n10540), .A2(n9789), .ZN(n5325) );
  INV_X1 U5383 ( .A(n5380), .ZN(n5379) );
  OAI21_X1 U5384 ( .B1(n6055), .B2(n5381), .A(n6087), .ZN(n5380) );
  INV_X1 U5385 ( .A(n6069), .ZN(n5381) );
  NAND2_X1 U5386 ( .A1(n5418), .A2(n6027), .ZN(n5417) );
  NAND2_X1 U5387 ( .A1(n5407), .A2(n5886), .ZN(n5404) );
  INV_X1 U5388 ( .A(n5574), .ZN(n5573) );
  OAI21_X1 U5389 ( .B1(n5576), .B2(n5575), .A(n9101), .ZN(n5574) );
  OR2_X1 U5390 ( .A1(n7331), .A2(n7359), .ZN(n5220) );
  NAND2_X1 U5391 ( .A1(n5220), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5217) );
  AND2_X1 U5392 ( .A1(n7331), .A2(n7359), .ZN(n7332) );
  AOI21_X1 U5393 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n9213), .A(n9208), .ZN(
        n9225) );
  INV_X1 U5394 ( .A(n5292), .ZN(n5291) );
  OAI21_X1 U5395 ( .B1(n5295), .B2(n5293), .A(n6636), .ZN(n5292) );
  INV_X1 U5396 ( .A(n6625), .ZN(n5293) );
  OR2_X1 U5397 ( .A1(n9406), .A2(n9415), .ZN(n8693) );
  AND2_X1 U5398 ( .A1(n9041), .A2(n5350), .ZN(n5349) );
  NAND2_X1 U5399 ( .A1(n5351), .A2(n8800), .ZN(n5350) );
  INV_X1 U5400 ( .A(n9501), .ZN(n5351) );
  INV_X1 U5401 ( .A(n8805), .ZN(n5348) );
  NAND3_X1 U5402 ( .A1(n6331), .A2(n5336), .A3(n10933), .ZN(n8721) );
  INV_X1 U5403 ( .A(n8836), .ZN(n8847) );
  NAND2_X1 U5404 ( .A1(n5302), .A2(n5364), .ZN(n6724) );
  INV_X1 U5405 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5303) );
  NOR2_X1 U5406 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n6257) );
  INV_X1 U5407 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8359) );
  NOR2_X1 U5408 ( .A1(n5465), .A2(n5469), .ZN(n5476) );
  INV_X1 U5409 ( .A(n8920), .ZN(n5465) );
  AOI21_X1 U5410 ( .B1(n8920), .B2(n5468), .A(n5466), .ZN(n8953) );
  INV_X1 U5411 ( .A(n10598), .ZN(n5708) );
  OR2_X1 U5412 ( .A1(n10299), .A2(n10310), .ZN(n10061) );
  NAND2_X1 U5413 ( .A1(n5333), .A2(n10562), .ZN(n5332) );
  NOR2_X1 U5414 ( .A1(n10553), .A2(n10556), .ZN(n5333) );
  OR2_X1 U5415 ( .A1(n10507), .A2(n10425), .ZN(n9899) );
  OR2_X1 U5416 ( .A1(n10432), .A2(n10449), .ZN(n10034) );
  OR2_X1 U5417 ( .A1(n10517), .A2(n10426), .ZN(n10029) );
  OR2_X1 U5418 ( .A1(n9864), .A2(n9799), .ZN(n10024) );
  NOR2_X1 U5419 ( .A1(n7675), .A2(n8029), .ZN(n7676) );
  NOR2_X1 U5420 ( .A1(n5513), .A2(n5509), .ZN(n5508) );
  INV_X1 U5421 ( .A(n5884), .ZN(n5513) );
  NAND2_X1 U5422 ( .A1(n5884), .A2(n5512), .ZN(n5511) );
  INV_X1 U5423 ( .A(n5868), .ZN(n5512) );
  NOR2_X1 U5424 ( .A1(n5814), .A2(n5813), .ZN(n5827) );
  NAND2_X1 U5425 ( .A1(n10056), .A2(n10057), .ZN(n10314) );
  AND2_X1 U5426 ( .A1(n5548), .A2(n6202), .ZN(n5547) );
  NAND2_X1 U5427 ( .A1(n5545), .A2(n5548), .ZN(n5544) );
  NAND2_X1 U5428 ( .A1(n6203), .A2(n5546), .ZN(n5545) );
  INV_X1 U5429 ( .A(n6129), .ZN(n5546) );
  AND2_X1 U5430 ( .A1(n10350), .A2(n10368), .ZN(n6129) );
  NAND2_X1 U5431 ( .A1(n6117), .A2(n6116), .ZN(n6131) );
  NAND2_X1 U5432 ( .A1(n6095), .A2(n6094), .ZN(n6112) );
  OR2_X1 U5433 ( .A1(n6035), .A2(n6034), .ZN(n6049) );
  NAND2_X1 U5434 ( .A1(n5485), .A2(n5560), .ZN(n5484) );
  AND2_X1 U5435 ( .A1(n5698), .A2(n5486), .ZN(n5485) );
  INV_X1 U5436 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5486) );
  AND2_X1 U5437 ( .A1(n5676), .A2(n5675), .ZN(n5962) );
  INV_X1 U5438 ( .A(n5667), .ZN(n5393) );
  INV_X1 U5439 ( .A(n5392), .ZN(n5391) );
  OAI21_X1 U5440 ( .B1(n5395), .B2(n5125), .A(n5672), .ZN(n5392) );
  XNOR2_X1 U5441 ( .A(n5657), .B(SI_13_), .ZN(n5903) );
  NAND2_X1 U5442 ( .A1(n5400), .A2(n5397), .ZN(n5904) );
  INV_X1 U5443 ( .A(n5398), .ZN(n5397) );
  NAND2_X1 U5444 ( .A1(n5647), .A2(n5401), .ZN(n5400) );
  OAI21_X1 U5445 ( .B1(n5404), .B2(n5399), .A(n5157), .ZN(n5398) );
  OR2_X1 U5446 ( .A1(n5645), .A2(n5644), .ZN(n5646) );
  NAND2_X1 U5447 ( .A1(n5638), .A2(n8224), .ZN(n5836) );
  XNOR2_X1 U5448 ( .A(n5635), .B(SI_7_), .ZN(n5805) );
  INV_X1 U5449 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5370) );
  AND2_X1 U5450 ( .A1(n7723), .A2(n7713), .ZN(n5191) );
  XNOR2_X1 U5451 ( .A(n9092), .B(n9196), .ZN(n9041) );
  OR2_X1 U5452 ( .A1(n6541), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6543) );
  OR2_X1 U5453 ( .A1(n7500), .A2(n7499), .ZN(n7712) );
  NOR2_X1 U5454 ( .A1(n5571), .A2(n5198), .ZN(n5197) );
  INV_X1 U5455 ( .A(n9042), .ZN(n5198) );
  INV_X1 U5456 ( .A(n5572), .ZN(n5569) );
  NOR2_X1 U5457 ( .A1(n5575), .A2(n5129), .ZN(n5572) );
  XNOR2_X1 U5458 ( .A(n9622), .B(n9050), .ZN(n9046) );
  INV_X1 U5459 ( .A(n7716), .ZN(n7723) );
  NAND2_X1 U5460 ( .A1(n5587), .A2(n5586), .ZN(n5585) );
  INV_X1 U5461 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8495) );
  INV_X1 U5462 ( .A(n8853), .ZN(n5375) );
  AOI211_X1 U5463 ( .C1(n8677), .C2(n8843), .A(n8848), .B(n8676), .ZN(n8689)
         );
  INV_X1 U5464 ( .A(n8882), .ZN(n8889) );
  NOR2_X1 U5465 ( .A1(n8886), .A2(n9658), .ZN(n8887) );
  OR2_X1 U5466 ( .A1(n6478), .A2(n6933), .ZN(n6309) );
  OAI21_X1 U5467 ( .B1(n6868), .B2(n6844), .A(n6874), .ZN(n6846) );
  NOR2_X1 U5468 ( .A1(n7366), .A2(n7367), .ZN(n7563) );
  NAND2_X1 U5469 ( .A1(n10845), .A2(n7345), .ZN(n7347) );
  NAND2_X1 U5470 ( .A1(n7347), .A2(n7346), .ZN(n7558) );
  NAND2_X1 U5471 ( .A1(n7780), .A2(n5603), .ZN(n7781) );
  NAND2_X1 U5472 ( .A1(n5209), .A2(n7783), .ZN(n7900) );
  NAND2_X1 U5473 ( .A1(n7803), .A2(n7804), .ZN(n7894) );
  XNOR2_X1 U5474 ( .A(n8060), .B(n7895), .ZN(n7896) );
  NAND2_X1 U5475 ( .A1(n8076), .A2(n8077), .ZN(n8078) );
  NAND2_X1 U5476 ( .A1(n8078), .A2(n8079), .ZN(n9215) );
  NAND2_X1 U5477 ( .A1(n7894), .A2(n5305), .ZN(n8060) );
  OR2_X1 U5478 ( .A1(n7898), .A2(n7792), .ZN(n5305) );
  NAND2_X1 U5479 ( .A1(n9234), .A2(n9235), .ZN(n9266) );
  XNOR2_X1 U5480 ( .A(n9225), .B(n9226), .ZN(n9209) );
  OR2_X1 U5481 ( .A1(n9209), .A2(n6477), .ZN(n5429) );
  NAND2_X1 U5482 ( .A1(n9274), .A2(n9257), .ZN(n9258) );
  AOI21_X1 U5483 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n9301), .A(n9298), .ZN(
        n9320) );
  INV_X1 U5484 ( .A(n9193), .ZN(n8675) );
  XNOR2_X1 U5485 ( .A(n9072), .B(n9380), .ZN(n9067) );
  NAND2_X1 U5486 ( .A1(n9380), .A2(n10926), .ZN(n9383) );
  INV_X1 U5487 ( .A(n5605), .ZN(n5341) );
  NOR2_X1 U5488 ( .A1(n5605), .A2(n5343), .ZN(n5342) );
  NOR2_X1 U5489 ( .A1(n5148), .A2(n5356), .ZN(n5355) );
  NOR2_X1 U5490 ( .A1(n5357), .A2(n8821), .ZN(n5356) );
  NOR2_X1 U5491 ( .A1(n8826), .A2(n5359), .ZN(n5358) );
  INV_X1 U5492 ( .A(n8822), .ZN(n5359) );
  OR2_X1 U5493 ( .A1(n9622), .A2(n9460), .ZN(n8822) );
  NAND2_X1 U5494 ( .A1(n9450), .A2(n8821), .ZN(n5360) );
  OR2_X1 U5495 ( .A1(n9510), .A2(n9487), .ZN(n8800) );
  NAND2_X1 U5496 ( .A1(n9497), .A2(n9501), .ZN(n9496) );
  OR2_X1 U5497 ( .A1(n9537), .A2(n9037), .ZN(n8787) );
  OAI21_X1 U5498 ( .B1(n9552), .B2(n9551), .A(n8777), .ZN(n9535) );
  OR2_X1 U5499 ( .A1(n9535), .A2(n9536), .ZN(n9533) );
  OR2_X1 U5500 ( .A1(n6492), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6505) );
  AND2_X1 U5501 ( .A1(n6699), .A2(n8769), .ZN(n5361) );
  AND2_X1 U5502 ( .A1(n6698), .A2(n8784), .ZN(n9570) );
  INV_X1 U5503 ( .A(n6462), .ZN(n6278) );
  INV_X1 U5504 ( .A(n6422), .ZN(n6277) );
  OR3_X1 U5505 ( .A1(n6928), .A2(n6711), .A3(n6712), .ZN(n9021) );
  INV_X1 U5506 ( .A(n6360), .ZN(n6555) );
  INV_X1 U5507 ( .A(n6313), .ZN(n6554) );
  INV_X1 U5508 ( .A(n9200), .ZN(n7738) );
  NAND2_X1 U5509 ( .A1(n7651), .A2(n6688), .ZN(n7733) );
  INV_X1 U5510 ( .A(n10926), .ZN(n9564) );
  INV_X1 U5511 ( .A(n10928), .ZN(n9559) );
  NAND2_X1 U5512 ( .A1(n6275), .A2(n8259), .ZN(n6368) );
  INV_X1 U5513 ( .A(n6350), .ZN(n6275) );
  NAND2_X1 U5514 ( .A1(n6912), .A2(n6680), .ZN(n7145) );
  OR2_X1 U5515 ( .A1(n6728), .A2(P2_D_REG_0__SCAN_IN), .ZN(n6727) );
  NAND2_X1 U5516 ( .A1(n8668), .A2(n8667), .ZN(n8885) );
  NOR2_X1 U5517 ( .A1(n6377), .A2(n8654), .ZN(n5373) );
  NOR2_X1 U5518 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n5363) );
  NAND2_X1 U5519 ( .A1(n6664), .A2(n5563), .ZN(n6714) );
  AND2_X1 U5520 ( .A1(n6269), .A2(n6260), .ZN(n6320) );
  INV_X1 U5521 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5181) );
  INV_X1 U5522 ( .A(n7766), .ZN(n7764) );
  NAND2_X1 U5523 ( .A1(n5451), .A2(n5599), .ZN(n5450) );
  INV_X1 U5524 ( .A(n7974), .ZN(n5451) );
  NOR2_X1 U5525 ( .A1(n8170), .A2(n8901), .ZN(n5445) );
  OR2_X1 U5526 ( .A1(n8171), .A2(n5444), .ZN(n5443) );
  INV_X1 U5527 ( .A(n8901), .ZN(n5444) );
  AOI21_X1 U5528 ( .B1(n9734), .B2(n8965), .A(n8962), .ZN(n8970) );
  NAND2_X1 U5529 ( .A1(n7033), .A2(n5601), .ZN(n7054) );
  NAND2_X1 U5530 ( .A1(n7030), .A2(n9905), .ZN(n5479) );
  NAND2_X1 U5531 ( .A1(n5111), .A2(n5449), .ZN(n5448) );
  INV_X1 U5532 ( .A(n5599), .ZN(n5449) );
  NAND2_X1 U5533 ( .A1(n5450), .A2(n5111), .ZN(n8032) );
  NAND2_X1 U5534 ( .A1(n5476), .A2(n5475), .ZN(n9856) );
  NAND2_X1 U5535 ( .A1(n7233), .A2(n5128), .ZN(n7242) );
  INV_X1 U5536 ( .A(n5457), .ZN(n9869) );
  AOI21_X1 U5537 ( .B1(n9810), .B2(n9807), .A(n5458), .ZN(n5457) );
  NAND2_X1 U5538 ( .A1(n9773), .A2(n5459), .ZN(n5458) );
  NAND2_X1 U5539 ( .A1(n9808), .A2(n9807), .ZN(n5459) );
  NAND2_X1 U5540 ( .A1(n9773), .A2(n5461), .ZN(n5460) );
  AND2_X1 U5541 ( .A1(n9872), .A2(n9868), .ZN(n5463) );
  NOR2_X1 U5542 ( .A1(n5113), .A2(n5456), .ZN(n5455) );
  INV_X1 U5543 ( .A(n8970), .ZN(n5456) );
  NOR2_X1 U5544 ( .A1(n5113), .A2(n5464), .ZN(n5453) );
  NAND2_X1 U5545 ( .A1(n8166), .A2(n8165), .ZN(n8172) );
  NAND2_X1 U5546 ( .A1(n10598), .A2(n5706), .ZN(n6079) );
  NAND2_X1 U5547 ( .A1(n5707), .A2(n10598), .ZN(n9889) );
  OAI22_X1 U5548 ( .A1(n7324), .A2(n6079), .B1(n9889), .B2(n5713), .ZN(n5250)
         );
  NAND2_X1 U5549 ( .A1(n10061), .A2(n10132), .ZN(n10102) );
  AND2_X1 U5550 ( .A1(n5541), .A2(n10314), .ZN(n5540) );
  NAND2_X1 U5551 ( .A1(n5544), .A2(n5542), .ZN(n5541) );
  INV_X1 U5552 ( .A(n5547), .ZN(n5542) );
  INV_X1 U5553 ( .A(n5544), .ZN(n5543) );
  NAND2_X1 U5554 ( .A1(n10360), .A2(n5331), .ZN(n10290) );
  NOR2_X1 U5555 ( .A1(n10299), .A2(n5332), .ZN(n5331) );
  AND2_X1 U5556 ( .A1(n10381), .A2(n10365), .ZN(n10360) );
  NAND2_X1 U5557 ( .A1(n10397), .A2(n10398), .ZN(n5490) );
  NAND2_X1 U5558 ( .A1(n5489), .A2(n5490), .ZN(n10373) );
  AND2_X1 U5559 ( .A1(n10379), .A2(n10037), .ZN(n5489) );
  AND2_X1 U5560 ( .A1(n10048), .A2(n10040), .ZN(n10379) );
  NOR2_X1 U5561 ( .A1(n10382), .A2(n10391), .ZN(n10381) );
  NAND2_X1 U5562 ( .A1(n5230), .A2(n5228), .ZN(n10397) );
  AOI21_X1 U5563 ( .B1(n5232), .B2(n5235), .A(n5229), .ZN(n5228) );
  NAND2_X1 U5564 ( .A1(n10445), .A2(n5232), .ZN(n5230) );
  INV_X1 U5565 ( .A(n9932), .ZN(n5235) );
  INV_X1 U5566 ( .A(n5525), .ZN(n5524) );
  OAI22_X1 U5567 ( .A1(n10415), .A2(n5531), .B1(n10399), .B2(n10507), .ZN(
        n5525) );
  AND2_X1 U5568 ( .A1(n10036), .A2(n10037), .ZN(n10398) );
  NOR2_X1 U5569 ( .A1(n10415), .A2(n5528), .ZN(n5527) );
  AND2_X1 U5570 ( .A1(n9899), .A2(n10124), .ZN(n10415) );
  INV_X1 U5571 ( .A(n5516), .ZN(n5514) );
  AOI22_X1 U5572 ( .A1(n8152), .A2(n5997), .B1(n8155), .B2(n10448), .ZN(n10436) );
  OAI21_X1 U5573 ( .B1(n7989), .B2(n10010), .A(n10006), .ZN(n8139) );
  NAND2_X1 U5574 ( .A1(n7994), .A2(n5602), .ZN(n8086) );
  OR2_X1 U5575 ( .A1(n8102), .A2(n9798), .ZN(n5602) );
  AND4_X1 U5576 ( .A1(n5947), .A2(n5946), .A3(n5945), .A4(n5944), .ZN(n9787)
         );
  INV_X1 U5577 ( .A(n5554), .ZN(n5553) );
  OAI22_X1 U5578 ( .A1(n10088), .A2(n5555), .B1(n10540), .B2(n10160), .ZN(
        n5554) );
  NAND2_X1 U5579 ( .A1(n5933), .A2(n5934), .ZN(n5555) );
  NAND2_X1 U5580 ( .A1(n5551), .A2(n5549), .ZN(n7994) );
  AND2_X1 U5581 ( .A1(n5553), .A2(n5550), .ZN(n5549) );
  AND2_X1 U5582 ( .A1(n10003), .A2(n10005), .ZN(n10088) );
  NOR2_X1 U5583 ( .A1(n11034), .A2(n7973), .ZN(n6212) );
  OR2_X1 U5584 ( .A1(n7636), .A2(n5900), .ZN(n5902) );
  AND4_X1 U5585 ( .A1(n5833), .A2(n5832), .A3(n5831), .A4(n5830), .ZN(n7627)
         );
  NAND2_X1 U5586 ( .A1(n7300), .A2(n9961), .ZN(n7302) );
  NAND2_X1 U5587 ( .A1(n5504), .A2(n5773), .ZN(n7471) );
  NOR2_X1 U5588 ( .A1(n5774), .A2(n5506), .ZN(n5505) );
  XNOR2_X1 U5589 ( .A(n10171), .B(n5247), .ZN(n10069) );
  AND3_X1 U5590 ( .A1(n7032), .A2(P1_STATE_REG_SCAN_IN), .A3(n7743), .ZN(
        n10584) );
  AND2_X1 U5591 ( .A1(n5684), .A2(n5561), .ZN(n5560) );
  INV_X1 U5592 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5561) );
  AND2_X1 U5593 ( .A1(n5691), .A2(n5698), .ZN(n5692) );
  XNOR2_X1 U5594 ( .A(n6228), .B(P1_IR_REG_22__SCAN_IN), .ZN(n10111) );
  NAND2_X1 U5595 ( .A1(n5414), .A2(n5418), .ZN(n6030) );
  NAND2_X1 U5596 ( .A1(n5112), .A2(n5167), .ZN(n5414) );
  NAND2_X1 U5597 ( .A1(n5112), .A2(n5978), .ZN(n5999) );
  NAND2_X1 U5598 ( .A1(n5937), .A2(n5698), .ZN(n5950) );
  NAND2_X1 U5599 ( .A1(n5394), .A2(n5667), .ZN(n5949) );
  NAND2_X1 U5600 ( .A1(n5921), .A2(n5395), .ZN(n5394) );
  NAND2_X1 U5601 ( .A1(n5921), .A2(n5665), .ZN(n5936) );
  INV_X1 U5602 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5684) );
  NOR2_X1 U5603 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5682) );
  NAND2_X1 U5604 ( .A1(n5405), .A2(n5407), .ZN(n5887) );
  OR2_X1 U5605 ( .A1(n5647), .A2(n5408), .ZN(n5405) );
  NOR2_X1 U5606 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5766) );
  INV_X1 U5607 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5679) );
  NAND2_X1 U5608 ( .A1(n9064), .A2(n5194), .ZN(n9077) );
  NOR2_X1 U5609 ( .A1(n9076), .A2(n5195), .ZN(n5194) );
  INV_X1 U5610 ( .A(n9063), .ZN(n5195) );
  NAND2_X1 U5611 ( .A1(n6638), .A2(n6637), .ZN(n9601) );
  NAND2_X1 U5612 ( .A1(n8134), .A2(n6416), .ZN(n6638) );
  NAND2_X1 U5613 ( .A1(n5200), .A2(n8001), .ZN(n9034) );
  INV_X1 U5614 ( .A(n5592), .ZN(n5590) );
  OR2_X1 U5615 ( .A1(n9117), .A2(n9037), .ZN(n5201) );
  NAND2_X1 U5616 ( .A1(n9117), .A2(n9037), .ZN(n5203) );
  INV_X1 U5617 ( .A(n9398), .ZN(n9425) );
  NAND2_X1 U5618 ( .A1(n9053), .A2(n9052), .ZN(n9054) );
  NAND2_X1 U5619 ( .A1(n6616), .A2(n6615), .ZN(n9421) );
  AND4_X1 U5620 ( .A1(n6535), .A2(n6534), .A3(n6533), .A4(n6532), .ZN(n9503)
         );
  NAND2_X1 U5621 ( .A1(n6299), .A2(n6298), .ZN(n9381) );
  XNOR2_X1 U5622 ( .A(n6358), .B(P2_IR_REG_4__SCAN_IN), .ZN(n10837) );
  NAND2_X1 U5623 ( .A1(n10862), .A2(n10861), .ZN(n10860) );
  OR2_X1 U5624 ( .A1(n10853), .A2(n7513), .ZN(n5424) );
  NAND2_X1 U5625 ( .A1(n5421), .A2(n5212), .ZN(n5211) );
  NAND2_X1 U5626 ( .A1(n7335), .A2(n5425), .ZN(n5421) );
  OR2_X1 U5627 ( .A1(n10853), .A2(n5422), .ZN(n5212) );
  NAND2_X1 U5628 ( .A1(n5425), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5422) );
  NAND2_X1 U5629 ( .A1(n8063), .A2(n8064), .ZN(n9205) );
  INV_X1 U5630 ( .A(n9274), .ZN(n9276) );
  NAND2_X1 U5631 ( .A1(n6514), .A2(n6513), .ZN(n6553) );
  NAND2_X1 U5632 ( .A1(n8674), .A2(n8673), .ZN(n9596) );
  XNOR2_X1 U5633 ( .A(n9018), .B(n9017), .ZN(n9593) );
  NAND2_X1 U5634 ( .A1(n5159), .A2(n6313), .ZN(n5298) );
  NAND2_X1 U5635 ( .A1(n5925), .A2(n5924), .ZN(n8128) );
  OAI21_X1 U5636 ( .B1(n10146), .B2(n10145), .A(n10153), .ZN(n5252) );
  NAND2_X1 U5637 ( .A1(n5255), .A2(n5254), .ZN(n5253) );
  AND2_X1 U5638 ( .A1(n10144), .A2(n10145), .ZN(n5254) );
  NAND2_X1 U5639 ( .A1(n10122), .A2(n5256), .ZN(n5255) );
  INV_X1 U5640 ( .A(n10111), .ZN(n10151) );
  NAND2_X1 U5641 ( .A1(n9204), .A2(n10938), .ZN(n8716) );
  NAND2_X1 U5642 ( .A1(n9975), .A2(n10075), .ZN(n5281) );
  NAND2_X1 U5643 ( .A1(n9970), .A2(n9969), .ZN(n5284) );
  NAND2_X1 U5644 ( .A1(n5277), .A2(n5274), .ZN(n9996) );
  NAND2_X1 U5645 ( .A1(n5278), .A2(n5141), .ZN(n5277) );
  NAND2_X1 U5646 ( .A1(n5276), .A2(n5275), .ZN(n5274) );
  OAI21_X1 U5647 ( .B1(n5260), .B2(n10039), .A(n5259), .ZN(n10047) );
  AND2_X1 U5648 ( .A1(n10379), .A2(n10038), .ZN(n5259) );
  AOI21_X1 U5649 ( .B1(n5262), .B2(n10035), .A(n5261), .ZN(n5260) );
  AND2_X1 U5650 ( .A1(n10049), .A2(n10060), .ZN(n5272) );
  INV_X1 U5651 ( .A(n6266), .ZN(n5365) );
  INV_X1 U5652 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6523) );
  INV_X1 U5653 ( .A(n9794), .ZN(n5469) );
  NOR2_X1 U5654 ( .A1(n5470), .A2(n5469), .ZN(n5468) );
  INV_X1 U5655 ( .A(n5471), .ZN(n5470) );
  NAND2_X1 U5656 ( .A1(n5145), .A2(n5467), .ZN(n5466) );
  NAND2_X1 U5657 ( .A1(n5471), .A2(n5474), .ZN(n5467) );
  NOR2_X1 U5658 ( .A1(n8942), .A2(n9857), .ZN(n5474) );
  NAND2_X1 U5659 ( .A1(n5269), .A2(n5147), .ZN(n10059) );
  NAND2_X1 U5660 ( .A1(n7603), .A2(n10969), .ZN(n5329) );
  NAND2_X1 U5661 ( .A1(n5383), .A2(n5382), .ZN(n8645) );
  AOI21_X1 U5662 ( .B1(n5384), .B2(n5386), .A(n5178), .ZN(n5382) );
  NAND2_X1 U5663 ( .A1(n6136), .A2(n5384), .ZN(n5383) );
  OAI22_X1 U5664 ( .A1(n5167), .A2(n5417), .B1(n6029), .B2(n8197), .ZN(n5416)
         );
  INV_X1 U5665 ( .A(n5962), .ZN(n5389) );
  NAND2_X1 U5666 ( .A1(n5669), .A2(n8206), .ZN(n5672) );
  INV_X1 U5667 ( .A(n5408), .ZN(n5399) );
  INV_X1 U5668 ( .A(n5404), .ZN(n5401) );
  INV_X1 U5669 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5368) );
  INV_X1 U5670 ( .A(n9142), .ZN(n5576) );
  INV_X1 U5671 ( .A(n9044), .ZN(n5575) );
  NAND2_X1 U5672 ( .A1(n9287), .A2(n9288), .ZN(n9289) );
  AND2_X1 U5673 ( .A1(n9324), .A2(n5187), .ZN(n9329) );
  NAND2_X1 U5674 ( .A1(n9326), .A2(n9325), .ZN(n5187) );
  NAND2_X1 U5675 ( .A1(n9312), .A2(n5307), .ZN(n9336) );
  NAND2_X1 U5676 ( .A1(n9301), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5307) );
  NAND2_X1 U5677 ( .A1(n9415), .A2(n9667), .ZN(n5296) );
  AND2_X1 U5678 ( .A1(n5296), .A2(n5294), .ZN(n5289) );
  INV_X1 U5679 ( .A(n5295), .ZN(n5294) );
  INV_X1 U5680 ( .A(n5358), .ZN(n5357) );
  AND2_X1 U5681 ( .A1(n6283), .A2(n8484), .ZN(n6586) );
  INV_X1 U5682 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8480) );
  INV_X1 U5683 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8447) );
  INV_X1 U5684 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8259) );
  OR2_X1 U5685 ( .A1(n5108), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6328) );
  OR2_X1 U5686 ( .A1(n5110), .A2(n6326), .ZN(n6330) );
  INV_X1 U5687 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5565) );
  AND2_X1 U5688 ( .A1(n5563), .A2(n5365), .ZN(n5304) );
  INV_X1 U5689 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6525) );
  OAI211_X1 U5690 ( .C1(n9905), .C2(n9001), .A(n7030), .B(n5478), .ZN(n7055)
         );
  INV_X1 U5691 ( .A(n9002), .ZN(n8974) );
  INV_X1 U5692 ( .A(n5226), .ZN(n5225) );
  OAI21_X1 U5693 ( .B1(n5487), .B2(n5227), .A(n10346), .ZN(n5226) );
  INV_X1 U5694 ( .A(n9898), .ZN(n5227) );
  NOR2_X1 U5695 ( .A1(n10358), .A2(n5488), .ZN(n5487) );
  INV_X1 U5696 ( .A(n10048), .ZN(n5488) );
  NAND2_X1 U5697 ( .A1(n5524), .A2(n5137), .ZN(n5523) );
  NAND2_X1 U5698 ( .A1(n10501), .A2(n10376), .ZN(n5530) );
  NOR2_X1 U5699 ( .A1(n5523), .A2(n5516), .ZN(n5515) );
  AOI21_X1 U5700 ( .B1(n5234), .B2(n9932), .A(n5233), .ZN(n5232) );
  INV_X1 U5701 ( .A(n9899), .ZN(n5233) );
  INV_X1 U5702 ( .A(n9930), .ZN(n5234) );
  NAND2_X1 U5703 ( .A1(n5318), .A2(n10409), .ZN(n5317) );
  NOR2_X1 U5704 ( .A1(n10517), .A2(n10156), .ZN(n5516) );
  AND2_X1 U5705 ( .A1(n8623), .A2(n5323), .ZN(n8147) );
  AND2_X1 U5706 ( .A1(n5119), .A2(n10580), .ZN(n5323) );
  NAND2_X1 U5707 ( .A1(n7474), .A2(n6189), .ZN(n7303) );
  INV_X1 U5708 ( .A(n7478), .ZN(n5328) );
  NOR2_X1 U5709 ( .A1(n5329), .A2(n7433), .ZN(n5327) );
  INV_X1 U5710 ( .A(n9950), .ZN(n5494) );
  NAND2_X1 U5711 ( .A1(n9820), .A2(n5245), .ZN(n9950) );
  OR2_X1 U5712 ( .A1(n10169), .A2(n10899), .ZN(n9951) );
  NAND2_X1 U5713 ( .A1(n7318), .A2(n6186), .ZN(n9949) );
  NAND2_X1 U5714 ( .A1(n10348), .A2(n10484), .ZN(n10334) );
  NAND2_X1 U5715 ( .A1(n8623), .A2(n5325), .ZN(n8088) );
  NAND2_X1 U5716 ( .A1(n8623), .A2(n8630), .ZN(n8624) );
  NOR2_X1 U5717 ( .A1(n7478), .A2(n5329), .ZN(n7311) );
  XNOR2_X1 U5718 ( .A(n8645), .B(n8644), .ZN(n8642) );
  NAND2_X1 U5719 ( .A1(n6112), .A2(n6111), .ZN(n6117) );
  NAND2_X1 U5720 ( .A1(n5378), .A2(n5376), .ZN(n6095) );
  AOI21_X1 U5721 ( .B1(n5379), .B2(n5381), .A(n5377), .ZN(n5376) );
  INV_X1 U5722 ( .A(n6089), .ZN(n5377) );
  OAI21_X1 U5723 ( .B1(n5980), .B2(n5412), .A(n5415), .ZN(n6035) );
  NAND2_X1 U5724 ( .A1(n5413), .A2(n5976), .ZN(n5412) );
  INV_X1 U5725 ( .A(n5416), .ZN(n5415) );
  INV_X1 U5726 ( .A(n5417), .ZN(n5413) );
  NAND2_X1 U5727 ( .A1(n5174), .A2(n6015), .ZN(n5418) );
  NAND2_X1 U5728 ( .A1(n5131), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5963) );
  INV_X1 U5729 ( .A(n5484), .ZN(n5482) );
  NOR2_X1 U5730 ( .A1(n5668), .A2(n5396), .ZN(n5395) );
  INV_X1 U5731 ( .A(n5665), .ZN(n5396) );
  NAND2_X1 U5732 ( .A1(n5660), .A2(n8422), .ZN(n5665) );
  NAND2_X1 U5733 ( .A1(n5659), .A2(n5658), .ZN(n5919) );
  NAND2_X1 U5734 ( .A1(n5904), .A2(n5656), .ZN(n5659) );
  OR2_X1 U5735 ( .A1(n5842), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5889) );
  NAND2_X1 U5736 ( .A1(n5403), .A2(n5402), .ZN(n5407) );
  NAND2_X1 U5737 ( .A1(n5408), .A2(n5654), .ZN(n5403) );
  NAND2_X1 U5738 ( .A1(n5641), .A2(SI_9_), .ZN(n5838) );
  NAND2_X1 U5739 ( .A1(n5836), .A2(n5640), .ZN(n5834) );
  OAI21_X1 U5740 ( .B1(n8662), .B2(n5627), .A(n5626), .ZN(n5628) );
  OAI21_X1 U5741 ( .B1(n6772), .B2(n5411), .A(n5410), .ZN(n5623) );
  NAND2_X1 U5742 ( .A1(n6772), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5410) );
  OAI21_X1 U5743 ( .B1(n5618), .B2(n5609), .A(n5608), .ZN(n5612) );
  AOI21_X1 U5744 ( .B1(n5584), .B2(n9039), .A(n5155), .ZN(n5582) );
  INV_X1 U5745 ( .A(n5584), .ZN(n5583) );
  XNOR2_X1 U5746 ( .A(n7152), .B(n7148), .ZN(n6952) );
  NOR2_X1 U5747 ( .A1(n7926), .A2(n9198), .ZN(n5595) );
  NAND2_X1 U5748 ( .A1(n5598), .A2(n5597), .ZN(n5596) );
  NAND2_X1 U5749 ( .A1(n5577), .A2(n5576), .ZN(n9139) );
  INV_X1 U5750 ( .A(n9141), .ZN(n5577) );
  NOR2_X1 U5751 ( .A1(n7927), .A2(n5153), .ZN(n5592) );
  OR2_X1 U5752 ( .A1(n6595), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6605) );
  NOR2_X1 U5753 ( .A1(n9158), .A2(n5589), .ZN(n5584) );
  INV_X1 U5754 ( .A(n6543), .ZN(n6281) );
  OR2_X1 U5755 ( .A1(n6531), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6558) );
  INV_X1 U5756 ( .A(n7176), .ZN(n5193) );
  NAND2_X1 U5757 ( .A1(n6280), .A2(n8500), .ZN(n6541) );
  INV_X1 U5758 ( .A(n6505), .ZN(n6280) );
  OR2_X1 U5759 ( .A1(n5219), .A2(n7332), .ZN(n10810) );
  INV_X1 U5760 ( .A(n5220), .ZN(n5219) );
  NOR2_X1 U5761 ( .A1(n5217), .A2(n7332), .ZN(n10809) );
  NAND2_X1 U5762 ( .A1(n10811), .A2(n7343), .ZN(n10828) );
  INV_X1 U5763 ( .A(n7332), .ZN(n5218) );
  XNOR2_X1 U5764 ( .A(n7344), .B(n10847), .ZN(n10846) );
  NAND2_X1 U5765 ( .A1(n10860), .A2(n7365), .ZN(n7366) );
  INV_X1 U5766 ( .A(n7337), .ZN(n5425) );
  NAND2_X1 U5767 ( .A1(n7558), .A2(n7559), .ZN(n7689) );
  NOR2_X1 U5768 ( .A1(n5211), .A2(n5210), .ZN(n7683) );
  NOR2_X1 U5769 ( .A1(n7352), .A2(n7349), .ZN(n5210) );
  OR2_X1 U5770 ( .A1(n7788), .A2(n7787), .ZN(n5183) );
  AND2_X1 U5771 ( .A1(n5183), .A2(n7790), .ZN(n7855) );
  OR2_X1 U5772 ( .A1(n7847), .A2(n7782), .ZN(n5209) );
  NAND2_X1 U5773 ( .A1(n7849), .A2(n7802), .ZN(n7803) );
  XNOR2_X1 U5774 ( .A(n8065), .B(n8074), .ZN(n7902) );
  NOR2_X1 U5775 ( .A1(n7855), .A2(n7791), .ZN(n7890) );
  NOR2_X1 U5776 ( .A1(n7902), .A2(n7965), .ZN(n8067) );
  OAI21_X1 U5777 ( .B1(n7902), .B2(n5432), .A(n5431), .ZN(n9208) );
  NAND2_X1 U5778 ( .A1(n5433), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5432) );
  NAND2_X1 U5779 ( .A1(n8066), .A2(n5433), .ZN(n5431) );
  INV_X1 U5780 ( .A(n8070), .ZN(n5433) );
  NAND2_X1 U5781 ( .A1(n9215), .A2(n9216), .ZN(n9217) );
  NAND2_X1 U5782 ( .A1(n9205), .A2(n5308), .ZN(n9241) );
  NAND2_X1 U5783 ( .A1(n9213), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5308) );
  NAND2_X1 U5784 ( .A1(n9266), .A2(n9267), .ZN(n9268) );
  NAND2_X1 U5785 ( .A1(n9268), .A2(n9269), .ZN(n9287) );
  NAND2_X1 U5786 ( .A1(n9281), .A2(n9282), .ZN(n9312) );
  XNOR2_X1 U5787 ( .A(n9336), .B(n9325), .ZN(n9314) );
  NAND2_X1 U5788 ( .A1(n9314), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n9338) );
  NAND2_X1 U5789 ( .A1(n5186), .A2(n9348), .ZN(n9332) );
  INV_X1 U5790 ( .A(n9347), .ZN(n5186) );
  INV_X1 U5791 ( .A(n9323), .ZN(n5439) );
  NOR2_X1 U5792 ( .A1(n9329), .A2(n9328), .ZN(n9347) );
  NAND2_X1 U5793 ( .A1(n8672), .A2(n8671), .ZN(n9018) );
  INV_X1 U5794 ( .A(n6670), .ZN(n9023) );
  INV_X1 U5795 ( .A(n9016), .ZN(n9017) );
  NAND2_X1 U5796 ( .A1(n5340), .A2(n5338), .ZN(n9388) );
  AOI21_X1 U5797 ( .B1(n5342), .B2(n8830), .A(n5339), .ZN(n5338) );
  INV_X1 U5798 ( .A(n8693), .ZN(n5339) );
  NAND2_X1 U5799 ( .A1(n9388), .A2(n9387), .ZN(n9386) );
  NAND2_X1 U5800 ( .A1(n5290), .A2(n5291), .ZN(n9396) );
  NAND2_X1 U5801 ( .A1(n9423), .A2(n5294), .ZN(n5290) );
  OR2_X1 U5802 ( .A1(n6605), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6617) );
  NAND2_X1 U5803 ( .A1(n6285), .A2(n8263), .ZN(n6628) );
  INV_X1 U5804 ( .A(n6617), .ZN(n6285) );
  NOR2_X1 U5805 ( .A1(n5606), .A2(n5130), .ZN(n6571) );
  AOI21_X1 U5806 ( .B1(n5349), .B2(n5352), .A(n5348), .ZN(n5347) );
  INV_X1 U5807 ( .A(n8800), .ZN(n5352) );
  OR2_X1 U5808 ( .A1(n6550), .A2(n6549), .ZN(n6551) );
  NAND2_X1 U5809 ( .A1(n9480), .A2(n9481), .ZN(n9528) );
  INV_X1 U5810 ( .A(n9529), .ZN(n9563) );
  INV_X1 U5811 ( .A(n9570), .ZN(n6699) );
  NAND2_X1 U5812 ( .A1(n6279), .A2(n8488), .ZN(n6492) );
  OR2_X1 U5813 ( .A1(n6448), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6462) );
  AND2_X1 U5814 ( .A1(n5366), .A2(n5124), .ZN(n8015) );
  AND2_X1 U5815 ( .A1(n8758), .A2(n8759), .ZN(n8869) );
  OR2_X1 U5816 ( .A1(n6435), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6448) );
  NAND2_X1 U5817 ( .A1(n6689), .A2(n8740), .ZN(n7816) );
  OR2_X1 U5818 ( .A1(n6405), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6422) );
  AND2_X1 U5819 ( .A1(n6276), .A2(n8495), .ZN(n6396) );
  INV_X1 U5820 ( .A(n6368), .ZN(n6276) );
  NAND2_X1 U5821 ( .A1(n6396), .A2(n8447), .ZN(n6405) );
  INV_X1 U5822 ( .A(n9201), .ZN(n7814) );
  NAND2_X1 U5823 ( .A1(n6687), .A2(n8861), .ZN(n7651) );
  AOI21_X1 U5824 ( .B1(n10930), .B2(n6686), .A(n6685), .ZN(n7509) );
  INV_X1 U5825 ( .A(n10951), .ZN(n5300) );
  NOR2_X1 U5826 ( .A1(n7154), .A2(n10951), .ZN(n5301) );
  NAND2_X1 U5827 ( .A1(n7163), .A2(n6274), .ZN(n6350) );
  INV_X1 U5828 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6274) );
  NAND2_X1 U5829 ( .A1(n8855), .A2(n8721), .ZN(n7388) );
  NOR2_X1 U5830 ( .A1(n6777), .A2(n8662), .ZN(n5299) );
  AND2_X1 U5831 ( .A1(n6960), .A2(n8836), .ZN(n10926) );
  AND2_X1 U5832 ( .A1(n6900), .A2(n6904), .ZN(n6908) );
  INV_X1 U5833 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6662) );
  OAI21_X1 U5834 ( .B1(n6502), .B2(n5204), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5206) );
  NAND2_X1 U5835 ( .A1(n6513), .A2(n5205), .ZN(n5204) );
  NOR2_X1 U5836 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n6259) );
  NOR2_X1 U5837 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n6258) );
  NAND2_X1 U5838 ( .A1(n6176), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6228) );
  OR2_X1 U5839 ( .A1(n5862), .A2(n5861), .ZN(n5878) );
  NOR3_X1 U5840 ( .A1(n5258), .A2(n5139), .A3(n5257), .ZN(n5256) );
  NOR2_X1 U5841 ( .A1(n10115), .A2(n10105), .ZN(n5258) );
  AND4_X1 U5842 ( .A1(n5796), .A2(n5795), .A3(n5794), .A4(n5793), .ZN(n7443)
         );
  OR2_X1 U5843 ( .A1(n6209), .A2(n6997), .ZN(n5780) );
  NAND2_X1 U5844 ( .A1(n10306), .A2(n10057), .ZN(n5503) );
  INV_X1 U5845 ( .A(n10102), .ZN(n5502) );
  INV_X1 U5846 ( .A(n5332), .ZN(n5330) );
  AND4_X1 U5847 ( .A1(n6147), .A2(n6146), .A3(n6145), .A4(n6144), .ZN(n10309)
         );
  INV_X1 U5848 ( .A(n10314), .ZN(n10308) );
  NAND2_X1 U5849 ( .A1(n10307), .A2(n10308), .ZN(n10306) );
  NAND2_X1 U5850 ( .A1(n5224), .A2(n5222), .ZN(n10324) );
  AOI21_X1 U5851 ( .B1(n5225), .B2(n5227), .A(n5223), .ZN(n5222) );
  NAND2_X1 U5852 ( .A1(n10373), .A2(n5225), .ZN(n5224) );
  INV_X1 U5853 ( .A(n10044), .ZN(n5223) );
  INV_X1 U5854 ( .A(n6203), .ZN(n10329) );
  AND4_X1 U5855 ( .A1(n6128), .A2(n6127), .A3(n6126), .A4(n6125), .ZN(n10325)
         );
  NAND2_X1 U5856 ( .A1(n10366), .A2(n9898), .ZN(n10341) );
  INV_X1 U5857 ( .A(n6202), .ZN(n10346) );
  OAI21_X1 U5858 ( .B1(n10373), .B2(n5227), .A(n5225), .ZN(n10340) );
  NAND2_X1 U5859 ( .A1(n10373), .A2(n5487), .ZN(n10366) );
  NAND2_X1 U5860 ( .A1(n5522), .A2(n5520), .ZN(n10380) );
  INV_X1 U5861 ( .A(n5521), .ZN(n5520) );
  NAND2_X1 U5862 ( .A1(n5517), .A2(n5515), .ZN(n5522) );
  OAI21_X1 U5863 ( .B1(n5523), .B2(n5527), .A(n5530), .ZN(n5521) );
  NOR3_X1 U5864 ( .A1(n10439), .A2(n5316), .A3(n10432), .ZN(n6213) );
  OR2_X1 U5865 ( .A1(n5317), .A2(n10501), .ZN(n5316) );
  NAND2_X1 U5866 ( .A1(n5231), .A2(n9932), .ZN(n10414) );
  NAND2_X1 U5867 ( .A1(n10445), .A2(n9930), .ZN(n5231) );
  NOR3_X1 U5868 ( .A1(n10439), .A2(n10432), .A3(n10517), .ZN(n10420) );
  INV_X1 U5869 ( .A(n6007), .ZN(n6008) );
  NOR2_X1 U5870 ( .A1(n10439), .A2(n10517), .ZN(n10437) );
  AND2_X1 U5871 ( .A1(n10029), .A2(n10026), .ZN(n10446) );
  AND2_X1 U5872 ( .A1(n5702), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5992) );
  AND4_X1 U5873 ( .A1(n6012), .A2(n6011), .A3(n6010), .A4(n6009), .ZN(n10426)
         );
  INV_X1 U5874 ( .A(n5243), .ZN(n8159) );
  OAI21_X1 U5875 ( .B1(n8139), .B2(n10091), .A(n6199), .ZN(n5243) );
  NAND2_X1 U5876 ( .A1(n8147), .A2(n8155), .ZN(n10439) );
  AND2_X1 U5877 ( .A1(n10019), .A2(n10027), .ZN(n10093) );
  AND2_X1 U5878 ( .A1(n10535), .A2(n10159), .ZN(n5975) );
  NAND2_X1 U5879 ( .A1(n6198), .A2(n10003), .ZN(n7989) );
  NOR2_X1 U5880 ( .A1(n5954), .A2(n7830), .ZN(n5970) );
  NOR2_X1 U5881 ( .A1(n5927), .A2(n5926), .ZN(n5941) );
  AND2_X1 U5882 ( .A1(n7676), .A2(n8056), .ZN(n8623) );
  NAND2_X1 U5883 ( .A1(n5908), .A2(n5907), .ZN(n8029) );
  NAND2_X1 U5884 ( .A1(n5498), .A2(n5496), .ZN(n7912) );
  NOR2_X1 U5885 ( .A1(n10085), .A2(n5497), .ZN(n5496) );
  INV_X1 U5886 ( .A(n9988), .ZN(n5497) );
  NAND2_X1 U5887 ( .A1(n5498), .A2(n9988), .ZN(n7670) );
  NAND2_X1 U5888 ( .A1(n5892), .A2(n5891), .ZN(n7973) );
  AND2_X1 U5889 ( .A1(n5511), .A2(n5885), .ZN(n5510) );
  NAND2_X1 U5890 ( .A1(n7450), .A2(n10079), .ZN(n7449) );
  NOR2_X1 U5891 ( .A1(n7451), .A2(n7773), .ZN(n11036) );
  NAND2_X1 U5892 ( .A1(n5532), .A2(n5535), .ZN(n7418) );
  AOI21_X1 U5893 ( .B1(n9968), .B2(n5536), .A(n5152), .ZN(n5535) );
  INV_X1 U5894 ( .A(n5820), .ZN(n5536) );
  OR2_X1 U5895 ( .A1(n7548), .A2(n10457), .ZN(n7451) );
  NAND2_X1 U5896 ( .A1(n5327), .A2(n5328), .ZN(n7546) );
  AND4_X1 U5897 ( .A1(n5852), .A2(n5851), .A3(n5850), .A4(n5849), .ZN(n7770)
         );
  AND4_X1 U5898 ( .A1(n5819), .A2(n5818), .A3(n5817), .A4(n5816), .ZN(n7539)
         );
  OAI21_X1 U5899 ( .B1(n7471), .B2(n9957), .A(n5790), .ZN(n7216) );
  NAND2_X1 U5900 ( .A1(n7216), .A2(n9964), .ZN(n7215) );
  NOR2_X1 U5901 ( .A1(n7478), .A2(n7482), .ZN(n7481) );
  OAI211_X1 U5902 ( .C1(n6188), .C2(n5494), .A(n5491), .B(n9957), .ZN(n7474)
         );
  NAND2_X1 U5903 ( .A1(n10907), .A2(n5492), .ZN(n5491) );
  NOR2_X1 U5904 ( .A1(n5494), .A2(n5495), .ZN(n5492) );
  INV_X1 U5905 ( .A(n9951), .ZN(n5495) );
  OR2_X1 U5906 ( .A1(n10897), .A2(n9820), .ZN(n7478) );
  NAND2_X1 U5907 ( .A1(n5493), .A2(n6188), .ZN(n7472) );
  NAND2_X1 U5908 ( .A1(n10907), .A2(n9951), .ZN(n5493) );
  NAND2_X1 U5909 ( .A1(n9953), .A2(n9950), .ZN(n10071) );
  NAND2_X1 U5910 ( .A1(n9949), .A2(n7285), .ZN(n10905) );
  NOR2_X1 U5911 ( .A1(n7325), .A2(n9848), .ZN(n10898) );
  NAND2_X1 U5912 ( .A1(n9951), .A2(n9947), .ZN(n10903) );
  OR2_X1 U5913 ( .A1(n10438), .A2(n10274), .ZN(n7038) );
  OR2_X1 U5914 ( .A1(n5247), .A2(n7382), .ZN(n7325) );
  NAND2_X1 U5915 ( .A1(n10069), .A2(n7319), .ZN(n7318) );
  OR2_X1 U5916 ( .A1(n7283), .A2(n7282), .ZN(n7292) );
  OAI21_X1 U5917 ( .B1(n10347), .B2(n5543), .A(n5540), .ZN(n10313) );
  NAND2_X1 U5918 ( .A1(n5539), .A2(n5544), .ZN(n10315) );
  NAND2_X1 U5919 ( .A1(n6120), .A2(n6119), .ZN(n10350) );
  NAND2_X1 U5920 ( .A1(n6098), .A2(n6097), .ZN(n10491) );
  NAND2_X1 U5921 ( .A1(n6038), .A2(n6037), .ZN(n10507) );
  AND2_X1 U5922 ( .A1(n7917), .A2(n8045), .ZN(n10543) );
  OAI22_X1 U5923 ( .A1(n6777), .A2(n6772), .B1(n6776), .B2(n8662), .ZN(n5320)
         );
  NAND2_X1 U5924 ( .A1(n8661), .A2(n8656), .ZN(n8658) );
  NAND2_X1 U5925 ( .A1(n5692), .A2(n5314), .ZN(n5696) );
  AND2_X1 U5926 ( .A1(n5123), .A2(n5558), .ZN(n5314) );
  AND2_X1 U5927 ( .A1(n5560), .A2(n5559), .ZN(n5558) );
  INV_X1 U5928 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5559) );
  NAND2_X1 U5929 ( .A1(n6131), .A2(n6130), .ZN(n6136) );
  NAND2_X1 U5930 ( .A1(n6136), .A2(n6135), .ZN(n6149) );
  OR2_X1 U5931 ( .A1(n6217), .A2(n6216), .ZN(n6221) );
  NAND2_X1 U5932 ( .A1(n5937), .A2(n5692), .ZN(n6219) );
  NAND2_X1 U5933 ( .A1(n6049), .A2(n6048), .ZN(n6056) );
  NAND2_X1 U5934 ( .A1(n6056), .A2(n6055), .ZN(n6070) );
  XNOR2_X1 U5935 ( .A(n6225), .B(P1_IR_REG_21__SCAN_IN), .ZN(n10107) );
  AND2_X1 U5936 ( .A1(n5483), .A2(n5123), .ZN(n6177) );
  NOR2_X1 U5937 ( .A1(n5484), .A2(n5151), .ZN(n5483) );
  NAND2_X1 U5938 ( .A1(n5112), .A2(n5419), .ZN(n6016) );
  NAND2_X1 U5939 ( .A1(n5387), .A2(n5391), .ZN(n5961) );
  OR2_X1 U5940 ( .A1(n5921), .A2(n5125), .ZN(n5387) );
  NAND2_X1 U5941 ( .A1(n5406), .A2(n5649), .ZN(n5870) );
  NAND2_X1 U5942 ( .A1(n5647), .A2(n5146), .ZN(n5406) );
  NAND2_X1 U5943 ( .A1(n5647), .A2(n5646), .ZN(n5855) );
  OR2_X1 U5944 ( .A1(n5821), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5842) );
  XNOR2_X1 U5945 ( .A(n5628), .B(n8431), .ZN(n5786) );
  NAND2_X1 U5946 ( .A1(n6490), .A2(n6489), .ZN(n8773) );
  XNOR2_X1 U5947 ( .A(n9041), .B(n9050), .ZN(n9094) );
  NAND2_X1 U5948 ( .A1(n5579), .A2(n5582), .ZN(n9095) );
  OR2_X1 U5949 ( .A1(n5587), .A2(n5583), .ZN(n5579) );
  NAND2_X1 U5950 ( .A1(n6585), .A2(n6584), .ZN(n9105) );
  NAND2_X1 U5951 ( .A1(n5596), .A2(n5593), .ZN(n7953) );
  INV_X1 U5952 ( .A(n5595), .ZN(n5593) );
  NAND2_X1 U5953 ( .A1(n6460), .A2(n6459), .ZN(n8018) );
  NAND2_X1 U5954 ( .A1(n6627), .A2(n6626), .ZN(n9411) );
  XNOR2_X1 U5955 ( .A(n9056), .B(n9194), .ZN(n9133) );
  NAND2_X1 U5956 ( .A1(n9093), .A2(n9042), .ZN(n9141) );
  NAND2_X1 U5957 ( .A1(n5591), .A2(n5114), .ZN(n8002) );
  NAND2_X1 U5958 ( .A1(n5598), .A2(n5592), .ZN(n5591) );
  AOI21_X1 U5959 ( .B1(n5570), .B2(n5569), .A(n5568), .ZN(n5567) );
  NAND2_X1 U5960 ( .A1(n9093), .A2(n5197), .ZN(n5199) );
  INV_X1 U5961 ( .A(n9150), .ZN(n5568) );
  NAND2_X1 U5962 ( .A1(n5566), .A2(n5570), .ZN(n9151) );
  NAND2_X1 U5963 ( .A1(n9141), .A2(n5572), .ZN(n5566) );
  NAND2_X1 U5964 ( .A1(n7723), .A2(n7722), .ZN(n7724) );
  NAND2_X1 U5965 ( .A1(n5585), .A2(n5588), .ZN(n9159) );
  NAND2_X1 U5966 ( .A1(n5585), .A2(n5584), .ZN(n9160) );
  NAND2_X1 U5967 ( .A1(n7175), .A2(n7174), .ZN(n5189) );
  NAND2_X1 U5968 ( .A1(n6504), .A2(n6503), .ZN(n9553) );
  AOI21_X1 U5969 ( .B1(n8889), .B2(n8888), .A(n8887), .ZN(n8890) );
  NAND2_X1 U5970 ( .A1(n6635), .A2(n6634), .ZN(n9398) );
  INV_X1 U5971 ( .A(n9426), .ZN(n9448) );
  NAND4_X1 U5972 ( .A1(n6427), .A2(n6426), .A3(n6425), .A4(n6424), .ZN(n9200)
         );
  OR2_X1 U5973 ( .A1(n5110), .A2(n7818), .ZN(n6424) );
  NAND4_X1 U5974 ( .A1(n6372), .A2(n6371), .A3(n6370), .A4(n6369), .ZN(n9203)
         );
  OR2_X1 U5975 ( .A1(n5110), .A2(n7513), .ZN(n6353) );
  INV_X1 U5976 ( .A(P2_U3893), .ZN(n9331) );
  OR2_X1 U5977 ( .A1(n6338), .A2(n6828), .ZN(n6308) );
  NAND2_X1 U5978 ( .A1(n6845), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6875) );
  INV_X1 U5979 ( .A(n6846), .ZN(n6845) );
  NAND2_X1 U5980 ( .A1(n10838), .A2(n5185), .ZN(n10862) );
  OR2_X1 U5981 ( .A1(n7363), .A2(n10837), .ZN(n5185) );
  INV_X1 U5982 ( .A(n5424), .ZN(n10852) );
  INV_X1 U5983 ( .A(n7335), .ZN(n5423) );
  XNOR2_X1 U5984 ( .A(n7689), .B(n5306), .ZN(n7560) );
  OR2_X1 U5985 ( .A1(n7688), .A2(n7687), .ZN(n7780) );
  NOR2_X1 U5986 ( .A1(n7848), .A2(n7818), .ZN(n7847) );
  INV_X1 U5987 ( .A(n7900), .ZN(n7899) );
  INV_X1 U5988 ( .A(n5209), .ZN(n7785) );
  NAND2_X1 U5989 ( .A1(n7893), .A2(n7892), .ZN(n8076) );
  NAND2_X1 U5990 ( .A1(n8061), .A2(n8062), .ZN(n8063) );
  INV_X1 U5991 ( .A(n5429), .ZN(n9228) );
  XNOR2_X1 U5992 ( .A(n9241), .B(n9226), .ZN(n9207) );
  OAI21_X1 U5993 ( .B1(n9209), .B2(n5427), .A(n5426), .ZN(n9255) );
  NAND2_X1 U5994 ( .A1(n5430), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5427) );
  INV_X1 U5995 ( .A(n9230), .ZN(n5430) );
  INV_X1 U5996 ( .A(n9227), .ZN(n5428) );
  NOR2_X1 U5997 ( .A1(n9258), .A2(n9554), .ZN(n9275) );
  OAI21_X1 U5998 ( .B1(n9258), .B2(n5435), .A(n5434), .ZN(n9298) );
  NAND2_X1 U5999 ( .A1(n5436), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5435) );
  INV_X1 U6000 ( .A(n9277), .ZN(n5436) );
  XNOR2_X1 U6001 ( .A(n9320), .B(n9325), .ZN(n9299) );
  NOR2_X1 U6002 ( .A1(n9299), .A2(n9300), .ZN(n9322) );
  NAND2_X1 U6003 ( .A1(n5216), .A2(n5437), .ZN(n9346) );
  NAND2_X1 U6004 ( .A1(n9321), .A2(n5439), .ZN(n5437) );
  OR2_X1 U6005 ( .A1(n9299), .A2(n5438), .ZN(n5216) );
  NAND2_X1 U6006 ( .A1(n5439), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5438) );
  XNOR2_X1 U6007 ( .A(n5214), .B(n9351), .ZN(n5213) );
  NOR2_X1 U6008 ( .A1(n9346), .A2(n5215), .ZN(n5214) );
  NOR2_X1 U6009 ( .A1(n9349), .A2(n9507), .ZN(n5215) );
  AOI21_X1 U6010 ( .B1(n6677), .B2(n9399), .A(n6676), .ZN(n6678) );
  NOR2_X1 U6011 ( .A1(n8675), .A2(n9564), .ZN(n6676) );
  NAND2_X1 U6012 ( .A1(n9383), .A2(n9382), .ZN(n9384) );
  NAND2_X1 U6013 ( .A1(n5344), .A2(n5342), .ZN(n9394) );
  NAND2_X1 U6014 ( .A1(n5345), .A2(n6710), .ZN(n5344) );
  NAND2_X1 U6015 ( .A1(n6273), .A2(n6272), .ZN(n9406) );
  OAI21_X1 U6016 ( .B1(n9423), .B2(n6625), .A(n5297), .ZN(n9413) );
  NAND2_X1 U6017 ( .A1(n5360), .A2(n5358), .ZN(n9430) );
  NAND2_X1 U6018 ( .A1(n5360), .A2(n8822), .ZN(n9439) );
  NAND2_X1 U6019 ( .A1(n6594), .A2(n6593), .ZN(n9622) );
  NAND2_X1 U6020 ( .A1(n9496), .A2(n8800), .ZN(n9490) );
  NAND2_X1 U6021 ( .A1(n6516), .A2(n6515), .ZN(n9510) );
  NAND2_X1 U6022 ( .A1(n9533), .A2(n8787), .ZN(n9520) );
  NAND2_X1 U6023 ( .A1(n6696), .A2(n8769), .ZN(n9569) );
  OR3_X1 U6024 ( .A1(n6394), .A2(n6393), .A3(n6392), .ZN(n7661) );
  AND2_X1 U6025 ( .A1(n10944), .A2(n9417), .ZN(n10941) );
  AND2_X1 U6026 ( .A1(n6748), .A2(n8836), .ZN(n6928) );
  INV_X1 U6027 ( .A(n8885), .ZN(n9658) );
  INV_X1 U6028 ( .A(n8691), .ZN(n9661) );
  AND2_X1 U6029 ( .A1(n9598), .A2(n9597), .ZN(n9599) );
  AND2_X1 U6030 ( .A1(n5363), .A2(n6290), .ZN(n5362) );
  OR2_X1 U6031 ( .A1(n6716), .A2(n6715), .ZN(n6717) );
  INV_X1 U6032 ( .A(n10837), .ZN(n7338) );
  INV_X1 U6033 ( .A(n10815), .ZN(n7359) );
  NAND2_X1 U6034 ( .A1(n6319), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n6322) );
  NOR2_X1 U6035 ( .A1(n6261), .A2(n6320), .ZN(n6321) );
  NAND2_X1 U6036 ( .A1(n6306), .A2(n5221), .ZN(n6868) );
  MUX2_X1 U6037 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6305), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n6306) );
  AND2_X1 U6038 ( .A1(n6232), .A2(n6248), .ZN(n6227) );
  AND2_X1 U6039 ( .A1(n7429), .A2(n7428), .ZN(n7520) );
  NAND2_X1 U6040 ( .A1(n9856), .A2(n9857), .ZN(n9751) );
  NAND2_X1 U6041 ( .A1(n5990), .A2(n5989), .ZN(n10522) );
  AND2_X1 U6042 ( .A1(n5450), .A2(n5133), .ZN(n7979) );
  NAND2_X1 U6043 ( .A1(n5134), .A2(n9807), .ZN(n9772) );
  OAI21_X1 U6044 ( .B1(n8172), .B2(n5445), .A(n5443), .ZN(n9781) );
  NAND2_X1 U6045 ( .A1(n6075), .A2(n6074), .ZN(n10382) );
  NAND2_X1 U6046 ( .A1(n5446), .A2(n5447), .ZN(n8122) );
  AND2_X1 U6047 ( .A1(n8031), .A2(n5448), .ZN(n5447) );
  NAND2_X1 U6048 ( .A1(n7974), .A2(n5111), .ZN(n5446) );
  NAND2_X1 U6049 ( .A1(n7242), .A2(n7241), .ZN(n7244) );
  NAND2_X1 U6050 ( .A1(n5454), .A2(n5452), .ZN(n9870) );
  NOR2_X1 U6051 ( .A1(n5150), .A2(n5453), .ZN(n5452) );
  NAND2_X1 U6052 ( .A1(n8172), .A2(n8171), .ZN(n8902) );
  AND2_X1 U6053 ( .A1(n5764), .A2(n5765), .ZN(n5246) );
  NAND2_X1 U6054 ( .A1(n9885), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5248) );
  INV_X1 U6055 ( .A(n5250), .ZN(n5249) );
  NAND2_X1 U6056 ( .A1(n5118), .A2(n11035), .ZN(n10470) );
  AOI21_X1 U6057 ( .B1(n5501), .B2(n10402), .A(n5499), .ZN(n10305) );
  OAI21_X1 U6058 ( .B1(n10326), .B2(n10900), .A(n5500), .ZN(n5499) );
  XNOR2_X1 U6059 ( .A(n5503), .B(n5502), .ZN(n5501) );
  NAND2_X1 U6060 ( .A1(n10286), .A2(n10155), .ZN(n5500) );
  AOI21_X1 U6061 ( .B1(n5540), .B2(n5543), .A(n5171), .ZN(n5538) );
  AND2_X1 U6062 ( .A1(n5490), .A2(n10037), .ZN(n10374) );
  NAND2_X1 U6063 ( .A1(n5526), .A2(n5524), .ZN(n10390) );
  NAND2_X1 U6064 ( .A1(n10427), .A2(n5527), .ZN(n5526) );
  AOI21_X1 U6065 ( .B1(n10427), .B2(n10428), .A(n5529), .ZN(n10406) );
  NAND2_X1 U6066 ( .A1(n5551), .A2(n5553), .ZN(n7992) );
  NAND2_X1 U6067 ( .A1(n5953), .A2(n5952), .ZN(n9789) );
  NAND2_X1 U6068 ( .A1(n5552), .A2(n5934), .ZN(n8619) );
  OR2_X1 U6069 ( .A1(n7911), .A2(n5933), .ZN(n5552) );
  NAND2_X1 U6070 ( .A1(n7538), .A2(n9968), .ZN(n7537) );
  NAND2_X1 U6071 ( .A1(n7302), .A2(n5820), .ZN(n7538) );
  INV_X1 U6072 ( .A(n11056), .ZN(n10440) );
  INV_X1 U6073 ( .A(n10335), .ZN(n11045) );
  INV_X1 U6074 ( .A(n8052), .ZN(n10532) );
  AND2_X1 U6075 ( .A1(n10470), .A2(n10469), .ZN(n10549) );
  INV_X1 U6076 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n5239) );
  NAND2_X1 U6077 ( .A1(n10472), .A2(n5241), .ZN(n10552) );
  INV_X1 U6078 ( .A(n5242), .ZN(n5241) );
  OAI21_X1 U6079 ( .B1(n10473), .B2(n10543), .A(n10471), .ZN(n5242) );
  NAND2_X1 U6080 ( .A1(n6151), .A2(n6150), .ZN(n10553) );
  INV_X1 U6081 ( .A(n10350), .ZN(n10562) );
  XNOR2_X1 U6082 ( .A(n8666), .B(n8665), .ZN(n10593) );
  NAND2_X1 U6083 ( .A1(n8661), .A2(n8660), .ZN(n8666) );
  INV_X1 U6084 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n10588) );
  AND2_X1 U6085 ( .A1(n5266), .A2(n5123), .ZN(n5265) );
  AND2_X1 U6086 ( .A1(n5162), .A2(n5115), .ZN(n5266) );
  NOR2_X1 U6087 ( .A1(n6772), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10592) );
  OR2_X1 U6088 ( .A1(n5705), .A2(n5905), .ZN(n5244) );
  NAND2_X1 U6089 ( .A1(n5692), .A2(n5115), .ZN(n5268) );
  XNOR2_X1 U6090 ( .A(n6161), .B(n6160), .ZN(n8609) );
  NAND2_X1 U6091 ( .A1(n6149), .A2(n6148), .ZN(n6161) );
  NAND2_X1 U6092 ( .A1(n6149), .A2(n6137), .ZN(n8134) );
  OR2_X1 U6093 ( .A1(n6136), .A2(n6135), .ZN(n6137) );
  NAND2_X1 U6094 ( .A1(n5123), .A2(n5684), .ZN(n5922) );
  AND2_X1 U6095 ( .A1(n5785), .A2(n5784), .ZN(n10242) );
  INV_X1 U6096 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7276) );
  XNOR2_X1 U6097 ( .A(n5196), .B(n9068), .ZN(n9074) );
  AOI21_X1 U6098 ( .B1(n5179), .B2(n7337), .A(n5211), .ZN(n7377) );
  OAI211_X1 U6099 ( .C1(n5313), .C2(n10833), .A(n5312), .B(n5311), .ZN(
        P2_U3201) );
  XNOR2_X1 U6100 ( .A(n9360), .B(n9359), .ZN(n5313) );
  AOI21_X1 U6101 ( .B1(n9362), .B2(n10859), .A(n9361), .ZN(n5312) );
  NAND2_X1 U6102 ( .A1(n5213), .A2(n6858), .ZN(n5311) );
  AOI21_X1 U6103 ( .B1(n5253), .B2(n5251), .A(n10152), .ZN(n10154) );
  INV_X1 U6104 ( .A(n5252), .ZN(n5251) );
  OAI21_X1 U6105 ( .B1(n10549), .B2(n11080), .A(n5321), .ZN(P1_U3552) );
  INV_X1 U6106 ( .A(n5322), .ZN(n5321) );
  OAI22_X1 U6107 ( .A1(n10551), .A2(n10532), .B1(n6208), .B2(n11081), .ZN(
        n5322) );
  NAND2_X1 U6108 ( .A1(n5240), .A2(n5237), .ZN(P1_U3518) );
  AOI21_X1 U6109 ( .B1(n10553), .B2(n10557), .A(n5238), .ZN(n5237) );
  NAND2_X1 U6110 ( .A1(n10552), .A2(n11085), .ZN(n5240) );
  NOR2_X1 U6111 ( .A1(n11085), .A2(n5239), .ZN(n5238) );
  BUF_X1 U6112 ( .A(n6338), .Z(n8680) );
  AND2_X1 U6113 ( .A1(n5133), .A2(n7980), .ZN(n5111) );
  AND4_X1 U6114 ( .A1(n6343), .A2(n6342), .A3(n6341), .A4(n6340), .ZN(n7156)
         );
  OR2_X1 U6115 ( .A1(n5980), .A2(n5979), .ZN(n5112) );
  INV_X1 U6116 ( .A(n6307), .ZN(n6518) );
  OR2_X1 U6117 ( .A1(n5462), .A2(n9808), .ZN(n5113) );
  OR2_X1 U6118 ( .A1(n5594), .A2(n5153), .ZN(n5114) );
  NOR2_X1 U6119 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n5115) );
  AND4_X1 U6120 ( .A1(n6382), .A2(n6259), .A3(n6258), .A4(n6257), .ZN(n5116)
         );
  INV_X1 U6121 ( .A(n7927), .ZN(n5597) );
  OR2_X1 U6122 ( .A1(n5476), .A2(n5475), .ZN(n5117) );
  INV_X1 U6123 ( .A(n9039), .ZN(n5586) );
  INV_X2 U6124 ( .A(n5618), .ZN(n6772) );
  XOR2_X1 U6125 ( .A(n10291), .B(n10290), .Z(n5118) );
  AND2_X1 U6126 ( .A1(n5325), .A2(n5324), .ZN(n5119) );
  NAND2_X1 U6127 ( .A1(n6059), .A2(n6058), .ZN(n10501) );
  AND2_X1 U6128 ( .A1(n5114), .A2(n5175), .ZN(n5120) );
  OR2_X1 U6129 ( .A1(n8172), .A2(n8171), .ZN(n5121) );
  AND2_X1 U6130 ( .A1(n8662), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5122) );
  NAND2_X1 U6131 ( .A1(n6955), .A2(n7043), .ZN(n6956) );
  INV_X1 U6132 ( .A(n9000), .ZN(n8991) );
  NAND2_X1 U6133 ( .A1(n5707), .A2(n5708), .ZN(n5776) );
  OR2_X1 U6134 ( .A1(n6690), .A2(n8750), .ZN(n5124) );
  OR2_X1 U6135 ( .A1(n5948), .A2(n5393), .ZN(n5125) );
  NAND2_X1 U6136 ( .A1(n8721), .A2(n5334), .ZN(n8855) );
  AND2_X1 U6137 ( .A1(n5218), .A2(n5217), .ZN(n5126) );
  OAI211_X1 U6138 ( .C1(n6313), .C2(n7359), .A(n6333), .B(n6332), .ZN(n10933)
         );
  NAND2_X1 U6139 ( .A1(n6664), .A2(n6267), .ZN(n5127) );
  NOR2_X1 U6140 ( .A1(n9816), .A2(n7240), .ZN(n5128) );
  AND2_X1 U6141 ( .A1(n9045), .A2(n9471), .ZN(n5129) );
  AND2_X1 U6142 ( .A1(n7032), .A2(n7021), .ZN(n7759) );
  NOR2_X1 U6143 ( .A1(n9092), .A2(n9196), .ZN(n5130) );
  NAND2_X1 U6144 ( .A1(n5482), .A2(n5123), .ZN(n5131) );
  INV_X1 U6145 ( .A(n10428), .ZN(n5528) );
  INV_X1 U6146 ( .A(n9195), .ZN(n9488) );
  AND2_X1 U6147 ( .A1(n6267), .A2(n6662), .ZN(n5132) );
  XNOR2_X1 U6148 ( .A(n5648), .B(n8427), .ZN(n5854) );
  NAND2_X1 U6149 ( .A1(n9139), .A2(n9044), .ZN(n9100) );
  XNOR2_X1 U6150 ( .A(n9051), .B(n9052), .ZN(n9085) );
  XNOR2_X1 U6151 ( .A(n5612), .B(n8441), .ZN(n5715) );
  NAND2_X1 U6152 ( .A1(n5517), .A2(n5514), .ZN(n10427) );
  INV_X1 U6153 ( .A(n10079), .ZN(n5509) );
  NAND2_X1 U6154 ( .A1(n7978), .A2(n7977), .ZN(n5133) );
  INV_X1 U6155 ( .A(n7352), .ZN(n7557) );
  NAND4_X1 U6156 ( .A1(n6311), .A2(n6310), .A3(n6309), .A4(n6308), .ZN(n6912)
         );
  AND2_X1 U6157 ( .A1(n5719), .A2(n5319), .ZN(n5729) );
  XNOR2_X1 U6158 ( .A(n5704), .B(n10588), .ZN(n5707) );
  NOR2_X1 U6159 ( .A1(n6442), .A2(n6266), .ZN(n6664) );
  OAI211_X1 U6160 ( .C1(n8656), .C2(n6377), .A(n8659), .B(n5372), .ZN(n8691)
         );
  OR2_X1 U6161 ( .A1(n9810), .A2(n9808), .ZN(n5134) );
  NAND2_X1 U6162 ( .A1(n9064), .A2(n9063), .ZN(n9075) );
  NAND2_X1 U6163 ( .A1(n10360), .A2(n5330), .ZN(n5135) );
  NAND2_X1 U6164 ( .A1(n9092), .A2(n9196), .ZN(n5136) );
  OR2_X1 U6165 ( .A1(n10501), .A2(n10376), .ZN(n5137) );
  NOR2_X1 U6166 ( .A1(n9322), .A2(n9321), .ZN(n5138) );
  NAND2_X1 U6167 ( .A1(n5940), .A2(n5939), .ZN(n10540) );
  NOR2_X1 U6168 ( .A1(n10119), .A2(n10118), .ZN(n5139) );
  NAND2_X1 U6169 ( .A1(n5304), .A2(n5364), .ZN(n6722) );
  NAND2_X1 U6170 ( .A1(n6664), .A2(n5132), .ZN(n6660) );
  AND2_X1 U6171 ( .A1(n10373), .A2(n10048), .ZN(n5140) );
  INV_X4 U6172 ( .A(n6772), .ZN(n8662) );
  NOR2_X1 U6173 ( .A1(n9981), .A2(n10060), .ZN(n5141) );
  INV_X1 U6174 ( .A(n10969), .ZN(n7482) );
  AND2_X1 U6175 ( .A1(n5789), .A2(n5788), .ZN(n10969) );
  AND2_X1 U6176 ( .A1(n7182), .A2(n7178), .ZN(n5142) );
  AND2_X1 U6177 ( .A1(n9036), .A2(n9529), .ZN(n5143) );
  XNOR2_X1 U6178 ( .A(n5655), .B(n8415), .ZN(n5886) );
  NAND2_X1 U6179 ( .A1(n9759), .A2(n8946), .ZN(n5144) );
  INV_X1 U6180 ( .A(n10556), .ZN(n10484) );
  NAND2_X1 U6181 ( .A1(n6139), .A2(n6138), .ZN(n10556) );
  OR2_X1 U6182 ( .A1(n5144), .A2(n9757), .ZN(n5145) );
  NAND2_X1 U6183 ( .A1(n6165), .A2(n6164), .ZN(n10299) );
  INV_X1 U6184 ( .A(n5571), .ZN(n5570) );
  NOR2_X1 U6185 ( .A1(n5573), .A2(n5129), .ZN(n5571) );
  AND2_X1 U6186 ( .A1(n5646), .A2(n5854), .ZN(n5146) );
  AND2_X1 U6187 ( .A1(n10308), .A2(n10054), .ZN(n5147) );
  NAND2_X1 U6188 ( .A1(n6708), .A2(n9429), .ZN(n5148) );
  INV_X1 U6189 ( .A(n5589), .ZN(n5588) );
  AND2_X1 U6190 ( .A1(n8693), .A2(n8694), .ZN(n9395) );
  INV_X1 U6191 ( .A(n9395), .ZN(n5343) );
  NAND2_X1 U6192 ( .A1(n9406), .A2(n9381), .ZN(n5149) );
  NAND2_X1 U6193 ( .A1(n5463), .A2(n5460), .ZN(n5150) );
  NAND3_X1 U6194 ( .A1(n6175), .A2(n6174), .A3(n8573), .ZN(n5151) );
  NOR2_X1 U6195 ( .A1(n7549), .A2(n10165), .ZN(n5152) );
  AND2_X1 U6196 ( .A1(n7930), .A2(n9578), .ZN(n5153) );
  INV_X1 U6197 ( .A(n5531), .ZN(n5529) );
  NAND2_X1 U6198 ( .A1(n10573), .A2(n10449), .ZN(n5531) );
  NOR2_X1 U6199 ( .A1(n8864), .A2(n6690), .ZN(n5154) );
  NOR2_X1 U6200 ( .A1(n9040), .A2(n9487), .ZN(n5155) );
  OR2_X1 U6201 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5156) );
  NAND2_X1 U6202 ( .A1(n5655), .A2(SI_12_), .ZN(n5157) );
  OR2_X1 U6203 ( .A1(n9411), .A2(n9398), .ZN(n5158) );
  OR2_X1 U6204 ( .A1(n5299), .A2(n5122), .ZN(n5159) );
  INV_X1 U6205 ( .A(n7175), .ZN(n5192) );
  NAND2_X1 U6206 ( .A1(n5291), .A2(n5149), .ZN(n5160) );
  AND2_X1 U6207 ( .A1(n5154), .A2(n8740), .ZN(n5161) );
  NOR2_X1 U6208 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n6382) );
  AND2_X1 U6209 ( .A1(n5560), .A2(n8369), .ZN(n5162) );
  NAND2_X1 U6210 ( .A1(n5701), .A2(n5700), .ZN(n9864) );
  AND2_X1 U6211 ( .A1(n7519), .A2(n7428), .ZN(n5163) );
  INV_X1 U6212 ( .A(n5337), .ZN(n5336) );
  AND2_X1 U6213 ( .A1(n5344), .A2(n5341), .ZN(n5164) );
  AND2_X1 U6214 ( .A1(n6691), .A2(n5124), .ZN(n5165) );
  INV_X1 U6215 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6260) );
  INV_X1 U6216 ( .A(n9961), .ZN(n5534) );
  INV_X1 U6217 ( .A(n7928), .ZN(n5598) );
  INV_X1 U6218 ( .A(n9126), .ZN(n5587) );
  INV_X1 U6219 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n5411) );
  INV_X1 U6220 ( .A(n8942), .ZN(n5475) );
  INV_X1 U6221 ( .A(n9399), .ZN(n9174) );
  NAND2_X1 U6222 ( .A1(n6649), .A2(n6648), .ZN(n9399) );
  AND2_X1 U6223 ( .A1(n8623), .A2(n5119), .ZN(n5166) );
  NAND2_X1 U6224 ( .A1(n6651), .A2(n6650), .ZN(n9072) );
  INV_X1 U6225 ( .A(n7690), .ZN(n5306) );
  AND2_X1 U6226 ( .A1(n5419), .A2(n6015), .ZN(n5167) );
  INV_X1 U6227 ( .A(n9807), .ZN(n5461) );
  NAND2_X1 U6228 ( .A1(n7449), .A2(n5868), .ZN(n11020) );
  AND2_X1 U6229 ( .A1(n10004), .A2(n10006), .ZN(n10089) );
  INV_X1 U6230 ( .A(n10089), .ZN(n5550) );
  NAND2_X1 U6231 ( .A1(n6502), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6514) );
  INV_X1 U6232 ( .A(n10124), .ZN(n5229) );
  INV_X1 U6233 ( .A(n5315), .ZN(n10407) );
  NOR3_X1 U6234 ( .A1(n10439), .A2(n10432), .A3(n5317), .ZN(n5315) );
  NOR2_X1 U6235 ( .A1(n8067), .A2(n8066), .ZN(n5168) );
  NOR2_X1 U6236 ( .A1(n9275), .A2(n9276), .ZN(n5169) );
  AND2_X1 U6237 ( .A1(n5596), .A2(n5594), .ZN(n5170) );
  AND2_X1 U6238 ( .A1(n10553), .A2(n6159), .ZN(n5171) );
  NOR2_X1 U6239 ( .A1(n8018), .A2(n9578), .ZN(n5172) );
  AND2_X1 U6240 ( .A1(n5429), .A2(n5428), .ZN(n5173) );
  INV_X1 U6241 ( .A(n5267), .ZN(n5937) );
  NAND2_X1 U6242 ( .A1(n5123), .A2(n5560), .ZN(n5267) );
  NAND2_X1 U6243 ( .A1(n6014), .A2(n6013), .ZN(n5174) );
  INV_X1 U6244 ( .A(n11080), .ZN(n11081) );
  NAND2_X1 U6245 ( .A1(n6005), .A2(n6004), .ZN(n10517) );
  INV_X1 U6246 ( .A(n10517), .ZN(n5318) );
  NAND2_X1 U6247 ( .A1(n5507), .A2(n5510), .ZN(n7636) );
  INV_X1 U6248 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5205) );
  OR2_X1 U6249 ( .A1(n7931), .A2(n9197), .ZN(n5175) );
  NAND2_X1 U6250 ( .A1(n5965), .A2(n5964), .ZN(n10535) );
  INV_X1 U6251 ( .A(n10535), .ZN(n5324) );
  INV_X1 U6252 ( .A(n8171), .ZN(n8170) );
  AND2_X1 U6253 ( .A1(n7411), .A2(n7410), .ZN(n7714) );
  NAND2_X1 U6254 ( .A1(n7193), .A2(n7178), .ZN(n7180) );
  AND2_X1 U6255 ( .A1(n9264), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5176) );
  NAND2_X1 U6256 ( .A1(n6664), .A2(n5564), .ZN(n5177) );
  AND2_X1 U6257 ( .A1(n6163), .A2(n8396), .ZN(n5178) );
  XNOR2_X1 U6258 ( .A(n5694), .B(n5693), .ZN(n6210) );
  OAI211_X1 U6259 ( .C1(n9887), .C2(n6977), .A(n5763), .B(n5246), .ZN(n9745)
         );
  INV_X1 U6260 ( .A(n9745), .ZN(n5245) );
  INV_X1 U6261 ( .A(n7549), .ZN(n5326) );
  AND2_X1 U6262 ( .A1(n5424), .A2(n5423), .ZN(n5179) );
  AND2_X1 U6263 ( .A1(n10138), .A2(n7066), .ZN(n11027) );
  AND2_X1 U6264 ( .A1(n7157), .A2(n7169), .ZN(n7159) );
  AND2_X1 U6265 ( .A1(n6772), .A2(P2_U3151), .ZN(n5180) );
  NAND2_X1 U6266 ( .A1(n5692), .A2(n5265), .ZN(n10587) );
  INV_X1 U6267 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5371) );
  INV_X2 U6268 ( .A(n5180), .ZN(n9719) );
  NAND2_X2 U6269 ( .A1(n6849), .A2(n6260), .ZN(n6386) );
  INV_X1 U6270 ( .A(n5183), .ZN(n7857) );
  NOR2_X1 U6271 ( .A1(n7701), .A2(n7700), .ZN(n7788) );
  NAND3_X1 U6272 ( .A1(n5189), .A2(n5188), .A3(n5142), .ZN(n7411) );
  NAND2_X1 U6273 ( .A1(n7176), .A2(n7174), .ZN(n5188) );
  NAND2_X1 U6274 ( .A1(n5190), .A2(n7174), .ZN(n7193) );
  NAND2_X1 U6275 ( .A1(n5193), .A2(n5192), .ZN(n5190) );
  NAND2_X1 U6276 ( .A1(n7714), .A2(n5191), .ZN(n7718) );
  NAND2_X1 U6277 ( .A1(n9077), .A2(n9066), .ZN(n5196) );
  OAI22_X2 U6278 ( .A1(n9034), .A2(n9033), .B1(n9032), .B2(n9577), .ZN(n9186)
         );
  AOI21_X2 U6279 ( .B1(n8633), .B2(n7962), .A(n7726), .ZN(n7928) );
  NOR2_X2 U6280 ( .A1(n9184), .A2(n5143), .ZN(n9117) );
  NAND3_X1 U6281 ( .A1(n6955), .A2(n7043), .A3(n6957), .ZN(n7044) );
  NAND2_X1 U6282 ( .A1(n7044), .A2(n7043), .ZN(n7045) );
  NAND2_X2 U6283 ( .A1(n5207), .A2(n6948), .ZN(n7152) );
  NAND2_X1 U6284 ( .A1(n9276), .A2(n5436), .ZN(n5434) );
  INV_X1 U6285 ( .A(n6849), .ZN(n5221) );
  NAND4_X1 U6286 ( .A1(n5683), .A2(n5682), .A3(n5680), .A4(n5681), .ZN(n5236)
         );
  NAND3_X1 U6287 ( .A1(n5766), .A2(n5739), .A3(n5679), .ZN(n5783) );
  INV_X1 U6288 ( .A(n10069), .ZN(n6184) );
  INV_X2 U6289 ( .A(n5729), .ZN(n5247) );
  NAND3_X1 U6291 ( .A1(n10123), .A2(n10140), .A3(n10121), .ZN(n5257) );
  NOR2_X1 U6292 ( .A1(n5267), .A2(n5268), .ZN(n5705) );
  NAND3_X1 U6293 ( .A1(n5273), .A2(n5270), .A3(n10329), .ZN(n5269) );
  NAND3_X1 U6294 ( .A1(n10051), .A2(n10055), .A3(n10050), .ZN(n5273) );
  AOI21_X2 U6295 ( .B1(n5285), .B2(n10928), .A(n9022), .ZN(n9600) );
  XNOR2_X1 U6296 ( .A(n5286), .B(n9017), .ZN(n5285) );
  OAI21_X1 U6297 ( .B1(n9015), .B2(n9014), .A(n9013), .ZN(n5286) );
  NAND2_X1 U6298 ( .A1(n9423), .A2(n5289), .ZN(n5287) );
  OR2_X1 U6299 ( .A1(n9421), .A2(n9194), .ZN(n5297) );
  NAND2_X1 U6300 ( .A1(n6313), .A2(n6772), .ZN(n6377) );
  NAND2_X2 U6301 ( .A1(n6313), .A2(n8662), .ZN(n6360) );
  NAND2_X1 U6302 ( .A1(n7511), .A2(n7171), .ZN(n6363) );
  OAI22_X2 U6303 ( .A1(n7390), .A2(n5301), .B1(n5300), .B2(n7156), .ZN(n7511)
         );
  NAND2_X4 U6304 ( .A1(n6210), .A2(n10660), .ZN(n6803) );
  NAND2_X1 U6305 ( .A1(n6803), .A2(n5320), .ZN(n5319) );
  NAND2_X2 U6306 ( .A1(n6803), .A2(n6772), .ZN(n9895) );
  NAND3_X1 U6307 ( .A1(n5328), .A2(n5327), .A3(n5326), .ZN(n7548) );
  AND2_X1 U6308 ( .A1(n10360), .A2(n10562), .ZN(n10348) );
  OAI21_X1 U6309 ( .B1(n5337), .B2(n5335), .A(n10938), .ZN(n5334) );
  INV_X1 U6310 ( .A(n6331), .ZN(n5335) );
  NAND3_X1 U6311 ( .A1(n6329), .A2(n6330), .A3(n6328), .ZN(n5337) );
  NAND2_X1 U6312 ( .A1(n9410), .A2(n5342), .ZN(n5340) );
  INV_X1 U6313 ( .A(n9410), .ZN(n5345) );
  NAND2_X1 U6314 ( .A1(n5346), .A2(n5347), .ZN(n9472) );
  NAND2_X1 U6315 ( .A1(n9497), .A2(n5349), .ZN(n5346) );
  NAND2_X1 U6316 ( .A1(n5353), .A2(n5354), .ZN(n6703) );
  NAND2_X1 U6317 ( .A1(n9535), .A2(n8787), .ZN(n5353) );
  OAI21_X1 U6318 ( .B1(n9450), .B2(n5357), .A(n5355), .ZN(n6709) );
  NAND2_X1 U6319 ( .A1(n6696), .A2(n5361), .ZN(n9567) );
  AND2_X1 U6320 ( .A1(n6271), .A2(n5363), .ZN(n6289) );
  NAND2_X1 U6321 ( .A1(n6271), .A2(n5362), .ZN(n9710) );
  NAND2_X1 U6322 ( .A1(n6271), .A2(n6268), .ZN(n5562) );
  NOR2_X2 U6323 ( .A1(n6442), .A2(n5156), .ZN(n5364) );
  NAND2_X1 U6324 ( .A1(n5366), .A2(n5165), .ZN(n6695) );
  NAND2_X1 U6325 ( .A1(n6689), .A2(n5161), .ZN(n5366) );
  NAND3_X1 U6326 ( .A1(n5368), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n5367) );
  NAND3_X1 U6327 ( .A1(n7276), .A2(n5371), .A3(n5370), .ZN(n5369) );
  NAND2_X1 U6328 ( .A1(n8653), .A2(n8652), .ZN(n8661) );
  NAND2_X1 U6329 ( .A1(n8653), .A2(n5373), .ZN(n5372) );
  NAND3_X1 U6330 ( .A1(n5374), .A2(n8890), .A3(n8891), .ZN(n8893) );
  NAND3_X1 U6331 ( .A1(n5375), .A2(n8850), .A3(n8849), .ZN(n5374) );
  NAND2_X1 U6332 ( .A1(n6056), .A2(n5379), .ZN(n5378) );
  NAND2_X1 U6333 ( .A1(n5921), .A2(n5391), .ZN(n5390) );
  NAND3_X1 U6334 ( .A1(n5646), .A2(n5854), .A3(n5654), .ZN(n5402) );
  MUX2_X1 U6335 ( .A(n7665), .B(n7668), .S(n6772), .Z(n6031) );
  MUX2_X1 U6336 ( .A(n8043), .B(n8617), .S(n6772), .Z(n6091) );
  MUX2_X1 U6337 ( .A(n8106), .B(n8105), .S(n6772), .Z(n6113) );
  MUX2_X1 U6338 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n6772), .Z(n6162) );
  MUX2_X1 U6339 ( .A(n9894), .B(n9030), .S(n6772), .Z(n8649) );
  XNOR2_X1 U6340 ( .A(n7334), .B(n10847), .ZN(n10853) );
  NAND2_X1 U6341 ( .A1(n9227), .A2(n5430), .ZN(n5426) );
  INV_X1 U6342 ( .A(n5440), .ZN(n9780) );
  AOI21_X1 U6343 ( .B1(n8971), .B2(n8970), .A(n8969), .ZN(n9810) );
  NAND2_X1 U6344 ( .A1(n8971), .A2(n5455), .ZN(n5454) );
  INV_X1 U6345 ( .A(n8969), .ZN(n5464) );
  NAND2_X1 U6346 ( .A1(n5479), .A2(n5477), .ZN(n7033) );
  NAND3_X1 U6347 ( .A1(n7030), .A2(n9001), .A3(n9002), .ZN(n5477) );
  NAND2_X2 U6348 ( .A1(n9001), .A2(n9002), .ZN(n9000) );
  NAND2_X1 U6349 ( .A1(n7429), .A2(n5163), .ZN(n7522) );
  NAND2_X1 U6350 ( .A1(n7638), .A2(n10083), .ZN(n5498) );
  NAND2_X1 U6351 ( .A1(n7912), .A2(n6196), .ZN(n6197) );
  NAND2_X1 U6352 ( .A1(n5761), .A2(n5760), .ZN(n7457) );
  NAND2_X1 U6353 ( .A1(n5761), .A2(n5505), .ZN(n5504) );
  INV_X1 U6354 ( .A(n5760), .ZN(n5506) );
  NAND2_X1 U6355 ( .A1(n7450), .A2(n5508), .ZN(n5507) );
  NAND2_X1 U6356 ( .A1(n7300), .A2(n5533), .ZN(n5532) );
  AND2_X1 U6357 ( .A1(n9961), .A2(n9968), .ZN(n5533) );
  NAND2_X1 U6358 ( .A1(n10347), .A2(n5540), .ZN(n5537) );
  NAND2_X1 U6359 ( .A1(n5537), .A2(n5538), .ZN(n6173) );
  NAND2_X1 U6360 ( .A1(n10347), .A2(n5547), .ZN(n5539) );
  AOI21_X1 U6361 ( .B1(n10347), .B2(n6202), .A(n6129), .ZN(n10330) );
  NAND2_X1 U6362 ( .A1(n7911), .A2(n5556), .ZN(n5551) );
  NAND2_X1 U6363 ( .A1(n5562), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6270) );
  OAI21_X2 U6364 ( .B1(n9126), .B2(n5578), .A(n5580), .ZN(n9093) );
  NOR2_X1 U6365 ( .A1(n9038), .A2(n9530), .ZN(n5589) );
  XNOR2_X1 U6366 ( .A(n8642), .B(SI_29_), .ZN(n9716) );
  INV_X1 U6367 ( .A(n8855), .ZN(n10932) );
  INV_X1 U6368 ( .A(n8857), .ZN(n6681) );
  OR2_X1 U6369 ( .A1(n9889), .A2(n5732), .ZN(n5733) );
  XNOR2_X1 U6370 ( .A(n7720), .B(n7719), .ZN(n8633) );
  NAND2_X1 U6371 ( .A1(n7718), .A2(n7717), .ZN(n7720) );
  XNOR2_X1 U6372 ( .A(n9015), .B(n9067), .ZN(n6679) );
  NOR2_X1 U6373 ( .A1(n7388), .A2(n6684), .ZN(n6685) );
  NAND2_X1 U6374 ( .A1(n7976), .A2(n7975), .ZN(n5599) );
  OR2_X1 U6375 ( .A1(n9875), .A2(n10365), .ZN(n5600) );
  OR2_X1 U6376 ( .A1(n7032), .A2(n7031), .ZN(n5601) );
  OR2_X1 U6377 ( .A1(n7799), .A2(n7779), .ZN(n5603) );
  INV_X1 U6378 ( .A(n8849), .ZN(n8888) );
  AND4_X1 U6379 ( .A1(n6158), .A2(n6157), .A3(n6156), .A4(n6155), .ZN(n10326)
         );
  OR2_X1 U6380 ( .A1(n6960), .A2(n8847), .ZN(n9562) );
  INV_X1 U6381 ( .A(n9562), .ZN(n6677) );
  INV_X1 U6382 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5609) );
  INV_X1 U6383 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n5627) );
  INV_X1 U6384 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5905) );
  INV_X1 U6385 ( .A(n10553), .ZN(n10477) );
  INV_X1 U6386 ( .A(n11093), .ZN(n11017) );
  OR2_X1 U6387 ( .A1(n6313), .A2(n6868), .ZN(n5604) );
  INV_X1 U6388 ( .A(n6213), .ZN(n10391) );
  NAND2_X1 U6389 ( .A1(n8843), .A2(n8842), .ZN(n9016) );
  AND2_X1 U6390 ( .A1(n9411), .A2(n9425), .ZN(n5605) );
  NAND2_X1 U6391 ( .A1(n7201), .A2(n7202), .ZN(n7200) );
  NOR2_X1 U6392 ( .A1(n6570), .A2(n9482), .ZN(n5606) );
  NOR3_X1 U6393 ( .A1(n10127), .A2(n10125), .A3(n9933), .ZN(n5607) );
  INV_X1 U6394 ( .A(n10529), .ZN(n11080) );
  INV_X1 U6395 ( .A(n9460), .ZN(n9047) );
  INV_X1 U6396 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n6262) );
  INV_X1 U6397 ( .A(n6575), .ZN(n6283) );
  INV_X1 U6398 ( .A(n9585), .ZN(n6483) );
  INV_X1 U6399 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6267) );
  INV_X1 U6400 ( .A(n10326), .ZN(n6159) );
  OR2_X1 U6401 ( .A1(n8645), .A2(n8644), .ZN(n8646) );
  INV_X1 U6402 ( .A(n5903), .ZN(n5656) );
  INV_X1 U6403 ( .A(n7181), .ZN(n7182) );
  AND2_X1 U6404 ( .A1(n6640), .A2(n9169), .ZN(n6641) );
  NOR2_X1 U6405 ( .A1(n10837), .A2(n7392), .ZN(n7333) );
  INV_X1 U6406 ( .A(n9536), .ZN(n6701) );
  INV_X1 U6407 ( .A(n6475), .ZN(n6279) );
  OR2_X1 U6408 ( .A1(n8680), .A2(n6337), .ZN(n6342) );
  NAND2_X1 U6409 ( .A1(n7054), .A2(n7053), .ZN(n7057) );
  OR2_X1 U6410 ( .A1(n8951), .A2(n8950), .ZN(n8952) );
  INV_X1 U6411 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5813) );
  NAND2_X1 U6412 ( .A1(n7452), .A2(n5509), .ZN(n11022) );
  INV_X1 U6413 ( .A(n8655), .ZN(n8653) );
  INV_X1 U6414 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5698) );
  AND2_X1 U6415 ( .A1(n5836), .A2(n5839), .ZN(n5644) );
  NAND2_X1 U6416 ( .A1(n5618), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5608) );
  INV_X1 U6417 ( .A(n6558), .ZN(n6282) );
  INV_X1 U6418 ( .A(n7722), .ZN(n7719) );
  OR2_X1 U6419 ( .A1(n6652), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6670) );
  NAND2_X1 U6420 ( .A1(n6586), .A2(n6284), .ZN(n6595) );
  NAND2_X1 U6421 ( .A1(n6281), .A2(n8476), .ZN(n6531) );
  NAND2_X1 U6422 ( .A1(n6278), .A2(n8255), .ZN(n6475) );
  NAND2_X1 U6423 ( .A1(n6277), .A2(n8480), .ZN(n6435) );
  NAND2_X1 U6424 ( .A1(n7758), .A2(n7757), .ZN(n7766) );
  NAND2_X1 U6425 ( .A1(n8966), .A2(n9733), .ZN(n8967) );
  NAND2_X1 U6426 ( .A1(n8953), .A2(n8952), .ZN(n9732) );
  OR2_X1 U6427 ( .A1(n5910), .A2(n5909), .ZN(n5927) );
  OR2_X1 U6428 ( .A1(n10789), .A2(n10788), .ZN(n10791) );
  NAND2_X1 U6429 ( .A1(n10567), .A2(n9775), .ZN(n6084) );
  NOR2_X1 U6430 ( .A1(n5878), .A2(n5877), .ZN(n5894) );
  OR2_X1 U6431 ( .A1(n5846), .A2(n5845), .ZN(n5862) );
  NAND2_X1 U6432 ( .A1(n5651), .A2(n8423), .ZN(n5654) );
  NAND2_X1 U6433 ( .A1(n8662), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5626) );
  NAND2_X1 U6434 ( .A1(n6282), .A2(n8247), .ZN(n6575) );
  INV_X1 U6435 ( .A(n9546), .ZN(n9037) );
  NAND2_X1 U6436 ( .A1(n6420), .A2(n6419), .ZN(n7494) );
  INV_X1 U6437 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n7163) );
  NAND2_X1 U6438 ( .A1(n9381), .A2(n6677), .ZN(n9382) );
  NAND2_X1 U6439 ( .A1(n6286), .A2(n8469), .ZN(n6639) );
  INV_X1 U6440 ( .A(n9194), .ZN(n9437) );
  INV_X1 U6441 ( .A(n9516), .ZN(n9487) );
  NAND2_X1 U6442 ( .A1(n8776), .A2(n8777), .ZN(n9551) );
  AND2_X1 U6443 ( .A1(n8770), .A2(n8769), .ZN(n9585) );
  NAND2_X1 U6444 ( .A1(n6951), .A2(n7148), .ZN(n6683) );
  NAND2_X1 U6445 ( .A1(n9596), .A2(n11017), .ZN(n9597) );
  AND2_X1 U6446 ( .A1(n9376), .A2(n11097), .ZN(n6713) );
  INV_X1 U6447 ( .A(n9197), .ZN(n9561) );
  NAND2_X1 U6448 ( .A1(n7764), .A2(n7763), .ZN(n7875) );
  AND3_X1 U6449 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5792) );
  NAND2_X1 U6450 ( .A1(n8968), .A2(n8967), .ZN(n8969) );
  OR2_X1 U6451 ( .A1(n7039), .A2(n10148), .ZN(n7037) );
  XNOR2_X1 U6452 ( .A(n6173), .B(n10102), .ZN(n10295) );
  INV_X1 U6453 ( .A(n10522), .ZN(n8155) );
  INV_X1 U6454 ( .A(n11027), .ZN(n10900) );
  NAND2_X1 U6455 ( .A1(n10587), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5704) );
  NAND2_X1 U6456 ( .A1(n5677), .A2(n5676), .ZN(n5980) );
  NAND2_X1 U6457 ( .A1(n5654), .A2(n5653), .ZN(n5869) );
  OAI211_X2 U6458 ( .C1(n6313), .C2(n7339), .A(n6324), .B(n6323), .ZN(n8710)
         );
  AND2_X1 U6459 ( .A1(n6612), .A2(n6611), .ZN(n9426) );
  NAND4_X1 U6460 ( .A1(n6356), .A2(n6355), .A3(n6354), .A4(n6353), .ZN(n7171)
         );
  INV_X1 U6461 ( .A(n7780), .ZN(n7686) );
  AND2_X1 U6462 ( .A1(n8800), .A2(n8801), .ZN(n9501) );
  OR2_X1 U6463 ( .A1(n6918), .A2(n7207), .ZN(n10937) );
  NAND2_X1 U6464 ( .A1(n6758), .A2(n8676), .ZN(n10928) );
  INV_X1 U6465 ( .A(n9655), .ZN(n6754) );
  INV_X1 U6466 ( .A(n9866), .ZN(n9871) );
  AND4_X1 U6467 ( .A1(n6047), .A2(n6046), .A3(n6045), .A4(n6044), .ZN(n10425)
         );
  AND4_X1 U6468 ( .A1(n5712), .A2(n5711), .A3(n5710), .A4(n5709), .ZN(n9799)
         );
  AND4_X1 U6469 ( .A1(n5867), .A2(n5866), .A3(n5865), .A4(n5864), .ZN(n7883)
         );
  OR2_X1 U6470 ( .A1(n7090), .A2(n10145), .ZN(n10438) );
  AND2_X1 U6471 ( .A1(n11081), .A2(n10541), .ZN(n8052) );
  AND2_X1 U6472 ( .A1(n11085), .A2(n10541), .ZN(n10557) );
  INV_X1 U6473 ( .A(n10543), .ZN(n11078) );
  OR2_X1 U6474 ( .A1(n7283), .A2(n6247), .ZN(n6252) );
  XNOR2_X1 U6475 ( .A(n5631), .B(n8436), .ZN(n5798) );
  INV_X1 U6476 ( .A(n7661), .ZN(n10988) );
  INV_X1 U6477 ( .A(n9171), .ZN(n9183) );
  NAND2_X1 U6478 ( .A1(n6659), .A2(n6658), .ZN(n9380) );
  INV_X1 U6479 ( .A(n9503), .ZN(n9530) );
  INV_X1 U6480 ( .A(n7962), .ZN(n9199) );
  INV_X1 U6481 ( .A(n10848), .ZN(n9330) );
  OR2_X1 U6482 ( .A1(n6932), .A2(n9583), .ZN(n10939) );
  NAND2_X1 U6483 ( .A1(n6932), .A2(n10937), .ZN(n10944) );
  INV_X1 U6484 ( .A(n10946), .ZN(n9589) );
  INV_X1 U6485 ( .A(n11100), .ZN(n11099) );
  INV_X1 U6486 ( .A(n11104), .ZN(n11101) );
  INV_X1 U6487 ( .A(n10491), .ZN(n10365) );
  INV_X1 U6488 ( .A(n9863), .ZN(n9882) );
  AND4_X1 U6489 ( .A1(n6172), .A2(n6171), .A3(n6170), .A4(n6169), .ZN(n10310)
         );
  AND4_X1 U6490 ( .A1(n6026), .A2(n6025), .A3(n6024), .A4(n6023), .ZN(n10449)
         );
  AND4_X1 U6491 ( .A1(n5960), .A2(n5959), .A3(n5958), .A4(n5957), .ZN(n9798)
         );
  OR2_X1 U6492 ( .A1(n6806), .A2(n6970), .ZN(n10808) );
  INV_X1 U6493 ( .A(n10458), .ZN(n10452) );
  NAND2_X1 U6494 ( .A1(n10299), .A2(n8052), .ZN(n6250) );
  INV_X1 U6495 ( .A(n10283), .ZN(n10547) );
  INV_X1 U6496 ( .A(n10432), .ZN(n10573) );
  INV_X1 U6497 ( .A(n10557), .ZN(n10579) );
  OR2_X1 U6498 ( .A1(n6252), .A2(n7020), .ZN(n11082) );
  INV_X1 U6499 ( .A(n10602), .ZN(n10603) );
  INV_X1 U6500 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n8539) );
  INV_X1 U6501 ( .A(SI_1_), .ZN(n8441) );
  AND2_X1 U6502 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5610) );
  NAND2_X1 U6503 ( .A1(n5618), .A2(n5610), .ZN(n5727) );
  NAND3_X1 U6504 ( .A1(n6772), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n5611) );
  NAND2_X1 U6505 ( .A1(n5727), .A2(n5611), .ZN(n5716) );
  NAND2_X1 U6506 ( .A1(n5715), .A2(n5716), .ZN(n5614) );
  NAND2_X1 U6507 ( .A1(n5612), .A2(SI_1_), .ZN(n5613) );
  NAND2_X1 U6508 ( .A1(n5614), .A2(n5613), .ZN(n5738) );
  MUX2_X1 U6509 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5618), .Z(n5615) );
  INV_X1 U6510 ( .A(SI_2_), .ZN(n8229) );
  XNOR2_X1 U6511 ( .A(n5615), .B(n8229), .ZN(n5737) );
  NAND2_X1 U6512 ( .A1(n5738), .A2(n5737), .ZN(n5617) );
  NAND2_X1 U6513 ( .A1(n5615), .A2(SI_2_), .ZN(n5616) );
  NAND2_X1 U6514 ( .A1(n5617), .A2(n5616), .ZN(n5752) );
  MUX2_X1 U6515 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n5618), .Z(n5619) );
  INV_X1 U6516 ( .A(SI_3_), .ZN(n8218) );
  XNOR2_X1 U6517 ( .A(n5619), .B(n8218), .ZN(n5751) );
  NAND2_X1 U6518 ( .A1(n5752), .A2(n5751), .ZN(n5621) );
  NAND2_X1 U6519 ( .A1(n5619), .A2(SI_3_), .ZN(n5620) );
  NAND2_X1 U6520 ( .A1(n5621), .A2(n5620), .ZN(n5770) );
  INV_X1 U6521 ( .A(SI_4_), .ZN(n5622) );
  XNOR2_X1 U6522 ( .A(n5623), .B(n5622), .ZN(n5769) );
  NAND2_X1 U6523 ( .A1(n5770), .A2(n5769), .ZN(n5625) );
  NAND2_X1 U6524 ( .A1(n5623), .A2(SI_4_), .ZN(n5624) );
  NAND2_X1 U6525 ( .A1(n5625), .A2(n5624), .ZN(n5787) );
  INV_X1 U6526 ( .A(SI_5_), .ZN(n8431) );
  NAND2_X1 U6527 ( .A1(n5787), .A2(n5786), .ZN(n5630) );
  NAND2_X1 U6528 ( .A1(n5628), .A2(SI_5_), .ZN(n5629) );
  NAND2_X1 U6529 ( .A1(n5630), .A2(n5629), .ZN(n5797) );
  MUX2_X1 U6530 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n8662), .Z(n5631) );
  INV_X1 U6531 ( .A(SI_6_), .ZN(n8436) );
  NAND2_X1 U6532 ( .A1(n5797), .A2(n5798), .ZN(n5633) );
  NAND2_X1 U6533 ( .A1(n5631), .A2(SI_6_), .ZN(n5632) );
  NAND2_X1 U6534 ( .A1(n5633), .A2(n5632), .ZN(n5804) );
  MUX2_X1 U6535 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n8662), .Z(n5635) );
  NAND2_X1 U6536 ( .A1(n5804), .A2(n5634), .ZN(n5637) );
  NAND2_X1 U6537 ( .A1(n5635), .A2(SI_7_), .ZN(n5636) );
  NAND2_X1 U6538 ( .A1(n5637), .A2(n5636), .ZN(n5835) );
  INV_X1 U6539 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6793) );
  INV_X1 U6540 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n8322) );
  MUX2_X1 U6541 ( .A(n6793), .B(n8322), .S(n8662), .Z(n5638) );
  INV_X1 U6542 ( .A(SI_8_), .ZN(n8224) );
  INV_X1 U6543 ( .A(n5638), .ZN(n5639) );
  NAND2_X1 U6544 ( .A1(n5639), .A2(SI_8_), .ZN(n5640) );
  INV_X1 U6545 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6798) );
  MUX2_X1 U6546 ( .A(n6798), .B(n8539), .S(n8662), .Z(n5643) );
  INV_X1 U6547 ( .A(n5643), .ZN(n5641) );
  INV_X1 U6548 ( .A(SI_9_), .ZN(n8219) );
  NAND2_X1 U6549 ( .A1(n5643), .A2(n8219), .ZN(n5839) );
  MUX2_X1 U6550 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n8662), .Z(n5648) );
  INV_X1 U6551 ( .A(SI_10_), .ZN(n8427) );
  NAND2_X1 U6552 ( .A1(n5648), .A2(SI_10_), .ZN(n5649) );
  INV_X1 U6553 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6808) );
  INV_X1 U6554 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5650) );
  MUX2_X1 U6555 ( .A(n6808), .B(n5650), .S(n8662), .Z(n5651) );
  INV_X1 U6556 ( .A(SI_11_), .ZN(n8423) );
  INV_X1 U6557 ( .A(n5651), .ZN(n5652) );
  NAND2_X1 U6558 ( .A1(n5652), .A2(SI_11_), .ZN(n5653) );
  MUX2_X1 U6559 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n8662), .Z(n5655) );
  INV_X1 U6560 ( .A(SI_12_), .ZN(n8415) );
  MUX2_X1 U6561 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n8662), .Z(n5657) );
  NAND2_X1 U6562 ( .A1(n5657), .A2(SI_13_), .ZN(n5658) );
  INV_X1 U6563 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6866) );
  INV_X1 U6564 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n8529) );
  MUX2_X1 U6565 ( .A(n6866), .B(n8529), .S(n8662), .Z(n5660) );
  INV_X1 U6566 ( .A(SI_14_), .ZN(n8422) );
  INV_X1 U6567 ( .A(n5660), .ZN(n5661) );
  NAND2_X1 U6568 ( .A1(n5661), .A2(SI_14_), .ZN(n5662) );
  NAND2_X1 U6569 ( .A1(n5665), .A2(n5662), .ZN(n5918) );
  MUX2_X1 U6570 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n8662), .Z(n5666) );
  INV_X1 U6571 ( .A(SI_15_), .ZN(n8418) );
  XNOR2_X1 U6572 ( .A(n5666), .B(n8418), .ZN(n5935) );
  INV_X1 U6573 ( .A(n5935), .ZN(n5668) );
  NAND2_X1 U6574 ( .A1(n5666), .A2(SI_15_), .ZN(n5667) );
  INV_X1 U6575 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7072) );
  INV_X1 U6576 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n8525) );
  MUX2_X1 U6577 ( .A(n7072), .B(n8525), .S(n8662), .Z(n5669) );
  INV_X1 U6578 ( .A(SI_16_), .ZN(n8206) );
  INV_X1 U6579 ( .A(n5669), .ZN(n5670) );
  NAND2_X1 U6580 ( .A1(n5670), .A2(SI_16_), .ZN(n5671) );
  NAND2_X1 U6581 ( .A1(n5672), .A2(n5671), .ZN(n5948) );
  INV_X1 U6582 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7086) );
  INV_X1 U6583 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n8309) );
  MUX2_X1 U6584 ( .A(n7086), .B(n8309), .S(n8662), .Z(n5673) );
  INV_X1 U6585 ( .A(SI_17_), .ZN(n8198) );
  NAND2_X1 U6586 ( .A1(n5673), .A2(n8198), .ZN(n5676) );
  INV_X1 U6587 ( .A(n5673), .ZN(n5674) );
  NAND2_X1 U6588 ( .A1(n5674), .A2(SI_17_), .ZN(n5675) );
  MUX2_X1 U6589 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n8662), .Z(n5977) );
  INV_X1 U6590 ( .A(SI_18_), .ZN(n5678) );
  XNOR2_X1 U6591 ( .A(n5977), .B(n5678), .ZN(n5976) );
  XNOR2_X1 U6592 ( .A(n5980), .B(n5976), .ZN(n7137) );
  NOR2_X1 U6593 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5683) );
  NOR2_X1 U6594 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n5688) );
  NOR2_X1 U6595 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5687) );
  NOR2_X1 U6596 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5686) );
  NOR2_X1 U6597 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n5685) );
  NAND4_X1 U6598 ( .A1(n5688), .A2(n5687), .A3(n5686), .A4(n5685), .ZN(n5690)
         );
  NOR2_X1 U6599 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5689) );
  INV_X1 U6600 ( .A(n6215), .ZN(n6223) );
  NOR2_X1 U6601 ( .A1(n5690), .A2(n6223), .ZN(n5691) );
  INV_X1 U6602 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5693) );
  NAND2_X1 U6603 ( .A1(n6219), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5695) );
  INV_X1 U6604 ( .A(n5799), .ZN(n5806) );
  NAND2_X1 U6605 ( .A1(n7137), .A2(n9893), .ZN(n5701) );
  INV_X2 U6606 ( .A(n9895), .ZN(n5988) );
  INV_X1 U6607 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6175) );
  NAND2_X1 U6608 ( .A1(n5963), .A2(n6175), .ZN(n5699) );
  NAND2_X1 U6609 ( .A1(n5699), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5984) );
  XNOR2_X1 U6610 ( .A(n5984), .B(P1_IR_REG_18__SCAN_IN), .ZN(n10271) );
  AOI22_X1 U6611 ( .A1(n5988), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5987), .B2(
        n10271), .ZN(n5700) );
  NAND2_X1 U6612 ( .A1(n5792), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5814) );
  NAND2_X1 U6613 ( .A1(n5827), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5846) );
  INV_X1 U6614 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5845) );
  INV_X1 U6615 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5861) );
  INV_X1 U6616 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5877) );
  NAND2_X1 U6617 ( .A1(n5894), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5910) );
  INV_X1 U6618 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5909) );
  INV_X1 U6619 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5926) );
  NAND2_X1 U6620 ( .A1(n5941), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5954) );
  INV_X1 U6621 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n7830) );
  NAND2_X1 U6622 ( .A1(n5970), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5969) );
  INV_X1 U6623 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5703) );
  INV_X1 U6624 ( .A(n5969), .ZN(n5702) );
  AOI21_X1 U6625 ( .B1(n5969), .B2(n5703), .A(n5992), .ZN(n8146) );
  INV_X1 U6626 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n8369) );
  INV_X1 U6627 ( .A(n5707), .ZN(n5706) );
  INV_X1 U6628 ( .A(n5791), .ZN(n5972) );
  NAND2_X1 U6629 ( .A1(n8146), .A2(n5972), .ZN(n5712) );
  INV_X1 U6630 ( .A(n6079), .ZN(n6205) );
  NAND2_X1 U6631 ( .A1(n6205), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5711) );
  NAND2_X1 U6632 ( .A1(n9885), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5710) );
  NAND2_X1 U6633 ( .A1(n5825), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5709) );
  INV_X1 U6634 ( .A(n9799), .ZN(n10158) );
  INV_X1 U6635 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n10178) );
  OR2_X1 U6636 ( .A1(n5791), .A2(n10178), .ZN(n5714) );
  INV_X1 U6637 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7324) );
  INV_X1 U6638 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5713) );
  XNOR2_X1 U6639 ( .A(n5715), .B(n5716), .ZN(n6777) );
  INV_X1 U6640 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6776) );
  INV_X1 U6641 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5718) );
  NAND2_X1 U6642 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5717) );
  XNOR2_X1 U6643 ( .A(n5718), .B(n5717), .ZN(n6990) );
  OR2_X1 U6644 ( .A1(n6803), .A2(n6990), .ZN(n5719) );
  NAND2_X1 U6645 ( .A1(n5825), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5724) );
  INV_X1 U6646 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n7031) );
  OR2_X1 U6647 ( .A1(n5776), .A2(n7031), .ZN(n5723) );
  INV_X1 U6648 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n5720) );
  OR2_X1 U6649 ( .A1(n5791), .A2(n5720), .ZN(n5722) );
  INV_X1 U6650 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10662) );
  OR2_X1 U6651 ( .A1(n6079), .A2(n10662), .ZN(n5721) );
  NAND2_X1 U6652 ( .A1(n8662), .A2(SI_0_), .ZN(n5726) );
  INV_X1 U6653 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5725) );
  NAND2_X1 U6654 ( .A1(n5726), .A2(n5725), .ZN(n5728) );
  AND2_X1 U6655 ( .A1(n5728), .A2(n5727), .ZN(n10599) );
  MUX2_X1 U6656 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10599), .S(n6803), .Z(n7382)
         );
  NAND2_X1 U6657 ( .A1(n9906), .A2(n7382), .ZN(n7317) );
  NAND2_X1 U6658 ( .A1(n6184), .A2(n7317), .ZN(n5731) );
  INV_X1 U6659 ( .A(n10171), .ZN(n6185) );
  NAND2_X1 U6660 ( .A1(n6185), .A2(n5729), .ZN(n5730) );
  NAND2_X1 U6661 ( .A1(n5731), .A2(n5730), .ZN(n7279) );
  NAND2_X1 U6662 ( .A1(n9885), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5736) );
  INV_X1 U6663 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10191) );
  OR2_X1 U6664 ( .A1(n5791), .A2(n10191), .ZN(n5735) );
  INV_X1 U6665 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7290) );
  OR2_X1 U6666 ( .A1(n6079), .A2(n7290), .ZN(n5734) );
  INV_X1 U6667 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5732) );
  INV_X1 U6668 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6774) );
  OR2_X1 U6669 ( .A1(n9895), .A2(n6774), .ZN(n5743) );
  XNOR2_X1 U6670 ( .A(n5738), .B(n5737), .ZN(n6775) );
  OR2_X1 U6671 ( .A1(n5799), .A2(n6775), .ZN(n5742) );
  OR2_X1 U6672 ( .A1(n5739), .A2(n5905), .ZN(n5753) );
  INV_X1 U6673 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5740) );
  XNOR2_X1 U6674 ( .A(n5753), .B(n5740), .ZN(n6989) );
  OR2_X1 U6675 ( .A1(n6803), .A2(n6989), .ZN(n5741) );
  OR2_X2 U6676 ( .A1(n10170), .A2(n10884), .ZN(n10904) );
  NAND2_X1 U6677 ( .A1(n10170), .A2(n10884), .ZN(n9948) );
  NAND2_X1 U6678 ( .A1(n10904), .A2(n9948), .ZN(n10065) );
  NAND2_X1 U6679 ( .A1(n7279), .A2(n10065), .ZN(n5745) );
  OR2_X1 U6680 ( .A1(n10170), .A2(n9848), .ZN(n5744) );
  NAND2_X1 U6681 ( .A1(n5745), .A2(n5744), .ZN(n10896) );
  NAND2_X1 U6682 ( .A1(n9885), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5750) );
  OR2_X1 U6683 ( .A1(n5791), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5749) );
  INV_X1 U6684 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10914) );
  OR2_X1 U6685 ( .A1(n6079), .A2(n10914), .ZN(n5748) );
  INV_X1 U6686 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5746) );
  OR2_X1 U6687 ( .A1(n9889), .A2(n5746), .ZN(n5747) );
  NAND4_X1 U6688 ( .A1(n5750), .A2(n5749), .A3(n5748), .A4(n5747), .ZN(n10169)
         );
  XNOR2_X1 U6689 ( .A(n5752), .B(n5751), .ZN(n6780) );
  OR2_X1 U6690 ( .A1(n5799), .A2(n6780), .ZN(n5758) );
  INV_X1 U6691 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6778) );
  OR2_X1 U6692 ( .A1(n9895), .A2(n6778), .ZN(n5757) );
  NAND2_X1 U6693 ( .A1(n5753), .A2(n5740), .ZN(n5754) );
  NAND2_X1 U6694 ( .A1(n5754), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5755) );
  INV_X1 U6695 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n8332) );
  XNOR2_X1 U6696 ( .A(n5755), .B(n8332), .ZN(n6993) );
  OR2_X1 U6697 ( .A1(n6803), .A2(n6993), .ZN(n5756) );
  NAND2_X1 U6698 ( .A1(n10169), .A2(n10899), .ZN(n9947) );
  NAND2_X1 U6699 ( .A1(n10896), .A2(n10903), .ZN(n5761) );
  INV_X1 U6700 ( .A(n10169), .ZN(n5759) );
  NAND2_X1 U6701 ( .A1(n5759), .A2(n10899), .ZN(n5760) );
  NAND2_X1 U6702 ( .A1(n9885), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5765) );
  INV_X1 U6703 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5762) );
  OR2_X1 U6704 ( .A1(n9889), .A2(n5762), .ZN(n5764) );
  XNOR2_X1 U6705 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n9821) );
  OR2_X1 U6706 ( .A1(n6167), .A2(n9821), .ZN(n5763) );
  INV_X1 U6707 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6977) );
  NAND2_X1 U6708 ( .A1(n5739), .A2(n5766), .ZN(n5767) );
  NAND2_X1 U6709 ( .A1(n5767), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5768) );
  XNOR2_X1 U6710 ( .A(n5768), .B(n5679), .ZN(n10217) );
  OR2_X1 U6711 ( .A1(n9895), .A2(n5411), .ZN(n5772) );
  XNOR2_X1 U6712 ( .A(n5770), .B(n5769), .ZN(n6773) );
  OR2_X1 U6713 ( .A1(n5799), .A2(n6773), .ZN(n5771) );
  OAI211_X1 U6714 ( .C1(n6803), .C2(n10217), .A(n5772), .B(n5771), .ZN(n9820)
         );
  NOR2_X1 U6715 ( .A1(n9745), .A2(n9820), .ZN(n5774) );
  NAND2_X1 U6716 ( .A1(n9745), .A2(n9820), .ZN(n5773) );
  AOI21_X1 U6717 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5775) );
  NOR2_X1 U6718 ( .A1(n5775), .A2(n5792), .ZN(n7483) );
  NAND2_X1 U6719 ( .A1(n5972), .A2(n7483), .ZN(n5781) );
  INV_X1 U6720 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6997) );
  INV_X1 U6721 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5777) );
  OR2_X1 U6722 ( .A1(n9889), .A2(n5777), .ZN(n5779) );
  INV_X1 U6723 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6979) );
  OR2_X1 U6724 ( .A1(n6079), .A2(n6979), .ZN(n5778) );
  NAND2_X1 U6725 ( .A1(n5783), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5782) );
  MUX2_X1 U6726 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5782), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5785) );
  NOR2_X1 U6727 ( .A1(n5783), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5808) );
  INV_X1 U6728 ( .A(n5808), .ZN(n5784) );
  AOI22_X1 U6729 ( .A1(n5988), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n5987), .B2(
        n10242), .ZN(n5789) );
  XNOR2_X1 U6730 ( .A(n5787), .B(n5786), .ZN(n6783) );
  OR2_X1 U6731 ( .A1(n6783), .A2(n5799), .ZN(n5788) );
  OR2_X1 U6732 ( .A1(n10168), .A2(n10969), .ZN(n9912) );
  NAND2_X1 U6733 ( .A1(n10168), .A2(n10969), .ZN(n9955) );
  NAND2_X1 U6734 ( .A1(n9912), .A2(n9955), .ZN(n10072) );
  INV_X1 U6735 ( .A(n10072), .ZN(n9957) );
  INV_X1 U6736 ( .A(n10168), .ZN(n7220) );
  NAND2_X1 U6737 ( .A1(n7220), .A2(n10969), .ZN(n5790) );
  NAND2_X1 U6738 ( .A1(n5825), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5796) );
  INV_X1 U6739 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6999) );
  OR2_X1 U6740 ( .A1(n6209), .A2(n6999), .ZN(n5795) );
  OAI21_X1 U6741 ( .B1(n5792), .B2(P1_REG3_REG_6__SCAN_IN), .A(n5814), .ZN(
        n7599) );
  OR2_X1 U6742 ( .A1(n6167), .A2(n7599), .ZN(n5794) );
  INV_X1 U6743 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6981) );
  OR2_X1 U6744 ( .A1(n9887), .A2(n6981), .ZN(n5793) );
  XNOR2_X1 U6745 ( .A(n5797), .B(n5798), .ZN(n6785) );
  OR2_X1 U6746 ( .A1(n6785), .A2(n5799), .ZN(n5802) );
  OR2_X1 U6747 ( .A1(n5808), .A2(n5905), .ZN(n5800) );
  XNOR2_X1 U6748 ( .A(n5800), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10253) );
  AOI22_X1 U6749 ( .A1(n5988), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5987), .B2(
        n10253), .ZN(n5801) );
  NAND2_X1 U6750 ( .A1(n5802), .A2(n5801), .ZN(n7747) );
  NAND2_X1 U6751 ( .A1(n7443), .A2(n7747), .ZN(n10070) );
  INV_X1 U6752 ( .A(n7747), .ZN(n7603) );
  INV_X1 U6753 ( .A(n7443), .ZN(n10167) );
  NAND2_X1 U6754 ( .A1(n7603), .A2(n10167), .ZN(n9962) );
  NAND2_X1 U6755 ( .A1(n10070), .A2(n9962), .ZN(n9964) );
  NAND2_X1 U6756 ( .A1(n7443), .A2(n7603), .ZN(n5803) );
  NAND2_X1 U6757 ( .A1(n7215), .A2(n5803), .ZN(n7300) );
  XNOR2_X1 U6758 ( .A(n5804), .B(n5805), .ZN(n6786) );
  NAND2_X1 U6759 ( .A1(n6786), .A2(n5806), .ZN(n5811) );
  INV_X1 U6760 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5807) );
  NAND2_X1 U6761 ( .A1(n5808), .A2(n5807), .ZN(n5821) );
  NAND2_X1 U6762 ( .A1(n5821), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5809) );
  XNOR2_X1 U6763 ( .A(n5809), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10678) );
  AOI22_X1 U6764 ( .A1(n5988), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5987), .B2(
        n10678), .ZN(n5810) );
  NAND2_X1 U6765 ( .A1(n5811), .A2(n5810), .ZN(n7433) );
  NAND2_X1 U6766 ( .A1(n5825), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5819) );
  INV_X1 U6767 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5812) );
  OR2_X1 U6768 ( .A1(n6209), .A2(n5812), .ZN(n5818) );
  AND2_X1 U6769 ( .A1(n5814), .A2(n5813), .ZN(n5815) );
  OR2_X1 U6770 ( .A1(n5815), .A2(n5827), .ZN(n7442) );
  OR2_X1 U6771 ( .A1(n6167), .A2(n7442), .ZN(n5817) );
  INV_X1 U6772 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7310) );
  OR2_X1 U6773 ( .A1(n9887), .A2(n7310), .ZN(n5816) );
  OR2_X1 U6774 ( .A1(n7433), .A2(n7539), .ZN(n9967) );
  NAND2_X1 U6775 ( .A1(n7433), .A2(n7539), .ZN(n9966) );
  NAND2_X1 U6776 ( .A1(n9967), .A2(n9966), .ZN(n9961) );
  INV_X1 U6777 ( .A(n7539), .ZN(n10166) );
  OR2_X1 U6778 ( .A1(n7433), .A2(n10166), .ZN(n5820) );
  XNOR2_X1 U6779 ( .A(n5835), .B(n5834), .ZN(n6790) );
  NAND2_X1 U6780 ( .A1(n6790), .A2(n5806), .ZN(n5824) );
  NAND2_X1 U6781 ( .A1(n5842), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5822) );
  XNOR2_X1 U6782 ( .A(n5822), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10692) );
  AOI22_X1 U6783 ( .A1(n5988), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5987), .B2(
        n10692), .ZN(n5823) );
  NAND2_X1 U6784 ( .A1(n5824), .A2(n5823), .ZN(n7549) );
  NAND2_X1 U6785 ( .A1(n5825), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5833) );
  INV_X1 U6786 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n5826) );
  OR2_X1 U6787 ( .A1(n6209), .A2(n5826), .ZN(n5832) );
  OR2_X1 U6788 ( .A1(n5827), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5828) );
  NAND2_X1 U6789 ( .A1(n5846), .A2(n5828), .ZN(n7529) );
  OR2_X1 U6790 ( .A1(n6167), .A2(n7529), .ZN(n5831) );
  INV_X1 U6791 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n5829) );
  OR2_X1 U6792 ( .A1(n9887), .A2(n5829), .ZN(n5830) );
  XNOR2_X1 U6793 ( .A(n7549), .B(n7627), .ZN(n9968) );
  INV_X1 U6794 ( .A(n7627), .ZN(n10165) );
  OR2_X1 U6795 ( .A1(n5835), .A2(n5834), .ZN(n5837) );
  NAND2_X1 U6796 ( .A1(n5837), .A2(n5836), .ZN(n5841) );
  AND2_X1 U6797 ( .A1(n5839), .A2(n5838), .ZN(n5840) );
  NAND2_X1 U6798 ( .A1(n6796), .A2(n5806), .ZN(n5844) );
  NAND2_X1 U6799 ( .A1(n5889), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5856) );
  XNOR2_X1 U6800 ( .A(n5856), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10798) );
  AOI22_X1 U6801 ( .A1(n5988), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5987), .B2(
        n10798), .ZN(n5843) );
  NAND2_X2 U6802 ( .A1(n5844), .A2(n5843), .ZN(n10457) );
  NAND2_X1 U6803 ( .A1(n5825), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5852) );
  INV_X1 U6804 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7003) );
  OR2_X1 U6805 ( .A1(n6209), .A2(n7003), .ZN(n5851) );
  NAND2_X1 U6806 ( .A1(n5846), .A2(n5845), .ZN(n5847) );
  NAND2_X1 U6807 ( .A1(n5862), .A2(n5847), .ZN(n10455) );
  OR2_X1 U6808 ( .A1(n6167), .A2(n10455), .ZN(n5850) );
  INV_X1 U6809 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n5848) );
  OR2_X1 U6810 ( .A1(n9887), .A2(n5848), .ZN(n5849) );
  OR2_X1 U6811 ( .A1(n10457), .A2(n7770), .ZN(n9977) );
  NAND2_X1 U6812 ( .A1(n10457), .A2(n7770), .ZN(n10075) );
  NAND2_X1 U6813 ( .A1(n9977), .A2(n10075), .ZN(n7425) );
  NAND2_X1 U6814 ( .A1(n7418), .A2(n7425), .ZN(n7417) );
  INV_X1 U6815 ( .A(n7770), .ZN(n10164) );
  OR2_X1 U6816 ( .A1(n10457), .A2(n10164), .ZN(n5853) );
  NAND2_X1 U6817 ( .A1(n7417), .A2(n5853), .ZN(n7450) );
  XNOR2_X1 U6818 ( .A(n5855), .B(n5854), .ZN(n6794) );
  NAND2_X1 U6819 ( .A1(n6794), .A2(n9893), .ZN(n5859) );
  INV_X1 U6820 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8342) );
  NAND2_X1 U6821 ( .A1(n5856), .A2(n8342), .ZN(n5857) );
  NAND2_X1 U6822 ( .A1(n5857), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5871) );
  XNOR2_X1 U6823 ( .A(n5871), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10774) );
  AOI22_X1 U6824 ( .A1(n5988), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5987), .B2(
        n10774), .ZN(n5858) );
  NAND2_X1 U6825 ( .A1(n9885), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5867) );
  INV_X1 U6826 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5860) );
  OR2_X1 U6827 ( .A1(n9889), .A2(n5860), .ZN(n5866) );
  NAND2_X1 U6828 ( .A1(n5862), .A2(n5861), .ZN(n5863) );
  NAND2_X1 U6829 ( .A1(n5878), .A2(n5863), .ZN(n7769) );
  OR2_X1 U6830 ( .A1(n6167), .A2(n7769), .ZN(n5865) );
  INV_X1 U6831 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7588) );
  OR2_X1 U6832 ( .A1(n9887), .A2(n7588), .ZN(n5864) );
  OR2_X1 U6833 ( .A1(n7773), .A2(n7883), .ZN(n9975) );
  NAND2_X1 U6834 ( .A1(n7773), .A2(n7883), .ZN(n11021) );
  NAND2_X1 U6835 ( .A1(n9975), .A2(n11021), .ZN(n10079) );
  INV_X1 U6836 ( .A(n7883), .ZN(n11028) );
  OR2_X1 U6837 ( .A1(n7773), .A2(n11028), .ZN(n5868) );
  XNOR2_X1 U6838 ( .A(n5870), .B(n5869), .ZN(n6801) );
  NAND2_X1 U6839 ( .A1(n6801), .A2(n9893), .ZN(n5875) );
  INV_X1 U6840 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n8558) );
  NAND2_X1 U6841 ( .A1(n5871), .A2(n8558), .ZN(n5872) );
  NAND2_X1 U6842 ( .A1(n5872), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5873) );
  XNOR2_X1 U6843 ( .A(n5873), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10709) );
  AOI22_X1 U6844 ( .A1(n5988), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5987), .B2(
        n10709), .ZN(n5874) );
  NAND2_X1 U6845 ( .A1(n5875), .A2(n5874), .ZN(n11055) );
  NAND2_X1 U6846 ( .A1(n5825), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5883) );
  INV_X1 U6847 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7006) );
  OR2_X1 U6848 ( .A1(n6209), .A2(n7006), .ZN(n5882) );
  INV_X1 U6849 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n5876) );
  OR2_X1 U6850 ( .A1(n9887), .A2(n5876), .ZN(n5881) );
  AND2_X1 U6851 ( .A1(n5878), .A2(n5877), .ZN(n5879) );
  OR2_X1 U6852 ( .A1(n5879), .A2(n5894), .ZN(n11049) );
  OR2_X1 U6853 ( .A1(n6167), .A2(n11049), .ZN(n5880) );
  NAND4_X1 U6854 ( .A1(n5883), .A2(n5882), .A3(n5881), .A4(n5880), .ZN(n10163)
         );
  NAND2_X1 U6855 ( .A1(n11055), .A2(n10163), .ZN(n5884) );
  OR2_X1 U6856 ( .A1(n11055), .A2(n10163), .ZN(n5885) );
  XNOR2_X1 U6857 ( .A(n5887), .B(n5886), .ZN(n6834) );
  NAND2_X1 U6858 ( .A1(n6834), .A2(n9893), .ZN(n5892) );
  INV_X1 U6859 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n8559) );
  NAND3_X1 U6860 ( .A1(n8559), .A2(n8342), .A3(n8558), .ZN(n5888) );
  OAI21_X1 U6861 ( .B1(n5889), .B2(n5888), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5890) );
  XNOR2_X1 U6862 ( .A(n5890), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7835) );
  AOI22_X1 U6863 ( .A1(n5988), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5987), .B2(
        n7835), .ZN(n5891) );
  NAND2_X1 U6864 ( .A1(n5825), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5899) );
  INV_X1 U6865 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n5893) );
  OR2_X1 U6866 ( .A1(n6209), .A2(n5893), .ZN(n5898) );
  OR2_X1 U6867 ( .A1(n5894), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5895) );
  NAND2_X1 U6868 ( .A1(n5910), .A2(n5895), .ZN(n7982) );
  OR2_X1 U6869 ( .A1(n6167), .A2(n7982), .ZN(n5897) );
  INV_X1 U6870 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7643) );
  OR2_X1 U6871 ( .A1(n9887), .A2(n7643), .ZN(n5896) );
  NAND4_X1 U6872 ( .A1(n5899), .A2(n5898), .A3(n5897), .A4(n5896), .ZN(n11025)
         );
  NOR2_X1 U6873 ( .A1(n7973), .A2(n11025), .ZN(n5900) );
  NAND2_X1 U6874 ( .A1(n7973), .A2(n11025), .ZN(n5901) );
  NAND2_X1 U6875 ( .A1(n5902), .A2(n5901), .ZN(n7669) );
  XNOR2_X1 U6876 ( .A(n5904), .B(n5903), .ZN(n6838) );
  NAND2_X1 U6877 ( .A1(n6838), .A2(n9893), .ZN(n5908) );
  OR2_X1 U6878 ( .A1(n5123), .A2(n5905), .ZN(n5906) );
  XNOR2_X1 U6879 ( .A(n5906), .B(P1_IR_REG_13__SCAN_IN), .ZN(n10767) );
  AOI22_X1 U6880 ( .A1(n5988), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5987), .B2(
        n10767), .ZN(n5907) );
  NAND2_X1 U6881 ( .A1(n5825), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5915) );
  INV_X1 U6882 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7823) );
  OR2_X1 U6883 ( .A1(n6209), .A2(n7823), .ZN(n5914) );
  NAND2_X1 U6884 ( .A1(n5910), .A2(n5909), .ZN(n5911) );
  NAND2_X1 U6885 ( .A1(n5927), .A2(n5911), .ZN(n8035) );
  OR2_X1 U6886 ( .A1(n6167), .A2(n8035), .ZN(n5913) );
  INV_X1 U6887 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7677) );
  OR2_X1 U6888 ( .A1(n9887), .A2(n7677), .ZN(n5912) );
  NAND4_X1 U6889 ( .A1(n5915), .A2(n5914), .A3(n5913), .A4(n5912), .ZN(n10162)
         );
  AND2_X1 U6890 ( .A1(n8029), .A2(n10162), .ZN(n5917) );
  OR2_X1 U6891 ( .A1(n8029), .A2(n10162), .ZN(n5916) );
  OAI21_X2 U6892 ( .B1(n7669), .B2(n5917), .A(n5916), .ZN(n7911) );
  NAND2_X1 U6893 ( .A1(n5919), .A2(n5918), .ZN(n5920) );
  NAND2_X1 U6894 ( .A1(n5921), .A2(n5920), .ZN(n6863) );
  NAND2_X1 U6895 ( .A1(n6863), .A2(n9893), .ZN(n5925) );
  NAND2_X1 U6896 ( .A1(n5922), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5923) );
  XNOR2_X1 U6897 ( .A(n5923), .B(P1_IR_REG_14__SCAN_IN), .ZN(n10726) );
  AOI22_X1 U6898 ( .A1(n5988), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5987), .B2(
        n10726), .ZN(n5924) );
  NAND2_X1 U6899 ( .A1(n5825), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5932) );
  INV_X1 U6900 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n8054) );
  OR2_X1 U6901 ( .A1(n6209), .A2(n8054), .ZN(n5931) );
  INV_X1 U6902 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7919) );
  OR2_X1 U6903 ( .A1(n6079), .A2(n7919), .ZN(n5930) );
  AND2_X1 U6904 ( .A1(n5927), .A2(n5926), .ZN(n5928) );
  OR2_X1 U6905 ( .A1(n5928), .A2(n5941), .ZN(n8124) );
  OR2_X1 U6906 ( .A1(n6167), .A2(n8124), .ZN(n5929) );
  NAND4_X1 U6907 ( .A1(n5932), .A2(n5931), .A3(n5930), .A4(n5929), .ZN(n10161)
         );
  NOR2_X1 U6908 ( .A1(n8128), .A2(n10161), .ZN(n5933) );
  NAND2_X1 U6909 ( .A1(n8128), .A2(n10161), .ZN(n5934) );
  XNOR2_X1 U6910 ( .A(n5936), .B(n5935), .ZN(n6942) );
  NAND2_X1 U6911 ( .A1(n6942), .A2(n9893), .ZN(n5940) );
  NAND2_X1 U6912 ( .A1(n5267), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5938) );
  XNOR2_X1 U6913 ( .A(n5938), .B(n5698), .ZN(n7837) );
  INV_X1 U6914 ( .A(n7837), .ZN(n10741) );
  AOI22_X1 U6915 ( .A1(n5988), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5987), .B2(
        n10741), .ZN(n5939) );
  NAND2_X1 U6916 ( .A1(n5825), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5947) );
  INV_X1 U6917 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10735) );
  OR2_X1 U6918 ( .A1(n6209), .A2(n10735), .ZN(n5946) );
  OR2_X1 U6919 ( .A1(n5941), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5942) );
  NAND2_X1 U6920 ( .A1(n5942), .A2(n5954), .ZN(n8175) );
  OR2_X1 U6921 ( .A1(n6167), .A2(n8175), .ZN(n5945) );
  INV_X1 U6922 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n5943) );
  OR2_X1 U6923 ( .A1(n9887), .A2(n5943), .ZN(n5944) );
  NAND2_X1 U6924 ( .A1(n10540), .A2(n9787), .ZN(n10005) );
  INV_X1 U6925 ( .A(n9787), .ZN(n10160) );
  XNOR2_X1 U6926 ( .A(n5949), .B(n5948), .ZN(n7071) );
  NAND2_X1 U6927 ( .A1(n7071), .A2(n9893), .ZN(n5953) );
  NAND2_X1 U6928 ( .A1(n5950), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5951) );
  XNOR2_X1 U6929 ( .A(n5951), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7866) );
  AOI22_X1 U6930 ( .A1(n5988), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5987), .B2(
        n7866), .ZN(n5952) );
  NAND2_X1 U6931 ( .A1(n5825), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5960) );
  INV_X1 U6932 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n8097) );
  OR2_X1 U6933 ( .A1(n6209), .A2(n8097), .ZN(n5959) );
  INV_X1 U6934 ( .A(n5954), .ZN(n5956) );
  INV_X1 U6935 ( .A(n5970), .ZN(n5955) );
  OAI21_X1 U6936 ( .B1(P1_REG3_REG_16__SCAN_IN), .B2(n5956), .A(n5955), .ZN(
        n9784) );
  OR2_X1 U6937 ( .A1(n5791), .A2(n9784), .ZN(n5958) );
  INV_X1 U6938 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7995) );
  OR2_X1 U6939 ( .A1(n9887), .A2(n7995), .ZN(n5957) );
  OR2_X1 U6940 ( .A1(n9789), .A2(n9798), .ZN(n10004) );
  NAND2_X1 U6941 ( .A1(n9789), .A2(n9798), .ZN(n10006) );
  INV_X1 U6942 ( .A(n9789), .ZN(n8102) );
  XNOR2_X1 U6943 ( .A(n5961), .B(n5962), .ZN(n7084) );
  NAND2_X1 U6944 ( .A1(n7084), .A2(n9893), .ZN(n5965) );
  XNOR2_X1 U6945 ( .A(n5963), .B(P1_IR_REG_17__SCAN_IN), .ZN(n7867) );
  AOI22_X1 U6946 ( .A1(n5988), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5987), .B2(
        n7867), .ZN(n5964) );
  INV_X1 U6947 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10268) );
  NAND2_X1 U6948 ( .A1(n5825), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5967) );
  INV_X1 U6949 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n10258) );
  OR2_X1 U6950 ( .A1(n6079), .A2(n10258), .ZN(n5966) );
  OAI211_X1 U6951 ( .C1(n10268), .C2(n6209), .A(n5967), .B(n5966), .ZN(n5968)
         );
  INV_X1 U6952 ( .A(n5968), .ZN(n5974) );
  OAI21_X1 U6953 ( .B1(n5970), .B2(P1_REG3_REG_17__SCAN_IN), .A(n5969), .ZN(
        n5971) );
  INV_X1 U6954 ( .A(n5971), .ZN(n9802) );
  NAND2_X1 U6955 ( .A1(n9802), .A2(n5972), .ZN(n5973) );
  AND2_X1 U6956 ( .A1(n5974), .A2(n5973), .ZN(n9860) );
  OR2_X1 U6957 ( .A1(n10535), .A2(n9860), .ZN(n8137) );
  NAND2_X1 U6958 ( .A1(n10535), .A2(n9860), .ZN(n8136) );
  NAND2_X1 U6959 ( .A1(n8137), .A2(n8136), .ZN(n10012) );
  INV_X1 U6960 ( .A(n9860), .ZN(n10159) );
  AOI21_X2 U6961 ( .B1(n8086), .B2(n10012), .A(n5975), .ZN(n8145) );
  NAND2_X1 U6962 ( .A1(n9864), .A2(n9799), .ZN(n10017) );
  NAND2_X1 U6963 ( .A1(n10024), .A2(n10017), .ZN(n8144) );
  INV_X1 U6964 ( .A(n5976), .ZN(n5979) );
  NAND2_X1 U6965 ( .A1(n5977), .A2(SI_18_), .ZN(n5978) );
  INV_X1 U6966 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7409) );
  INV_X1 U6967 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8304) );
  MUX2_X1 U6968 ( .A(n7409), .B(n8304), .S(n8662), .Z(n5981) );
  INV_X1 U6969 ( .A(SI_19_), .ZN(n8407) );
  NAND2_X1 U6970 ( .A1(n5981), .A2(n8407), .ZN(n6014) );
  INV_X1 U6971 ( .A(n5981), .ZN(n5982) );
  NAND2_X1 U6972 ( .A1(n5982), .A2(SI_19_), .ZN(n5983) );
  NAND2_X1 U6973 ( .A1(n6014), .A2(n5983), .ZN(n5998) );
  XNOR2_X1 U6974 ( .A(n5999), .B(n5998), .ZN(n7407) );
  NAND2_X1 U6975 ( .A1(n7407), .A2(n9893), .ZN(n5990) );
  INV_X1 U6976 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n8573) );
  NAND2_X1 U6977 ( .A1(n5984), .A2(n8573), .ZN(n5985) );
  NAND2_X1 U6978 ( .A1(n5985), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5986) );
  INV_X1 U6979 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6174) );
  XNOR2_X2 U6980 ( .A(n5986), .B(n6174), .ZN(n10274) );
  INV_X1 U6981 ( .A(n10274), .ZN(n10280) );
  AOI22_X1 U6982 ( .A1(n5988), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10280), 
        .B2(n5987), .ZN(n5989) );
  NAND2_X1 U6983 ( .A1(n5825), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5996) );
  INV_X1 U6984 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n5991) );
  OR2_X1 U6985 ( .A1(n6209), .A2(n5991), .ZN(n5995) );
  NAND2_X1 U6986 ( .A1(n5992), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6007) );
  OAI21_X1 U6987 ( .B1(P1_REG3_REG_19__SCAN_IN), .B2(n5992), .A(n6007), .ZN(
        n9752) );
  OR2_X1 U6988 ( .A1(n6167), .A2(n9752), .ZN(n5994) );
  INV_X1 U6989 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n8156) );
  OR2_X1 U6990 ( .A1(n6079), .A2(n8156), .ZN(n5993) );
  NAND4_X1 U6991 ( .A1(n5996), .A2(n5995), .A3(n5994), .A4(n5993), .ZN(n10157)
         );
  NAND2_X1 U6992 ( .A1(n10522), .A2(n10157), .ZN(n5997) );
  INV_X1 U6993 ( .A(n10157), .ZN(n10448) );
  NAND2_X1 U6994 ( .A1(n6016), .A2(n6014), .ZN(n6003) );
  INV_X1 U6995 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7555) );
  INV_X1 U6996 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7535) );
  MUX2_X1 U6997 ( .A(n7555), .B(n7535), .S(n8662), .Z(n6000) );
  INV_X1 U6998 ( .A(SI_20_), .ZN(n8406) );
  NAND2_X1 U6999 ( .A1(n6000), .A2(n8406), .ZN(n6013) );
  INV_X1 U7000 ( .A(n6000), .ZN(n6001) );
  NAND2_X1 U7001 ( .A1(n6001), .A2(SI_20_), .ZN(n6015) );
  AND2_X1 U7002 ( .A1(n6013), .A2(n6015), .ZN(n6002) );
  NAND2_X1 U7003 ( .A1(n7534), .A2(n9893), .ZN(n6005) );
  OR2_X1 U7004 ( .A1(n9895), .A2(n7535), .ZN(n6004) );
  NAND2_X1 U7005 ( .A1(n5825), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6012) );
  INV_X1 U7006 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n6006) );
  OR2_X1 U7007 ( .A1(n6209), .A2(n6006), .ZN(n6011) );
  NAND2_X1 U7008 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(n6008), .ZN(n6021) );
  OAI21_X1 U7009 ( .B1(P1_REG3_REG_20__SCAN_IN), .B2(n6008), .A(n6021), .ZN(
        n10441) );
  OR2_X1 U7010 ( .A1(n6167), .A2(n10441), .ZN(n6010) );
  INV_X1 U7011 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n10442) );
  OR2_X1 U7012 ( .A1(n9887), .A2(n10442), .ZN(n6009) );
  NAND2_X1 U7013 ( .A1(n10517), .A2(n10426), .ZN(n10026) );
  INV_X1 U7014 ( .A(n10426), .ZN(n10156) );
  MUX2_X1 U7015 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n8662), .Z(n6028) );
  INV_X1 U7016 ( .A(SI_21_), .ZN(n8197) );
  XNOR2_X1 U7017 ( .A(n6028), .B(n8197), .ZN(n6027) );
  XNOR2_X1 U7018 ( .A(n6030), .B(n6027), .ZN(n7595) );
  NAND2_X1 U7019 ( .A1(n7595), .A2(n9893), .ZN(n6018) );
  INV_X1 U7020 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7596) );
  OR2_X1 U7021 ( .A1(n9895), .A2(n7596), .ZN(n6017) );
  NAND2_X1 U7022 ( .A1(n5825), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6026) );
  INV_X1 U7023 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n10513) );
  OR2_X1 U7024 ( .A1(n6209), .A2(n10513), .ZN(n6025) );
  INV_X1 U7025 ( .A(n6021), .ZN(n6019) );
  NAND2_X1 U7026 ( .A1(n6019), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6042) );
  INV_X1 U7027 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n6020) );
  NAND2_X1 U7028 ( .A1(n6021), .A2(n6020), .ZN(n6022) );
  NAND2_X1 U7029 ( .A1(n6042), .A2(n6022), .ZN(n10429) );
  OR2_X1 U7030 ( .A1(n5791), .A2(n10429), .ZN(n6024) );
  INV_X1 U7031 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n10430) );
  OR2_X1 U7032 ( .A1(n6079), .A2(n10430), .ZN(n6023) );
  NAND2_X1 U7033 ( .A1(n10432), .A2(n10449), .ZN(n10033) );
  NAND2_X1 U7034 ( .A1(n10034), .A2(n10033), .ZN(n10428) );
  INV_X1 U7035 ( .A(n6028), .ZN(n6029) );
  INV_X1 U7036 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7668) );
  INV_X1 U7037 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7665) );
  INV_X1 U7038 ( .A(SI_22_), .ZN(n8400) );
  NAND2_X1 U7039 ( .A1(n6031), .A2(n8400), .ZN(n6048) );
  INV_X1 U7040 ( .A(n6031), .ZN(n6032) );
  NAND2_X1 U7041 ( .A1(n6032), .A2(SI_22_), .ZN(n6033) );
  NAND2_X1 U7042 ( .A1(n6048), .A2(n6033), .ZN(n6034) );
  NAND2_X1 U7043 ( .A1(n6035), .A2(n6034), .ZN(n6036) );
  NAND2_X1 U7044 ( .A1(n6049), .A2(n6036), .ZN(n7664) );
  NAND2_X1 U7045 ( .A1(n7664), .A2(n9893), .ZN(n6038) );
  OR2_X1 U7046 ( .A1(n9895), .A2(n7665), .ZN(n6037) );
  NAND2_X1 U7047 ( .A1(n5825), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6047) );
  INV_X1 U7048 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n6039) );
  OR2_X1 U7049 ( .A1(n6209), .A2(n6039), .ZN(n6046) );
  INV_X1 U7050 ( .A(n6042), .ZN(n6040) );
  NAND2_X1 U7051 ( .A1(n6040), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6062) );
  INV_X1 U7052 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n6041) );
  NAND2_X1 U7053 ( .A1(n6042), .A2(n6041), .ZN(n6043) );
  NAND2_X1 U7054 ( .A1(n6062), .A2(n6043), .ZN(n10410) );
  OR2_X1 U7055 ( .A1(n6167), .A2(n10410), .ZN(n6045) );
  INV_X1 U7056 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n10411) );
  OR2_X1 U7057 ( .A1(n9887), .A2(n10411), .ZN(n6044) );
  NAND2_X1 U7058 ( .A1(n10507), .A2(n10425), .ZN(n10124) );
  INV_X1 U7059 ( .A(n10425), .ZN(n10399) );
  INV_X1 U7060 ( .A(n6056), .ZN(n6053) );
  INV_X1 U7061 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7778) );
  INV_X1 U7062 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8294) );
  MUX2_X1 U7063 ( .A(n7778), .B(n8294), .S(n8662), .Z(n6050) );
  INV_X1 U7064 ( .A(SI_23_), .ZN(n8401) );
  NAND2_X1 U7065 ( .A1(n6050), .A2(n8401), .ZN(n6069) );
  INV_X1 U7066 ( .A(n6050), .ZN(n6051) );
  NAND2_X1 U7067 ( .A1(n6051), .A2(SI_23_), .ZN(n6052) );
  NAND2_X1 U7068 ( .A1(n6069), .A2(n6052), .ZN(n6054) );
  NAND2_X1 U7069 ( .A1(n6053), .A2(n6054), .ZN(n6057) );
  INV_X1 U7070 ( .A(n6054), .ZN(n6055) );
  NAND2_X1 U7071 ( .A1(n6057), .A2(n6070), .ZN(n7776) );
  NAND2_X1 U7072 ( .A1(n7776), .A2(n9893), .ZN(n6059) );
  OR2_X1 U7073 ( .A1(n9895), .A2(n8294), .ZN(n6058) );
  NAND2_X1 U7074 ( .A1(n9885), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6068) );
  INV_X1 U7075 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n6060) );
  OR2_X1 U7076 ( .A1(n9889), .A2(n6060), .ZN(n6067) );
  INV_X1 U7077 ( .A(n6062), .ZN(n6061) );
  NAND2_X1 U7078 ( .A1(n6061), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6077) );
  INV_X1 U7079 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9736) );
  NAND2_X1 U7080 ( .A1(n6062), .A2(n9736), .ZN(n6063) );
  NAND2_X1 U7081 ( .A1(n6077), .A2(n6063), .ZN(n10392) );
  OR2_X1 U7082 ( .A1(n6167), .A2(n10392), .ZN(n6066) );
  INV_X1 U7083 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n6064) );
  OR2_X1 U7084 ( .A1(n9887), .A2(n6064), .ZN(n6065) );
  NAND4_X1 U7085 ( .A1(n6068), .A2(n6067), .A3(n6066), .A4(n6065), .ZN(n10376)
         );
  INV_X1 U7086 ( .A(n10501), .ZN(n10396) );
  INV_X1 U7087 ( .A(n10376), .ZN(n10417) );
  INV_X1 U7088 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8059) );
  INV_X1 U7089 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8508) );
  MUX2_X1 U7090 ( .A(n8059), .B(n8508), .S(n8662), .Z(n6071) );
  INV_X1 U7091 ( .A(SI_24_), .ZN(n8388) );
  NAND2_X1 U7092 ( .A1(n6071), .A2(n8388), .ZN(n6089) );
  INV_X1 U7093 ( .A(n6071), .ZN(n6072) );
  NAND2_X1 U7094 ( .A1(n6072), .A2(SI_24_), .ZN(n6073) );
  AND2_X1 U7095 ( .A1(n6089), .A2(n6073), .ZN(n6087) );
  NAND2_X1 U7096 ( .A1(n7958), .A2(n9893), .ZN(n6075) );
  OR2_X1 U7097 ( .A1(n9895), .A2(n8508), .ZN(n6074) );
  NAND2_X1 U7098 ( .A1(n5825), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6083) );
  INV_X1 U7099 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n10498) );
  OR2_X1 U7100 ( .A1(n6209), .A2(n10498), .ZN(n6082) );
  INV_X1 U7101 ( .A(n6077), .ZN(n6076) );
  NAND2_X1 U7102 ( .A1(n6076), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6102) );
  INV_X1 U7103 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9811) );
  NAND2_X1 U7104 ( .A1(n6077), .A2(n9811), .ZN(n6078) );
  NAND2_X1 U7105 ( .A1(n6102), .A2(n6078), .ZN(n10383) );
  OR2_X1 U7106 ( .A1(n5791), .A2(n10383), .ZN(n6081) );
  INV_X1 U7107 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n10384) );
  OR2_X1 U7108 ( .A1(n6079), .A2(n10384), .ZN(n6080) );
  NAND4_X1 U7109 ( .A1(n6083), .A2(n6082), .A3(n6081), .A4(n6080), .ZN(n10400)
         );
  INV_X1 U7110 ( .A(n10382), .ZN(n10567) );
  INV_X1 U7111 ( .A(n10400), .ZN(n9775) );
  OAI21_X1 U7112 ( .B1(n10380), .B2(n6085), .A(n6084), .ZN(n6086) );
  INV_X1 U7113 ( .A(n6086), .ZN(n10359) );
  INV_X1 U7114 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8617) );
  INV_X1 U7115 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8043) );
  INV_X1 U7116 ( .A(SI_25_), .ZN(n6090) );
  NAND2_X1 U7117 ( .A1(n6091), .A2(n6090), .ZN(n6111) );
  INV_X1 U7118 ( .A(n6091), .ZN(n6092) );
  NAND2_X1 U7119 ( .A1(n6092), .A2(SI_25_), .ZN(n6093) );
  AND2_X1 U7120 ( .A1(n6111), .A2(n6093), .ZN(n6094) );
  OR2_X1 U7121 ( .A1(n6095), .A2(n6094), .ZN(n6096) );
  NAND2_X1 U7122 ( .A1(n6112), .A2(n6096), .ZN(n8042) );
  NAND2_X1 U7123 ( .A1(n8042), .A2(n9893), .ZN(n6098) );
  OR2_X1 U7124 ( .A1(n9895), .A2(n8043), .ZN(n6097) );
  NAND2_X1 U7125 ( .A1(n5825), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6108) );
  INV_X1 U7126 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n6099) );
  OR2_X1 U7127 ( .A1(n6209), .A2(n6099), .ZN(n6107) );
  INV_X1 U7128 ( .A(n6102), .ZN(n6100) );
  NAND2_X1 U7129 ( .A1(n6100), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6123) );
  INV_X1 U7130 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6101) );
  NAND2_X1 U7131 ( .A1(n6102), .A2(n6101), .ZN(n6103) );
  NAND2_X1 U7132 ( .A1(n6123), .A2(n6103), .ZN(n10362) );
  OR2_X1 U7133 ( .A1(n6167), .A2(n10362), .ZN(n6106) );
  INV_X1 U7134 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n6104) );
  OR2_X1 U7135 ( .A1(n9887), .A2(n6104), .ZN(n6105) );
  NAND4_X1 U7136 ( .A1(n6108), .A2(n6107), .A3(n6106), .A4(n6105), .ZN(n10375)
         );
  NAND2_X1 U7137 ( .A1(n10359), .A2(n6109), .ZN(n6110) );
  INV_X1 U7138 ( .A(n10375), .ZN(n9875) );
  NAND2_X1 U7139 ( .A1(n6110), .A2(n5600), .ZN(n10347) );
  INV_X1 U7140 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8105) );
  INV_X1 U7141 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8106) );
  INV_X1 U7142 ( .A(SI_26_), .ZN(n8386) );
  NAND2_X1 U7143 ( .A1(n6113), .A2(n8386), .ZN(n6130) );
  INV_X1 U7144 ( .A(n6113), .ZN(n6114) );
  NAND2_X1 U7145 ( .A1(n6114), .A2(SI_26_), .ZN(n6115) );
  AND2_X1 U7146 ( .A1(n6130), .A2(n6115), .ZN(n6116) );
  OR2_X1 U7147 ( .A1(n6117), .A2(n6116), .ZN(n6118) );
  NAND2_X1 U7148 ( .A1(n6131), .A2(n6118), .ZN(n8103) );
  NAND2_X1 U7149 ( .A1(n8103), .A2(n9893), .ZN(n6120) );
  OR2_X1 U7150 ( .A1(n9895), .A2(n8106), .ZN(n6119) );
  NAND2_X1 U7151 ( .A1(n5825), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6128) );
  INV_X1 U7152 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n10488) );
  OR2_X1 U7153 ( .A1(n6209), .A2(n10488), .ZN(n6127) );
  INV_X1 U7154 ( .A(n6123), .ZN(n6121) );
  NAND2_X1 U7155 ( .A1(n6121), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6142) );
  INV_X1 U7156 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6122) );
  NAND2_X1 U7157 ( .A1(n6123), .A2(n6122), .ZN(n6124) );
  NAND2_X1 U7158 ( .A1(n6142), .A2(n6124), .ZN(n10351) );
  OR2_X1 U7159 ( .A1(n6167), .A2(n10351), .ZN(n6126) );
  INV_X1 U7160 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n10352) );
  OR2_X1 U7161 ( .A1(n9887), .A2(n10352), .ZN(n6125) );
  NAND2_X1 U7162 ( .A1(n10350), .A2(n10325), .ZN(n10044) );
  NAND2_X1 U7163 ( .A1(n10049), .A2(n10044), .ZN(n6202) );
  INV_X1 U7164 ( .A(n10325), .ZN(n10368) );
  INV_X1 U7165 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8133) );
  INV_X1 U7166 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8290) );
  MUX2_X1 U7167 ( .A(n8133), .B(n8290), .S(n8662), .Z(n6132) );
  INV_X1 U7168 ( .A(SI_27_), .ZN(n8387) );
  NAND2_X1 U7169 ( .A1(n6132), .A2(n8387), .ZN(n6148) );
  INV_X1 U7170 ( .A(n6132), .ZN(n6133) );
  NAND2_X1 U7171 ( .A1(n6133), .A2(SI_27_), .ZN(n6134) );
  AND2_X1 U7172 ( .A1(n6148), .A2(n6134), .ZN(n6135) );
  NAND2_X1 U7173 ( .A1(n8134), .A2(n5806), .ZN(n6139) );
  OR2_X1 U7174 ( .A1(n9895), .A2(n8290), .ZN(n6138) );
  NAND2_X1 U7175 ( .A1(n5825), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6147) );
  INV_X1 U7176 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n10482) );
  OR2_X1 U7177 ( .A1(n6209), .A2(n10482), .ZN(n6146) );
  INV_X1 U7178 ( .A(n6142), .ZN(n6140) );
  NAND2_X1 U7179 ( .A1(n6140), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n6153) );
  INV_X1 U7180 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6141) );
  NAND2_X1 U7181 ( .A1(n6142), .A2(n6141), .ZN(n6143) );
  NAND2_X1 U7182 ( .A1(n6153), .A2(n6143), .ZN(n10332) );
  OR2_X1 U7183 ( .A1(n5791), .A2(n10332), .ZN(n6145) );
  INV_X1 U7184 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n10333) );
  OR2_X1 U7185 ( .A1(n9887), .A2(n10333), .ZN(n6144) );
  OR2_X1 U7186 ( .A1(n10556), .A2(n10309), .ZN(n10053) );
  NAND2_X1 U7187 ( .A1(n10556), .A2(n10309), .ZN(n10052) );
  NAND2_X1 U7188 ( .A1(n10053), .A2(n10052), .ZN(n6203) );
  INV_X1 U7189 ( .A(SI_28_), .ZN(n8396) );
  XNOR2_X1 U7190 ( .A(n6162), .B(n8396), .ZN(n6160) );
  NAND2_X1 U7191 ( .A1(n8609), .A2(n9893), .ZN(n6151) );
  INV_X1 U7192 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8181) );
  OR2_X1 U7193 ( .A1(n9895), .A2(n8181), .ZN(n6150) );
  NAND2_X1 U7194 ( .A1(n5825), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6158) );
  INV_X1 U7195 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n10475) );
  OR2_X1 U7196 ( .A1(n6209), .A2(n10475), .ZN(n6157) );
  INV_X1 U7197 ( .A(n6153), .ZN(n6152) );
  NAND2_X1 U7198 ( .A1(n6152), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n10297) );
  INV_X1 U7199 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9008) );
  NAND2_X1 U7200 ( .A1(n6153), .A2(n9008), .ZN(n6154) );
  NAND2_X1 U7201 ( .A1(n10297), .A2(n6154), .ZN(n10317) );
  OR2_X1 U7202 ( .A1(n6167), .A2(n10317), .ZN(n6156) );
  INV_X1 U7203 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n10318) );
  OR2_X1 U7204 ( .A1(n9887), .A2(n10318), .ZN(n6155) );
  NAND2_X1 U7205 ( .A1(n10553), .A2(n10326), .ZN(n10057) );
  INV_X1 U7206 ( .A(n6162), .ZN(n6163) );
  INV_X1 U7207 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9717) );
  INV_X1 U7208 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10596) );
  MUX2_X1 U7209 ( .A(n9717), .B(n10596), .S(n8662), .Z(n8644) );
  NAND2_X1 U7210 ( .A1(n9716), .A2(n9893), .ZN(n6165) );
  OR2_X1 U7211 ( .A1(n9895), .A2(n10596), .ZN(n6164) );
  NAND2_X1 U7212 ( .A1(n5825), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6172) );
  INV_X1 U7213 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6166) );
  OR2_X1 U7214 ( .A1(n6209), .A2(n6166), .ZN(n6171) );
  OR2_X1 U7215 ( .A1(n6167), .A2(n10297), .ZN(n6170) );
  INV_X1 U7216 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n6168) );
  OR2_X1 U7217 ( .A1(n9887), .A2(n6168), .ZN(n6169) );
  NAND2_X1 U7218 ( .A1(n10299), .A2(n10310), .ZN(n10132) );
  INV_X1 U7219 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8577) );
  NAND2_X1 U7220 ( .A1(n6177), .A2(n8577), .ZN(n6217) );
  NAND2_X1 U7221 ( .A1(n6217), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6225) );
  NAND2_X1 U7222 ( .A1(n6225), .A2(n8359), .ZN(n6176) );
  NAND2_X1 U7223 ( .A1(n10111), .A2(n10274), .ZN(n7028) );
  INV_X1 U7224 ( .A(n6177), .ZN(n6178) );
  NAND2_X1 U7225 ( .A1(n6178), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6179) );
  XNOR2_X1 U7226 ( .A(n6179), .B(n8577), .ZN(n7536) );
  NAND2_X1 U7227 ( .A1(n10107), .A2(n7536), .ZN(n7027) );
  OR2_X1 U7228 ( .A1(n7028), .A2(n7027), .ZN(n10147) );
  INV_X1 U7229 ( .A(n10107), .ZN(n10117) );
  NAND2_X1 U7230 ( .A1(n10151), .A2(n10117), .ZN(n7090) );
  AND2_X1 U7231 ( .A1(n10274), .A2(n7536), .ZN(n7022) );
  INV_X1 U7232 ( .A(n7022), .ZN(n6180) );
  NAND2_X1 U7233 ( .A1(n7028), .A2(n6180), .ZN(n6181) );
  NAND3_X1 U7234 ( .A1(n10147), .A2(n7090), .A3(n6181), .ZN(n7917) );
  NAND2_X1 U7235 ( .A1(n10151), .A2(n10280), .ZN(n10060) );
  INV_X1 U7236 ( .A(n7536), .ZN(n10145) );
  OR2_X1 U7237 ( .A1(n10060), .A2(n10145), .ZN(n8045) );
  NAND2_X1 U7238 ( .A1(n10111), .A2(n10280), .ZN(n6183) );
  NAND2_X1 U7239 ( .A1(n10107), .A2(n10145), .ZN(n6182) );
  NAND2_X1 U7240 ( .A1(n6183), .A2(n6182), .ZN(n10402) );
  OR2_X1 U7241 ( .A1(n10382), .A2(n9775), .ZN(n10048) );
  NAND2_X1 U7242 ( .A1(n10382), .A2(n9775), .ZN(n10040) );
  OR2_X1 U7243 ( .A1(n10501), .A2(n10417), .ZN(n10036) );
  NAND2_X1 U7244 ( .A1(n10501), .A2(n10417), .ZN(n10037) );
  AND2_X1 U7245 ( .A1(n10034), .A2(n10029), .ZN(n9930) );
  OR2_X1 U7246 ( .A1(n10522), .A2(n10448), .ZN(n10019) );
  NAND2_X1 U7247 ( .A1(n10522), .A2(n10448), .ZN(n10027) );
  INV_X1 U7248 ( .A(n7382), .ZN(n9905) );
  NOR2_X1 U7249 ( .A1(n9906), .A2(n9905), .ZN(n7319) );
  NAND2_X1 U7250 ( .A1(n6185), .A2(n5247), .ZN(n6186) );
  INV_X1 U7251 ( .A(n10065), .ZN(n7285) );
  NAND2_X1 U7252 ( .A1(n10905), .A2(n10904), .ZN(n6187) );
  INV_X1 U7253 ( .A(n10903), .ZN(n10066) );
  NAND2_X1 U7254 ( .A1(n6187), .A2(n10066), .ZN(n10907) );
  INV_X1 U7255 ( .A(n9820), .ZN(n10955) );
  NAND2_X1 U7256 ( .A1(n9745), .A2(n10955), .ZN(n9953) );
  INV_X1 U7257 ( .A(n10071), .ZN(n6188) );
  AND2_X1 U7258 ( .A1(n9912), .A2(n10070), .ZN(n6189) );
  OR2_X1 U7259 ( .A1(n7549), .A2(n7627), .ZN(n7422) );
  NAND2_X1 U7260 ( .A1(n9977), .A2(n7422), .ZN(n9973) );
  NAND2_X1 U7261 ( .A1(n9967), .A2(n9962), .ZN(n6190) );
  NOR2_X1 U7262 ( .A1(n9973), .A2(n6190), .ZN(n10078) );
  NAND2_X1 U7263 ( .A1(n7303), .A2(n10078), .ZN(n6192) );
  NAND2_X1 U7264 ( .A1(n7549), .A2(n7627), .ZN(n9971) );
  AND2_X1 U7265 ( .A1(n9971), .A2(n9966), .ZN(n10077) );
  OR2_X1 U7266 ( .A1(n9973), .A2(n10077), .ZN(n6191) );
  AND2_X1 U7267 ( .A1(n6191), .A2(n10075), .ZN(n9916) );
  NAND2_X1 U7268 ( .A1(n6192), .A2(n9916), .ZN(n7452) );
  INV_X1 U7269 ( .A(n10163), .ZN(n7983) );
  OR2_X1 U7270 ( .A1(n11055), .A2(n7983), .ZN(n9976) );
  NAND2_X1 U7271 ( .A1(n11055), .A2(n7983), .ZN(n9983) );
  NAND2_X1 U7272 ( .A1(n9976), .A2(n9983), .ZN(n11023) );
  INV_X1 U7273 ( .A(n11021), .ZN(n9978) );
  NOR2_X1 U7274 ( .A1(n11023), .A2(n9978), .ZN(n6193) );
  NAND2_X1 U7275 ( .A1(n11022), .A2(n6193), .ZN(n6194) );
  NAND2_X1 U7276 ( .A1(n6194), .A2(n9976), .ZN(n7638) );
  INV_X1 U7277 ( .A(n11025), .ZN(n8036) );
  OR2_X1 U7278 ( .A1(n7973), .A2(n8036), .ZN(n9988) );
  NAND2_X1 U7279 ( .A1(n7973), .A2(n8036), .ZN(n9980) );
  AND2_X1 U7280 ( .A1(n9988), .A2(n9980), .ZN(n10083) );
  INV_X1 U7281 ( .A(n10162), .ZN(n8125) );
  OR2_X1 U7282 ( .A1(n8029), .A2(n8125), .ZN(n9994) );
  NAND2_X1 U7283 ( .A1(n8029), .A2(n8125), .ZN(n9989) );
  NAND2_X1 U7284 ( .A1(n9994), .A2(n9989), .ZN(n10085) );
  INV_X1 U7285 ( .A(n10161), .ZN(n8622) );
  OR2_X1 U7286 ( .A1(n8128), .A2(n8622), .ZN(n9997) );
  NAND2_X1 U7287 ( .A1(n8128), .A2(n8622), .ZN(n9999) );
  NAND2_X1 U7288 ( .A1(n9997), .A2(n9999), .ZN(n10086) );
  INV_X1 U7289 ( .A(n9989), .ZN(n6195) );
  NOR2_X1 U7290 ( .A1(n10086), .A2(n6195), .ZN(n6196) );
  NAND2_X1 U7291 ( .A1(n6197), .A2(n9997), .ZN(n8620) );
  NAND2_X1 U7292 ( .A1(n8620), .A2(n10005), .ZN(n6198) );
  INV_X1 U7293 ( .A(n10004), .ZN(n10010) );
  NAND2_X1 U7294 ( .A1(n10017), .A2(n8136), .ZN(n10091) );
  NAND2_X1 U7295 ( .A1(n10024), .A2(n8137), .ZN(n10016) );
  NAND2_X1 U7296 ( .A1(n10016), .A2(n10017), .ZN(n6199) );
  NAND2_X1 U7297 ( .A1(n10093), .A2(n8159), .ZN(n6200) );
  NAND2_X1 U7298 ( .A1(n6200), .A2(n10027), .ZN(n10445) );
  INV_X1 U7299 ( .A(n10026), .ZN(n10422) );
  NAND2_X1 U7300 ( .A1(n10034), .A2(n10422), .ZN(n6201) );
  AND2_X1 U7301 ( .A1(n6201), .A2(n10033), .ZN(n9932) );
  OR2_X1 U7302 ( .A1(n10491), .A2(n9875), .ZN(n10042) );
  NAND2_X1 U7303 ( .A1(n10491), .A2(n9875), .ZN(n9898) );
  NAND2_X1 U7304 ( .A1(n10042), .A2(n9898), .ZN(n10358) );
  NAND2_X1 U7305 ( .A1(n10324), .A2(n10329), .ZN(n6204) );
  NAND2_X1 U7306 ( .A1(n6204), .A2(n10052), .ZN(n10307) );
  INV_X1 U7307 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n6208) );
  NAND2_X1 U7308 ( .A1(n6205), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6207) );
  NAND2_X1 U7309 ( .A1(n5825), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6206) );
  OAI211_X1 U7310 ( .C1(n6209), .C2(n6208), .A(n6207), .B(n6206), .ZN(n10155)
         );
  NAND2_X1 U7311 ( .A1(n10111), .A2(n10107), .ZN(n10106) );
  INV_X1 U7312 ( .A(n6210), .ZN(n7066) );
  OR2_X1 U7313 ( .A1(n10106), .A2(n7066), .ZN(n10902) );
  INV_X1 U7314 ( .A(P1_B_REG_SCAN_IN), .ZN(n10150) );
  NOR2_X1 U7315 ( .A1(n10660), .A2(n10150), .ZN(n6211) );
  NOR2_X1 U7316 ( .A1(n10902), .A2(n6211), .ZN(n10286) );
  INV_X1 U7317 ( .A(n10106), .ZN(n10138) );
  INV_X1 U7318 ( .A(n10507), .ZN(n10409) );
  INV_X1 U7319 ( .A(n9864), .ZN(n10580) );
  NAND2_X1 U7320 ( .A1(n10898), .A2(n10899), .ZN(n10897) );
  INV_X1 U7321 ( .A(n7433), .ZN(n10983) );
  INV_X1 U7322 ( .A(n11055), .ZN(n11037) );
  NAND2_X1 U7323 ( .A1(n11036), .A2(n11037), .ZN(n11034) );
  INV_X1 U7324 ( .A(n6212), .ZN(n7675) );
  INV_X1 U7325 ( .A(n8128), .ZN(n8056) );
  INV_X1 U7326 ( .A(n10540), .ZN(n8630) );
  AOI21_X1 U7327 ( .B1(n10299), .B2(n5135), .A(n10438), .ZN(n6214) );
  NAND2_X1 U7328 ( .A1(n6214), .A2(n10290), .ZN(n10301) );
  OAI211_X1 U7329 ( .C1(n10295), .C2(n10543), .A(n10305), .B(n10301), .ZN(
        n6253) );
  INV_X1 U7330 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n8582) );
  NAND2_X1 U7331 ( .A1(n6215), .A2(n8582), .ZN(n6216) );
  OAI21_X1 U7332 ( .B1(n6221), .B2(P1_IR_REG_25__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6218) );
  MUX2_X1 U7333 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6218), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n6220) );
  NAND2_X1 U7334 ( .A1(n6220), .A2(n6219), .ZN(n8108) );
  NAND2_X1 U7335 ( .A1(n6221), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6222) );
  XNOR2_X1 U7336 ( .A(n6222), .B(P1_IR_REG_25__SCAN_IN), .ZN(n6232) );
  NAND2_X1 U7337 ( .A1(n6223), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6224) );
  NAND2_X1 U7338 ( .A1(n6225), .A2(n6224), .ZN(n6226) );
  XNOR2_X1 U7339 ( .A(n6226), .B(n8582), .ZN(n6248) );
  INV_X1 U7340 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n8581) );
  NAND2_X1 U7341 ( .A1(n6228), .A2(n8581), .ZN(n6229) );
  NAND2_X1 U7342 ( .A1(n6229), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6231) );
  INV_X1 U7343 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6230) );
  XNOR2_X1 U7344 ( .A(n6231), .B(n6230), .ZN(n7743) );
  OAI211_X1 U7345 ( .C1(n10106), .C2(n7022), .A(n7032), .B(n7743), .ZN(n7128)
         );
  NOR2_X1 U7346 ( .A1(n7128), .A2(P1_U3086), .ZN(n7040) );
  INV_X1 U7347 ( .A(n6232), .ZN(n8044) );
  NAND2_X1 U7348 ( .A1(n8044), .A2(P1_B_REG_SCAN_IN), .ZN(n6233) );
  MUX2_X1 U7349 ( .A(n6233), .B(P1_B_REG_SCAN_IN), .S(n6248), .Z(n6235) );
  NAND2_X1 U7350 ( .A1(n6235), .A2(n6234), .ZN(n10583) );
  INV_X1 U7351 ( .A(n10583), .ZN(n6246) );
  NOR4_X1 U7352 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_27__SCAN_IN), .ZN(n6244) );
  NOR4_X1 U7353 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n6243) );
  OR4_X1 U7354 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6241) );
  NOR4_X1 U7355 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n6239) );
  NOR4_X1 U7356 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n6238) );
  NOR4_X1 U7357 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n6237) );
  NOR4_X1 U7358 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n6236) );
  NAND4_X1 U7359 ( .A1(n6239), .A2(n6238), .A3(n6237), .A4(n6236), .ZN(n6240)
         );
  NOR4_X1 U7360 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        n6241), .A4(n6240), .ZN(n6242) );
  NAND3_X1 U7361 ( .A1(n6244), .A2(n6243), .A3(n6242), .ZN(n6245) );
  NAND2_X1 U7362 ( .A1(n6246), .A2(n6245), .ZN(n7019) );
  NAND2_X1 U7363 ( .A1(n7040), .A2(n7019), .ZN(n7283) );
  NAND2_X1 U7364 ( .A1(n8108), .A2(n8044), .ZN(n10585) );
  OAI21_X1 U7365 ( .B1(n10583), .B2(P1_D_REG_1__SCAN_IN), .A(n10585), .ZN(
        n7018) );
  NAND2_X1 U7366 ( .A1(n7018), .A2(n7038), .ZN(n6247) );
  INV_X1 U7367 ( .A(n6248), .ZN(n7959) );
  NAND2_X1 U7368 ( .A1(n8108), .A2(n7959), .ZN(n10586) );
  OAI21_X1 U7369 ( .B1(n10583), .B2(P1_D_REG_0__SCAN_IN), .A(n10586), .ZN(
        n7280) );
  NOR2_X2 U7370 ( .A1(n6252), .A2(n7280), .ZN(n10529) );
  MUX2_X1 U7371 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n6253), .S(n11081), .Z(n6249) );
  INV_X1 U7372 ( .A(n6249), .ZN(n6251) );
  OR2_X1 U7373 ( .A1(n7090), .A2(n7022), .ZN(n11074) );
  INV_X1 U7374 ( .A(n11074), .ZN(n10541) );
  NAND2_X1 U7375 ( .A1(n6251), .A2(n6250), .ZN(P1_U3551) );
  INV_X1 U7376 ( .A(n7280), .ZN(n7020) );
  INV_X2 U7377 ( .A(n11082), .ZN(n11085) );
  MUX2_X1 U7378 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n6253), .S(n11085), .Z(n6254) );
  INV_X1 U7379 ( .A(n6254), .ZN(n6256) );
  NAND2_X1 U7380 ( .A1(n10299), .A2(n10557), .ZN(n6255) );
  NAND2_X1 U7381 ( .A1(n6256), .A2(n6255), .ZN(P1_U3519) );
  INV_X1 U7382 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6753) );
  NOR2_X1 U7383 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n6265) );
  NOR2_X1 U7384 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n6264) );
  NOR2_X1 U7385 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n6263) );
  INV_X1 U7386 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6268) );
  INV_X1 U7387 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6269) );
  INV_X1 U7388 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6287) );
  NAND2_X1 U7389 ( .A1(n8103), .A2(n6416), .ZN(n6273) );
  OR2_X1 U7390 ( .A1(n6360), .A2(n8105), .ZN(n6272) );
  INV_X1 U7391 ( .A(n9406), .ZN(n9667) );
  INV_X1 U7392 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8255) );
  INV_X1 U7393 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8488) );
  INV_X1 U7394 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8500) );
  INV_X1 U7395 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8476) );
  INV_X1 U7396 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8247) );
  INV_X1 U7397 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8484) );
  INV_X1 U7398 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n6284) );
  INV_X1 U7399 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8263) );
  INV_X1 U7400 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8469) );
  XNOR2_X1 U7401 ( .A(n6639), .B(P2_REG3_REG_26__SCAN_IN), .ZN(n9402) );
  INV_X1 U7402 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6290) );
  INV_X1 U7403 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9711) );
  XNOR2_X2 U7404 ( .A(n6291), .B(n6290), .ZN(n9718) );
  NAND2_X1 U7405 ( .A1(n9402), .A2(n6671), .ZN(n6299) );
  INV_X1 U7406 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n9403) );
  NAND2_X2 U7407 ( .A1(n6293), .A2(n6294), .ZN(n6338) );
  NAND2_X1 U7408 ( .A1(n6300), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6296) );
  AND2_X2 U7409 ( .A1(n6293), .A2(n9718), .ZN(n6307) );
  NAND2_X1 U7410 ( .A1(n8678), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6295) );
  OAI211_X1 U7411 ( .C1(n9403), .C2(n5110), .A(n6296), .B(n6295), .ZN(n6297)
         );
  INV_X1 U7412 ( .A(n6297), .ZN(n6298) );
  NAND2_X1 U7413 ( .A1(n5109), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6304) );
  INV_X1 U7414 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7147) );
  OR2_X1 U7415 ( .A1(n6478), .A2(n7147), .ZN(n6303) );
  INV_X1 U7416 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6964) );
  NAND2_X1 U7417 ( .A1(n6307), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6301) );
  NAND2_X1 U7418 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6305) );
  NAND2_X2 U7419 ( .A1(n8706), .A2(n6683), .ZN(n8857) );
  NAND2_X1 U7420 ( .A1(n6307), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6311) );
  INV_X1 U7421 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6929) );
  OR2_X1 U7422 ( .A1(n5108), .A2(n6929), .ZN(n6310) );
  INV_X1 U7423 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6933) );
  INV_X1 U7424 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6828) );
  NAND2_X1 U7425 ( .A1(n6772), .A2(SI_0_), .ZN(n6312) );
  XNOR2_X1 U7426 ( .A(n6312), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9720) );
  MUX2_X1 U7427 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9720), .S(n6313), .Z(n6680) );
  NAND2_X1 U7428 ( .A1(n8857), .A2(n7145), .ZN(n7144) );
  CLKBUF_X1 U7429 ( .A(n6951), .Z(n7048) );
  INV_X1 U7430 ( .A(n7148), .ZN(n10869) );
  NAND2_X1 U7431 ( .A1(n7048), .A2(n10869), .ZN(n6314) );
  NAND2_X1 U7432 ( .A1(n7144), .A2(n6314), .ZN(n7201) );
  NAND2_X1 U7433 ( .A1(n6307), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6318) );
  INV_X1 U7434 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7341) );
  OR2_X1 U7435 ( .A1(n6338), .A2(n7341), .ZN(n6317) );
  INV_X1 U7436 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6873) );
  OR2_X1 U7437 ( .A1(n6478), .A2(n6873), .ZN(n6316) );
  INV_X1 U7438 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7208) );
  OR2_X1 U7439 ( .A1(n5108), .A2(n7208), .ZN(n6315) );
  NOR2_X1 U7440 ( .A1(n6849), .A2(n6269), .ZN(n6319) );
  INV_X1 U7441 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6771) );
  OR2_X1 U7442 ( .A1(n6360), .A2(n6771), .ZN(n6324) );
  OR2_X1 U7443 ( .A1(n6377), .A2(n6775), .ZN(n6323) );
  OR2_X1 U7444 ( .A1(n10925), .A2(n8710), .ZN(n6325) );
  NAND2_X1 U7445 ( .A1(n7200), .A2(n6325), .ZN(n10924) );
  NAND2_X1 U7446 ( .A1(n6307), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6331) );
  INV_X1 U7447 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6326) );
  INV_X1 U7448 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6327) );
  OR2_X1 U7449 ( .A1(n8680), .A2(n6327), .ZN(n6329) );
  NAND2_X1 U7450 ( .A1(n6386), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6344) );
  XNOR2_X1 U7451 ( .A(n6344), .B(P2_IR_REG_3__SCAN_IN), .ZN(n10815) );
  OR2_X1 U7452 ( .A1(n6377), .A2(n6780), .ZN(n6333) );
  INV_X1 U7453 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6781) );
  OR2_X1 U7454 ( .A1(n6360), .A2(n6781), .ZN(n6332) );
  NAND2_X1 U7455 ( .A1(n9204), .A2(n10933), .ZN(n6334) );
  NAND2_X1 U7456 ( .A1(n10924), .A2(n6334), .ZN(n6336) );
  OR2_X1 U7457 ( .A1(n9204), .A2(n10933), .ZN(n6335) );
  NAND2_X1 U7458 ( .A1(n6307), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6343) );
  INV_X1 U7459 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6337) );
  NAND2_X1 U7460 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6339) );
  AND2_X1 U7461 ( .A1(n6350), .A2(n6339), .ZN(n7393) );
  OR2_X1 U7462 ( .A1(n5108), .A2(n7393), .ZN(n6341) );
  INV_X1 U7463 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7392) );
  OR2_X1 U7464 ( .A1(n5110), .A2(n7392), .ZN(n6340) );
  INV_X1 U7465 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n6383) );
  NAND2_X1 U7466 ( .A1(n6344), .A2(n6383), .ZN(n6345) );
  NAND2_X1 U7467 ( .A1(n6345), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6358) );
  INV_X1 U7468 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6346) );
  OR2_X1 U7469 ( .A1(n6360), .A2(n6346), .ZN(n6348) );
  OR2_X1 U7470 ( .A1(n6377), .A2(n6773), .ZN(n6347) );
  NAND2_X1 U7471 ( .A1(n6307), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6356) );
  INV_X1 U7472 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6349) );
  OR2_X1 U7473 ( .A1(n8680), .A2(n6349), .ZN(n6355) );
  NAND2_X1 U7474 ( .A1(n6350), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6351) );
  AND2_X1 U7475 ( .A1(n6368), .A2(n6351), .ZN(n7514) );
  OR2_X1 U7476 ( .A1(n5108), .A2(n7514), .ZN(n6354) );
  INV_X1 U7477 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7513) );
  INV_X1 U7478 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6357) );
  NAND2_X1 U7479 ( .A1(n6358), .A2(n6357), .ZN(n6359) );
  NAND2_X1 U7480 ( .A1(n6359), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6374) );
  XNOR2_X1 U7481 ( .A(n6374), .B(P2_IR_REG_5__SCAN_IN), .ZN(n10847) );
  INV_X1 U7482 ( .A(n10847), .ZN(n7353) );
  OR2_X1 U7483 ( .A1(n6377), .A2(n6783), .ZN(n6362) );
  OR2_X1 U7484 ( .A1(n6360), .A2(n5627), .ZN(n6361) );
  OAI211_X1 U7485 ( .C1(n6313), .C2(n7353), .A(n6362), .B(n6361), .ZN(n7516)
         );
  INV_X1 U7486 ( .A(n7516), .ZN(n10961) );
  NAND2_X1 U7487 ( .A1(n6363), .A2(n10961), .ZN(n6367) );
  INV_X1 U7488 ( .A(n7511), .ZN(n6365) );
  INV_X1 U7489 ( .A(n7171), .ZN(n6364) );
  NAND2_X1 U7490 ( .A1(n6365), .A2(n6364), .ZN(n6366) );
  NAND2_X1 U7491 ( .A1(n6367), .A2(n6366), .ZN(n7575) );
  NAND2_X1 U7492 ( .A1(n8678), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6372) );
  INV_X1 U7493 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7349) );
  OR2_X1 U7494 ( .A1(n5110), .A2(n7349), .ZN(n6371) );
  XNOR2_X1 U7495 ( .A(n6368), .B(n8495), .ZN(n7580) );
  OR2_X1 U7496 ( .A1(n5108), .A2(n7580), .ZN(n6370) );
  INV_X1 U7497 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7348) );
  OR2_X1 U7498 ( .A1(n8680), .A2(n7348), .ZN(n6369) );
  INV_X1 U7499 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6373) );
  NAND2_X1 U7500 ( .A1(n6374), .A2(n6373), .ZN(n6375) );
  NAND2_X1 U7501 ( .A1(n6375), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6376) );
  XNOR2_X1 U7502 ( .A(n6376), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7352) );
  OR2_X1 U7503 ( .A1(n6377), .A2(n6785), .ZN(n6379) );
  INV_X1 U7504 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6782) );
  OR2_X1 U7505 ( .A1(n6360), .A2(n6782), .ZN(n6378) );
  OAI211_X1 U7506 ( .C1(n6313), .C2(n7557), .A(n6379), .B(n6378), .ZN(n7179)
         );
  INV_X1 U7507 ( .A(n7179), .ZN(n10974) );
  NAND2_X1 U7508 ( .A1(n9203), .A2(n10974), .ZN(n8726) );
  NAND2_X1 U7509 ( .A1(n8745), .A2(n8726), .ZN(n7577) );
  NAND2_X1 U7510 ( .A1(n7575), .A2(n7577), .ZN(n6381) );
  OR2_X1 U7511 ( .A1(n9203), .A2(n7179), .ZN(n6380) );
  NAND2_X1 U7512 ( .A1(n6381), .A2(n6380), .ZN(n7655) );
  AND2_X1 U7513 ( .A1(n6786), .A2(n6416), .ZN(n6394) );
  INV_X1 U7514 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6384) );
  NAND3_X1 U7515 ( .A1(n6382), .A2(n6384), .A3(n6383), .ZN(n6385) );
  OR2_X1 U7516 ( .A1(n6386), .A2(n6385), .ZN(n6388) );
  NAND2_X1 U7517 ( .A1(n6388), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6387) );
  MUX2_X1 U7518 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6387), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n6391) );
  INV_X1 U7519 ( .A(n6388), .ZN(n6390) );
  INV_X1 U7520 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6389) );
  NAND2_X1 U7521 ( .A1(n6390), .A2(n6389), .ZN(n6417) );
  NAND2_X1 U7522 ( .A1(n6391), .A2(n6417), .ZN(n7690) );
  NOR2_X1 U7523 ( .A1(n6313), .A2(n7690), .ZN(n6393) );
  INV_X1 U7524 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6789) );
  NOR2_X1 U7525 ( .A1(n6360), .A2(n6789), .ZN(n6392) );
  NAND2_X1 U7526 ( .A1(n6307), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6402) );
  INV_X1 U7527 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6395) );
  OR2_X1 U7528 ( .A1(n8680), .A2(n6395), .ZN(n6401) );
  INV_X1 U7529 ( .A(n6396), .ZN(n6397) );
  NAND2_X1 U7530 ( .A1(n6397), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6398) );
  AND2_X1 U7531 ( .A1(n6405), .A2(n6398), .ZN(n7658) );
  OR2_X1 U7532 ( .A1(n5108), .A2(n7658), .ZN(n6400) );
  INV_X1 U7533 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7659) );
  OR2_X1 U7534 ( .A1(n5110), .A2(n7659), .ZN(n6399) );
  NAND4_X1 U7535 ( .A1(n6402), .A2(n6401), .A3(n6400), .A4(n6399), .ZN(n9202)
         );
  OR2_X1 U7536 ( .A1(n10988), .A2(n9202), .ZN(n8739) );
  NAND2_X1 U7537 ( .A1(n9202), .A2(n10988), .ZN(n7732) );
  NAND2_X1 U7538 ( .A1(n8739), .A2(n7732), .ZN(n8865) );
  NAND2_X1 U7539 ( .A1(n7655), .A2(n8865), .ZN(n6404) );
  OR2_X1 U7540 ( .A1(n9202), .A2(n7661), .ZN(n6403) );
  NAND2_X1 U7541 ( .A1(n6404), .A2(n6403), .ZN(n7735) );
  NAND2_X1 U7542 ( .A1(n6307), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6410) );
  INV_X1 U7543 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7698) );
  OR2_X1 U7544 ( .A1(n8680), .A2(n7698), .ZN(n6409) );
  NAND2_X1 U7545 ( .A1(n6405), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6406) );
  AND2_X1 U7546 ( .A1(n6422), .A2(n6406), .ZN(n7739) );
  OR2_X1 U7547 ( .A1(n5108), .A2(n7739), .ZN(n6408) );
  INV_X1 U7548 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7779) );
  OR2_X1 U7549 ( .A1(n5110), .A2(n7779), .ZN(n6407) );
  NAND4_X1 U7550 ( .A1(n6410), .A2(n6409), .A3(n6408), .A4(n6407), .ZN(n9201)
         );
  NAND2_X1 U7551 ( .A1(n6790), .A2(n6416), .ZN(n6413) );
  NAND2_X1 U7552 ( .A1(n6417), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6411) );
  XNOR2_X1 U7553 ( .A(n6411), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7799) );
  AOI22_X1 U7554 ( .A1(n6555), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6554), .B2(
        n7799), .ZN(n6412) );
  OR2_X1 U7555 ( .A1(n7814), .A2(n10997), .ZN(n8732) );
  NAND2_X1 U7556 ( .A1(n7814), .A2(n10997), .ZN(n8740) );
  NAND2_X1 U7557 ( .A1(n8732), .A2(n8740), .ZN(n8863) );
  NAND2_X1 U7558 ( .A1(n7735), .A2(n8863), .ZN(n6415) );
  OR2_X1 U7559 ( .A1(n9201), .A2(n10997), .ZN(n6414) );
  NAND2_X1 U7560 ( .A1(n6415), .A2(n6414), .ZN(n7812) );
  NAND2_X1 U7561 ( .A1(n6796), .A2(n6416), .ZN(n6420) );
  OR2_X1 U7562 ( .A1(n6417), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n6430) );
  NAND2_X1 U7563 ( .A1(n6430), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6418) );
  XNOR2_X1 U7564 ( .A(n6418), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7861) );
  AOI22_X1 U7565 ( .A1(n6555), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6554), .B2(
        n7861), .ZN(n6419) );
  NAND2_X1 U7566 ( .A1(n6307), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6427) );
  INV_X1 U7567 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6421) );
  OR2_X1 U7568 ( .A1(n8680), .A2(n6421), .ZN(n6426) );
  NAND2_X1 U7569 ( .A1(n6422), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6423) );
  AND2_X1 U7570 ( .A1(n6435), .A2(n6423), .ZN(n7817) );
  OR2_X1 U7571 ( .A1(n5108), .A2(n7817), .ZN(n6425) );
  INV_X1 U7572 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7818) );
  NAND2_X1 U7573 ( .A1(n7494), .A2(n7738), .ZN(n8741) );
  NAND2_X1 U7574 ( .A1(n8733), .A2(n8741), .ZN(n8864) );
  NAND2_X1 U7575 ( .A1(n7812), .A2(n8864), .ZN(n6429) );
  OR2_X1 U7576 ( .A1(n7494), .A2(n9200), .ZN(n6428) );
  NAND2_X1 U7577 ( .A1(n6429), .A2(n6428), .ZN(n7943) );
  NAND2_X1 U7578 ( .A1(n6794), .A2(n6416), .ZN(n6433) );
  OAI21_X1 U7579 ( .B1(n6430), .B2(P2_IR_REG_9__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6431) );
  XNOR2_X1 U7580 ( .A(n6431), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7898) );
  AOI22_X1 U7581 ( .A1(n6555), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6554), .B2(
        n7898), .ZN(n6432) );
  NAND2_X1 U7582 ( .A1(n6433), .A2(n6432), .ZN(n11010) );
  NAND2_X1 U7583 ( .A1(n6300), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6440) );
  INV_X1 U7584 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n6434) );
  OR2_X1 U7585 ( .A1(n6518), .A2(n6434), .ZN(n6439) );
  NAND2_X1 U7586 ( .A1(n6435), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6436) );
  AND2_X1 U7587 ( .A1(n6448), .A2(n6436), .ZN(n8638) );
  OR2_X1 U7588 ( .A1(n5108), .A2(n8638), .ZN(n6438) );
  INV_X1 U7589 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7947) );
  OR2_X1 U7590 ( .A1(n5110), .A2(n7947), .ZN(n6437) );
  NAND2_X1 U7591 ( .A1(n11010), .A2(n9199), .ZN(n7939) );
  NAND2_X1 U7592 ( .A1(n7943), .A2(n7939), .ZN(n6441) );
  OR2_X1 U7593 ( .A1(n11010), .A2(n9199), .ZN(n7940) );
  NAND2_X1 U7594 ( .A1(n6441), .A2(n7940), .ZN(n7960) );
  NAND2_X1 U7595 ( .A1(n6801), .A2(n6416), .ZN(n6447) );
  NAND2_X1 U7596 ( .A1(n6442), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6443) );
  MUX2_X1 U7597 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6443), .S(
        P2_IR_REG_11__SCAN_IN), .Z(n6445) );
  INV_X1 U7598 ( .A(n6470), .ZN(n6444) );
  NAND2_X1 U7599 ( .A1(n6445), .A2(n6444), .ZN(n8074) );
  INV_X1 U7600 ( .A(n8074), .ZN(n7895) );
  AOI22_X1 U7601 ( .A1(n6555), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6554), .B2(
        n7895), .ZN(n6446) );
  NAND2_X1 U7602 ( .A1(n6447), .A2(n6446), .ZN(n11016) );
  NAND2_X1 U7603 ( .A1(n8678), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6454) );
  INV_X1 U7604 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7965) );
  OR2_X1 U7605 ( .A1(n5110), .A2(n7965), .ZN(n6453) );
  NAND2_X1 U7606 ( .A1(n6448), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6449) );
  AND2_X1 U7607 ( .A1(n6462), .A2(n6449), .ZN(n7964) );
  OR2_X1 U7608 ( .A1(n5108), .A2(n7964), .ZN(n6452) );
  INV_X1 U7609 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6450) );
  OR2_X1 U7610 ( .A1(n8680), .A2(n6450), .ZN(n6451) );
  NAND4_X1 U7611 ( .A1(n6454), .A2(n6453), .A3(n6452), .A4(n6451), .ZN(n9198)
         );
  NAND2_X1 U7612 ( .A1(n11016), .A2(n9198), .ZN(n6455) );
  NAND2_X1 U7613 ( .A1(n7960), .A2(n6455), .ZN(n6457) );
  OR2_X1 U7614 ( .A1(n11016), .A2(n9198), .ZN(n6456) );
  NAND2_X1 U7615 ( .A1(n6834), .A2(n6416), .ZN(n6460) );
  OR2_X1 U7616 ( .A1(n6470), .A2(n6269), .ZN(n6458) );
  XNOR2_X1 U7617 ( .A(n6458), .B(P2_IR_REG_12__SCAN_IN), .ZN(n9206) );
  AOI22_X1 U7618 ( .A1(n6555), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6554), .B2(
        n9206), .ZN(n6459) );
  NAND2_X1 U7619 ( .A1(n8678), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6467) );
  INV_X1 U7620 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6461) );
  OR2_X1 U7621 ( .A1(n8680), .A2(n6461), .ZN(n6466) );
  NAND2_X1 U7622 ( .A1(n6462), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6463) );
  AND2_X1 U7623 ( .A1(n6475), .A2(n6463), .ZN(n8008) );
  OR2_X1 U7624 ( .A1(n5108), .A2(n8008), .ZN(n6465) );
  INV_X1 U7625 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8068) );
  OR2_X1 U7626 ( .A1(n5110), .A2(n8068), .ZN(n6464) );
  NAND4_X1 U7627 ( .A1(n6467), .A2(n6466), .A3(n6465), .A4(n6464), .ZN(n9578)
         );
  NAND2_X1 U7628 ( .A1(n8018), .A2(n9578), .ZN(n6468) );
  INV_X1 U7629 ( .A(n9574), .ZN(n6484) );
  NAND2_X1 U7630 ( .A1(n6838), .A2(n6416), .ZN(n6473) );
  INV_X1 U7631 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6469) );
  OR2_X1 U7632 ( .A1(n6487), .A2(n6269), .ZN(n6471) );
  XNOR2_X1 U7633 ( .A(n6471), .B(P2_IR_REG_13__SCAN_IN), .ZN(n9226) );
  AOI22_X1 U7634 ( .A1(n6555), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6554), .B2(
        n9226), .ZN(n6472) );
  NAND2_X1 U7635 ( .A1(n6473), .A2(n6472), .ZN(n9581) );
  NAND2_X1 U7636 ( .A1(n8678), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6482) );
  INV_X1 U7637 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6474) );
  OR2_X1 U7638 ( .A1(n8680), .A2(n6474), .ZN(n6481) );
  NAND2_X1 U7639 ( .A1(n6475), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6476) );
  AND2_X1 U7640 ( .A1(n6492), .A2(n6476), .ZN(n9582) );
  OR2_X1 U7641 ( .A1(n5108), .A2(n9582), .ZN(n6480) );
  INV_X1 U7642 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6477) );
  OR2_X1 U7643 ( .A1(n5110), .A2(n6477), .ZN(n6479) );
  NAND4_X1 U7644 ( .A1(n6482), .A2(n6481), .A3(n6480), .A4(n6479), .ZN(n9197)
         );
  OR2_X1 U7645 ( .A1(n9581), .A2(n9561), .ZN(n8770) );
  NAND2_X1 U7646 ( .A1(n9581), .A2(n9561), .ZN(n8769) );
  NAND2_X1 U7647 ( .A1(n6484), .A2(n6483), .ZN(n9573) );
  OR2_X1 U7648 ( .A1(n9581), .A2(n9197), .ZN(n6485) );
  NAND2_X1 U7649 ( .A1(n6863), .A2(n6416), .ZN(n6490) );
  INV_X1 U7650 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6486) );
  NAND2_X1 U7651 ( .A1(n6487), .A2(n6486), .ZN(n6499) );
  NAND2_X1 U7652 ( .A1(n6499), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6488) );
  XNOR2_X1 U7653 ( .A(n6488), .B(P2_IR_REG_14__SCAN_IN), .ZN(n9240) );
  AOI22_X1 U7654 ( .A1(n6555), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6554), .B2(
        n9240), .ZN(n6489) );
  NAND2_X1 U7655 ( .A1(n8678), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6498) );
  INV_X1 U7656 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n6491) );
  OR2_X1 U7657 ( .A1(n8680), .A2(n6491), .ZN(n6497) );
  NAND2_X1 U7658 ( .A1(n6492), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6493) );
  AND2_X1 U7659 ( .A1(n6505), .A2(n6493), .ZN(n9565) );
  OR2_X1 U7660 ( .A1(n5108), .A2(n9565), .ZN(n6496) );
  INV_X1 U7661 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6494) );
  OR2_X1 U7662 ( .A1(n5110), .A2(n6494), .ZN(n6495) );
  NAND4_X1 U7663 ( .A1(n6498), .A2(n6497), .A3(n6496), .A4(n6495), .ZN(n9577)
         );
  NOR2_X1 U7664 ( .A1(n8773), .A2(n9577), .ZN(n6697) );
  NAND2_X1 U7665 ( .A1(n8773), .A2(n9577), .ZN(n8784) );
  NAND2_X1 U7666 ( .A1(n6942), .A2(n6416), .ZN(n6504) );
  INV_X1 U7667 ( .A(n6499), .ZN(n6501) );
  INV_X1 U7668 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6500) );
  NAND2_X1 U7669 ( .A1(n6501), .A2(n6500), .ZN(n6502) );
  XNOR2_X1 U7670 ( .A(n6514), .B(P2_IR_REG_15__SCAN_IN), .ZN(n9263) );
  AOI22_X1 U7671 ( .A1(n6555), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6554), .B2(
        n9263), .ZN(n6503) );
  NAND2_X1 U7672 ( .A1(n8678), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6510) );
  INV_X1 U7673 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9653) );
  OR2_X1 U7674 ( .A1(n8680), .A2(n9653), .ZN(n6509) );
  NAND2_X1 U7675 ( .A1(n6505), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6506) );
  AND2_X1 U7676 ( .A1(n6541), .A2(n6506), .ZN(n9544) );
  OR2_X1 U7677 ( .A1(n5108), .A2(n9544), .ZN(n6508) );
  INV_X1 U7678 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9554) );
  OR2_X1 U7679 ( .A1(n5110), .A2(n9554), .ZN(n6507) );
  NAND4_X1 U7680 ( .A1(n6510), .A2(n6509), .A3(n6508), .A4(n6507), .ZN(n9529)
         );
  OR2_X1 U7681 ( .A1(n9553), .A2(n9563), .ZN(n8776) );
  NAND2_X1 U7682 ( .A1(n9553), .A2(n9563), .ZN(n8777) );
  NAND2_X1 U7683 ( .A1(n9553), .A2(n9529), .ZN(n9481) );
  NAND2_X1 U7684 ( .A1(n7137), .A2(n6416), .ZN(n6516) );
  INV_X1 U7685 ( .A(n6511), .ZN(n6512) );
  NAND2_X1 U7686 ( .A1(n6512), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6513) );
  XNOR2_X1 U7687 ( .A(n6553), .B(n5205), .ZN(n9349) );
  AOI22_X1 U7688 ( .A1(n6555), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6554), .B2(
        n9349), .ZN(n6515) );
  NAND2_X1 U7689 ( .A1(n6531), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6517) );
  NAND2_X1 U7690 ( .A1(n6558), .A2(n6517), .ZN(n9505) );
  NAND2_X1 U7691 ( .A1(n6671), .A2(n9505), .ZN(n6522) );
  INV_X1 U7692 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9641) );
  OR2_X1 U7693 ( .A1(n8680), .A2(n9641), .ZN(n6521) );
  INV_X1 U7694 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9694) );
  OR2_X1 U7695 ( .A1(n6518), .A2(n9694), .ZN(n6520) );
  INV_X1 U7696 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9507) );
  OR2_X1 U7697 ( .A1(n5110), .A2(n9507), .ZN(n6519) );
  NAND4_X1 U7698 ( .A1(n6522), .A2(n6521), .A3(n6520), .A4(n6519), .ZN(n9516)
         );
  OR2_X1 U7699 ( .A1(n9510), .A2(n9516), .ZN(n6568) );
  INV_X1 U7700 ( .A(n6568), .ZN(n6552) );
  NAND2_X1 U7701 ( .A1(n7084), .A2(n6416), .ZN(n6529) );
  NAND2_X1 U7702 ( .A1(n6514), .A2(n6523), .ZN(n6524) );
  NAND2_X1 U7703 ( .A1(n6524), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6538) );
  NAND2_X1 U7704 ( .A1(n6538), .A2(n6525), .ZN(n6526) );
  NAND2_X1 U7705 ( .A1(n6526), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6527) );
  XNOR2_X1 U7706 ( .A(n6527), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9325) );
  AOI22_X1 U7707 ( .A1(n6555), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6554), .B2(
        n9325), .ZN(n6528) );
  NAND2_X1 U7708 ( .A1(n8678), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6535) );
  OR2_X1 U7709 ( .A1(n5110), .A2(n9300), .ZN(n6534) );
  NAND2_X1 U7710 ( .A1(n6543), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6530) );
  AND2_X1 U7711 ( .A1(n6531), .A2(n6530), .ZN(n9522) );
  OR2_X1 U7712 ( .A1(n5108), .A2(n9522), .ZN(n6533) );
  INV_X1 U7713 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9645) );
  OR2_X1 U7714 ( .A1(n8680), .A2(n9645), .ZN(n6532) );
  NAND2_X1 U7715 ( .A1(n9521), .A2(n9530), .ZN(n9499) );
  NAND2_X1 U7716 ( .A1(n9510), .A2(n9516), .ZN(n6536) );
  AND2_X1 U7717 ( .A1(n9499), .A2(n6536), .ZN(n6548) );
  INV_X1 U7718 ( .A(n6548), .ZN(n6537) );
  OR2_X1 U7719 ( .A1(n6537), .A2(n9519), .ZN(n6567) );
  INV_X1 U7720 ( .A(n6567), .ZN(n6550) );
  NAND2_X1 U7721 ( .A1(n7071), .A2(n6416), .ZN(n6540) );
  XNOR2_X1 U7722 ( .A(n6538), .B(P2_IR_REG_16__SCAN_IN), .ZN(n9313) );
  AOI22_X1 U7723 ( .A1(n6555), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6554), .B2(
        n9313), .ZN(n6539) );
  NAND2_X1 U7724 ( .A1(n8678), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6547) );
  INV_X1 U7725 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9649) );
  OR2_X1 U7726 ( .A1(n8680), .A2(n9649), .ZN(n6546) );
  NAND2_X1 U7727 ( .A1(n6541), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6542) );
  AND2_X1 U7728 ( .A1(n6543), .A2(n6542), .ZN(n9538) );
  OR2_X1 U7729 ( .A1(n5108), .A2(n9538), .ZN(n6545) );
  INV_X1 U7730 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n9539) );
  OR2_X1 U7731 ( .A1(n5110), .A2(n9539), .ZN(n6544) );
  NAND4_X1 U7732 ( .A1(n6547), .A2(n6546), .A3(n6545), .A4(n6544), .ZN(n9546)
         );
  NAND2_X1 U7733 ( .A1(n9537), .A2(n9546), .ZN(n9498) );
  AND2_X1 U7734 ( .A1(n9498), .A2(n6548), .ZN(n6549) );
  NAND2_X1 U7735 ( .A1(n7407), .A2(n6416), .ZN(n6557) );
  AOI22_X1 U7736 ( .A1(n6555), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6711), .B2(
        n6554), .ZN(n6556) );
  NAND2_X1 U7737 ( .A1(n6558), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6559) );
  NAND2_X1 U7738 ( .A1(n6575), .A2(n6559), .ZN(n9491) );
  NAND2_X1 U7739 ( .A1(n9491), .A2(n6671), .ZN(n6564) );
  NAND2_X1 U7740 ( .A1(n6300), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6563) );
  NAND2_X1 U7741 ( .A1(n8678), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6562) );
  INV_X1 U7742 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n6560) );
  OR2_X1 U7743 ( .A1(n5110), .A2(n6560), .ZN(n6561) );
  NAND4_X1 U7744 ( .A1(n6564), .A2(n6563), .A3(n6562), .A4(n6561), .ZN(n9196)
         );
  AND2_X1 U7745 ( .A1(n9481), .A2(n6566), .ZN(n6565) );
  NAND2_X1 U7746 ( .A1(n9480), .A2(n6565), .ZN(n6572) );
  INV_X1 U7747 ( .A(n6566), .ZN(n6570) );
  NAND2_X1 U7748 ( .A1(n9537), .A2(n9037), .ZN(n8788) );
  NAND2_X1 U7749 ( .A1(n8787), .A2(n8788), .ZN(n9536) );
  AND2_X1 U7750 ( .A1(n9536), .A2(n6567), .ZN(n6569) );
  AND2_X1 U7751 ( .A1(n6569), .A2(n6568), .ZN(n9482) );
  NAND2_X1 U7752 ( .A1(n6572), .A2(n6571), .ZN(n9468) );
  NAND2_X1 U7753 ( .A1(n7534), .A2(n6416), .ZN(n6574) );
  OR2_X1 U7754 ( .A1(n6360), .A2(n7555), .ZN(n6573) );
  XNOR2_X1 U7755 ( .A(n6575), .B(P2_REG3_REG_20__SCAN_IN), .ZN(n9475) );
  NAND2_X1 U7756 ( .A1(n9475), .A2(n6671), .ZN(n6581) );
  INV_X1 U7757 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n6578) );
  NAND2_X1 U7758 ( .A1(n6300), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6577) );
  NAND2_X1 U7759 ( .A1(n8678), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6576) );
  OAI211_X1 U7760 ( .C1(n6578), .C2(n5110), .A(n6577), .B(n6576), .ZN(n6579)
         );
  INV_X1 U7761 ( .A(n6579), .ZN(n6580) );
  NAND2_X1 U7762 ( .A1(n6581), .A2(n6580), .ZN(n9195) );
  XNOR2_X1 U7763 ( .A(n9474), .B(n9488), .ZN(n9473) );
  NAND2_X1 U7764 ( .A1(n9468), .A2(n9473), .ZN(n6583) );
  OR2_X1 U7765 ( .A1(n9474), .A2(n9195), .ZN(n6582) );
  NAND2_X1 U7766 ( .A1(n6583), .A2(n6582), .ZN(n9458) );
  NAND2_X1 U7767 ( .A1(n7595), .A2(n6416), .ZN(n6585) );
  INV_X1 U7768 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7635) );
  OR2_X1 U7769 ( .A1(n6360), .A2(n7635), .ZN(n6584) );
  INV_X1 U7770 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n6591) );
  INV_X1 U7771 ( .A(n6586), .ZN(n6587) );
  NAND2_X1 U7772 ( .A1(n6587), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6588) );
  NAND2_X1 U7773 ( .A1(n6595), .A2(n6588), .ZN(n9463) );
  NAND2_X1 U7774 ( .A1(n9463), .A2(n6671), .ZN(n6590) );
  AOI22_X1 U7775 ( .A1(n8678), .A2(P2_REG0_REG_21__SCAN_IN), .B1(n6300), .B2(
        P2_REG1_REG_21__SCAN_IN), .ZN(n6589) );
  OAI211_X1 U7776 ( .C1(n5110), .C2(n6591), .A(n6590), .B(n6589), .ZN(n9447)
         );
  INV_X1 U7777 ( .A(n9447), .ZN(n9471) );
  XNOR2_X1 U7778 ( .A(n9105), .B(n9471), .ZN(n9462) );
  NAND2_X1 U7779 ( .A1(n9458), .A2(n9462), .ZN(n6592) );
  OR2_X1 U7780 ( .A1(n9105), .A2(n9447), .ZN(n8812) );
  NAND2_X1 U7781 ( .A1(n6592), .A2(n8812), .ZN(n9446) );
  NAND2_X1 U7782 ( .A1(n7664), .A2(n6416), .ZN(n6594) );
  OR2_X1 U7783 ( .A1(n6360), .A2(n7668), .ZN(n6593) );
  NAND2_X1 U7784 ( .A1(n6595), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6596) );
  NAND2_X1 U7785 ( .A1(n6605), .A2(n6596), .ZN(n9452) );
  INV_X1 U7786 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n6599) );
  NAND2_X1 U7787 ( .A1(n8678), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6598) );
  NAND2_X1 U7788 ( .A1(n6300), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6597) );
  OAI211_X1 U7789 ( .C1(n5110), .C2(n6599), .A(n6598), .B(n6597), .ZN(n6600)
         );
  AOI21_X1 U7790 ( .B1(n9452), .B2(n6671), .A(n6600), .ZN(n9460) );
  NAND2_X1 U7791 ( .A1(n9622), .A2(n9460), .ZN(n8821) );
  NAND2_X1 U7792 ( .A1(n8822), .A2(n8821), .ZN(n9451) );
  NAND2_X1 U7793 ( .A1(n9446), .A2(n9451), .ZN(n6602) );
  OR2_X1 U7794 ( .A1(n9622), .A2(n9047), .ZN(n6601) );
  NAND2_X1 U7795 ( .A1(n7776), .A2(n6416), .ZN(n6604) );
  OR2_X1 U7796 ( .A1(n6360), .A2(n7778), .ZN(n6603) );
  NAND2_X1 U7797 ( .A1(n6605), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6606) );
  NAND2_X1 U7798 ( .A1(n6617), .A2(n6606), .ZN(n9441) );
  NAND2_X1 U7799 ( .A1(n9441), .A2(n6671), .ZN(n6612) );
  INV_X1 U7800 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n6609) );
  NAND2_X1 U7801 ( .A1(n6300), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6608) );
  NAND2_X1 U7802 ( .A1(n8678), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6607) );
  OAI211_X1 U7803 ( .C1(n6609), .C2(n5110), .A(n6608), .B(n6607), .ZN(n6610)
         );
  INV_X1 U7804 ( .A(n6610), .ZN(n6611) );
  NOR2_X1 U7805 ( .A1(n9440), .A2(n9448), .ZN(n6614) );
  NAND2_X1 U7806 ( .A1(n9440), .A2(n9448), .ZN(n6613) );
  OAI21_X2 U7807 ( .B1(n9435), .B2(n6614), .A(n6613), .ZN(n9423) );
  NAND2_X1 U7808 ( .A1(n7958), .A2(n6416), .ZN(n6616) );
  OR2_X1 U7809 ( .A1(n6360), .A2(n8059), .ZN(n6615) );
  NAND2_X1 U7810 ( .A1(n6617), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6618) );
  NAND2_X1 U7811 ( .A1(n6628), .A2(n6618), .ZN(n9428) );
  NAND2_X1 U7812 ( .A1(n9428), .A2(n6671), .ZN(n6624) );
  INV_X1 U7813 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6621) );
  NAND2_X1 U7814 ( .A1(n6300), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6620) );
  NAND2_X1 U7815 ( .A1(n8678), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6619) );
  OAI211_X1 U7816 ( .C1(n6621), .C2(n5110), .A(n6620), .B(n6619), .ZN(n6622)
         );
  INV_X1 U7817 ( .A(n6622), .ZN(n6623) );
  NAND2_X1 U7818 ( .A1(n6624), .A2(n6623), .ZN(n9194) );
  AND2_X1 U7819 ( .A1(n9421), .A2(n9194), .ZN(n6625) );
  NAND2_X1 U7820 ( .A1(n8042), .A2(n6416), .ZN(n6627) );
  OR2_X1 U7821 ( .A1(n6360), .A2(n8617), .ZN(n6626) );
  NAND2_X1 U7822 ( .A1(n6628), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6629) );
  NAND2_X1 U7823 ( .A1(n6639), .A2(n6629), .ZN(n9418) );
  NAND2_X1 U7824 ( .A1(n9418), .A2(n6671), .ZN(n6635) );
  INV_X1 U7825 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n6632) );
  NAND2_X1 U7826 ( .A1(n6300), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6631) );
  NAND2_X1 U7827 ( .A1(n8678), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6630) );
  OAI211_X1 U7828 ( .C1(n6632), .C2(n5110), .A(n6631), .B(n6630), .ZN(n6633)
         );
  INV_X1 U7829 ( .A(n6633), .ZN(n6634) );
  NAND2_X1 U7830 ( .A1(n9411), .A2(n9398), .ZN(n6636) );
  OR2_X1 U7831 ( .A1(n6360), .A2(n8133), .ZN(n6637) );
  INV_X1 U7832 ( .A(n6639), .ZN(n6640) );
  INV_X1 U7833 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9169) );
  INV_X1 U7834 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8454) );
  NAND2_X1 U7835 ( .A1(n6641), .A2(n8454), .ZN(n6652) );
  INV_X1 U7836 ( .A(n6641), .ZN(n6642) );
  NAND2_X1 U7837 ( .A1(n6642), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6643) );
  NAND2_X1 U7838 ( .A1(n6652), .A2(n6643), .ZN(n9389) );
  NAND2_X1 U7839 ( .A1(n9389), .A2(n6671), .ZN(n6649) );
  INV_X1 U7840 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n6646) );
  NAND2_X1 U7841 ( .A1(n8678), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6645) );
  NAND2_X1 U7842 ( .A1(n6300), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6644) );
  OAI211_X1 U7843 ( .C1(n6646), .C2(n5110), .A(n6645), .B(n6644), .ZN(n6647)
         );
  INV_X1 U7844 ( .A(n6647), .ZN(n6648) );
  NAND2_X1 U7845 ( .A1(n8609), .A2(n6416), .ZN(n6651) );
  INV_X1 U7846 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8612) );
  OR2_X1 U7847 ( .A1(n6360), .A2(n8612), .ZN(n6650) );
  NAND2_X1 U7848 ( .A1(n6652), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6653) );
  NAND2_X1 U7849 ( .A1(n6670), .A2(n6653), .ZN(n9372) );
  NAND2_X1 U7850 ( .A1(n9372), .A2(n6671), .ZN(n6659) );
  INV_X1 U7851 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n6656) );
  NAND2_X1 U7852 ( .A1(n6300), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6655) );
  NAND2_X1 U7853 ( .A1(n8678), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6654) );
  OAI211_X1 U7854 ( .C1(n6656), .C2(n5110), .A(n6655), .B(n6654), .ZN(n6657)
         );
  INV_X1 U7855 ( .A(n6657), .ZN(n6658) );
  NAND2_X1 U7856 ( .A1(n6660), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6661) );
  XNOR2_X1 U7857 ( .A(n6661), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8897) );
  NAND2_X1 U7858 ( .A1(n6711), .A2(n8897), .ZN(n6758) );
  NAND2_X1 U7859 ( .A1(n5127), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6663) );
  XNOR2_X1 U7860 ( .A(n6663), .B(n6662), .ZN(n8879) );
  INV_X1 U7861 ( .A(n6664), .ZN(n6665) );
  NAND2_X1 U7862 ( .A1(n6665), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6666) );
  MUX2_X1 U7863 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6666), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n6667) );
  NAND2_X1 U7864 ( .A1(n6667), .A2(n5127), .ZN(n8849) );
  OR2_X1 U7865 ( .A1(n8879), .A2(n8849), .ZN(n8676) );
  INV_X1 U7866 ( .A(n6668), .ZN(n8894) );
  XNOR2_X1 U7867 ( .A(n8894), .B(n6859), .ZN(n6960) );
  INV_X1 U7868 ( .A(n8879), .ZN(n6947) );
  AND2_X2 U7869 ( .A1(n8897), .A2(n6947), .ZN(n8836) );
  NAND2_X1 U7870 ( .A1(n9023), .A2(n6671), .ZN(n8686) );
  INV_X1 U7871 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n9024) );
  NAND2_X1 U7872 ( .A1(n8678), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6673) );
  NAND2_X1 U7873 ( .A1(n6300), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6672) );
  OAI211_X1 U7874 ( .C1(n9024), .C2(n5110), .A(n6673), .B(n6672), .ZN(n6674)
         );
  INV_X1 U7875 ( .A(n6674), .ZN(n6675) );
  NAND2_X1 U7876 ( .A1(n8686), .A2(n6675), .ZN(n9193) );
  OAI21_X2 U7877 ( .B1(n6679), .B2(n9559), .A(n6678), .ZN(n9371) );
  INV_X1 U7878 ( .A(n6680), .ZN(n6949) );
  OR2_X1 U7879 ( .A1(n6912), .A2(n6949), .ZN(n8699) );
  INV_X1 U7880 ( .A(n8699), .ZN(n6682) );
  NAND2_X1 U7881 ( .A1(n6682), .A2(n6681), .ZN(n7141) );
  NAND2_X1 U7882 ( .A1(n7141), .A2(n6683), .ZN(n7212) );
  INV_X1 U7883 ( .A(n7202), .ZN(n8859) );
  NAND2_X1 U7884 ( .A1(n7212), .A2(n8859), .ZN(n10930) );
  INV_X1 U7885 ( .A(n10933), .ZN(n10938) );
  OR2_X1 U7886 ( .A1(n10925), .A2(n7206), .ZN(n10929) );
  AND2_X1 U7887 ( .A1(n8721), .A2(n10929), .ZN(n7386) );
  AND2_X1 U7888 ( .A1(n7156), .A2(n10951), .ZN(n6684) );
  INV_X1 U7889 ( .A(n6684), .ZN(n8717) );
  AND2_X1 U7890 ( .A1(n7386), .A2(n8717), .ZN(n6686) );
  OR2_X1 U7891 ( .A1(n7156), .A2(n10951), .ZN(n7508) );
  NAND2_X1 U7892 ( .A1(n7171), .A2(n10961), .ZN(n8719) );
  AND2_X1 U7893 ( .A1(n7508), .A2(n8719), .ZN(n8722) );
  NAND2_X1 U7894 ( .A1(n7509), .A2(n8722), .ZN(n7578) );
  OR2_X1 U7895 ( .A1(n7171), .A2(n10961), .ZN(n8725) );
  NAND2_X1 U7896 ( .A1(n7578), .A2(n8725), .ZN(n6687) );
  INV_X1 U7897 ( .A(n7577), .ZN(n8861) );
  INV_X1 U7898 ( .A(n8745), .ZN(n7652) );
  NOR2_X1 U7899 ( .A1(n8865), .A2(n7652), .ZN(n6688) );
  AND2_X1 U7900 ( .A1(n8732), .A2(n7732), .ZN(n8751) );
  NAND2_X1 U7901 ( .A1(n7733), .A2(n8751), .ZN(n6689) );
  NAND2_X1 U7902 ( .A1(n11010), .A2(n7962), .ZN(n8753) );
  INV_X1 U7903 ( .A(n8753), .ZN(n6690) );
  OR2_X1 U7904 ( .A1(n11010), .A2(n7962), .ZN(n8757) );
  AND2_X1 U7905 ( .A1(n8757), .A2(n8733), .ZN(n8750) );
  INV_X1 U7906 ( .A(n9198), .ZN(n8635) );
  OR2_X1 U7907 ( .A1(n11016), .A2(n8635), .ZN(n8758) );
  NAND2_X1 U7908 ( .A1(n11016), .A2(n8635), .ZN(n8759) );
  INV_X1 U7909 ( .A(n9578), .ZN(n7963) );
  OR2_X1 U7910 ( .A1(n8018), .A2(n7963), .ZN(n8766) );
  AND2_X1 U7911 ( .A1(n8869), .A2(n8766), .ZN(n6691) );
  NAND2_X1 U7912 ( .A1(n8018), .A2(n7963), .ZN(n8765) );
  INV_X1 U7913 ( .A(n8766), .ZN(n6692) );
  OR2_X1 U7914 ( .A1(n6692), .A2(n8759), .ZN(n6693) );
  AND2_X1 U7915 ( .A1(n8765), .A2(n6693), .ZN(n6694) );
  NAND2_X1 U7916 ( .A1(n6695), .A2(n6694), .ZN(n9586) );
  NAND2_X1 U7917 ( .A1(n9586), .A2(n9585), .ZN(n6696) );
  INV_X1 U7918 ( .A(n6697), .ZN(n6698) );
  INV_X1 U7919 ( .A(n9577), .ZN(n9179) );
  OR2_X1 U7920 ( .A1(n8773), .A2(n9179), .ZN(n6700) );
  INV_X1 U7921 ( .A(n9519), .ZN(n8872) );
  OR2_X1 U7922 ( .A1(n9521), .A2(n9503), .ZN(n6702) );
  NAND2_X1 U7923 ( .A1(n6703), .A2(n6702), .ZN(n9497) );
  NAND2_X1 U7924 ( .A1(n9510), .A2(n9487), .ZN(n8801) );
  INV_X1 U7925 ( .A(n9196), .ZN(n9504) );
  OR2_X1 U7926 ( .A1(n9092), .A2(n9504), .ZN(n8805) );
  INV_X1 U7927 ( .A(n9473), .ZN(n9469) );
  NAND2_X1 U7928 ( .A1(n9472), .A2(n9469), .ZN(n6705) );
  OR2_X1 U7929 ( .A1(n9474), .A2(n9488), .ZN(n6704) );
  NAND2_X1 U7930 ( .A1(n6705), .A2(n6704), .ZN(n9461) );
  INV_X1 U7931 ( .A(n9462), .ZN(n9457) );
  NAND2_X1 U7932 ( .A1(n9461), .A2(n9457), .ZN(n6707) );
  OR2_X1 U7933 ( .A1(n9105), .A2(n9471), .ZN(n6706) );
  NAND2_X1 U7934 ( .A1(n6707), .A2(n6706), .ZN(n9450) );
  NOR2_X1 U7935 ( .A1(n9440), .A2(n9426), .ZN(n8826) );
  XNOR2_X1 U7936 ( .A(n9421), .B(n9437), .ZN(n9422) );
  INV_X1 U7937 ( .A(n9422), .ZN(n6708) );
  NAND2_X1 U7938 ( .A1(n9440), .A2(n9426), .ZN(n9429) );
  OR2_X1 U7939 ( .A1(n9421), .A2(n9437), .ZN(n8696) );
  NAND2_X1 U7940 ( .A1(n6709), .A2(n8696), .ZN(n9410) );
  NOR2_X1 U7941 ( .A1(n9411), .A2(n9425), .ZN(n8830) );
  INV_X1 U7942 ( .A(n8830), .ZN(n6710) );
  NAND2_X1 U7943 ( .A1(n9406), .A2(n9415), .ZN(n8694) );
  NAND2_X1 U7944 ( .A1(n9386), .A2(n8838), .ZN(n8670) );
  XOR2_X1 U7945 ( .A(n9067), .B(n8670), .Z(n9376) );
  NOR2_X1 U7946 ( .A1(n7207), .A2(n8897), .ZN(n9594) );
  INV_X1 U7947 ( .A(n9594), .ZN(n11006) );
  INV_X1 U7948 ( .A(n6711), .ZN(n8892) );
  AND2_X1 U7949 ( .A1(n8892), .A2(n8849), .ZN(n6748) );
  INV_X1 U7950 ( .A(n8897), .ZN(n7666) );
  NAND2_X1 U7951 ( .A1(n7666), .A2(n8879), .ZN(n11093) );
  OAI21_X1 U7952 ( .B1(n8897), .B2(n8849), .A(n11093), .ZN(n6712) );
  NAND2_X1 U7953 ( .A1(n11006), .A2(n9021), .ZN(n11097) );
  NOR2_X1 U7954 ( .A1(n9371), .A2(n6713), .ZN(n6764) );
  NAND2_X1 U7955 ( .A1(n6714), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6716) );
  INV_X1 U7956 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6715) );
  NAND2_X1 U7957 ( .A1(n6716), .A2(n6715), .ZN(n6718) );
  XNOR2_X1 U7958 ( .A(n8058), .B(P2_B_REG_SCAN_IN), .ZN(n6721) );
  NAND2_X1 U7959 ( .A1(n6718), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6720) );
  INV_X1 U7960 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6719) );
  NAND2_X1 U7961 ( .A1(n6721), .A2(n8615), .ZN(n6726) );
  NAND2_X1 U7962 ( .A1(n6722), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6723) );
  MUX2_X1 U7963 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6723), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6725) );
  AND2_X1 U7964 ( .A1(n6725), .A2(n6724), .ZN(n6733) );
  NAND2_X1 U7965 ( .A1(n6726), .A2(n6733), .ZN(n6728) );
  INV_X1 U7966 ( .A(n6733), .ZN(n8104) );
  NAND2_X1 U7967 ( .A1(n8104), .A2(n8058), .ZN(n6810) );
  OR2_X1 U7968 ( .A1(n6728), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6729) );
  NAND2_X1 U7969 ( .A1(n8615), .A2(n8104), .ZN(n6813) );
  NAND2_X1 U7970 ( .A1(n6729), .A2(n6813), .ZN(n6923) );
  INV_X1 U7971 ( .A(n6923), .ZN(n6730) );
  AND2_X1 U7972 ( .A1(n6946), .A2(n6730), .ZN(n6757) );
  INV_X1 U7973 ( .A(n8615), .ZN(n6732) );
  INV_X1 U7974 ( .A(n8058), .ZN(n6731) );
  NAND3_X1 U7975 ( .A1(n6733), .A2(n6732), .A3(n6731), .ZN(n6900) );
  NAND2_X1 U7976 ( .A1(n5177), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6735) );
  INV_X1 U7977 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6734) );
  XNOR2_X1 U7978 ( .A(n6735), .B(n6734), .ZN(n6820) );
  AND2_X1 U7979 ( .A1(n6820), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6904) );
  NOR2_X1 U7980 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6739) );
  NOR4_X1 U7981 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6738) );
  NOR4_X1 U7982 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6737) );
  NOR4_X1 U7983 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6736) );
  NAND4_X1 U7984 ( .A1(n6739), .A2(n6738), .A3(n6737), .A4(n6736), .ZN(n6745)
         );
  NOR4_X1 U7985 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6743) );
  NOR4_X1 U7986 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6742) );
  NOR4_X1 U7987 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6741) );
  NOR4_X1 U7988 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6740) );
  NAND4_X1 U7989 ( .A1(n6743), .A2(n6742), .A3(n6741), .A4(n6740), .ZN(n6744)
         );
  NOR2_X1 U7990 ( .A1(n6745), .A2(n6744), .ZN(n6746) );
  OR2_X1 U7991 ( .A1(n6728), .A2(n6746), .ZN(n6759) );
  NAND2_X1 U7992 ( .A1(n6908), .A2(n6759), .ZN(n6747) );
  NOR2_X1 U7993 ( .A1(n6757), .A2(n6747), .ZN(n6927) );
  OAI21_X1 U7994 ( .B1(n7207), .B2(n11093), .A(n6946), .ZN(n6751) );
  INV_X1 U7995 ( .A(n6748), .ZN(n6749) );
  NAND2_X1 U7996 ( .A1(n6749), .A2(n8836), .ZN(n6899) );
  OR3_X1 U7997 ( .A1(n6711), .A2(n8849), .A3(n7666), .ZN(n6750) );
  NAND2_X1 U7998 ( .A1(n6750), .A2(n8847), .ZN(n6924) );
  NAND2_X1 U7999 ( .A1(n6899), .A2(n6924), .ZN(n6922) );
  AOI22_X1 U8000 ( .A1(n6751), .A2(n6922), .B1(n6923), .B2(n6924), .ZN(n6752)
         );
  AND2_X2 U8001 ( .A1(n6927), .A2(n6752), .ZN(n11100) );
  MUX2_X1 U8002 ( .A(n6753), .B(n6764), .S(n11100), .Z(n6756) );
  INV_X1 U8003 ( .A(n9072), .ZN(n9374) );
  NAND2_X1 U8004 ( .A1(n11100), .A2(n11017), .ZN(n9655) );
  NAND2_X1 U8005 ( .A1(n9072), .A2(n6754), .ZN(n6755) );
  NAND2_X1 U8006 ( .A1(n6756), .A2(n6755), .ZN(P2_U3487) );
  INV_X1 U8007 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6765) );
  NAND2_X1 U8008 ( .A1(n6757), .A2(n6759), .ZN(n6915) );
  OR3_X1 U8009 ( .A1(n6758), .A2(n6947), .A3(n8849), .ZN(n6906) );
  INV_X1 U8010 ( .A(n6906), .ZN(n6898) );
  NOR2_X1 U8011 ( .A1(n6928), .A2(n6898), .ZN(n6763) );
  INV_X1 U8012 ( .A(n6946), .ZN(n6925) );
  NAND3_X1 U8013 ( .A1(n6925), .A2(n6923), .A3(n6759), .ZN(n6914) );
  INV_X1 U8014 ( .A(n6914), .ZN(n6761) );
  AND2_X1 U8015 ( .A1(n8847), .A2(n11093), .ZN(n6905) );
  NAND2_X1 U8016 ( .A1(n6906), .A2(n6905), .ZN(n6760) );
  NAND2_X1 U8017 ( .A1(n7207), .A2(n11017), .ZN(n9583) );
  NAND2_X1 U8018 ( .A1(n6760), .A2(n9583), .ZN(n6897) );
  NAND2_X1 U8019 ( .A1(n6761), .A2(n6897), .ZN(n6762) );
  OAI21_X1 U8020 ( .B1(n6915), .B2(n6763), .A(n6762), .ZN(n6766) );
  AND2_X2 U8021 ( .A1(n6766), .A2(n6908), .ZN(n11104) );
  MUX2_X1 U8022 ( .A(n6765), .B(n6764), .S(n11104), .Z(n6769) );
  AND2_X1 U8023 ( .A1(n6908), .A2(n11017), .ZN(n6917) );
  NAND2_X1 U8024 ( .A1(n6766), .A2(n6917), .ZN(n9708) );
  INV_X1 U8025 ( .A(n9708), .ZN(n6767) );
  NAND2_X1 U8026 ( .A1(n9072), .A2(n6767), .ZN(n6768) );
  NAND2_X1 U8027 ( .A1(n6769), .A2(n6768), .ZN(P2_U3455) );
  NOR2_X1 U8028 ( .A1(n7032), .A2(P1_U3086), .ZN(n6770) );
  AND2_X2 U8029 ( .A1(n6770), .A2(n7743), .ZN(P1_U3973) );
  INV_X1 U8030 ( .A(n6820), .ZN(n7074) );
  OR2_X1 U8031 ( .A1(n6900), .A2(n7074), .ZN(n6825) );
  NOR2_X2 U8032 ( .A1(n6825), .A2(P2_U3151), .ZN(P2_U3893) );
  OAI222_X1 U8033 ( .A1(P2_U3151), .A2(n6868), .B1(n9719), .B2(n6777), .C1(
        n5609), .C2(n8618), .ZN(P2_U3294) );
  OAI222_X1 U8034 ( .A1(P2_U3151), .A2(n7338), .B1(n9719), .B2(n6773), .C1(
        n8618), .C2(n6346), .ZN(P2_U3291) );
  OAI222_X1 U8035 ( .A1(P2_U3151), .A2(n7339), .B1(n9719), .B2(n6775), .C1(
        n6771), .C2(n8618), .ZN(P2_U3293) );
  NAND2_X1 U8036 ( .A1(n6772), .A2(P1_U3086), .ZN(n10595) );
  OAI222_X1 U8037 ( .A1(n10217), .A2(P1_U3086), .B1(n8657), .B2(n6773), .C1(
        n10595), .C2(n5411), .ZN(P1_U3351) );
  OAI222_X1 U8038 ( .A1(n6989), .A2(P1_U3086), .B1(n8657), .B2(n6775), .C1(
        n6774), .C2(n10595), .ZN(P1_U3353) );
  OAI222_X1 U8039 ( .A1(n6990), .A2(P1_U3086), .B1(n8657), .B2(n6777), .C1(
        n6776), .C2(n10595), .ZN(P1_U3354) );
  OAI222_X1 U8040 ( .A1(n6993), .A2(P1_U3086), .B1(n8657), .B2(n6780), .C1(
        n6778), .C2(n10595), .ZN(P1_U3352) );
  INV_X1 U8041 ( .A(n10595), .ZN(n7744) );
  AOI22_X1 U8042 ( .A1(n10242), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n7744), .ZN(n6779) );
  OAI21_X1 U8043 ( .B1(n6783), .B2(n8657), .A(n6779), .ZN(P1_U3350) );
  OAI222_X1 U8044 ( .A1(n8618), .A2(n6781), .B1(n9719), .B2(n6780), .C1(
        P2_U3151), .C2(n7359), .ZN(P2_U3292) );
  OAI222_X1 U8045 ( .A1(n8618), .A2(n6782), .B1(n9719), .B2(n6785), .C1(
        P2_U3151), .C2(n7557), .ZN(P2_U3289) );
  OAI222_X1 U8046 ( .A1(n8618), .A2(n5627), .B1(n9719), .B2(n6783), .C1(
        P2_U3151), .C2(n7353), .ZN(P2_U3290) );
  AOI22_X1 U8047 ( .A1(n10253), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n7744), .ZN(n6784) );
  OAI21_X1 U8048 ( .B1(n6785), .B2(n8657), .A(n6784), .ZN(P1_U3349) );
  INV_X1 U8049 ( .A(n6786), .ZN(n6788) );
  AOI22_X1 U8050 ( .A1(n10678), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n7744), .ZN(n6787) );
  OAI21_X1 U8051 ( .B1(n6788), .B2(n8657), .A(n6787), .ZN(P1_U3348) );
  OAI222_X1 U8052 ( .A1(n8618), .A2(n6789), .B1(n9719), .B2(n6788), .C1(
        P2_U3151), .C2(n7690), .ZN(P2_U3288) );
  INV_X1 U8053 ( .A(n6790), .ZN(n6792) );
  AOI22_X1 U8054 ( .A1(n10692), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n7744), .ZN(n6791) );
  OAI21_X1 U8055 ( .B1(n6792), .B2(n8657), .A(n6791), .ZN(P1_U3347) );
  NAND2_X1 U8056 ( .A1(n6908), .A2(n6728), .ZN(n6809) );
  AND2_X1 U8057 ( .A1(n6809), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8058 ( .A1(n6809), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8059 ( .A1(n6809), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8060 ( .A1(n6809), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8061 ( .A1(n6809), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8062 ( .A1(n6809), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8063 ( .A1(n6809), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8064 ( .A1(n6809), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8065 ( .A1(n6809), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8066 ( .A1(n6809), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8067 ( .A1(n6809), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8068 ( .A1(n6809), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8069 ( .A1(n6809), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  INV_X1 U8070 ( .A(n7799), .ZN(n7695) );
  OAI222_X1 U8071 ( .A1(n8618), .A2(n6793), .B1(n9719), .B2(n6792), .C1(
        P2_U3151), .C2(n7695), .ZN(P2_U3287) );
  INV_X1 U8072 ( .A(n6794), .ZN(n6799) );
  AOI22_X1 U8073 ( .A1(n10774), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n7744), .ZN(n6795) );
  OAI21_X1 U8074 ( .B1(n6799), .B2(n8657), .A(n6795), .ZN(P1_U3345) );
  INV_X1 U8075 ( .A(n10798), .ZN(n7004) );
  INV_X1 U8076 ( .A(n6796), .ZN(n6797) );
  OAI222_X1 U8077 ( .A1(P1_U3086), .A2(n7004), .B1(n8657), .B2(n6797), .C1(
        n8539), .C2(n10595), .ZN(P1_U3346) );
  INV_X1 U8078 ( .A(n7861), .ZN(n7800) );
  OAI222_X1 U8079 ( .A1(n8618), .A2(n6798), .B1(n9719), .B2(n6797), .C1(n7800), 
        .C2(P2_U3151), .ZN(P2_U3286) );
  INV_X1 U8080 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6800) );
  INV_X1 U8081 ( .A(n7898), .ZN(n7806) );
  OAI222_X1 U8082 ( .A1(n8618), .A2(n6800), .B1(n9719), .B2(n6799), .C1(n7806), 
        .C2(P2_U3151), .ZN(P2_U3285) );
  INV_X1 U8083 ( .A(n6801), .ZN(n6807) );
  AOI22_X1 U8084 ( .A1(n10709), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n7744), .ZN(n6802) );
  OAI21_X1 U8085 ( .B1(n6807), .B2(n8657), .A(n6802), .ZN(P1_U3344) );
  NAND2_X1 U8086 ( .A1(n10138), .A2(n7743), .ZN(n6804) );
  NAND2_X1 U8087 ( .A1(n6804), .A2(n6803), .ZN(n6969) );
  INV_X1 U8088 ( .A(n6969), .ZN(n6806) );
  INV_X1 U8089 ( .A(n7743), .ZN(n6805) );
  OAI21_X1 U8090 ( .B1(n6805), .B2(n7032), .A(P1_STATE_REG_SCAN_IN), .ZN(n6970) );
  INV_X1 U8091 ( .A(n10808), .ZN(n10666) );
  NOR2_X1 U8092 ( .A1(n10666), .A2(P1_U3973), .ZN(P1_U3085) );
  OAI222_X1 U8093 ( .A1(n8618), .A2(n6808), .B1(n9719), .B2(n6807), .C1(
        P2_U3151), .C2(n8074), .ZN(P2_U3284) );
  INV_X1 U8094 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6812) );
  INV_X1 U8095 ( .A(n6810), .ZN(n6811) );
  AOI22_X1 U8096 ( .A1(n6809), .A2(n6812), .B1(n6811), .B2(n6904), .ZN(
        P2_U3376) );
  INV_X1 U8097 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6815) );
  INV_X1 U8098 ( .A(n6813), .ZN(n6814) );
  AOI22_X1 U8099 ( .A1(n6809), .A2(n6815), .B1(n6814), .B2(n6904), .ZN(
        P2_U3377) );
  AND2_X1 U8100 ( .A1(n6809), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8101 ( .A1(n6809), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8102 ( .A1(n6809), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8103 ( .A1(n6809), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8104 ( .A1(n6809), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8105 ( .A1(n6809), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8106 ( .A1(n6809), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8107 ( .A1(n6809), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8108 ( .A1(n6809), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8109 ( .A1(n6809), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8110 ( .A1(n6809), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8111 ( .A1(n6809), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8112 ( .A1(n6809), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8113 ( .A1(n6809), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8114 ( .A1(n6809), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8115 ( .A1(n6809), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8116 ( .A1(n6809), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  NAND2_X1 U8117 ( .A1(P1_U3973), .A2(n9745), .ZN(n6816) );
  OAI21_X1 U8118 ( .B1(P1_U3973), .B2(n6346), .A(n6816), .ZN(P1_U3558) );
  INV_X1 U8119 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6818) );
  NAND2_X1 U8120 ( .A1(P1_U3973), .A2(n9906), .ZN(n6817) );
  OAI21_X1 U8121 ( .B1(P1_U3973), .B2(n6818), .A(n6817), .ZN(P1_U3554) );
  NAND2_X1 U8122 ( .A1(n7154), .A2(P2_U3893), .ZN(n6819) );
  OAI21_X1 U8123 ( .B1(P2_U3893), .B2(n5411), .A(n6819), .ZN(P2_U3495) );
  NAND2_X1 U8124 ( .A1(n8836), .A2(n6820), .ZN(n6821) );
  NAND2_X1 U8125 ( .A1(n6825), .A2(n6821), .ZN(n6827) );
  INV_X1 U8126 ( .A(n6827), .ZN(n6822) );
  NAND2_X1 U8127 ( .A1(n6822), .A2(n6313), .ZN(n6823) );
  NAND2_X1 U8128 ( .A1(n6823), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  OR2_X1 U8129 ( .A1(n9327), .A2(P2_U3151), .ZN(n8131) );
  NOR2_X1 U8130 ( .A1(n6827), .A2(n8131), .ZN(n6824) );
  MUX2_X1 U8131 ( .A(n6824), .B(P2_U3893), .S(n8894), .Z(n10848) );
  INV_X1 U8132 ( .A(P2_U3150), .ZN(n6826) );
  NAND2_X1 U8133 ( .A1(n6826), .A2(n6825), .ZN(n10843) );
  INV_X1 U8134 ( .A(n10843), .ZN(n10858) );
  AND2_X1 U8135 ( .A1(P2_U3893), .A2(n6668), .ZN(n10859) );
  OR2_X1 U8136 ( .A1(n6668), .A2(P2_U3151), .ZN(n8610) );
  NOR2_X1 U8137 ( .A1(n6827), .A2(n8610), .ZN(n6848) );
  MUX2_X1 U8138 ( .A(n6933), .B(n6828), .S(n9327), .Z(n6829) );
  NAND2_X1 U8139 ( .A1(n6829), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6870) );
  OAI21_X1 U8140 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n6829), .A(n6870), .ZN(n6830) );
  OAI21_X1 U8141 ( .B1(n10859), .B2(n6848), .A(n6830), .ZN(n6831) );
  OAI21_X1 U8142 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n6929), .A(n6831), .ZN(n6832) );
  AOI21_X1 U8143 ( .B1(n10858), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n6832), .ZN(
        n6833) );
  OAI21_X1 U8144 ( .B1(n5182), .B2(n9330), .A(n6833), .ZN(P2_U3182) );
  INV_X1 U8145 ( .A(n7835), .ZN(n7014) );
  INV_X1 U8146 ( .A(n6834), .ZN(n6836) );
  INV_X1 U8147 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6835) );
  OAI222_X1 U8148 ( .A1(P1_U3086), .A2(n7014), .B1(n8657), .B2(n6836), .C1(
        n6835), .C2(n10595), .ZN(P1_U3343) );
  INV_X1 U8149 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6837) );
  INV_X1 U8150 ( .A(n9206), .ZN(n9213) );
  OAI222_X1 U8151 ( .A1(n8618), .A2(n6837), .B1(n9719), .B2(n6836), .C1(n9213), 
        .C2(P2_U3151), .ZN(P2_U3283) );
  INV_X1 U8152 ( .A(n6838), .ZN(n6842) );
  AOI22_X1 U8153 ( .A1(n10767), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n7744), .ZN(n6839) );
  OAI21_X1 U8154 ( .B1(n6842), .B2(n8657), .A(n6839), .ZN(P1_U3342) );
  INV_X1 U8155 ( .A(P1_U3973), .ZN(n7088) );
  NAND2_X1 U8156 ( .A1(n7088), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n6840) );
  OAI21_X1 U8157 ( .B1(n7088), .B2(n9798), .A(n6840), .ZN(P1_U3570) );
  NAND2_X1 U8158 ( .A1(n7088), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6841) );
  OAI21_X1 U8159 ( .B1(n7088), .B2(n10449), .A(n6841), .ZN(P1_U3575) );
  INV_X1 U8160 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6843) );
  INV_X1 U8161 ( .A(n9226), .ZN(n9242) );
  OAI222_X1 U8162 ( .A1(n8618), .A2(n6843), .B1(n9719), .B2(n6842), .C1(
        P2_U3151), .C2(n9242), .ZN(P2_U3282) );
  NAND2_X1 U8163 ( .A1(n6848), .A2(n6859), .ZN(n10854) );
  INV_X1 U8164 ( .A(n10854), .ZN(n6858) );
  NOR2_X1 U8165 ( .A1(n6933), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6844) );
  NAND2_X1 U8166 ( .A1(n6849), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6874) );
  NAND2_X1 U8167 ( .A1(n6846), .A2(n7147), .ZN(n6847) );
  NAND2_X1 U8168 ( .A1(n6875), .A2(n6847), .ZN(n6857) );
  NAND2_X1 U8169 ( .A1(n6848), .A2(n9327), .ZN(n10833) );
  NAND2_X1 U8170 ( .A1(n6849), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6883) );
  NAND2_X1 U8171 ( .A1(n6868), .A2(n6883), .ZN(n6852) );
  NAND2_X1 U8172 ( .A1(n5182), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6850) );
  OR2_X1 U8173 ( .A1(n6850), .A2(n6849), .ZN(n6851) );
  NAND2_X1 U8174 ( .A1(n6852), .A2(n6851), .ZN(n6882) );
  INV_X1 U8175 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6853) );
  XNOR2_X1 U8176 ( .A(n6882), .B(n6853), .ZN(n6854) );
  OAI22_X1 U8177 ( .A1(n10833), .A2(n6854), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6964), .ZN(n6856) );
  INV_X1 U8178 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10608) );
  NOR2_X1 U8179 ( .A1(n10843), .A2(n10608), .ZN(n6855) );
  AOI211_X1 U8180 ( .C1(n6858), .C2(n6857), .A(n6856), .B(n6855), .ZN(n6862)
         );
  MUX2_X1 U8181 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n9327), .Z(n6869) );
  XOR2_X1 U8182 ( .A(n6868), .B(n6869), .Z(n6871) );
  XOR2_X1 U8183 ( .A(n6870), .B(n6871), .Z(n6860) );
  NAND2_X1 U8184 ( .A1(n6860), .A2(n10859), .ZN(n6861) );
  OAI211_X1 U8185 ( .C1(n9330), .C2(n6868), .A(n6862), .B(n6861), .ZN(P2_U3183) );
  INV_X1 U8186 ( .A(n6863), .ZN(n6865) );
  AOI22_X1 U8187 ( .A1(n10726), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n7744), .ZN(n6864) );
  OAI21_X1 U8188 ( .B1(n6865), .B2(n8657), .A(n6864), .ZN(P1_U3341) );
  INV_X1 U8189 ( .A(n9240), .ZN(n9264) );
  OAI222_X1 U8190 ( .A1(n8618), .A2(n6866), .B1(n9719), .B2(n6865), .C1(
        P2_U3151), .C2(n9264), .ZN(P2_U3281) );
  NAND2_X1 U8191 ( .A1(P1_U3973), .A2(n10376), .ZN(n6867) );
  OAI21_X1 U8192 ( .B1(P1_U3973), .B2(n7778), .A(n6867), .ZN(P1_U3577) );
  INV_X1 U8193 ( .A(n10859), .ZN(n10823) );
  AOI22_X1 U8194 ( .A1(n6871), .A2(n6870), .B1(n6869), .B2(n6868), .ZN(n7358)
         );
  MUX2_X1 U8195 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n9327), .Z(n7354) );
  XNOR2_X1 U8196 ( .A(n7354), .B(n7339), .ZN(n7357) );
  XNOR2_X1 U8197 ( .A(n7358), .B(n7357), .ZN(n6896) );
  NOR2_X1 U8198 ( .A1(n9330), .A2(n7339), .ZN(n6894) );
  INV_X1 U8199 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n6872) );
  NOR2_X1 U8200 ( .A1(n10843), .A2(n6872), .ZN(n6893) );
  XNOR2_X1 U8201 ( .A(n7339), .B(n6873), .ZN(n6876) );
  NAND2_X1 U8202 ( .A1(n6875), .A2(n6874), .ZN(n6877) );
  NAND2_X1 U8203 ( .A1(n6876), .A2(n6877), .ZN(n7330) );
  INV_X1 U8204 ( .A(n6876), .ZN(n6879) );
  INV_X1 U8205 ( .A(n6877), .ZN(n6878) );
  NAND2_X1 U8206 ( .A1(n6879), .A2(n6878), .ZN(n6880) );
  AND2_X1 U8207 ( .A1(n7330), .A2(n6880), .ZN(n6881) );
  NOR2_X1 U8208 ( .A1(n10854), .A2(n6881), .ZN(n6892) );
  MUX2_X1 U8209 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n7341), .S(n7339), .Z(n6885)
         );
  NAND2_X1 U8210 ( .A1(n6882), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6884) );
  NAND2_X1 U8211 ( .A1(n6884), .A2(n6883), .ZN(n6886) );
  NAND2_X1 U8212 ( .A1(n6885), .A2(n6886), .ZN(n7340) );
  INV_X1 U8213 ( .A(n6885), .ZN(n6888) );
  INV_X1 U8214 ( .A(n6886), .ZN(n6887) );
  NAND2_X1 U8215 ( .A1(n6888), .A2(n6887), .ZN(n6889) );
  AND2_X1 U8216 ( .A1(n7340), .A2(n6889), .ZN(n6890) );
  OAI22_X1 U8217 ( .A1(n10833), .A2(n6890), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7208), .ZN(n6891) );
  NOR4_X1 U8218 ( .A1(n6894), .A2(n6893), .A3(n6892), .A4(n6891), .ZN(n6895)
         );
  OAI21_X1 U8219 ( .B1(n10823), .B2(n6896), .A(n6895), .ZN(P2_U3184) );
  NAND2_X1 U8220 ( .A1(n6915), .A2(n6897), .ZN(n6901) );
  NAND2_X1 U8221 ( .A1(n6914), .A2(n6898), .ZN(n6909) );
  NAND4_X1 U8222 ( .A1(n6901), .A2(n6900), .A3(n6909), .A4(n6899), .ZN(n6903)
         );
  NAND2_X1 U8223 ( .A1(n6908), .A2(n6928), .ZN(n6913) );
  INV_X1 U8224 ( .A(n6913), .ZN(n8895) );
  AND2_X1 U8225 ( .A1(n6914), .A2(n8895), .ZN(n6902) );
  AOI21_X1 U8226 ( .B1(n6903), .B2(P2_STATE_REG_SCAN_IN), .A(n6902), .ZN(n7075) );
  AND2_X1 U8227 ( .A1(n7075), .A2(n6904), .ZN(n7052) );
  INV_X1 U8228 ( .A(n6905), .ZN(n6907) );
  OAI21_X1 U8229 ( .B1(n6915), .B2(n6907), .A(n6906), .ZN(n6911) );
  AND2_X1 U8230 ( .A1(n6909), .A2(n6908), .ZN(n6910) );
  NAND2_X1 U8231 ( .A1(n6911), .A2(n6910), .ZN(n9185) );
  INV_X1 U8232 ( .A(n9185), .ZN(n9148) );
  AND2_X1 U8233 ( .A1(n6912), .A2(n6949), .ZN(n8705) );
  INV_X1 U8234 ( .A(n8705), .ZN(n8700) );
  NAND2_X1 U8235 ( .A1(n8699), .A2(n8700), .ZN(n8856) );
  NOR2_X1 U8236 ( .A1(n6914), .A2(n6913), .ZN(n6962) );
  AND2_X1 U8237 ( .A1(n6962), .A2(n6960), .ZN(n9181) );
  INV_X1 U8238 ( .A(n9181), .ZN(n9173) );
  INV_X1 U8239 ( .A(n6915), .ZN(n6916) );
  NAND2_X1 U8240 ( .A1(n6916), .A2(n6917), .ZN(n6919) );
  INV_X1 U8241 ( .A(n6917), .ZN(n6918) );
  NAND2_X1 U8242 ( .A1(n6919), .A2(n10937), .ZN(n9190) );
  INV_X1 U8243 ( .A(n9190), .ZN(n9166) );
  OAI22_X1 U8244 ( .A1(n7048), .A2(n9173), .B1(n9166), .B2(n6949), .ZN(n6920)
         );
  AOI21_X1 U8245 ( .B1(n9148), .B2(n8856), .A(n6920), .ZN(n6921) );
  OAI21_X1 U8246 ( .B1(n7052), .B2(n6929), .A(n6921), .ZN(P2_U3172) );
  AOI22_X1 U8247 ( .A1(n6925), .A2(n6924), .B1(n6923), .B2(n6922), .ZN(n6926)
         );
  NAND2_X1 U8248 ( .A1(n6927), .A2(n6926), .ZN(n6932) );
  NOR3_X1 U8249 ( .A1(n6932), .A2(n11017), .A3(n6928), .ZN(n6931) );
  OAI22_X1 U8250 ( .A1(n10939), .A2(n6949), .B1(n6929), .B2(n10937), .ZN(n6930) );
  AOI21_X1 U8251 ( .B1(n6931), .B2(n8856), .A(n6930), .ZN(n6935) );
  NAND2_X1 U8252 ( .A1(n6953), .A2(n10926), .ZN(n6936) );
  MUX2_X1 U8253 ( .A(n6933), .B(n6936), .S(n10944), .Z(n6934) );
  NAND2_X1 U8254 ( .A1(n6935), .A2(n6934), .ZN(P2_U3233) );
  OAI21_X1 U8255 ( .B1(n10928), .B2(n11097), .A(n8856), .ZN(n6937) );
  OAI211_X1 U8256 ( .C1(n11093), .C2(n6949), .A(n6937), .B(n6936), .ZN(n6939)
         );
  NAND2_X1 U8257 ( .A1(n6939), .A2(n11100), .ZN(n6938) );
  OAI21_X1 U8258 ( .B1(n11100), .B2(n6828), .A(n6938), .ZN(P2_U3459) );
  INV_X1 U8259 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6941) );
  NAND2_X1 U8260 ( .A1(n6939), .A2(n11104), .ZN(n6940) );
  OAI21_X1 U8261 ( .B1(n11104), .B2(n6941), .A(n6940), .ZN(P2_U3390) );
  INV_X1 U8262 ( .A(n6942), .ZN(n6944) );
  INV_X1 U8263 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6943) );
  OAI222_X1 U8264 ( .A1(P1_U3086), .A2(n7837), .B1(n8657), .B2(n6944), .C1(
        n6943), .C2(n10595), .ZN(P1_U3340) );
  INV_X1 U8265 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6945) );
  INV_X1 U8266 ( .A(n9263), .ZN(n9285) );
  OAI222_X1 U8267 ( .A1(n8618), .A2(n6945), .B1(n9719), .B2(n6944), .C1(n9285), 
        .C2(P2_U3151), .ZN(P2_U3280) );
  NAND2_X1 U8268 ( .A1(n6947), .A2(n8849), .ZN(n6948) );
  NAND2_X1 U8269 ( .A1(n6949), .A2(n7152), .ZN(n6950) );
  NAND2_X1 U8270 ( .A1(n6950), .A2(n7145), .ZN(n6959) );
  NAND2_X1 U8271 ( .A1(n6951), .A2(n6952), .ZN(n7043) );
  INV_X1 U8272 ( .A(n6952), .ZN(n6954) );
  NAND2_X1 U8273 ( .A1(n6954), .A2(n6953), .ZN(n6955) );
  INV_X1 U8274 ( .A(n6959), .ZN(n6957) );
  INV_X1 U8275 ( .A(n7044), .ZN(n6958) );
  AOI21_X1 U8276 ( .B1(n6959), .B2(n6956), .A(n6958), .ZN(n6968) );
  INV_X1 U8277 ( .A(n10925), .ZN(n8711) );
  INV_X1 U8278 ( .A(n6912), .ZN(n6963) );
  INV_X1 U8279 ( .A(n6960), .ZN(n6961) );
  NAND2_X1 U8280 ( .A1(n6962), .A2(n6961), .ZN(n9178) );
  OAI22_X1 U8281 ( .A1(n8711), .A2(n9173), .B1(n6963), .B2(n9178), .ZN(n6966)
         );
  NOR2_X1 U8282 ( .A1(n7052), .A2(n6964), .ZN(n6965) );
  AOI211_X1 U8283 ( .C1(n7148), .C2(n9190), .A(n6966), .B(n6965), .ZN(n6967)
         );
  OAI21_X1 U8284 ( .B1(n6968), .B2(n9185), .A(n6967), .ZN(P2_U3162) );
  OR2_X1 U8285 ( .A1(n6970), .A2(n6969), .ZN(n10669) );
  INV_X1 U8286 ( .A(n10669), .ZN(n7009) );
  OR2_X1 U8287 ( .A1(n6210), .A2(n10660), .ZN(n10663) );
  INV_X1 U8288 ( .A(n10663), .ZN(n6971) );
  NAND2_X1 U8289 ( .A1(n7009), .A2(n6971), .ZN(n10797) );
  INV_X1 U8290 ( .A(n10797), .ZN(n10776) );
  NOR2_X1 U8291 ( .A1(n7835), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6972) );
  AOI21_X1 U8292 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7835), .A(n6972), .ZN(
        n6987) );
  NAND2_X1 U8293 ( .A1(n10774), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6973) );
  OAI21_X1 U8294 ( .B1(n10774), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6973), .ZN(
        n10773) );
  AOI22_X1 U8295 ( .A1(n10798), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n5848), .B2(
        n7004), .ZN(n10793) );
  MUX2_X1 U8296 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n5829), .S(n10692), .Z(n10688) );
  MUX2_X1 U8297 ( .A(n7290), .B(P1_REG2_REG_2__SCAN_IN), .S(n6989), .Z(n10200)
         );
  MUX2_X1 U8298 ( .A(n7324), .B(P1_REG2_REG_1__SCAN_IN), .S(n6990), .Z(n10174)
         );
  AND2_X1 U8299 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n10173) );
  NAND2_X1 U8300 ( .A1(n10174), .A2(n10173), .ZN(n10172) );
  INV_X1 U8301 ( .A(n6990), .ZN(n10181) );
  NAND2_X1 U8302 ( .A1(n10181), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6974) );
  NAND2_X1 U8303 ( .A1(n10172), .A2(n6974), .ZN(n10199) );
  NAND2_X1 U8304 ( .A1(n10200), .A2(n10199), .ZN(n10198) );
  INV_X1 U8305 ( .A(n6989), .ZN(n10194) );
  NAND2_X1 U8306 ( .A1(n10194), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6975) );
  NAND2_X1 U8307 ( .A1(n10198), .A2(n6975), .ZN(n10205) );
  XNOR2_X1 U8308 ( .A(n6993), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n10206) );
  NAND2_X1 U8309 ( .A1(n10205), .A2(n10206), .ZN(n10204) );
  INV_X1 U8310 ( .A(n6993), .ZN(n10213) );
  NAND2_X1 U8311 ( .A1(n10213), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6976) );
  NAND2_X1 U8312 ( .A1(n10204), .A2(n6976), .ZN(n10224) );
  XNOR2_X1 U8313 ( .A(n10217), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n10225) );
  NAND2_X1 U8314 ( .A1(n10224), .A2(n10225), .ZN(n10223) );
  OR2_X1 U8315 ( .A1(n10217), .A2(n6977), .ZN(n6978) );
  NAND2_X1 U8316 ( .A1(n10223), .A2(n6978), .ZN(n10234) );
  XNOR2_X1 U8317 ( .A(n10242), .B(n6979), .ZN(n10235) );
  NAND2_X1 U8318 ( .A1(n10234), .A2(n10235), .ZN(n10233) );
  NAND2_X1 U8319 ( .A1(n10242), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6980) );
  NAND2_X1 U8320 ( .A1(n10233), .A2(n6980), .ZN(n10247) );
  XNOR2_X1 U8321 ( .A(n10253), .B(n6981), .ZN(n10248) );
  NAND2_X1 U8322 ( .A1(n10247), .A2(n10248), .ZN(n10246) );
  NAND2_X1 U8323 ( .A1(n10253), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6982) );
  NAND2_X1 U8324 ( .A1(n10246), .A2(n6982), .ZN(n10674) );
  MUX2_X1 U8325 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n7310), .S(n10678), .Z(n10673) );
  AND2_X1 U8326 ( .A1(n10674), .A2(n10673), .ZN(n10676) );
  AOI21_X1 U8327 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n10678), .A(n10676), .ZN(
        n6983) );
  INV_X1 U8328 ( .A(n6983), .ZN(n10687) );
  NAND2_X1 U8329 ( .A1(n10688), .A2(n10687), .ZN(n10686) );
  NAND2_X1 U8330 ( .A1(n10692), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6984) );
  AND2_X1 U8331 ( .A1(n10686), .A2(n6984), .ZN(n10792) );
  NAND2_X1 U8332 ( .A1(n10793), .A2(n10792), .ZN(n10794) );
  OAI21_X1 U8333 ( .B1(n10798), .B2(P1_REG2_REG_9__SCAN_IN), .A(n10794), .ZN(
        n10772) );
  NOR2_X1 U8334 ( .A1(n10773), .A2(n10772), .ZN(n10771) );
  AOI21_X1 U8335 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n10774), .A(n10771), .ZN(
        n10700) );
  NAND2_X1 U8336 ( .A1(n10709), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6985) );
  OAI21_X1 U8337 ( .B1(n10709), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6985), .ZN(
        n10701) );
  NOR2_X1 U8338 ( .A1(n10700), .A2(n10701), .ZN(n10702) );
  AOI21_X1 U8339 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n10709), .A(n10702), .ZN(
        n6986) );
  NAND2_X1 U8340 ( .A1(n6987), .A2(n6986), .ZN(n7834) );
  OAI21_X1 U8341 ( .B1(n6987), .B2(n6986), .A(n7834), .ZN(n7016) );
  NOR2_X2 U8342 ( .A1(n10669), .A2(n7066), .ZN(n10799) );
  INV_X1 U8343 ( .A(n10799), .ZN(n10754) );
  AOI22_X1 U8344 ( .A1(n7835), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n5893), .B2(
        n7014), .ZN(n7008) );
  INV_X1 U8345 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6988) );
  MUX2_X1 U8346 ( .A(n6988), .B(P1_REG1_REG_10__SCAN_IN), .S(n10774), .Z(
        n10777) );
  INV_X1 U8347 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10889) );
  MUX2_X1 U8348 ( .A(n10889), .B(P1_REG1_REG_2__SCAN_IN), .S(n6989), .Z(n10197) );
  INV_X1 U8349 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10881) );
  MUX2_X1 U8350 ( .A(n10881), .B(P1_REG1_REG_1__SCAN_IN), .S(n6990), .Z(n10177) );
  AND2_X1 U8351 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n10176) );
  NAND2_X1 U8352 ( .A1(n10177), .A2(n10176), .ZN(n10175) );
  NAND2_X1 U8353 ( .A1(n10181), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6991) );
  NAND2_X1 U8354 ( .A1(n10175), .A2(n6991), .ZN(n10196) );
  NAND2_X1 U8355 ( .A1(n10197), .A2(n10196), .ZN(n10195) );
  NAND2_X1 U8356 ( .A1(n10194), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6992) );
  NAND2_X1 U8357 ( .A1(n10195), .A2(n6992), .ZN(n10208) );
  XNOR2_X1 U8358 ( .A(n6993), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n10209) );
  NAND2_X1 U8359 ( .A1(n10208), .A2(n10209), .ZN(n10207) );
  NAND2_X1 U8360 ( .A1(n10213), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6994) );
  NAND2_X1 U8361 ( .A1(n10207), .A2(n6994), .ZN(n10227) );
  XNOR2_X1 U8362 ( .A(n10217), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n10228) );
  NAND2_X1 U8363 ( .A1(n10227), .A2(n10228), .ZN(n10226) );
  INV_X1 U8364 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6995) );
  OR2_X1 U8365 ( .A1(n10217), .A2(n6995), .ZN(n6996) );
  NAND2_X1 U8366 ( .A1(n10226), .A2(n6996), .ZN(n10237) );
  XNOR2_X1 U8367 ( .A(n10242), .B(n6997), .ZN(n10238) );
  NAND2_X1 U8368 ( .A1(n10237), .A2(n10238), .ZN(n10236) );
  NAND2_X1 U8369 ( .A1(n10242), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6998) );
  NAND2_X1 U8370 ( .A1(n10236), .A2(n6998), .ZN(n10250) );
  XNOR2_X1 U8371 ( .A(n10253), .B(n6999), .ZN(n10251) );
  NAND2_X1 U8372 ( .A1(n10250), .A2(n10251), .ZN(n10249) );
  NAND2_X1 U8373 ( .A1(n10253), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7000) );
  NAND2_X1 U8374 ( .A1(n10249), .A2(n7000), .ZN(n10671) );
  MUX2_X1 U8375 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n5812), .S(n10678), .Z(n10672) );
  NAND2_X1 U8376 ( .A1(n10671), .A2(n10672), .ZN(n10670) );
  NAND2_X1 U8377 ( .A1(n10678), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7001) );
  NAND2_X1 U8378 ( .A1(n10670), .A2(n7001), .ZN(n10690) );
  MUX2_X1 U8379 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n5826), .S(n10692), .Z(n10691) );
  NAND2_X1 U8380 ( .A1(n10690), .A2(n10691), .ZN(n10689) );
  NAND2_X1 U8381 ( .A1(n10692), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7002) );
  NAND2_X1 U8382 ( .A1(n10689), .A2(n7002), .ZN(n10789) );
  MUX2_X1 U8383 ( .A(n7003), .B(P1_REG1_REG_9__SCAN_IN), .S(n10798), .Z(n10788) );
  NAND2_X1 U8384 ( .A1(n7004), .A2(n7003), .ZN(n7005) );
  NAND2_X1 U8385 ( .A1(n10791), .A2(n7005), .ZN(n10778) );
  NOR2_X1 U8386 ( .A1(n10777), .A2(n10778), .ZN(n10779) );
  AOI21_X1 U8387 ( .B1(n10774), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10779), .ZN(
        n10706) );
  MUX2_X1 U8388 ( .A(n7006), .B(P1_REG1_REG_11__SCAN_IN), .S(n10709), .Z(
        n10707) );
  NOR2_X1 U8389 ( .A1(n10706), .A2(n10707), .ZN(n10705) );
  AOI21_X1 U8390 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n10709), .A(n10705), .ZN(
        n7007) );
  NAND2_X1 U8391 ( .A1(n7008), .A2(n7007), .ZN(n7825) );
  OAI21_X1 U8392 ( .B1(n7008), .B2(n7007), .A(n7825), .ZN(n7010) );
  NAND2_X1 U8393 ( .A1(n7009), .A2(n10660), .ZN(n10803) );
  INV_X1 U8394 ( .A(n10803), .ZN(n10782) );
  NAND2_X1 U8395 ( .A1(n7010), .A2(n10782), .ZN(n7013) );
  INV_X1 U8396 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7011) );
  NOR2_X1 U8397 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7011), .ZN(n7985) );
  AOI21_X1 U8398 ( .B1(n10666), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n7985), .ZN(
        n7012) );
  OAI211_X1 U8399 ( .C1(n10754), .C2(n7014), .A(n7013), .B(n7012), .ZN(n7015)
         );
  AOI21_X1 U8400 ( .B1(n10776), .B2(n7016), .A(n7015), .ZN(n7017) );
  INV_X1 U8401 ( .A(n7017), .ZN(P1_U3255) );
  INV_X1 U8402 ( .A(n7018), .ZN(n7281) );
  NAND3_X1 U8403 ( .A1(n7020), .A2(n7281), .A3(n7019), .ZN(n7039) );
  INV_X1 U8404 ( .A(n10584), .ZN(n10148) );
  NOR2_X1 U8405 ( .A1(n7037), .A2(n10147), .ZN(n7067) );
  NAND2_X1 U8406 ( .A1(n7067), .A2(n6210), .ZN(n9877) );
  INV_X1 U8407 ( .A(n9877), .ZN(n9845) );
  INV_X1 U8408 ( .A(n7027), .ZN(n7021) );
  OR2_X1 U8409 ( .A1(n7027), .A2(n10274), .ZN(n7458) );
  NAND2_X1 U8410 ( .A1(n10151), .A2(n7022), .ZN(n7023) );
  NAND2_X1 U8411 ( .A1(n8976), .A2(n9906), .ZN(n7026) );
  INV_X1 U8412 ( .A(n7032), .ZN(n7024) );
  NAND2_X1 U8413 ( .A1(n7024), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n7025) );
  OAI211_X1 U8414 ( .C1(n7115), .C2(n9905), .A(n7026), .B(n7025), .ZN(n7053)
         );
  NAND2_X1 U8415 ( .A1(n7759), .A2(n9906), .ZN(n7030) );
  XOR2_X1 U8416 ( .A(n7053), .B(n7054), .Z(n10190) );
  INV_X1 U8417 ( .A(n7037), .ZN(n7035) );
  AND2_X1 U8418 ( .A1(n11074), .A2(n10106), .ZN(n7034) );
  NAND2_X1 U8419 ( .A1(n7035), .A2(n7034), .ZN(n9866) );
  AOI22_X1 U8420 ( .A1(n9845), .A2(n10171), .B1(n10190), .B2(n9871), .ZN(n7042) );
  OR2_X1 U8421 ( .A1(n7090), .A2(n7536), .ZN(n7291) );
  INV_X1 U8422 ( .A(n7038), .ZN(n7036) );
  NAND2_X2 U8423 ( .A1(n7036), .A2(n10584), .ZN(n11050) );
  OAI21_X2 U8424 ( .B1(n7037), .B2(n7291), .A(n11050), .ZN(n9863) );
  NAND2_X1 U8425 ( .A1(n7039), .A2(n7038), .ZN(n7130) );
  NAND2_X1 U8426 ( .A1(n7130), .A2(n7040), .ZN(n9847) );
  AOI22_X1 U8427 ( .A1(n9863), .A2(n7382), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n9847), .ZN(n7041) );
  NAND2_X1 U8428 ( .A1(n7042), .A2(n7041), .ZN(P1_U3232) );
  XNOR2_X1 U8429 ( .A(n8710), .B(n7152), .ZN(n7076) );
  XNOR2_X1 U8430 ( .A(n7076), .B(n10925), .ZN(n7046) );
  NAND2_X1 U8431 ( .A1(n7045), .A2(n7046), .ZN(n7078) );
  OAI21_X1 U8432 ( .B1(n7046), .B2(n7045), .A(n7078), .ZN(n7047) );
  NAND2_X1 U8433 ( .A1(n7047), .A2(n9148), .ZN(n7051) );
  INV_X1 U8434 ( .A(n9204), .ZN(n7165) );
  OAI22_X1 U8435 ( .A1(n7165), .A2(n9173), .B1(n7048), .B2(n9178), .ZN(n7049)
         );
  AOI21_X1 U8436 ( .B1(n8710), .B2(n9190), .A(n7049), .ZN(n7050) );
  OAI211_X1 U8437 ( .C1(n7052), .C2(n7208), .A(n7051), .B(n7050), .ZN(P2_U3177) );
  OR2_X1 U8438 ( .A1(n7055), .A2(n9002), .ZN(n7056) );
  NAND2_X1 U8439 ( .A1(n7057), .A2(n7056), .ZN(n7064) );
  INV_X1 U8440 ( .A(n7064), .ZN(n7062) );
  NAND2_X1 U8441 ( .A1(n9000), .A2(n5247), .ZN(n7059) );
  NAND2_X1 U8442 ( .A1(n7759), .A2(n10171), .ZN(n7058) );
  NAND2_X1 U8443 ( .A1(n7059), .A2(n7058), .ZN(n7060) );
  XNOR2_X1 U8444 ( .A(n7060), .B(n9002), .ZN(n7063) );
  INV_X1 U8445 ( .A(n7063), .ZN(n7061) );
  NAND2_X1 U8446 ( .A1(n7062), .A2(n7061), .ZN(n7097) );
  NAND2_X1 U8447 ( .A1(n7064), .A2(n7063), .ZN(n7096) );
  NAND2_X1 U8448 ( .A1(n7097), .A2(n7096), .ZN(n7065) );
  AOI22_X1 U8449 ( .A1(n8976), .A2(n10171), .B1(n8961), .B2(n5247), .ZN(n7095)
         );
  XNOR2_X1 U8450 ( .A(n7065), .B(n7095), .ZN(n7070) );
  NAND2_X1 U8451 ( .A1(n7067), .A2(n7066), .ZN(n9876) );
  INV_X1 U8452 ( .A(n9876), .ZN(n9846) );
  AOI22_X1 U8453 ( .A1(n9846), .A2(n9906), .B1(n9845), .B2(n10170), .ZN(n7069)
         );
  AOI22_X1 U8454 ( .A1(n9863), .A2(n5247), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n9847), .ZN(n7068) );
  OAI211_X1 U8455 ( .C1(n7070), .C2(n9866), .A(n7069), .B(n7068), .ZN(P1_U3222) );
  INV_X1 U8456 ( .A(n7071), .ZN(n7073) );
  INV_X1 U8457 ( .A(n9313), .ZN(n9301) );
  OAI222_X1 U8458 ( .A1(n8618), .A2(n7072), .B1(n9719), .B2(n7073), .C1(
        P2_U3151), .C2(n9301), .ZN(P2_U3279) );
  INV_X1 U8459 ( .A(n7866), .ZN(n7832) );
  OAI222_X1 U8460 ( .A1(n7832), .A2(P1_U3086), .B1(n8657), .B2(n7073), .C1(
        n8525), .C2(n10595), .ZN(P1_U3339) );
  NAND2_X1 U8461 ( .A1(n7074), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8899) );
  NAND2_X1 U8462 ( .A1(n7075), .A2(n8899), .ZN(n9171) );
  NAND2_X1 U8463 ( .A1(n8711), .A2(n7076), .ZN(n7077) );
  NAND2_X1 U8464 ( .A1(n7078), .A2(n7077), .ZN(n7176) );
  XNOR2_X1 U8465 ( .A(n10933), .B(n7079), .ZN(n7151) );
  XNOR2_X1 U8466 ( .A(n7151), .B(n9204), .ZN(n7170) );
  AOI21_X1 U8467 ( .B1(n7176), .B2(n7170), .A(n9185), .ZN(n7080) );
  OR2_X1 U8468 ( .A1(n7176), .A2(n7170), .ZN(n7160) );
  NAND2_X1 U8469 ( .A1(n7080), .A2(n7160), .ZN(n7083) );
  AND2_X1 U8470 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n10813) );
  OAI22_X1 U8471 ( .A1(n10938), .A2(n9166), .B1(n8711), .B2(n9178), .ZN(n7081)
         );
  AOI211_X1 U8472 ( .C1(n9181), .C2(n7154), .A(n10813), .B(n7081), .ZN(n7082)
         );
  OAI211_X1 U8473 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n9183), .A(n7083), .B(
        n7082), .ZN(P2_U3158) );
  INV_X1 U8474 ( .A(n7867), .ZN(n10267) );
  INV_X1 U8475 ( .A(n7084), .ZN(n7085) );
  OAI222_X1 U8476 ( .A1(P1_U3086), .A2(n10267), .B1(n8657), .B2(n7085), .C1(
        n8309), .C2(n10595), .ZN(P1_U3338) );
  INV_X1 U8477 ( .A(n9325), .ZN(n9337) );
  OAI222_X1 U8478 ( .A1(n8618), .A2(n7086), .B1(n9719), .B2(n7085), .C1(n9337), 
        .C2(P2_U3151), .ZN(P2_U3278) );
  NAND2_X1 U8479 ( .A1(n7088), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7087) );
  OAI21_X1 U8480 ( .B1(n7088), .B2(n10310), .A(n7087), .ZN(P1_U3583) );
  XNOR2_X1 U8481 ( .A(n9906), .B(n7382), .ZN(n10067) );
  INV_X1 U8482 ( .A(n10402), .ZN(n11030) );
  AND2_X1 U8483 ( .A1(n10543), .A2(n11030), .ZN(n7089) );
  OR2_X1 U8484 ( .A1(n10067), .A2(n7089), .ZN(n7093) );
  INV_X1 U8485 ( .A(n10902), .ZN(n11026) );
  AND2_X1 U8486 ( .A1(n10171), .A2(n11026), .ZN(n7381) );
  INV_X1 U8487 ( .A(n7090), .ZN(n7378) );
  AND2_X1 U8488 ( .A1(n7378), .A2(n7382), .ZN(n7091) );
  NOR2_X1 U8489 ( .A1(n7381), .A2(n7091), .ZN(n7092) );
  AND2_X1 U8490 ( .A1(n7093), .A2(n7092), .ZN(n10867) );
  NAND2_X1 U8491 ( .A1(n11080), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7094) );
  OAI21_X1 U8492 ( .B1(n11080), .B2(n10867), .A(n7094), .ZN(P1_U3522) );
  NAND2_X1 U8493 ( .A1(n7096), .A2(n7095), .ZN(n7098) );
  NAND2_X1 U8494 ( .A1(n7098), .A2(n7097), .ZN(n9850) );
  NAND2_X1 U8495 ( .A1(n9000), .A2(n9848), .ZN(n7100) );
  NAND2_X1 U8496 ( .A1(n7759), .A2(n10170), .ZN(n7099) );
  NAND2_X1 U8497 ( .A1(n7100), .A2(n7099), .ZN(n7101) );
  XNOR2_X1 U8498 ( .A(n7101), .B(n8974), .ZN(n7103) );
  AOI22_X1 U8499 ( .A1(n8976), .A2(n10170), .B1(n8961), .B2(n9848), .ZN(n7102)
         );
  NAND2_X1 U8500 ( .A1(n7103), .A2(n7102), .ZN(n7105) );
  OR2_X1 U8501 ( .A1(n7103), .A2(n7102), .ZN(n7104) );
  AND2_X1 U8502 ( .A1(n7105), .A2(n7104), .ZN(n9851) );
  NAND2_X1 U8503 ( .A1(n9850), .A2(n9851), .ZN(n9849) );
  NAND2_X1 U8504 ( .A1(n9849), .A2(n7105), .ZN(n9742) );
  INV_X1 U8505 ( .A(n10899), .ZN(n10917) );
  NAND2_X1 U8506 ( .A1(n9000), .A2(n10917), .ZN(n7107) );
  NAND2_X1 U8507 ( .A1(n8961), .A2(n10169), .ZN(n7106) );
  NAND2_X1 U8508 ( .A1(n7107), .A2(n7106), .ZN(n7108) );
  XNOR2_X1 U8509 ( .A(n7108), .B(n8974), .ZN(n7113) );
  NAND2_X1 U8510 ( .A1(n8976), .A2(n10169), .ZN(n7110) );
  NAND2_X1 U8511 ( .A1(n8961), .A2(n10917), .ZN(n7109) );
  NAND2_X1 U8512 ( .A1(n7110), .A2(n7109), .ZN(n7111) );
  XNOR2_X1 U8513 ( .A(n7113), .B(n7111), .ZN(n9743) );
  NAND2_X1 U8514 ( .A1(n9742), .A2(n9743), .ZN(n9741) );
  INV_X1 U8515 ( .A(n7111), .ZN(n7112) );
  NAND2_X1 U8516 ( .A1(n7113), .A2(n7112), .ZN(n7114) );
  NAND2_X1 U8517 ( .A1(n9741), .A2(n7114), .ZN(n9817) );
  NAND2_X1 U8518 ( .A1(n9000), .A2(n9820), .ZN(n7117) );
  NAND2_X1 U8519 ( .A1(n8938), .A2(n9745), .ZN(n7116) );
  NAND2_X1 U8520 ( .A1(n7117), .A2(n7116), .ZN(n7118) );
  XNOR2_X1 U8521 ( .A(n7118), .B(n8974), .ZN(n7120) );
  AOI22_X1 U8522 ( .A1(n8976), .A2(n9745), .B1(n8938), .B2(n9820), .ZN(n7119)
         );
  XNOR2_X1 U8523 ( .A(n7120), .B(n7119), .ZN(n9816) );
  OR2_X1 U8524 ( .A1(n9817), .A2(n9816), .ZN(n9818) );
  OR2_X1 U8525 ( .A1(n7120), .A2(n7119), .ZN(n7238) );
  NAND2_X1 U8526 ( .A1(n9818), .A2(n7238), .ZN(n7127) );
  NAND2_X1 U8527 ( .A1(n9000), .A2(n7482), .ZN(n7122) );
  NAND2_X1 U8528 ( .A1(n8938), .A2(n10168), .ZN(n7121) );
  NAND2_X1 U8529 ( .A1(n7122), .A2(n7121), .ZN(n7123) );
  XNOR2_X1 U8530 ( .A(n7123), .B(n8974), .ZN(n7234) );
  NAND2_X1 U8531 ( .A1(n8976), .A2(n10168), .ZN(n7125) );
  NAND2_X1 U8532 ( .A1(n8938), .A2(n7482), .ZN(n7124) );
  AND2_X1 U8533 ( .A1(n7125), .A2(n7124), .ZN(n7232) );
  INV_X1 U8534 ( .A(n7232), .ZN(n7235) );
  XNOR2_X1 U8535 ( .A(n7234), .B(n7235), .ZN(n7126) );
  XNOR2_X1 U8536 ( .A(n7127), .B(n7126), .ZN(n7136) );
  AOI22_X1 U8537 ( .A1(n9845), .A2(n10167), .B1(n7482), .B2(n9863), .ZN(n7135)
         );
  INV_X1 U8538 ( .A(n7128), .ZN(n7129) );
  NAND2_X1 U8539 ( .A1(n7130), .A2(n7129), .ZN(n7131) );
  NAND2_X1 U8540 ( .A1(n7131), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9874) );
  INV_X1 U8541 ( .A(n9874), .ZN(n9803) );
  NAND2_X1 U8542 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10239) );
  INV_X1 U8543 ( .A(n10239), .ZN(n7133) );
  NOR2_X1 U8544 ( .A1(n9876), .A2(n5245), .ZN(n7132) );
  AOI211_X1 U8545 ( .C1(n9803), .C2(n7483), .A(n7133), .B(n7132), .ZN(n7134)
         );
  OAI211_X1 U8546 ( .C1(n7136), .C2(n9866), .A(n7135), .B(n7134), .ZN(P1_U3227) );
  INV_X1 U8547 ( .A(n10271), .ZN(n10753) );
  INV_X1 U8548 ( .A(n7137), .ZN(n7139) );
  INV_X1 U8549 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7138) );
  OAI222_X1 U8550 ( .A1(P1_U3086), .A2(n10753), .B1(n8657), .B2(n7139), .C1(
        n7138), .C2(n10595), .ZN(P1_U3337) );
  INV_X1 U8551 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7140) );
  INV_X1 U8552 ( .A(n9349), .ZN(n9356) );
  OAI222_X1 U8553 ( .A1(n8618), .A2(n7140), .B1(P2_U3151), .B2(n9356), .C1(
        n7139), .C2(n9719), .ZN(P2_U3277) );
  INV_X1 U8554 ( .A(n7141), .ZN(n7142) );
  AOI21_X1 U8555 ( .B1(n8699), .B2(n8857), .A(n7142), .ZN(n10870) );
  NOR2_X1 U8556 ( .A1(n7207), .A2(n8879), .ZN(n7942) );
  INV_X1 U8557 ( .A(n7942), .ZN(n7143) );
  NAND2_X1 U8558 ( .A1(n9021), .A2(n7143), .ZN(n9417) );
  INV_X1 U8559 ( .A(n10941), .ZN(n9513) );
  OAI21_X1 U8560 ( .B1(n8857), .B2(n7145), .A(n7144), .ZN(n7146) );
  AOI222_X1 U8561 ( .A1(n10928), .A2(n7146), .B1(n10925), .B2(n10926), .C1(
        n6912), .C2(n6677), .ZN(n10868) );
  MUX2_X1 U8562 ( .A(n7147), .B(n10868), .S(n10944), .Z(n7150) );
  INV_X1 U8563 ( .A(n10939), .ZN(n9509) );
  INV_X1 U8564 ( .A(n10937), .ZN(n9550) );
  AOI22_X1 U8565 ( .A1(n9509), .A2(n7148), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n9550), .ZN(n7149) );
  OAI211_X1 U8566 ( .C1(n10870), .C2(n9513), .A(n7150), .B(n7149), .ZN(
        P2_U3232) );
  NAND2_X1 U8567 ( .A1(n7151), .A2(n9204), .ZN(n7158) );
  AND2_X1 U8568 ( .A1(n7160), .A2(n7158), .ZN(n7161) );
  INV_X1 U8569 ( .A(n7156), .ZN(n7154) );
  XNOR2_X1 U8570 ( .A(n10951), .B(n7152), .ZN(n7155) );
  INV_X1 U8571 ( .A(n7155), .ZN(n7153) );
  NAND2_X1 U8572 ( .A1(n7154), .A2(n7153), .ZN(n7157) );
  NAND2_X1 U8573 ( .A1(n7156), .A2(n7155), .ZN(n7169) );
  AND2_X1 U8574 ( .A1(n7159), .A2(n7158), .ZN(n7172) );
  NAND2_X1 U8575 ( .A1(n7160), .A2(n7172), .ZN(n7189) );
  OAI21_X1 U8576 ( .B1(n7161), .B2(n7159), .A(n7189), .ZN(n7162) );
  NAND2_X1 U8577 ( .A1(n7162), .A2(n9148), .ZN(n7168) );
  NOR2_X1 U8578 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7163), .ZN(n10836) );
  AOI21_X1 U8579 ( .B1(n9181), .B2(n7171), .A(n10836), .ZN(n7164) );
  OAI21_X1 U8580 ( .B1(n7165), .B2(n9178), .A(n7164), .ZN(n7166) );
  AOI21_X1 U8581 ( .B1(n10951), .B2(n9190), .A(n7166), .ZN(n7167) );
  OAI211_X1 U8582 ( .C1(n7393), .C2(n9183), .A(n7168), .B(n7167), .ZN(P2_U3170) );
  INV_X1 U8583 ( .A(n7169), .ZN(n7190) );
  OR2_X1 U8584 ( .A1(n7170), .A2(n7190), .ZN(n7175) );
  XNOR2_X1 U8585 ( .A(n7516), .B(n7152), .ZN(n7177) );
  XNOR2_X1 U8586 ( .A(n7177), .B(n7171), .ZN(n7191) );
  OAI21_X1 U8587 ( .B1(n7172), .B2(n7190), .A(n7191), .ZN(n7173) );
  INV_X1 U8588 ( .A(n7173), .ZN(n7174) );
  NAND2_X1 U8589 ( .A1(n6364), .A2(n7177), .ZN(n7178) );
  XNOR2_X1 U8590 ( .A(n7179), .B(n7079), .ZN(n7397) );
  XNOR2_X1 U8591 ( .A(n7397), .B(n9203), .ZN(n7181) );
  AOI21_X1 U8592 ( .B1(n7180), .B2(n7181), .A(n9185), .ZN(n7183) );
  NAND2_X1 U8593 ( .A1(n7183), .A2(n7411), .ZN(n7188) );
  INV_X1 U8594 ( .A(n7580), .ZN(n7186) );
  INV_X1 U8595 ( .A(n9202), .ZN(n7737) );
  INV_X1 U8596 ( .A(n9178), .ZN(n9152) );
  NOR2_X1 U8597 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8495), .ZN(n7368) );
  AOI21_X1 U8598 ( .B1(n9152), .B2(n7171), .A(n7368), .ZN(n7184) );
  OAI21_X1 U8599 ( .B1(n7737), .B2(n9173), .A(n7184), .ZN(n7185) );
  AOI21_X1 U8600 ( .B1(n7186), .B2(n9171), .A(n7185), .ZN(n7187) );
  OAI211_X1 U8601 ( .C1(n10974), .C2(n9166), .A(n7188), .B(n7187), .ZN(
        P2_U3179) );
  INV_X1 U8602 ( .A(n7189), .ZN(n7192) );
  NOR3_X1 U8603 ( .A1(n7192), .A2(n7190), .A3(n7191), .ZN(n7195) );
  INV_X1 U8604 ( .A(n7193), .ZN(n7194) );
  OAI21_X1 U8605 ( .B1(n7195), .B2(n7194), .A(n9148), .ZN(n7199) );
  NAND2_X1 U8606 ( .A1(n9181), .A2(n9203), .ZN(n7196) );
  NAND2_X1 U8607 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n10851) );
  OAI211_X1 U8608 ( .C1(n7156), .C2(n9178), .A(n7196), .B(n10851), .ZN(n7197)
         );
  AOI21_X1 U8609 ( .B1(n7516), .B2(n9190), .A(n7197), .ZN(n7198) );
  OAI211_X1 U8610 ( .C1(n7514), .C2(n9183), .A(n7199), .B(n7198), .ZN(P2_U3167) );
  INV_X2 U8611 ( .A(n10944), .ZN(n10946) );
  OAI21_X1 U8612 ( .B1(n7202), .B2(n7201), .A(n7200), .ZN(n7203) );
  NAND2_X1 U8613 ( .A1(n7203), .A2(n10928), .ZN(n7205) );
  AOI22_X1 U8614 ( .A1(n6953), .A2(n6677), .B1(n10926), .B2(n9204), .ZN(n7204)
         );
  NAND2_X1 U8615 ( .A1(n7205), .A2(n7204), .ZN(n10891) );
  NOR2_X1 U8616 ( .A1(n7206), .A2(n11093), .ZN(n10892) );
  INV_X1 U8617 ( .A(n10892), .ZN(n7210) );
  INV_X1 U8618 ( .A(n7207), .ZN(n7209) );
  OAI22_X1 U8619 ( .A1(n7210), .A2(n7209), .B1(n10937), .B2(n7208), .ZN(n7211)
         );
  OAI21_X1 U8620 ( .B1(n10891), .B2(n7211), .A(n9589), .ZN(n7214) );
  XNOR2_X1 U8621 ( .A(n7212), .B(n8859), .ZN(n10893) );
  NAND2_X1 U8622 ( .A1(n10893), .A2(n10941), .ZN(n7213) );
  OAI211_X1 U8623 ( .C1(n6873), .C2(n9589), .A(n7214), .B(n7213), .ZN(P2_U3231) );
  OAI21_X1 U8624 ( .B1(n7216), .B2(n9964), .A(n7215), .ZN(n7605) );
  INV_X1 U8625 ( .A(n7481), .ZN(n7217) );
  AOI211_X1 U8626 ( .C1(n7747), .C2(n7217), .A(n10438), .B(n7311), .ZN(n7598)
         );
  NAND2_X1 U8627 ( .A1(n7474), .A2(n9912), .ZN(n7218) );
  XNOR2_X1 U8628 ( .A(n7218), .B(n9964), .ZN(n7219) );
  OAI222_X1 U8629 ( .A1(n10902), .A2(n7539), .B1(n10900), .B2(n7220), .C1(
        n7219), .C2(n11030), .ZN(n7597) );
  AOI211_X1 U8630 ( .C1(n11078), .C2(n7605), .A(n7598), .B(n7597), .ZN(n7749)
         );
  AOI22_X1 U8631 ( .A1(n10557), .A2(n7747), .B1(n11082), .B2(
        P1_REG0_REG_6__SCAN_IN), .ZN(n7221) );
  OAI21_X1 U8632 ( .B1(n7749), .B2(n11082), .A(n7221), .ZN(P1_U3471) );
  NAND2_X1 U8633 ( .A1(n9000), .A2(n7747), .ZN(n7223) );
  OR2_X1 U8634 ( .A1(n7443), .A2(n7115), .ZN(n7222) );
  NAND2_X1 U8635 ( .A1(n7223), .A2(n7222), .ZN(n7224) );
  XNOR2_X1 U8636 ( .A(n7224), .B(n8974), .ZN(n7227) );
  OR2_X1 U8637 ( .A1(n9001), .A2(n7443), .ZN(n7226) );
  NAND2_X1 U8638 ( .A1(n8961), .A2(n7747), .ZN(n7225) );
  AND2_X1 U8639 ( .A1(n7226), .A2(n7225), .ZN(n7228) );
  NAND2_X1 U8640 ( .A1(n7227), .A2(n7228), .ZN(n7428) );
  INV_X1 U8641 ( .A(n7227), .ZN(n7230) );
  INV_X1 U8642 ( .A(n7228), .ZN(n7229) );
  NAND2_X1 U8643 ( .A1(n7230), .A2(n7229), .ZN(n7231) );
  NAND2_X1 U8644 ( .A1(n7428), .A2(n7231), .ZN(n7245) );
  INV_X1 U8645 ( .A(n9817), .ZN(n7233) );
  AND2_X1 U8646 ( .A1(n7234), .A2(n7232), .ZN(n7240) );
  INV_X1 U8647 ( .A(n7234), .ZN(n7236) );
  NAND2_X1 U8648 ( .A1(n7236), .A2(n7235), .ZN(n7237) );
  AND2_X1 U8649 ( .A1(n7238), .A2(n7237), .ZN(n7239) );
  OR2_X1 U8650 ( .A1(n7240), .A2(n7239), .ZN(n7241) );
  INV_X1 U8651 ( .A(n7429), .ZN(n7243) );
  AOI21_X1 U8652 ( .B1(n7245), .B2(n7244), .A(n7243), .ZN(n7250) );
  AOI22_X1 U8653 ( .A1(n9846), .A2(n10168), .B1(n7747), .B2(n9863), .ZN(n7249)
         );
  INV_X1 U8654 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7246) );
  NOR2_X1 U8655 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7246), .ZN(n10252) );
  NOR2_X1 U8656 ( .A1(n9874), .A2(n7599), .ZN(n7247) );
  AOI211_X1 U8657 ( .C1(n9845), .C2(n10166), .A(n10252), .B(n7247), .ZN(n7248)
         );
  OAI211_X1 U8658 ( .C1(n7250), .C2(n9866), .A(n7249), .B(n7248), .ZN(P1_U3239) );
  INV_X1 U8659 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n7254) );
  NAND2_X1 U8660 ( .A1(n8678), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7253) );
  INV_X1 U8661 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n7251) );
  OR2_X1 U8662 ( .A1(n6338), .A2(n7251), .ZN(n7252) );
  OAI211_X1 U8663 ( .C1(n7254), .C2(n5110), .A(n7253), .B(n7252), .ZN(n7255)
         );
  INV_X1 U8664 ( .A(n7255), .ZN(n7256) );
  AND2_X1 U8665 ( .A1(n8686), .A2(n7256), .ZN(n9365) );
  NAND2_X1 U8666 ( .A1(n9331), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n7257) );
  OAI21_X1 U8667 ( .B1(n9365), .B2(n9331), .A(n7257), .ZN(P2_U3522) );
  NOR2_X1 U8668 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n7258) );
  AOI21_X1 U8669 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(P2_ADDR_REG_18__SCAN_IN), 
        .A(n7258), .ZN(n10659) );
  NOR2_X1 U8670 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7259) );
  AOI21_X1 U8671 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7259), .ZN(n10656) );
  NOR2_X1 U8672 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7260) );
  AOI21_X1 U8673 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7260), .ZN(n10653) );
  NOR2_X1 U8674 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7261) );
  AOI21_X1 U8675 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7261), .ZN(n10650) );
  NOR2_X1 U8676 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7262) );
  AOI21_X1 U8677 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7262), .ZN(n10647) );
  NOR2_X1 U8678 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7263) );
  AOI21_X1 U8679 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7263), .ZN(n10644) );
  NOR2_X1 U8680 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7264) );
  AOI21_X1 U8681 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7264), .ZN(n10641) );
  NOR2_X1 U8682 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7265) );
  AOI21_X1 U8683 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7265), .ZN(n10638) );
  NOR2_X1 U8684 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7266) );
  AOI21_X1 U8685 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7266), .ZN(n10635) );
  NOR2_X1 U8686 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7267) );
  AOI21_X1 U8687 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7267), .ZN(n10632) );
  NOR2_X1 U8688 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7268) );
  AOI21_X1 U8689 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7268), .ZN(n10629) );
  NOR2_X1 U8690 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7269) );
  AOI21_X1 U8691 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7269), .ZN(n10626) );
  NOR2_X1 U8692 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7270) );
  AOI21_X1 U8693 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7270), .ZN(n10623) );
  NOR2_X1 U8694 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7271) );
  AOI21_X1 U8695 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n7271), .ZN(n10620) );
  AND2_X1 U8696 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .ZN(n7272) );
  NOR2_X1 U8697 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7272), .ZN(n10605) );
  INV_X1 U8698 ( .A(n10605), .ZN(n10606) );
  NAND3_X1 U8699 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10607) );
  NAND2_X1 U8700 ( .A1(n10608), .A2(n10607), .ZN(n10604) );
  NAND2_X1 U8701 ( .A1(n10606), .A2(n10604), .ZN(n10611) );
  NAND2_X1 U8702 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7273) );
  OAI21_X1 U8703 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7273), .ZN(n10610) );
  NOR2_X1 U8704 ( .A1(n10611), .A2(n10610), .ZN(n10609) );
  AOI21_X1 U8705 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10609), .ZN(n10614) );
  NAND2_X1 U8706 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n7274) );
  OAI21_X1 U8707 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n7274), .ZN(n10613) );
  NOR2_X1 U8708 ( .A1(n10614), .A2(n10613), .ZN(n10612) );
  AOI21_X1 U8709 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10612), .ZN(n10617) );
  NOR2_X1 U8710 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7275) );
  AOI21_X1 U8711 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7275), .ZN(n10616) );
  NAND2_X1 U8712 ( .A1(n10617), .A2(n10616), .ZN(n10615) );
  OAI21_X1 U8713 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10615), .ZN(n10619) );
  NAND2_X1 U8714 ( .A1(n10620), .A2(n10619), .ZN(n10618) );
  OAI21_X1 U8715 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10618), .ZN(n10622) );
  NAND2_X1 U8716 ( .A1(n10623), .A2(n10622), .ZN(n10621) );
  OAI21_X1 U8717 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10621), .ZN(n10625) );
  NAND2_X1 U8718 ( .A1(n10626), .A2(n10625), .ZN(n10624) );
  OAI21_X1 U8719 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10624), .ZN(n10628) );
  NAND2_X1 U8720 ( .A1(n10629), .A2(n10628), .ZN(n10627) );
  OAI21_X1 U8721 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10627), .ZN(n10631) );
  NAND2_X1 U8722 ( .A1(n10632), .A2(n10631), .ZN(n10630) );
  OAI21_X1 U8723 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10630), .ZN(n10634) );
  NAND2_X1 U8724 ( .A1(n10635), .A2(n10634), .ZN(n10633) );
  OAI21_X1 U8725 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10633), .ZN(n10637) );
  NAND2_X1 U8726 ( .A1(n10638), .A2(n10637), .ZN(n10636) );
  OAI21_X1 U8727 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10636), .ZN(n10640) );
  NAND2_X1 U8728 ( .A1(n10641), .A2(n10640), .ZN(n10639) );
  OAI21_X1 U8729 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10639), .ZN(n10643) );
  NAND2_X1 U8730 ( .A1(n10644), .A2(n10643), .ZN(n10642) );
  OAI21_X1 U8731 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10642), .ZN(n10646) );
  NAND2_X1 U8732 ( .A1(n10647), .A2(n10646), .ZN(n10645) );
  OAI21_X1 U8733 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10645), .ZN(n10649) );
  NAND2_X1 U8734 ( .A1(n10650), .A2(n10649), .ZN(n10648) );
  OAI21_X1 U8735 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10648), .ZN(n10652) );
  NAND2_X1 U8736 ( .A1(n10653), .A2(n10652), .ZN(n10651) );
  OAI21_X1 U8737 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10651), .ZN(n10655) );
  NAND2_X1 U8738 ( .A1(n10656), .A2(n10655), .ZN(n10654) );
  OAI21_X1 U8739 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10654), .ZN(n10658) );
  NAND2_X1 U8740 ( .A1(n10659), .A2(n10658), .ZN(n10657) );
  OAI21_X1 U8741 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(P1_ADDR_REG_18__SCAN_IN), 
        .A(n10657), .ZN(n7278) );
  XNOR2_X1 U8742 ( .A(n7276), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7277) );
  XNOR2_X1 U8743 ( .A(n7278), .B(n7277), .ZN(ADD_1068_U4) );
  XNOR2_X1 U8744 ( .A(n10065), .B(n7279), .ZN(n10888) );
  INV_X1 U8745 ( .A(n10888), .ZN(n7299) );
  NAND2_X1 U8746 ( .A1(n7281), .A2(n7280), .ZN(n7282) );
  NAND2_X2 U8747 ( .A1(n7292), .A2(n11050), .ZN(n10915) );
  INV_X1 U8748 ( .A(n7458), .ZN(n7284) );
  NAND2_X1 U8749 ( .A1(n10915), .A2(n7284), .ZN(n7924) );
  INV_X1 U8750 ( .A(n7917), .ZN(n11033) );
  NAND2_X1 U8751 ( .A1(n10888), .A2(n11033), .ZN(n7289) );
  OAI21_X1 U8752 ( .B1(n7285), .B2(n9949), .A(n10905), .ZN(n7286) );
  NAND2_X1 U8753 ( .A1(n7286), .A2(n10402), .ZN(n7288) );
  AOI22_X1 U8754 ( .A1(n11027), .A2(n10171), .B1(n10169), .B2(n11026), .ZN(
        n7287) );
  AND3_X1 U8755 ( .A1(n7289), .A2(n7288), .A3(n7287), .ZN(n10885) );
  MUX2_X1 U8756 ( .A(n7290), .B(n10885), .S(n10915), .Z(n7298) );
  INV_X2 U8757 ( .A(n10915), .ZN(n11051) );
  NOR2_X2 U8758 ( .A1(n11051), .A2(n7291), .ZN(n11056) );
  INV_X1 U8759 ( .A(n7292), .ZN(n7293) );
  NAND2_X1 U8760 ( .A1(n7293), .A2(n10274), .ZN(n10335) );
  NAND2_X1 U8761 ( .A1(n9848), .A2(n7325), .ZN(n7294) );
  INV_X1 U8762 ( .A(n10438), .ZN(n11035) );
  NAND2_X1 U8763 ( .A1(n7294), .A2(n11035), .ZN(n7295) );
  OR2_X1 U8764 ( .A1(n7295), .A2(n10898), .ZN(n10883) );
  OAI22_X1 U8765 ( .A1(n10335), .A2(n10883), .B1(n10191), .B2(n11050), .ZN(
        n7296) );
  AOI21_X1 U8766 ( .B1(n11056), .B2(n9848), .A(n7296), .ZN(n7297) );
  OAI211_X1 U8767 ( .C1(n7299), .C2(n7924), .A(n7298), .B(n7297), .ZN(P1_U3291) );
  OR2_X1 U8768 ( .A1(n7300), .A2(n9961), .ZN(n7301) );
  NAND2_X1 U8769 ( .A1(n7302), .A2(n7301), .ZN(n10980) );
  INV_X1 U8770 ( .A(n10980), .ZN(n7316) );
  NAND2_X1 U8771 ( .A1(n7303), .A2(n9962), .ZN(n7304) );
  NOR2_X1 U8772 ( .A1(n7304), .A2(n9961), .ZN(n7541) );
  AND2_X1 U8773 ( .A1(n7304), .A2(n9961), .ZN(n7305) );
  OAI21_X1 U8774 ( .B1(n7541), .B2(n7305), .A(n10402), .ZN(n7309) );
  OAI22_X1 U8775 ( .A1(n7443), .A2(n10900), .B1(n7627), .B2(n10902), .ZN(n7306) );
  INV_X1 U8776 ( .A(n7306), .ZN(n7308) );
  NAND2_X1 U8777 ( .A1(n10980), .A2(n11033), .ZN(n7307) );
  NAND3_X1 U8778 ( .A1(n7309), .A2(n7308), .A3(n7307), .ZN(n10985) );
  NAND2_X1 U8779 ( .A1(n10985), .A2(n10915), .ZN(n7315) );
  OAI22_X1 U8780 ( .A1(n10915), .A2(n7310), .B1(n7442), .B2(n11050), .ZN(n7313) );
  OAI211_X1 U8781 ( .C1(n7311), .C2(n10983), .A(n11035), .B(n7546), .ZN(n10981) );
  NOR2_X1 U8782 ( .A1(n10981), .A2(n10335), .ZN(n7312) );
  AOI211_X1 U8783 ( .C1(n11056), .C2(n7433), .A(n7313), .B(n7312), .ZN(n7314)
         );
  OAI211_X1 U8784 ( .C1(n7316), .C2(n7924), .A(n7315), .B(n7314), .ZN(P1_U3286) );
  XNOR2_X1 U8785 ( .A(n7317), .B(n10069), .ZN(n10875) );
  OAI21_X1 U8786 ( .B1(n10069), .B2(n7319), .A(n7318), .ZN(n7323) );
  INV_X1 U8787 ( .A(n9906), .ZN(n7320) );
  INV_X1 U8788 ( .A(n10170), .ZN(n10901) );
  OAI22_X1 U8789 ( .A1(n7320), .A2(n10900), .B1(n10901), .B2(n10902), .ZN(
        n7322) );
  NOR2_X1 U8790 ( .A1(n10875), .A2(n7917), .ZN(n7321) );
  AOI211_X1 U8791 ( .C1(n10402), .C2(n7323), .A(n7322), .B(n7321), .ZN(n10877)
         );
  MUX2_X1 U8792 ( .A(n7324), .B(n10877), .S(n10915), .Z(n7328) );
  OAI211_X1 U8793 ( .C1(n9905), .C2(n5729), .A(n11035), .B(n7325), .ZN(n10876)
         );
  OAI22_X1 U8794 ( .A1(n10335), .A2(n10876), .B1(n10178), .B2(n11050), .ZN(
        n7326) );
  AOI21_X1 U8795 ( .B1(n11056), .B2(n5247), .A(n7326), .ZN(n7327) );
  OAI211_X1 U8796 ( .C1(n10875), .C2(n7924), .A(n7328), .B(n7327), .ZN(
        P1_U3292) );
  NAND2_X1 U8797 ( .A1(n7339), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7329) );
  NAND2_X1 U8798 ( .A1(n7330), .A2(n7329), .ZN(n7331) );
  AOI22_X1 U8799 ( .A1(P2_REG2_REG_4__SCAN_IN), .A2(n10837), .B1(n7338), .B2(
        n7392), .ZN(n10831) );
  NOR2_X1 U8800 ( .A1(n5126), .A2(n10831), .ZN(n10830) );
  NOR2_X1 U8801 ( .A1(n10830), .A2(n7333), .ZN(n7334) );
  NOR2_X1 U8802 ( .A1(n10847), .A2(n7334), .ZN(n7335) );
  NAND2_X1 U8803 ( .A1(P2_REG2_REG_6__SCAN_IN), .A2(n7557), .ZN(n7336) );
  OAI21_X1 U8804 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n7557), .A(n7336), .ZN(
        n7337) );
  AOI22_X1 U8805 ( .A1(P2_REG1_REG_4__SCAN_IN), .A2(n7338), .B1(n10837), .B2(
        n6337), .ZN(n10829) );
  INV_X1 U8806 ( .A(n7339), .ZN(n7356) );
  OAI21_X1 U8807 ( .B1(n7356), .B2(n7341), .A(n7340), .ZN(n7342) );
  NAND2_X1 U8808 ( .A1(n7359), .A2(n7342), .ZN(n7343) );
  XNOR2_X1 U8809 ( .A(n7342), .B(n10815), .ZN(n10812) );
  NAND2_X1 U8810 ( .A1(P2_REG1_REG_3__SCAN_IN), .A2(n10812), .ZN(n10811) );
  NAND2_X1 U8811 ( .A1(n7353), .A2(n7344), .ZN(n7345) );
  NAND2_X1 U8812 ( .A1(P2_REG1_REG_5__SCAN_IN), .A2(n10846), .ZN(n10845) );
  AOI22_X1 U8813 ( .A1(n7352), .A2(n7348), .B1(P2_REG1_REG_6__SCAN_IN), .B2(
        n7557), .ZN(n7346) );
  OAI21_X1 U8814 ( .B1(n7347), .B2(n7346), .A(n7558), .ZN(n7375) );
  INV_X1 U8815 ( .A(n10833), .ZN(n10849) );
  NOR2_X1 U8816 ( .A1(n9330), .A2(n7557), .ZN(n7374) );
  MUX2_X1 U8817 ( .A(n7349), .B(n7348), .S(n9327), .Z(n7351) );
  AND2_X1 U8818 ( .A1(n7351), .A2(n7352), .ZN(n7564) );
  INV_X1 U8819 ( .A(n7564), .ZN(n7350) );
  OAI21_X1 U8820 ( .B1(n7352), .B2(n7351), .A(n7350), .ZN(n7367) );
  MUX2_X1 U8821 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n9327), .Z(n7364) );
  NAND2_X1 U8822 ( .A1(n7364), .A2(n7353), .ZN(n7365) );
  MUX2_X1 U8823 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n9327), .Z(n7362) );
  INV_X1 U8824 ( .A(n7362), .ZN(n7363) );
  MUX2_X1 U8825 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n9327), .Z(n7360) );
  INV_X1 U8826 ( .A(n7360), .ZN(n7361) );
  INV_X1 U8827 ( .A(n7354), .ZN(n7355) );
  OAI22_X1 U8828 ( .A1(n7358), .A2(n7357), .B1(n7356), .B2(n7355), .ZN(n10821)
         );
  XNOR2_X1 U8829 ( .A(n7360), .B(n7359), .ZN(n10822) );
  NOR2_X1 U8830 ( .A1(n10821), .A2(n10822), .ZN(n10820) );
  AOI21_X1 U8831 ( .B1(n10815), .B2(n7361), .A(n10820), .ZN(n10840) );
  XNOR2_X1 U8832 ( .A(n7362), .B(n10837), .ZN(n10839) );
  NAND2_X1 U8833 ( .A1(n10840), .A2(n10839), .ZN(n10838) );
  XNOR2_X1 U8834 ( .A(n7364), .B(n10847), .ZN(n10861) );
  AOI21_X1 U8835 ( .B1(n7367), .B2(n7366), .A(n7563), .ZN(n7372) );
  INV_X1 U8836 ( .A(n7368), .ZN(n7371) );
  INV_X1 U8837 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7369) );
  OR2_X1 U8838 ( .A1(n10843), .A2(n7369), .ZN(n7370) );
  OAI211_X1 U8839 ( .C1(n7372), .C2(n10823), .A(n7371), .B(n7370), .ZN(n7373)
         );
  AOI211_X1 U8840 ( .C1(n7375), .C2(n10849), .A(n7374), .B(n7373), .ZN(n7376)
         );
  OAI21_X1 U8841 ( .B1(n7377), .B2(n10854), .A(n7376), .ZN(P2_U3188) );
  INV_X1 U8842 ( .A(n11050), .ZN(n10393) );
  INV_X1 U8843 ( .A(n10147), .ZN(n7379) );
  NOR3_X1 U8844 ( .A1(n10067), .A2(n7379), .A3(n7378), .ZN(n7380) );
  AOI211_X1 U8845 ( .C1(n10393), .C2(P1_REG3_REG_0__SCAN_IN), .A(n7381), .B(
        n7380), .ZN(n7385) );
  NOR2_X1 U8846 ( .A1(n10335), .A2(n10438), .ZN(n10285) );
  OAI21_X1 U8847 ( .B1(n10285), .B2(n11056), .A(n7382), .ZN(n7384) );
  NAND2_X1 U8848 ( .A1(n11051), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n7383) );
  OAI211_X1 U8849 ( .C1(n11051), .C2(n7385), .A(n7384), .B(n7383), .ZN(
        P1_U3293) );
  NAND2_X1 U8850 ( .A1(n10930), .A2(n7386), .ZN(n7387) );
  AND2_X1 U8851 ( .A1(n7388), .A2(n7387), .ZN(n7389) );
  AND2_X1 U8852 ( .A1(n8717), .A2(n7508), .ZN(n8714) );
  INV_X1 U8853 ( .A(n8714), .ZN(n8858) );
  XNOR2_X1 U8854 ( .A(n7389), .B(n8858), .ZN(n10947) );
  XNOR2_X1 U8855 ( .A(n7390), .B(n8858), .ZN(n7391) );
  AOI222_X1 U8856 ( .A1(n10928), .A2(n7391), .B1(n7171), .B2(n10926), .C1(
        n9204), .C2(n6677), .ZN(n10948) );
  MUX2_X1 U8857 ( .A(n7392), .B(n10948), .S(n10944), .Z(n7396) );
  INV_X1 U8858 ( .A(n7393), .ZN(n7394) );
  AOI22_X1 U8859 ( .A1(n9509), .A2(n10951), .B1(n9550), .B2(n7394), .ZN(n7395)
         );
  OAI211_X1 U8860 ( .C1(n9513), .C2(n10947), .A(n7396), .B(n7395), .ZN(
        P2_U3229) );
  XNOR2_X1 U8861 ( .A(n7661), .B(n9050), .ZN(n7399) );
  XNOR2_X1 U8862 ( .A(n7399), .B(n9202), .ZN(n7713) );
  NAND2_X1 U8863 ( .A1(n7397), .A2(n9203), .ZN(n7410) );
  AND2_X1 U8864 ( .A1(n7713), .A2(n7410), .ZN(n7398) );
  NAND2_X1 U8865 ( .A1(n7411), .A2(n7398), .ZN(n7498) );
  NAND2_X1 U8866 ( .A1(n7399), .A2(n7737), .ZN(n7491) );
  NAND2_X1 U8867 ( .A1(n7498), .A2(n7491), .ZN(n7401) );
  XNOR2_X1 U8868 ( .A(n10997), .B(n7079), .ZN(n7492) );
  XNOR2_X1 U8869 ( .A(n7492), .B(n9201), .ZN(n7400) );
  XNOR2_X1 U8870 ( .A(n7401), .B(n7400), .ZN(n7406) );
  NAND2_X1 U8871 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7703) );
  OAI21_X1 U8872 ( .B1(n9173), .B2(n7738), .A(n7703), .ZN(n7402) );
  AOI21_X1 U8873 ( .B1(n9152), .B2(n9202), .A(n7402), .ZN(n7403) );
  OAI21_X1 U8874 ( .B1(n7739), .B2(n9183), .A(n7403), .ZN(n7404) );
  AOI21_X1 U8875 ( .B1(n10997), .B2(n9190), .A(n7404), .ZN(n7405) );
  OAI21_X1 U8876 ( .B1(n7406), .B2(n9185), .A(n7405), .ZN(P2_U3161) );
  INV_X1 U8877 ( .A(n7407), .ZN(n7408) );
  OAI222_X1 U8878 ( .A1(n10274), .A2(P1_U3086), .B1(n8657), .B2(n7408), .C1(
        n8304), .C2(n10595), .ZN(P1_U3336) );
  OAI222_X1 U8879 ( .A1(n8618), .A2(n7409), .B1(n9719), .B2(n7408), .C1(n8892), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  OAI21_X1 U8880 ( .B1(n7714), .B2(n7713), .A(n7498), .ZN(n7412) );
  NAND2_X1 U8881 ( .A1(n7412), .A2(n9148), .ZN(n7416) );
  NAND2_X1 U8882 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7568) );
  OAI21_X1 U8883 ( .B1(n9173), .B2(n7814), .A(n7568), .ZN(n7414) );
  NOR2_X1 U8884 ( .A1(n9183), .A2(n7658), .ZN(n7413) );
  AOI211_X1 U8885 ( .C1(n9152), .C2(n9203), .A(n7414), .B(n7413), .ZN(n7415)
         );
  OAI211_X1 U8886 ( .C1(n10988), .C2(n9166), .A(n7416), .B(n7415), .ZN(
        P2_U3153) );
  OAI21_X1 U8887 ( .B1(n7418), .B2(n7425), .A(n7417), .ZN(n10459) );
  AOI21_X1 U8888 ( .B1(n7548), .B2(n10457), .A(n10438), .ZN(n7419) );
  NAND2_X1 U8889 ( .A1(n7419), .A2(n7451), .ZN(n7421) );
  OR2_X1 U8890 ( .A1(n7883), .A2(n10902), .ZN(n7420) );
  NAND2_X1 U8891 ( .A1(n7421), .A2(n7420), .ZN(n10460) );
  INV_X1 U8892 ( .A(n10077), .ZN(n7423) );
  OAI21_X1 U8893 ( .B1(n7541), .B2(n7423), .A(n7422), .ZN(n7424) );
  XOR2_X1 U8894 ( .A(n7425), .B(n7424), .Z(n7426) );
  OAI22_X1 U8895 ( .A1(n7426), .A2(n11030), .B1(n7627), .B2(n10900), .ZN(
        n10453) );
  AOI211_X1 U8896 ( .C1(n11078), .C2(n10459), .A(n10460), .B(n10453), .ZN(
        n7753) );
  AOI22_X1 U8897 ( .A1(n10557), .A2(n10457), .B1(n11082), .B2(
        P1_REG0_REG_9__SCAN_IN), .ZN(n7427) );
  OAI21_X1 U8898 ( .B1(n7753), .B2(n11082), .A(n7427), .ZN(P1_U3480) );
  NAND2_X1 U8899 ( .A1(n7433), .A2(n9000), .ZN(n7431) );
  OR2_X1 U8900 ( .A1(n7539), .A2(n7115), .ZN(n7430) );
  NAND2_X1 U8901 ( .A1(n7431), .A2(n7430), .ZN(n7432) );
  XNOR2_X1 U8902 ( .A(n7432), .B(n8974), .ZN(n7439) );
  INV_X1 U8903 ( .A(n7439), .ZN(n7437) );
  NAND2_X1 U8904 ( .A1(n7433), .A2(n8961), .ZN(n7435) );
  OR2_X1 U8905 ( .A1(n9001), .A2(n7539), .ZN(n7434) );
  AND2_X1 U8906 ( .A1(n7435), .A2(n7434), .ZN(n7438) );
  INV_X1 U8907 ( .A(n7438), .ZN(n7436) );
  NAND2_X1 U8908 ( .A1(n7437), .A2(n7436), .ZN(n7521) );
  NAND2_X1 U8909 ( .A1(n7439), .A2(n7438), .ZN(n7519) );
  NAND2_X1 U8910 ( .A1(n7521), .A2(n7519), .ZN(n7440) );
  XNOR2_X1 U8911 ( .A(n7520), .B(n7440), .ZN(n7441) );
  NAND2_X1 U8912 ( .A1(n7441), .A2(n9871), .ZN(n7448) );
  INV_X1 U8913 ( .A(n7442), .ZN(n7446) );
  NAND2_X1 U8914 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n10683) );
  INV_X1 U8915 ( .A(n10683), .ZN(n7445) );
  OAI22_X1 U8916 ( .A1(n7443), .A2(n9876), .B1(n9877), .B2(n7627), .ZN(n7444)
         );
  AOI211_X1 U8917 ( .C1(n9803), .C2(n7446), .A(n7445), .B(n7444), .ZN(n7447)
         );
  OAI211_X1 U8918 ( .C1(n10983), .C2(n9882), .A(n7448), .B(n7447), .ZN(
        P1_U3213) );
  OAI21_X1 U8919 ( .B1(n7450), .B2(n10079), .A(n7449), .ZN(n7586) );
  AOI211_X1 U8920 ( .C1(n7773), .C2(n7451), .A(n10438), .B(n11036), .ZN(n7591)
         );
  OAI21_X1 U8921 ( .B1(n5509), .B2(n7452), .A(n11022), .ZN(n7453) );
  NAND2_X1 U8922 ( .A1(n7453), .A2(n10402), .ZN(n7455) );
  AOI22_X1 U8923 ( .A1(n10164), .A2(n11027), .B1(n11026), .B2(n10163), .ZN(
        n7454) );
  NAND2_X1 U8924 ( .A1(n7455), .A2(n7454), .ZN(n7585) );
  AOI211_X1 U8925 ( .C1(n7586), .C2(n11078), .A(n7591), .B(n7585), .ZN(n7751)
         );
  AOI22_X1 U8926 ( .A1(n10557), .A2(n7773), .B1(n11082), .B2(
        P1_REG0_REG_10__SCAN_IN), .ZN(n7456) );
  OAI21_X1 U8927 ( .B1(n7751), .B2(n11082), .A(n7456), .ZN(P1_U3483) );
  XNOR2_X1 U8928 ( .A(n7457), .B(n10071), .ZN(n10958) );
  INV_X1 U8929 ( .A(n10958), .ZN(n7470) );
  AND2_X1 U8930 ( .A1(n7917), .A2(n7458), .ZN(n7459) );
  NAND3_X1 U8931 ( .A1(n10907), .A2(n9951), .A3(n10071), .ZN(n7460) );
  NAND2_X1 U8932 ( .A1(n7472), .A2(n7460), .ZN(n7461) );
  NAND2_X1 U8933 ( .A1(n7461), .A2(n10402), .ZN(n7463) );
  AOI22_X1 U8934 ( .A1(n11027), .A2(n10169), .B1(n10168), .B2(n11026), .ZN(
        n7462) );
  NAND2_X1 U8935 ( .A1(n7463), .A2(n7462), .ZN(n10956) );
  INV_X1 U8936 ( .A(n10897), .ZN(n7464) );
  OAI211_X1 U8937 ( .C1(n7464), .C2(n10955), .A(n11035), .B(n7478), .ZN(n10954) );
  NAND2_X1 U8938 ( .A1(n11056), .A2(n9820), .ZN(n7467) );
  INV_X1 U8939 ( .A(n9821), .ZN(n7465) );
  AOI22_X1 U8940 ( .A1(n11051), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7465), .B2(
        n10393), .ZN(n7466) );
  OAI211_X1 U8941 ( .C1(n10335), .C2(n10954), .A(n7467), .B(n7466), .ZN(n7468)
         );
  AOI21_X1 U8942 ( .B1(n10956), .B2(n10915), .A(n7468), .ZN(n7469) );
  OAI21_X1 U8943 ( .B1(n7470), .B2(n10452), .A(n7469), .ZN(P1_U3289) );
  XNOR2_X1 U8944 ( .A(n7471), .B(n9957), .ZN(n10967) );
  INV_X1 U8945 ( .A(n10967), .ZN(n7488) );
  NAND3_X1 U8946 ( .A1(n7472), .A2(n9950), .A3(n10072), .ZN(n7473) );
  NAND2_X1 U8947 ( .A1(n7474), .A2(n7473), .ZN(n7475) );
  NAND2_X1 U8948 ( .A1(n7475), .A2(n10402), .ZN(n7477) );
  AOI22_X1 U8949 ( .A1(n10167), .A2(n11026), .B1(n11027), .B2(n9745), .ZN(
        n7476) );
  NAND2_X1 U8950 ( .A1(n7477), .A2(n7476), .ZN(n10971) );
  NAND2_X1 U8951 ( .A1(n7478), .A2(n7482), .ZN(n7479) );
  NAND2_X1 U8952 ( .A1(n7479), .A2(n11035), .ZN(n7480) );
  OR2_X1 U8953 ( .A1(n7481), .A2(n7480), .ZN(n10968) );
  NAND2_X1 U8954 ( .A1(n11056), .A2(n7482), .ZN(n7485) );
  AOI22_X1 U8955 ( .A1(n11051), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7483), .B2(
        n10393), .ZN(n7484) );
  OAI211_X1 U8956 ( .C1(n10968), .C2(n10335), .A(n7485), .B(n7484), .ZN(n7486)
         );
  AOI21_X1 U8957 ( .B1(n10971), .B2(n10915), .A(n7486), .ZN(n7487) );
  OAI21_X1 U8958 ( .B1(n10452), .B2(n7488), .A(n7487), .ZN(P1_U3288) );
  INV_X1 U8959 ( .A(n7494), .ZN(n11000) );
  INV_X1 U8960 ( .A(n7492), .ZN(n7489) );
  NAND2_X1 U8961 ( .A1(n7489), .A2(n7814), .ZN(n7490) );
  AND2_X1 U8962 ( .A1(n7491), .A2(n7490), .ZN(n7497) );
  NAND2_X1 U8963 ( .A1(n7498), .A2(n7497), .ZN(n7493) );
  NAND2_X1 U8964 ( .A1(n7492), .A2(n9201), .ZN(n7499) );
  AND2_X1 U8965 ( .A1(n7493), .A2(n7499), .ZN(n7495) );
  XNOR2_X1 U8966 ( .A(n7494), .B(n7079), .ZN(n7710) );
  XNOR2_X1 U8967 ( .A(n7710), .B(n9200), .ZN(n7500) );
  AOI21_X1 U8968 ( .B1(n7495), .B2(n7500), .A(n9185), .ZN(n7502) );
  INV_X1 U8969 ( .A(n7500), .ZN(n7496) );
  AND2_X1 U8970 ( .A1(n7497), .A2(n7496), .ZN(n7715) );
  NAND2_X1 U8971 ( .A1(n7498), .A2(n7715), .ZN(n7721) );
  AND2_X1 U8972 ( .A1(n7721), .A2(n7712), .ZN(n7501) );
  NAND2_X1 U8973 ( .A1(n7502), .A2(n7501), .ZN(n7507) );
  INV_X1 U8974 ( .A(n7817), .ZN(n7505) );
  NOR2_X1 U8975 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8480), .ZN(n7851) );
  AOI21_X1 U8976 ( .B1(n9152), .B2(n9201), .A(n7851), .ZN(n7503) );
  OAI21_X1 U8977 ( .B1(n7962), .B2(n9173), .A(n7503), .ZN(n7504) );
  AOI21_X1 U8978 ( .B1(n7505), .B2(n9171), .A(n7504), .ZN(n7506) );
  OAI211_X1 U8979 ( .C1(n11000), .C2(n9166), .A(n7507), .B(n7506), .ZN(
        P2_U3171) );
  NAND2_X1 U8980 ( .A1(n7509), .A2(n7508), .ZN(n7510) );
  AND2_X1 U8981 ( .A1(n8725), .A2(n8719), .ZN(n8860) );
  XNOR2_X1 U8982 ( .A(n7510), .B(n8860), .ZN(n10962) );
  XNOR2_X1 U8983 ( .A(n7511), .B(n8860), .ZN(n7512) );
  AOI222_X1 U8984 ( .A1(n10928), .A2(n7512), .B1(n9203), .B2(n10926), .C1(
        n7154), .C2(n6677), .ZN(n10960) );
  MUX2_X1 U8985 ( .A(n7513), .B(n10960), .S(n10944), .Z(n7518) );
  INV_X1 U8986 ( .A(n7514), .ZN(n7515) );
  AOI22_X1 U8987 ( .A1(n9509), .A2(n7516), .B1(n9550), .B2(n7515), .ZN(n7517)
         );
  OAI211_X1 U8988 ( .C1(n9513), .C2(n10962), .A(n7518), .B(n7517), .ZN(
        P2_U3228) );
  NAND2_X1 U8989 ( .A1(n7522), .A2(n7521), .ZN(n7528) );
  NAND2_X1 U8990 ( .A1(n7549), .A2(n9000), .ZN(n7524) );
  OR2_X1 U8991 ( .A1(n7627), .A2(n7115), .ZN(n7523) );
  NAND2_X1 U8992 ( .A1(n7524), .A2(n7523), .ZN(n7525) );
  XNOR2_X1 U8993 ( .A(n7525), .B(n9002), .ZN(n7616) );
  NOR2_X1 U8994 ( .A1(n7627), .A2(n9001), .ZN(n7526) );
  AOI21_X1 U8995 ( .B1(n7549), .B2(n8938), .A(n7526), .ZN(n7617) );
  XNOR2_X1 U8996 ( .A(n7616), .B(n7617), .ZN(n7527) );
  NAND2_X1 U8997 ( .A1(n7528), .A2(n7527), .ZN(n7620) );
  OAI211_X1 U8998 ( .C1(n7528), .C2(n7527), .A(n7620), .B(n9871), .ZN(n7533)
         );
  INV_X1 U8999 ( .A(n7529), .ZN(n7609) );
  NAND2_X1 U9000 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n10697) );
  INV_X1 U9001 ( .A(n10697), .ZN(n7531) );
  OAI22_X1 U9002 ( .A1(n7539), .A2(n9876), .B1(n9877), .B2(n7770), .ZN(n7530)
         );
  AOI211_X1 U9003 ( .C1(n7609), .C2(n9803), .A(n7531), .B(n7530), .ZN(n7532)
         );
  OAI211_X1 U9004 ( .C1(n5326), .C2(n9882), .A(n7533), .B(n7532), .ZN(P1_U3221) );
  INV_X1 U9005 ( .A(n7534), .ZN(n7554) );
  OAI222_X1 U9006 ( .A1(P1_U3086), .A2(n7536), .B1(n8657), .B2(n7554), .C1(
        n7535), .C2(n10595), .ZN(P1_U3335) );
  INV_X1 U9007 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7553) );
  OAI21_X1 U9008 ( .B1(n7538), .B2(n9968), .A(n7537), .ZN(n7613) );
  INV_X1 U9009 ( .A(n7613), .ZN(n7551) );
  OAI22_X1 U9010 ( .A1(n7539), .A2(n10900), .B1(n7770), .B2(n10902), .ZN(n7545) );
  INV_X1 U9011 ( .A(n9966), .ZN(n7540) );
  NOR2_X1 U9012 ( .A1(n7541), .A2(n7540), .ZN(n7542) );
  XOR2_X1 U9013 ( .A(n9968), .B(n7542), .Z(n7543) );
  NOR2_X1 U9014 ( .A1(n7543), .A2(n11030), .ZN(n7544) );
  AOI211_X1 U9015 ( .C1(n11033), .C2(n7613), .A(n7545), .B(n7544), .ZN(n7615)
         );
  NAND2_X1 U9016 ( .A1(n7546), .A2(n7549), .ZN(n7547) );
  AND2_X1 U9017 ( .A1(n7548), .A2(n7547), .ZN(n7608) );
  AOI22_X1 U9018 ( .A1(n7608), .A2(n11035), .B1(n10541), .B2(n7549), .ZN(n7550) );
  OAI211_X1 U9019 ( .C1(n7551), .C2(n8045), .A(n7615), .B(n7550), .ZN(n7649)
         );
  NAND2_X1 U9020 ( .A1(n7649), .A2(n11085), .ZN(n7552) );
  OAI21_X1 U9021 ( .B1(n11085), .B2(n7553), .A(n7552), .ZN(P1_U3477) );
  OAI222_X1 U9022 ( .A1(n8618), .A2(n7555), .B1(P2_U3151), .B2(n8849), .C1(
        n9719), .C2(n7554), .ZN(P2_U3275) );
  XNOR2_X1 U9023 ( .A(n5306), .B(n7683), .ZN(n7556) );
  NOR2_X1 U9024 ( .A1(n7659), .A2(n7556), .ZN(n7685) );
  AOI21_X1 U9025 ( .B1(n7659), .B2(n7556), .A(n7685), .ZN(n7574) );
  NAND2_X1 U9026 ( .A1(P2_REG1_REG_6__SCAN_IN), .A2(n7557), .ZN(n7559) );
  NAND2_X1 U9027 ( .A1(P2_REG1_REG_7__SCAN_IN), .A2(n7560), .ZN(n7691) );
  OAI21_X1 U9028 ( .B1(P2_REG1_REG_7__SCAN_IN), .B2(n7560), .A(n7691), .ZN(
        n7572) );
  NOR2_X1 U9029 ( .A1(n9330), .A2(n7690), .ZN(n7571) );
  MUX2_X1 U9030 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n9327), .Z(n7561) );
  NOR2_X1 U9031 ( .A1(n7561), .A2(n7690), .ZN(n7697) );
  AOI21_X1 U9032 ( .B1(n7561), .B2(n7690), .A(n7697), .ZN(n7562) );
  INV_X1 U9033 ( .A(n7562), .ZN(n7566) );
  NOR2_X1 U9034 ( .A1(n7564), .A2(n7563), .ZN(n7565) );
  NOR2_X1 U9035 ( .A1(n7565), .A2(n7566), .ZN(n7696) );
  AOI21_X1 U9036 ( .B1(n7566), .B2(n7565), .A(n7696), .ZN(n7569) );
  NAND2_X1 U9037 ( .A1(n10858), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7567) );
  OAI211_X1 U9038 ( .C1(n7569), .C2(n10823), .A(n7568), .B(n7567), .ZN(n7570)
         );
  AOI211_X1 U9039 ( .C1(n7572), .C2(n10849), .A(n7571), .B(n7570), .ZN(n7573)
         );
  OAI21_X1 U9040 ( .B1(n7574), .B2(n10854), .A(n7573), .ZN(P2_U3189) );
  XNOR2_X1 U9041 ( .A(n7575), .B(n8861), .ZN(n7576) );
  OAI222_X1 U9042 ( .A1(n9564), .A2(n7737), .B1(n9562), .B2(n6364), .C1(n9559), 
        .C2(n7576), .ZN(n10975) );
  INV_X1 U9043 ( .A(n10975), .ZN(n7584) );
  NAND3_X1 U9044 ( .A1(n7578), .A2(n8725), .A3(n7577), .ZN(n7579) );
  NAND2_X1 U9045 ( .A1(n7651), .A2(n7579), .ZN(n10977) );
  NOR2_X1 U9046 ( .A1(n10939), .A2(n10974), .ZN(n7582) );
  OAI22_X1 U9047 ( .A1(n9589), .A2(n7349), .B1(n7580), .B2(n10937), .ZN(n7581)
         );
  AOI211_X1 U9048 ( .C1(n10977), .C2(n10941), .A(n7582), .B(n7581), .ZN(n7583)
         );
  OAI21_X1 U9049 ( .B1(n7584), .B2(n10946), .A(n7583), .ZN(P2_U3227) );
  INV_X1 U9050 ( .A(n7585), .ZN(n7594) );
  NAND2_X1 U9051 ( .A1(n7586), .A2(n10458), .ZN(n7593) );
  INV_X1 U9052 ( .A(n7773), .ZN(n7587) );
  NOR2_X1 U9053 ( .A1(n10440), .A2(n7587), .ZN(n7590) );
  OAI22_X1 U9054 ( .A1(n10915), .A2(n7588), .B1(n7769), .B2(n11050), .ZN(n7589) );
  AOI211_X1 U9055 ( .C1(n7591), .C2(n11045), .A(n7590), .B(n7589), .ZN(n7592)
         );
  OAI211_X1 U9056 ( .C1(n11051), .C2(n7594), .A(n7593), .B(n7592), .ZN(
        P1_U3283) );
  INV_X1 U9057 ( .A(n7595), .ZN(n7634) );
  OAI222_X1 U9058 ( .A1(P1_U3086), .A2(n10117), .B1(n8657), .B2(n7634), .C1(
        n7596), .C2(n10595), .ZN(P1_U3334) );
  INV_X1 U9059 ( .A(n7597), .ZN(n7607) );
  NAND2_X1 U9060 ( .A1(n7598), .A2(n11045), .ZN(n7602) );
  INV_X1 U9061 ( .A(n7599), .ZN(n7600) );
  AOI22_X1 U9062 ( .A1(n11051), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7600), .B2(
        n10393), .ZN(n7601) );
  OAI211_X1 U9063 ( .C1(n7603), .C2(n10440), .A(n7602), .B(n7601), .ZN(n7604)
         );
  AOI21_X1 U9064 ( .B1(n7605), .B2(n10458), .A(n7604), .ZN(n7606) );
  OAI21_X1 U9065 ( .B1(n7607), .B2(n11051), .A(n7606), .ZN(P1_U3287) );
  INV_X1 U9066 ( .A(n7924), .ZN(n11046) );
  NAND2_X1 U9067 ( .A1(n7608), .A2(n10285), .ZN(n7611) );
  AOI22_X1 U9068 ( .A1(n11051), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7609), .B2(
        n10393), .ZN(n7610) );
  OAI211_X1 U9069 ( .C1(n5326), .C2(n10440), .A(n7611), .B(n7610), .ZN(n7612)
         );
  AOI21_X1 U9070 ( .B1(n7613), .B2(n11046), .A(n7612), .ZN(n7614) );
  OAI21_X1 U9071 ( .B1(n7615), .B2(n11051), .A(n7614), .ZN(P1_U3285) );
  INV_X1 U9072 ( .A(n10457), .ZN(n7633) );
  INV_X1 U9073 ( .A(n7616), .ZN(n7618) );
  OR2_X1 U9074 ( .A1(n7618), .A2(n7617), .ZN(n7619) );
  NAND2_X1 U9075 ( .A1(n7620), .A2(n7619), .ZN(n7626) );
  NAND2_X1 U9076 ( .A1(n10457), .A2(n9000), .ZN(n7622) );
  OR2_X1 U9077 ( .A1(n7770), .A2(n7115), .ZN(n7621) );
  NAND2_X1 U9078 ( .A1(n7622), .A2(n7621), .ZN(n7623) );
  XNOR2_X1 U9079 ( .A(n7623), .B(n9002), .ZN(n7754) );
  NOR2_X1 U9080 ( .A1(n7770), .A2(n9001), .ZN(n7624) );
  AOI21_X1 U9081 ( .B1(n10457), .B2(n8938), .A(n7624), .ZN(n7755) );
  XNOR2_X1 U9082 ( .A(n7754), .B(n7755), .ZN(n7625) );
  NAND2_X1 U9083 ( .A1(n7626), .A2(n7625), .ZN(n7758) );
  OAI211_X1 U9084 ( .C1(n7626), .C2(n7625), .A(n7758), .B(n9871), .ZN(n7632)
         );
  INV_X1 U9085 ( .A(n10455), .ZN(n7630) );
  NAND2_X1 U9086 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n10805) );
  INV_X1 U9087 ( .A(n10805), .ZN(n7629) );
  OAI22_X1 U9088 ( .A1(n7627), .A2(n9876), .B1(n9877), .B2(n7883), .ZN(n7628)
         );
  AOI211_X1 U9089 ( .C1(n7630), .C2(n9803), .A(n7629), .B(n7628), .ZN(n7631)
         );
  OAI211_X1 U9090 ( .C1(n7633), .C2(n9882), .A(n7632), .B(n7631), .ZN(P1_U3231) );
  OAI222_X1 U9091 ( .A1(n8618), .A2(n7635), .B1(P2_U3151), .B2(n8879), .C1(
        n9719), .C2(n7634), .ZN(P2_U3274) );
  XOR2_X1 U9092 ( .A(n7636), .B(n10083), .Z(n11070) );
  INV_X1 U9093 ( .A(n11070), .ZN(n7648) );
  INV_X1 U9094 ( .A(n10083), .ZN(n7637) );
  XNOR2_X1 U9095 ( .A(n7638), .B(n7637), .ZN(n7639) );
  NAND2_X1 U9096 ( .A1(n7639), .A2(n10402), .ZN(n7641) );
  AOI22_X1 U9097 ( .A1(n11026), .A2(n10162), .B1(n10163), .B2(n11027), .ZN(
        n7640) );
  NAND2_X1 U9098 ( .A1(n7641), .A2(n7640), .ZN(n11069) );
  INV_X1 U9099 ( .A(n11034), .ZN(n7642) );
  INV_X1 U9100 ( .A(n7973), .ZN(n11067) );
  OAI211_X1 U9101 ( .C1(n7642), .C2(n11067), .A(n11035), .B(n7675), .ZN(n11066) );
  OAI22_X1 U9102 ( .A1(n10915), .A2(n7643), .B1(n7982), .B2(n11050), .ZN(n7644) );
  AOI21_X1 U9103 ( .B1(n7973), .B2(n11056), .A(n7644), .ZN(n7645) );
  OAI21_X1 U9104 ( .B1(n11066), .B2(n10335), .A(n7645), .ZN(n7646) );
  AOI21_X1 U9105 ( .B1(n11069), .B2(n10915), .A(n7646), .ZN(n7647) );
  OAI21_X1 U9106 ( .B1(n7648), .B2(n10452), .A(n7647), .ZN(P1_U3281) );
  NAND2_X1 U9107 ( .A1(n7649), .A2(n11081), .ZN(n7650) );
  OAI21_X1 U9108 ( .B1(n11081), .B2(n5826), .A(n7650), .ZN(P1_U3530) );
  INV_X1 U9109 ( .A(n7651), .ZN(n7653) );
  OAI21_X1 U9110 ( .B1(n7653), .B2(n7652), .A(n8865), .ZN(n7654) );
  NAND2_X1 U9111 ( .A1(n7654), .A2(n7733), .ZN(n10989) );
  INV_X1 U9112 ( .A(n9203), .ZN(n7657) );
  INV_X1 U9113 ( .A(n8865), .ZN(n8737) );
  XNOR2_X1 U9114 ( .A(n7655), .B(n8737), .ZN(n7656) );
  OAI222_X1 U9115 ( .A1(n9562), .A2(n7657), .B1(n9564), .B2(n7814), .C1(n9559), 
        .C2(n7656), .ZN(n10991) );
  NAND2_X1 U9116 ( .A1(n10991), .A2(n10944), .ZN(n7663) );
  OAI22_X1 U9117 ( .A1(n9589), .A2(n7659), .B1(n7658), .B2(n10937), .ZN(n7660)
         );
  AOI21_X1 U9118 ( .B1(n9509), .B2(n7661), .A(n7660), .ZN(n7662) );
  OAI211_X1 U9119 ( .C1(n9513), .C2(n10989), .A(n7663), .B(n7662), .ZN(
        P2_U3226) );
  INV_X1 U9120 ( .A(n7664), .ZN(n7667) );
  OAI222_X1 U9121 ( .A1(n10151), .A2(P1_U3086), .B1(n8657), .B2(n7667), .C1(
        n7665), .C2(n10595), .ZN(P1_U3333) );
  OAI222_X1 U9122 ( .A1(n8618), .A2(n7668), .B1(n9719), .B2(n7667), .C1(
        P2_U3151), .C2(n7666), .ZN(P2_U3273) );
  XOR2_X1 U9123 ( .A(n10085), .B(n7669), .Z(n11079) );
  INV_X1 U9124 ( .A(n11079), .ZN(n7682) );
  NAND2_X1 U9125 ( .A1(n7670), .A2(n10085), .ZN(n7671) );
  NAND2_X1 U9126 ( .A1(n7912), .A2(n7671), .ZN(n7672) );
  NAND2_X1 U9127 ( .A1(n7672), .A2(n10402), .ZN(n7674) );
  AOI22_X1 U9128 ( .A1(n11026), .A2(n10161), .B1(n11025), .B2(n11027), .ZN(
        n7673) );
  NAND2_X1 U9129 ( .A1(n7674), .A2(n7673), .ZN(n11077) );
  INV_X1 U9130 ( .A(n8029), .ZN(n11075) );
  INV_X1 U9131 ( .A(n7676), .ZN(n7918) );
  OAI211_X1 U9132 ( .C1(n11075), .C2(n6212), .A(n7918), .B(n11035), .ZN(n11073) );
  OAI22_X1 U9133 ( .A1(n10915), .A2(n7677), .B1(n8035), .B2(n11050), .ZN(n7678) );
  AOI21_X1 U9134 ( .B1(n8029), .B2(n11056), .A(n7678), .ZN(n7679) );
  OAI21_X1 U9135 ( .B1(n11073), .B2(n10335), .A(n7679), .ZN(n7680) );
  AOI21_X1 U9136 ( .B1(n11077), .B2(n10915), .A(n7680), .ZN(n7681) );
  OAI21_X1 U9137 ( .B1(n7682), .B2(n10452), .A(n7681), .ZN(P1_U3280) );
  NOR2_X1 U9138 ( .A1(n5306), .A2(n7683), .ZN(n7684) );
  NOR2_X1 U9139 ( .A1(n7685), .A2(n7684), .ZN(n7688) );
  AOI22_X1 U9140 ( .A1(n7799), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n7779), .B2(
        n7695), .ZN(n7687) );
  AOI21_X1 U9141 ( .B1(n7688), .B2(n7687), .A(n7686), .ZN(n7709) );
  NAND2_X1 U9142 ( .A1(n7690), .A2(n7689), .ZN(n7692) );
  NAND2_X1 U9143 ( .A1(n7692), .A2(n7691), .ZN(n7694) );
  MUX2_X1 U9144 ( .A(n7698), .B(P2_REG1_REG_8__SCAN_IN), .S(n7799), .Z(n7693)
         );
  NAND2_X1 U9145 ( .A1(n7693), .A2(n7694), .ZN(n7798) );
  OAI21_X1 U9146 ( .B1(n7694), .B2(n7693), .A(n7798), .ZN(n7707) );
  NOR2_X1 U9147 ( .A1(n9330), .A2(n7695), .ZN(n7706) );
  NOR2_X1 U9148 ( .A1(n7697), .A2(n7696), .ZN(n7701) );
  MUX2_X1 U9149 ( .A(n7779), .B(n7698), .S(n9327), .Z(n7699) );
  NAND2_X1 U9150 ( .A1(n7699), .A2(n7799), .ZN(n7786) );
  OAI21_X1 U9151 ( .B1(n7699), .B2(n7799), .A(n7786), .ZN(n7700) );
  AOI21_X1 U9152 ( .B1(n7701), .B2(n7700), .A(n7788), .ZN(n7704) );
  NAND2_X1 U9153 ( .A1(n10858), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7702) );
  OAI211_X1 U9154 ( .C1(n7704), .C2(n10823), .A(n7703), .B(n7702), .ZN(n7705)
         );
  AOI211_X1 U9155 ( .C1(n7707), .C2(n10849), .A(n7706), .B(n7705), .ZN(n7708)
         );
  OAI21_X1 U9156 ( .B1(n7709), .B2(n10854), .A(n7708), .ZN(P2_U3190) );
  NAND2_X1 U9157 ( .A1(n7710), .A2(n9200), .ZN(n7711) );
  OR2_X1 U9158 ( .A1(n7716), .A2(n7715), .ZN(n7717) );
  XNOR2_X1 U9159 ( .A(n11010), .B(n9050), .ZN(n7722) );
  INV_X1 U9160 ( .A(n7721), .ZN(n7725) );
  NOR2_X1 U9161 ( .A1(n7725), .A2(n7724), .ZN(n7726) );
  XNOR2_X1 U9162 ( .A(n11016), .B(n9050), .ZN(n7925) );
  XOR2_X1 U9163 ( .A(n9198), .B(n7925), .Z(n7927) );
  XOR2_X1 U9164 ( .A(n7928), .B(n7927), .Z(n7731) );
  NAND2_X1 U9165 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7903) );
  OAI21_X1 U9166 ( .B1(n9173), .B2(n7963), .A(n7903), .ZN(n7727) );
  AOI21_X1 U9167 ( .B1(n9152), .B2(n9199), .A(n7727), .ZN(n7728) );
  OAI21_X1 U9168 ( .B1(n7964), .B2(n9183), .A(n7728), .ZN(n7729) );
  AOI21_X1 U9169 ( .B1(n11016), .B2(n9190), .A(n7729), .ZN(n7730) );
  OAI21_X1 U9170 ( .B1(n7731), .B2(n9185), .A(n7730), .ZN(P2_U3176) );
  NAND2_X1 U9171 ( .A1(n7733), .A2(n7732), .ZN(n7734) );
  XOR2_X1 U9172 ( .A(n8863), .B(n7734), .Z(n10994) );
  XOR2_X1 U9173 ( .A(n7735), .B(n8863), .Z(n7736) );
  OAI222_X1 U9174 ( .A1(n9564), .A2(n7738), .B1(n9562), .B2(n7737), .C1(n9559), 
        .C2(n7736), .ZN(n10995) );
  NAND2_X1 U9175 ( .A1(n10995), .A2(n10944), .ZN(n7742) );
  OAI22_X1 U9176 ( .A1(n9589), .A2(n7779), .B1(n7739), .B2(n10937), .ZN(n7740)
         );
  AOI21_X1 U9177 ( .B1(n9509), .B2(n10997), .A(n7740), .ZN(n7741) );
  OAI211_X1 U9178 ( .C1(n10994), .C2(n9513), .A(n7742), .B(n7741), .ZN(
        P2_U3225) );
  INV_X1 U9179 ( .A(n7776), .ZN(n7746) );
  NOR2_X1 U9180 ( .A1(n7743), .A2(P1_U3086), .ZN(n10153) );
  AOI21_X1 U9181 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n7744), .A(n10153), .ZN(
        n7745) );
  OAI21_X1 U9182 ( .B1(n7746), .B2(n8657), .A(n7745), .ZN(P1_U3332) );
  AOI22_X1 U9183 ( .A1(n8052), .A2(n7747), .B1(n11080), .B2(
        P1_REG1_REG_6__SCAN_IN), .ZN(n7748) );
  OAI21_X1 U9184 ( .B1(n7749), .B2(n11080), .A(n7748), .ZN(P1_U3528) );
  AOI22_X1 U9185 ( .A1(n8052), .A2(n7773), .B1(n11080), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7750) );
  OAI21_X1 U9186 ( .B1(n7751), .B2(n11080), .A(n7750), .ZN(P1_U3532) );
  AOI22_X1 U9187 ( .A1(n8052), .A2(n10457), .B1(n11080), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n7752) );
  OAI21_X1 U9188 ( .B1(n7753), .B2(n11080), .A(n7752), .ZN(P1_U3531) );
  INV_X1 U9189 ( .A(n7754), .ZN(n7756) );
  OR2_X1 U9190 ( .A1(n7756), .A2(n7755), .ZN(n7757) );
  NAND2_X1 U9191 ( .A1(n7773), .A2(n9000), .ZN(n7761) );
  OR2_X1 U9192 ( .A1(n7883), .A2(n7115), .ZN(n7760) );
  NAND2_X1 U9193 ( .A1(n7761), .A2(n7760), .ZN(n7762) );
  XNOR2_X1 U9194 ( .A(n7762), .B(n9002), .ZN(n7765) );
  INV_X1 U9195 ( .A(n7765), .ZN(n7763) );
  NAND2_X1 U9196 ( .A1(n7766), .A2(n7765), .ZN(n7874) );
  NAND2_X1 U9197 ( .A1(n7875), .A2(n7874), .ZN(n7768) );
  NOR2_X1 U9198 ( .A1(n7883), .A2(n9001), .ZN(n7767) );
  AOI21_X1 U9199 ( .B1(n7773), .B2(n8938), .A(n7767), .ZN(n7873) );
  XNOR2_X1 U9200 ( .A(n7768), .B(n7873), .ZN(n7775) );
  NAND2_X1 U9201 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n10785) );
  OAI21_X1 U9202 ( .B1(n9874), .B2(n7769), .A(n10785), .ZN(n7772) );
  OAI22_X1 U9203 ( .A1(n7770), .A2(n9876), .B1(n9877), .B2(n7983), .ZN(n7771)
         );
  AOI211_X1 U9204 ( .C1(n7773), .C2(n9863), .A(n7772), .B(n7771), .ZN(n7774)
         );
  OAI21_X1 U9205 ( .B1(n7775), .B2(n9866), .A(n7774), .ZN(P1_U3217) );
  NAND2_X1 U9206 ( .A1(n7776), .A2(n5180), .ZN(n7777) );
  OAI211_X1 U9207 ( .C1(n7778), .C2(n8618), .A(n7777), .B(n8899), .ZN(P2_U3272) );
  XNOR2_X1 U9208 ( .A(n7781), .B(n7800), .ZN(n7848) );
  AND2_X1 U9209 ( .A1(n7781), .A2(n7800), .ZN(n7782) );
  MUX2_X1 U9210 ( .A(n7947), .B(P2_REG2_REG_10__SCAN_IN), .S(n7898), .Z(n7783)
         );
  INV_X1 U9211 ( .A(n7783), .ZN(n7784) );
  AOI21_X1 U9212 ( .B1(n7785), .B2(n7784), .A(n7899), .ZN(n7811) );
  MUX2_X1 U9213 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n9327), .Z(n7789) );
  NOR2_X1 U9214 ( .A1(n7789), .A2(n7800), .ZN(n7791) );
  INV_X1 U9215 ( .A(n7786), .ZN(n7787) );
  AOI21_X1 U9216 ( .B1(n7789), .B2(n7800), .A(n7791), .ZN(n7790) );
  INV_X1 U9217 ( .A(n7790), .ZN(n7856) );
  INV_X1 U9218 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7792) );
  MUX2_X1 U9219 ( .A(n7947), .B(n7792), .S(n9327), .Z(n7793) );
  NAND2_X1 U9220 ( .A1(n7793), .A2(n7898), .ZN(n7889) );
  MUX2_X1 U9221 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n9327), .Z(n7794) );
  AND2_X1 U9222 ( .A1(n7794), .A2(n7806), .ZN(n7891) );
  INV_X1 U9223 ( .A(n7891), .ZN(n7795) );
  NAND2_X1 U9224 ( .A1(n7889), .A2(n7795), .ZN(n7796) );
  XNOR2_X1 U9225 ( .A(n7890), .B(n7796), .ZN(n7797) );
  NAND2_X1 U9226 ( .A1(n7797), .A2(n10859), .ZN(n7810) );
  AOI22_X1 U9227 ( .A1(n7898), .A2(n7792), .B1(P2_REG1_REG_10__SCAN_IN), .B2(
        n7806), .ZN(n7804) );
  OAI21_X1 U9228 ( .B1(n7799), .B2(n7698), .A(n7798), .ZN(n7801) );
  NAND2_X1 U9229 ( .A1(n7801), .A2(n7800), .ZN(n7802) );
  XNOR2_X1 U9230 ( .A(n7801), .B(n7861), .ZN(n7850) );
  NAND2_X1 U9231 ( .A1(P2_REG1_REG_9__SCAN_IN), .A2(n7850), .ZN(n7849) );
  OAI21_X1 U9232 ( .B1(n7804), .B2(n7803), .A(n7894), .ZN(n7808) );
  NAND2_X1 U9233 ( .A1(n10858), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n7805) );
  NAND2_X1 U9234 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8634) );
  OAI211_X1 U9235 ( .C1(n9330), .C2(n7806), .A(n7805), .B(n8634), .ZN(n7807)
         );
  AOI21_X1 U9236 ( .B1(n7808), .B2(n10849), .A(n7807), .ZN(n7809) );
  OAI211_X1 U9237 ( .C1(n7811), .C2(n10854), .A(n7810), .B(n7809), .ZN(
        P2_U3192) );
  XOR2_X1 U9238 ( .A(n7812), .B(n8864), .Z(n7813) );
  OAI222_X1 U9239 ( .A1(n9564), .A2(n7962), .B1(n9562), .B2(n7814), .C1(n9559), 
        .C2(n7813), .ZN(n11001) );
  INV_X1 U9240 ( .A(n11001), .ZN(n7822) );
  OR2_X1 U9241 ( .A1(n7816), .A2(n8864), .ZN(n7938) );
  INV_X1 U9242 ( .A(n7938), .ZN(n7815) );
  AOI21_X1 U9243 ( .B1(n8864), .B2(n7816), .A(n7815), .ZN(n11003) );
  NOR2_X1 U9244 ( .A1(n11000), .A2(n10939), .ZN(n7820) );
  OAI22_X1 U9245 ( .A1(n9589), .A2(n7818), .B1(n7817), .B2(n10937), .ZN(n7819)
         );
  AOI211_X1 U9246 ( .C1(n11003), .C2(n10941), .A(n7820), .B(n7819), .ZN(n7821)
         );
  OAI21_X1 U9247 ( .B1(n7822), .B2(n10946), .A(n7821), .ZN(P2_U3224) );
  NOR2_X1 U9248 ( .A1(n10767), .A2(n7823), .ZN(n7824) );
  AOI21_X1 U9249 ( .B1(n10767), .B2(n7823), .A(n7824), .ZN(n10760) );
  OAI21_X1 U9250 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n7835), .A(n7825), .ZN(
        n10761) );
  NOR2_X1 U9251 ( .A1(n10760), .A2(n10761), .ZN(n10759) );
  AOI21_X1 U9252 ( .B1(n10767), .B2(P1_REG1_REG_13__SCAN_IN), .A(n10759), .ZN(
        n10723) );
  XNOR2_X1 U9253 ( .A(n10726), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n10724) );
  NOR2_X1 U9254 ( .A1(n10723), .A2(n10724), .ZN(n10722) );
  AOI21_X1 U9255 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n10726), .A(n10722), .ZN(
        n7826) );
  NOR2_X1 U9256 ( .A1(n7826), .A2(n7837), .ZN(n7827) );
  XNOR2_X1 U9257 ( .A(n7837), .B(n7826), .ZN(n10736) );
  NOR2_X1 U9258 ( .A1(n10735), .A2(n10736), .ZN(n10734) );
  NOR2_X1 U9259 ( .A1(n7827), .A2(n10734), .ZN(n7829) );
  AOI22_X1 U9260 ( .A1(n7866), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n8097), .B2(
        n7832), .ZN(n7828) );
  NAND2_X1 U9261 ( .A1(n7828), .A2(n7829), .ZN(n7865) );
  OAI21_X1 U9262 ( .B1(n7829), .B2(n7828), .A(n7865), .ZN(n7845) );
  NOR2_X1 U9263 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7830), .ZN(n9785) );
  AOI21_X1 U9264 ( .B1(n10666), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n9785), .ZN(
        n7831) );
  OAI21_X1 U9265 ( .B1(n10754), .B2(n7832), .A(n7831), .ZN(n7844) );
  NAND2_X1 U9266 ( .A1(n10767), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7833) );
  OAI21_X1 U9267 ( .B1(n10767), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7833), .ZN(
        n10763) );
  OAI21_X1 U9268 ( .B1(n7835), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7834), .ZN(
        n10764) );
  NOR2_X1 U9269 ( .A1(n10763), .A2(n10764), .ZN(n10762) );
  AOI21_X1 U9270 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n10767), .A(n10762), .ZN(
        n10717) );
  NAND2_X1 U9271 ( .A1(n10726), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7836) );
  OAI21_X1 U9272 ( .B1(n10726), .B2(P1_REG2_REG_14__SCAN_IN), .A(n7836), .ZN(
        n10718) );
  NOR2_X1 U9273 ( .A1(n10717), .A2(n10718), .ZN(n10719) );
  AOI21_X1 U9274 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n10726), .A(n10719), .ZN(
        n7838) );
  NOR2_X1 U9275 ( .A1(n7838), .A2(n7837), .ZN(n7839) );
  XNOR2_X1 U9276 ( .A(n7838), .B(n7837), .ZN(n10738) );
  NOR2_X1 U9277 ( .A1(n5943), .A2(n10738), .ZN(n10737) );
  NOR2_X1 U9278 ( .A1(n7839), .A2(n10737), .ZN(n7842) );
  NAND2_X1 U9279 ( .A1(n7866), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7840) );
  OAI21_X1 U9280 ( .B1(n7866), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7840), .ZN(
        n7841) );
  NOR2_X1 U9281 ( .A1(n7842), .A2(n7841), .ZN(n7864) );
  AOI211_X1 U9282 ( .C1(n7842), .C2(n7841), .A(n7864), .B(n10797), .ZN(n7843)
         );
  AOI211_X1 U9283 ( .C1(n10782), .C2(n7845), .A(n7844), .B(n7843), .ZN(n7846)
         );
  INV_X1 U9284 ( .A(n7846), .ZN(P1_U3259) );
  AOI21_X1 U9285 ( .B1(n7848), .B2(n7818), .A(n7847), .ZN(n7863) );
  INV_X1 U9286 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7854) );
  OAI21_X1 U9287 ( .B1(n7850), .B2(P2_REG1_REG_9__SCAN_IN), .A(n7849), .ZN(
        n7852) );
  AOI21_X1 U9288 ( .B1(n10849), .B2(n7852), .A(n7851), .ZN(n7853) );
  OAI21_X1 U9289 ( .B1(n7854), .B2(n10843), .A(n7853), .ZN(n7860) );
  AOI21_X1 U9290 ( .B1(n7857), .B2(n7856), .A(n7855), .ZN(n7858) );
  NOR2_X1 U9291 ( .A1(n7858), .A2(n10823), .ZN(n7859) );
  AOI211_X1 U9292 ( .C1(n10848), .C2(n7861), .A(n7860), .B(n7859), .ZN(n7862)
         );
  OAI21_X1 U9293 ( .B1(n7863), .B2(n10854), .A(n7862), .ZN(P2_U3191) );
  XNOR2_X1 U9294 ( .A(n7867), .B(n10258), .ZN(n10259) );
  AOI21_X1 U9295 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n7866), .A(n7864), .ZN(
        n10260) );
  XOR2_X1 U9296 ( .A(n10259), .B(n10260), .Z(n7872) );
  OAI21_X1 U9297 ( .B1(n7866), .B2(P1_REG1_REG_16__SCAN_IN), .A(n7865), .ZN(
        n10270) );
  XNOR2_X1 U9298 ( .A(n7867), .B(n10268), .ZN(n10269) );
  XNOR2_X1 U9299 ( .A(n10270), .B(n10269), .ZN(n7870) );
  AND2_X1 U9300 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9801) );
  AOI21_X1 U9301 ( .B1(n10666), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n9801), .ZN(
        n7868) );
  OAI21_X1 U9302 ( .B1(n10754), .B2(n10267), .A(n7868), .ZN(n7869) );
  AOI21_X1 U9303 ( .B1(n7870), .B2(n10782), .A(n7869), .ZN(n7871) );
  OAI21_X1 U9304 ( .B1(n7872), .B2(n10797), .A(n7871), .ZN(P1_U3260) );
  NAND2_X1 U9305 ( .A1(n7874), .A2(n7873), .ZN(n7876) );
  NAND2_X1 U9306 ( .A1(n7876), .A2(n7875), .ZN(n7974) );
  NAND2_X1 U9307 ( .A1(n11055), .A2(n9000), .ZN(n7878) );
  NAND2_X1 U9308 ( .A1(n8961), .A2(n10163), .ZN(n7877) );
  NAND2_X1 U9309 ( .A1(n7878), .A2(n7877), .ZN(n7879) );
  XNOR2_X1 U9310 ( .A(n7879), .B(n8974), .ZN(n7976) );
  AND2_X1 U9311 ( .A1(n8976), .A2(n10163), .ZN(n7880) );
  AOI21_X1 U9312 ( .B1(n11055), .B2(n8938), .A(n7880), .ZN(n7975) );
  INV_X1 U9313 ( .A(n7975), .ZN(n7977) );
  XNOR2_X1 U9314 ( .A(n7976), .B(n7977), .ZN(n7881) );
  XNOR2_X1 U9315 ( .A(n7974), .B(n7881), .ZN(n7882) );
  NAND2_X1 U9316 ( .A1(n7882), .A2(n9871), .ZN(n7888) );
  INV_X1 U9317 ( .A(n11049), .ZN(n7886) );
  NAND2_X1 U9318 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n10714) );
  INV_X1 U9319 ( .A(n10714), .ZN(n7885) );
  OAI22_X1 U9320 ( .A1(n8036), .A2(n9877), .B1(n9876), .B2(n7883), .ZN(n7884)
         );
  AOI211_X1 U9321 ( .C1(n9803), .C2(n7886), .A(n7885), .B(n7884), .ZN(n7887)
         );
  OAI211_X1 U9322 ( .C1(n11037), .C2(n9882), .A(n7888), .B(n7887), .ZN(
        P1_U3236) );
  OAI21_X1 U9323 ( .B1(n7891), .B2(n7890), .A(n7889), .ZN(n7893) );
  MUX2_X1 U9324 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n9327), .Z(n8075) );
  XNOR2_X1 U9325 ( .A(n8075), .B(n7895), .ZN(n7892) );
  OAI21_X1 U9326 ( .B1(n7893), .B2(n7892), .A(n8076), .ZN(n7909) );
  NAND2_X1 U9327 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(n7896), .ZN(n8061) );
  OAI21_X1 U9328 ( .B1(n7896), .B2(P2_REG1_REG_11__SCAN_IN), .A(n8061), .ZN(
        n7897) );
  NAND2_X1 U9329 ( .A1(n7897), .A2(n10849), .ZN(n7907) );
  OR2_X1 U9330 ( .A1(n7898), .A2(n7947), .ZN(n7901) );
  NAND2_X1 U9331 ( .A1(n7901), .A2(n7900), .ZN(n8065) );
  AOI21_X1 U9332 ( .B1(n7965), .B2(n7902), .A(n8067), .ZN(n7904) );
  OAI21_X1 U9333 ( .B1(n10854), .B2(n7904), .A(n7903), .ZN(n7905) );
  AOI21_X1 U9334 ( .B1(n10858), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n7905), .ZN(
        n7906) );
  OAI211_X1 U9335 ( .C1(n9330), .C2(n8074), .A(n7907), .B(n7906), .ZN(n7908)
         );
  AOI21_X1 U9336 ( .B1(n7909), .B2(n10859), .A(n7908), .ZN(n7910) );
  INV_X1 U9337 ( .A(n7910), .ZN(P2_U3193) );
  INV_X1 U9338 ( .A(n10086), .ZN(n9992) );
  XNOR2_X1 U9339 ( .A(n7911), .B(n9992), .ZN(n8046) );
  AOI22_X1 U9340 ( .A1(n10160), .A2(n11026), .B1(n11027), .B2(n10162), .ZN(
        n7916) );
  NAND2_X1 U9341 ( .A1(n7912), .A2(n9989), .ZN(n7913) );
  XNOR2_X1 U9342 ( .A(n7913), .B(n9992), .ZN(n7914) );
  NAND2_X1 U9343 ( .A1(n7914), .A2(n10402), .ZN(n7915) );
  OAI211_X1 U9344 ( .C1(n8046), .C2(n7917), .A(n7916), .B(n7915), .ZN(n8047)
         );
  NAND2_X1 U9345 ( .A1(n8047), .A2(n10915), .ZN(n7923) );
  AOI211_X1 U9346 ( .C1(n8128), .C2(n7918), .A(n10438), .B(n8623), .ZN(n8048)
         );
  NOR2_X1 U9347 ( .A1(n8056), .A2(n10440), .ZN(n7921) );
  OAI22_X1 U9348 ( .A1(n10915), .A2(n7919), .B1(n8124), .B2(n11050), .ZN(n7920) );
  AOI211_X1 U9349 ( .C1(n8048), .C2(n11045), .A(n7921), .B(n7920), .ZN(n7922)
         );
  OAI211_X1 U9350 ( .C1(n8046), .C2(n7924), .A(n7923), .B(n7922), .ZN(P1_U3279) );
  INV_X1 U9351 ( .A(n7925), .ZN(n7926) );
  XNOR2_X1 U9352 ( .A(n8018), .B(n9050), .ZN(n7929) );
  XOR2_X1 U9353 ( .A(n9578), .B(n7929), .Z(n7954) );
  INV_X1 U9354 ( .A(n7929), .ZN(n7930) );
  XNOR2_X1 U9355 ( .A(n9581), .B(n7079), .ZN(n7931) );
  NAND2_X1 U9356 ( .A1(n7931), .A2(n9197), .ZN(n8001) );
  NAND2_X1 U9357 ( .A1(n5175), .A2(n8001), .ZN(n7932) );
  XNOR2_X1 U9358 ( .A(n8002), .B(n7932), .ZN(n7937) );
  NAND2_X1 U9359 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n9210) );
  OAI21_X1 U9360 ( .B1(n9173), .B2(n9179), .A(n9210), .ZN(n7933) );
  AOI21_X1 U9361 ( .B1(n9152), .B2(n9578), .A(n7933), .ZN(n7934) );
  OAI21_X1 U9362 ( .B1(n9582), .B2(n9183), .A(n7934), .ZN(n7935) );
  AOI21_X1 U9363 ( .B1(n9581), .B2(n9190), .A(n7935), .ZN(n7936) );
  OAI21_X1 U9364 ( .B1(n7937), .B2(n9185), .A(n7936), .ZN(P2_U3174) );
  NAND2_X1 U9365 ( .A1(n7938), .A2(n8733), .ZN(n7941) );
  NAND2_X1 U9366 ( .A1(n7940), .A2(n7939), .ZN(n8867) );
  XNOR2_X1 U9367 ( .A(n7941), .B(n8867), .ZN(n11007) );
  NAND2_X1 U9368 ( .A1(n9589), .A2(n7942), .ZN(n9025) );
  XOR2_X1 U9369 ( .A(n7943), .B(n8867), .Z(n7944) );
  NAND2_X1 U9370 ( .A1(n7944), .A2(n10928), .ZN(n7946) );
  AOI22_X1 U9371 ( .A1(n10926), .A2(n9198), .B1(n9200), .B2(n6677), .ZN(n7945)
         );
  OAI211_X1 U9372 ( .C1(n9021), .C2(n11007), .A(n7946), .B(n7945), .ZN(n11008)
         );
  NAND2_X1 U9373 ( .A1(n11008), .A2(n10944), .ZN(n7950) );
  OAI22_X1 U9374 ( .A1(n9589), .A2(n7947), .B1(n8638), .B2(n10937), .ZN(n7948)
         );
  AOI21_X1 U9375 ( .B1(n11010), .B2(n9509), .A(n7948), .ZN(n7949) );
  OAI211_X1 U9376 ( .C1(n11007), .C2(n9025), .A(n7950), .B(n7949), .ZN(
        P2_U3223) );
  NAND2_X1 U9377 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8071) );
  OAI21_X1 U9378 ( .B1(n9173), .B2(n9561), .A(n8071), .ZN(n7951) );
  AOI21_X1 U9379 ( .B1(n9152), .B2(n9198), .A(n7951), .ZN(n7952) );
  OAI21_X1 U9380 ( .B1(n8008), .B2(n9183), .A(n7952), .ZN(n7956) );
  AOI211_X1 U9381 ( .C1(n7954), .C2(n7953), .A(n9185), .B(n5170), .ZN(n7955)
         );
  AOI211_X1 U9382 ( .C1(n8018), .C2(n9190), .A(n7956), .B(n7955), .ZN(n7957)
         );
  INV_X1 U9383 ( .A(n7957), .ZN(P2_U3164) );
  INV_X1 U9384 ( .A(n7958), .ZN(n8057) );
  OAI222_X1 U9385 ( .A1(n10595), .A2(n8508), .B1(P1_U3086), .B2(n7959), .C1(
        n8057), .C2(n8657), .ZN(P1_U3331) );
  XOR2_X1 U9386 ( .A(n8015), .B(n8869), .Z(n11013) );
  XNOR2_X1 U9387 ( .A(n7960), .B(n8869), .ZN(n7961) );
  OAI222_X1 U9388 ( .A1(n9564), .A2(n7963), .B1(n9562), .B2(n7962), .C1(n9559), 
        .C2(n7961), .ZN(n11014) );
  NAND2_X1 U9389 ( .A1(n11014), .A2(n10944), .ZN(n7968) );
  OAI22_X1 U9390 ( .A1(n9589), .A2(n7965), .B1(n7964), .B2(n10937), .ZN(n7966)
         );
  AOI21_X1 U9391 ( .B1(n11016), .B2(n9509), .A(n7966), .ZN(n7967) );
  OAI211_X1 U9392 ( .C1(n9513), .C2(n11013), .A(n7968), .B(n7967), .ZN(
        P2_U3222) );
  NAND2_X1 U9393 ( .A1(n7973), .A2(n9000), .ZN(n7970) );
  NAND2_X1 U9394 ( .A1(n8961), .A2(n11025), .ZN(n7969) );
  NAND2_X1 U9395 ( .A1(n7970), .A2(n7969), .ZN(n7971) );
  XNOR2_X1 U9396 ( .A(n7971), .B(n9002), .ZN(n8022) );
  AND2_X1 U9397 ( .A1(n8976), .A2(n11025), .ZN(n7972) );
  AOI21_X1 U9398 ( .B1(n7973), .B2(n8938), .A(n7972), .ZN(n8023) );
  XNOR2_X1 U9399 ( .A(n8022), .B(n8023), .ZN(n7980) );
  INV_X1 U9400 ( .A(n7976), .ZN(n7978) );
  OAI21_X1 U9401 ( .B1(n7980), .B2(n7979), .A(n8032), .ZN(n7981) );
  NAND2_X1 U9402 ( .A1(n7981), .A2(n9871), .ZN(n7988) );
  INV_X1 U9403 ( .A(n7982), .ZN(n7986) );
  OAI22_X1 U9404 ( .A1(n8125), .A2(n9877), .B1(n9876), .B2(n7983), .ZN(n7984)
         );
  AOI211_X1 U9405 ( .C1(n9803), .C2(n7986), .A(n7985), .B(n7984), .ZN(n7987)
         );
  OAI211_X1 U9406 ( .C1(n11067), .C2(n9882), .A(n7988), .B(n7987), .ZN(
        P1_U3224) );
  XNOR2_X1 U9407 ( .A(n7989), .B(n5550), .ZN(n7991) );
  OAI22_X1 U9408 ( .A1(n9860), .A2(n10902), .B1(n9787), .B2(n10900), .ZN(n7990) );
  AOI21_X1 U9409 ( .B1(n7991), .B2(n10402), .A(n7990), .ZN(n8094) );
  NAND2_X1 U9410 ( .A1(n7992), .A2(n10089), .ZN(n7993) );
  AND2_X1 U9411 ( .A1(n7994), .A2(n7993), .ZN(n8096) );
  NAND2_X1 U9412 ( .A1(n8096), .A2(n10458), .ZN(n8000) );
  OAI22_X1 U9413 ( .A1(n10915), .A2(n7995), .B1(n9784), .B2(n11050), .ZN(n7998) );
  AOI21_X1 U9414 ( .B1(n8624), .B2(n9789), .A(n10438), .ZN(n7996) );
  NAND2_X1 U9415 ( .A1(n7996), .A2(n8088), .ZN(n8093) );
  NOR2_X1 U9416 ( .A1(n8093), .A2(n10335), .ZN(n7997) );
  AOI211_X1 U9417 ( .C1(n11056), .C2(n9789), .A(n7998), .B(n7997), .ZN(n7999)
         );
  OAI211_X1 U9418 ( .C1(n11051), .C2(n8094), .A(n8000), .B(n7999), .ZN(
        P1_U3277) );
  XNOR2_X1 U9419 ( .A(n8773), .B(n9050), .ZN(n9031) );
  XOR2_X1 U9420 ( .A(n9577), .B(n9031), .Z(n9033) );
  XOR2_X1 U9421 ( .A(n9033), .B(n9034), .Z(n8007) );
  NAND2_X1 U9422 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n9236) );
  OAI21_X1 U9423 ( .B1(n9173), .B2(n9563), .A(n9236), .ZN(n8003) );
  AOI21_X1 U9424 ( .B1(n9152), .B2(n9197), .A(n8003), .ZN(n8004) );
  OAI21_X1 U9425 ( .B1(n9565), .B2(n9183), .A(n8004), .ZN(n8005) );
  AOI21_X1 U9426 ( .B1(n8773), .B2(n9190), .A(n8005), .ZN(n8006) );
  OAI21_X1 U9427 ( .B1(n8007), .B2(n9185), .A(n8006), .ZN(P2_U3155) );
  INV_X1 U9428 ( .A(n8008), .ZN(n8014) );
  AND2_X1 U9429 ( .A1(n8766), .A2(n8765), .ZN(n8868) );
  INV_X1 U9430 ( .A(n8868), .ZN(n8009) );
  XNOR2_X1 U9431 ( .A(n8010), .B(n8009), .ZN(n8011) );
  NAND2_X1 U9432 ( .A1(n8011), .A2(n10928), .ZN(n8013) );
  AOI22_X1 U9433 ( .A1(n6677), .A2(n9198), .B1(n9197), .B2(n10926), .ZN(n8012)
         );
  NAND2_X1 U9434 ( .A1(n8013), .A2(n8012), .ZN(n11063) );
  AOI21_X1 U9435 ( .B1(n9550), .B2(n8014), .A(n11063), .ZN(n8021) );
  NAND2_X1 U9436 ( .A1(n8015), .A2(n8869), .ZN(n8016) );
  NAND2_X1 U9437 ( .A1(n8016), .A2(n8759), .ZN(n8017) );
  XNOR2_X1 U9438 ( .A(n8017), .B(n8868), .ZN(n11059) );
  INV_X1 U9439 ( .A(n8018), .ZN(n11061) );
  OAI22_X1 U9440 ( .A1(n11061), .A2(n10939), .B1(n8068), .B2(n10944), .ZN(
        n8019) );
  AOI21_X1 U9441 ( .B1(n11059), .B2(n10941), .A(n8019), .ZN(n8020) );
  OAI21_X1 U9442 ( .B1(n8021), .B2(n10946), .A(n8020), .ZN(P2_U3221) );
  INV_X1 U9443 ( .A(n8022), .ZN(n8024) );
  NAND2_X1 U9444 ( .A1(n8024), .A2(n8023), .ZN(n8030) );
  AND2_X1 U9445 ( .A1(n8032), .A2(n8030), .ZN(n8034) );
  NAND2_X1 U9446 ( .A1(n8029), .A2(n9000), .ZN(n8026) );
  NAND2_X1 U9447 ( .A1(n8938), .A2(n10162), .ZN(n8025) );
  NAND2_X1 U9448 ( .A1(n8026), .A2(n8025), .ZN(n8027) );
  XNOR2_X1 U9449 ( .A(n8027), .B(n9002), .ZN(n8113) );
  AND2_X1 U9450 ( .A1(n8976), .A2(n10162), .ZN(n8028) );
  AOI21_X1 U9451 ( .B1(n8029), .B2(n8938), .A(n8028), .ZN(n8111) );
  XNOR2_X1 U9452 ( .A(n8113), .B(n8111), .ZN(n8033) );
  AND2_X1 U9453 ( .A1(n8033), .A2(n8030), .ZN(n8031) );
  OAI211_X1 U9454 ( .C1(n8034), .C2(n8033), .A(n9871), .B(n8122), .ZN(n8041)
         );
  INV_X1 U9455 ( .A(n8035), .ZN(n8039) );
  NAND2_X1 U9456 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n10768) );
  INV_X1 U9457 ( .A(n10768), .ZN(n8038) );
  OAI22_X1 U9458 ( .A1(n8622), .A2(n9877), .B1(n9876), .B2(n8036), .ZN(n8037)
         );
  AOI211_X1 U9459 ( .C1(n9803), .C2(n8039), .A(n8038), .B(n8037), .ZN(n8040)
         );
  OAI211_X1 U9460 ( .C1(n11075), .C2(n9882), .A(n8041), .B(n8040), .ZN(
        P1_U3234) );
  INV_X1 U9461 ( .A(n8042), .ZN(n8616) );
  OAI222_X1 U9462 ( .A1(n8044), .A2(P1_U3086), .B1(n8657), .B2(n8616), .C1(
        n8043), .C2(n10595), .ZN(P1_U3330) );
  INV_X1 U9463 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n8050) );
  INV_X1 U9464 ( .A(n8045), .ZN(n11039) );
  INV_X1 U9465 ( .A(n8046), .ZN(n8049) );
  AOI211_X1 U9466 ( .C1(n11039), .C2(n8049), .A(n8048), .B(n8047), .ZN(n8053)
         );
  MUX2_X1 U9467 ( .A(n8050), .B(n8053), .S(n11085), .Z(n8051) );
  OAI21_X1 U9468 ( .B1(n8056), .B2(n10579), .A(n8051), .ZN(P1_U3495) );
  MUX2_X1 U9469 ( .A(n8054), .B(n8053), .S(n10529), .Z(n8055) );
  OAI21_X1 U9470 ( .B1(n8056), .B2(n10532), .A(n8055), .ZN(P1_U3536) );
  OAI222_X1 U9471 ( .A1(n8618), .A2(n8059), .B1(P2_U3151), .B2(n8058), .C1(
        n9719), .C2(n8057), .ZN(P2_U3271) );
  AOI22_X1 U9472 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n9213), .B1(n9206), .B2(
        n6461), .ZN(n8064) );
  NAND2_X1 U9473 ( .A1(n8060), .A2(n8074), .ZN(n8062) );
  OAI21_X1 U9474 ( .B1(n8064), .B2(n8063), .A(n9205), .ZN(n8084) );
  AND2_X1 U9475 ( .A1(n8065), .A2(n8074), .ZN(n8066) );
  NOR2_X1 U9476 ( .A1(n9213), .A2(n8068), .ZN(n8069) );
  AOI21_X1 U9477 ( .B1(n8068), .B2(n9213), .A(n8069), .ZN(n8070) );
  AOI21_X1 U9478 ( .B1(n5168), .B2(n8070), .A(n9208), .ZN(n8072) );
  OAI21_X1 U9479 ( .B1(n10854), .B2(n8072), .A(n8071), .ZN(n8073) );
  AOI21_X1 U9480 ( .B1(n10858), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n8073), .ZN(
        n8082) );
  MUX2_X1 U9481 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n9327), .Z(n9214) );
  XNOR2_X1 U9482 ( .A(n9214), .B(n9206), .ZN(n8079) );
  OR2_X1 U9483 ( .A1(n8075), .A2(n8074), .ZN(n8077) );
  OAI21_X1 U9484 ( .B1(n8079), .B2(n8078), .A(n9215), .ZN(n8080) );
  NAND2_X1 U9485 ( .A1(n8080), .A2(n10859), .ZN(n8081) );
  OAI211_X1 U9486 ( .C1(n9330), .C2(n9213), .A(n8082), .B(n8081), .ZN(n8083)
         );
  AOI21_X1 U9487 ( .B1(n8084), .B2(n10849), .A(n8083), .ZN(n8085) );
  INV_X1 U9488 ( .A(n8085), .ZN(P2_U3194) );
  XNOR2_X1 U9489 ( .A(n8086), .B(n10012), .ZN(n10537) );
  XNOR2_X1 U9490 ( .A(n8139), .B(n10012), .ZN(n8087) );
  OAI222_X1 U9491 ( .A1(n10900), .A2(n9798), .B1(n10902), .B2(n9799), .C1(
        n8087), .C2(n11030), .ZN(n10533) );
  AOI211_X1 U9492 ( .C1(n10535), .C2(n8088), .A(n10438), .B(n5166), .ZN(n10534) );
  NAND2_X1 U9493 ( .A1(n10534), .A2(n11045), .ZN(n8090) );
  AOI22_X1 U9494 ( .A1(n11051), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n10393), 
        .B2(n9802), .ZN(n8089) );
  OAI211_X1 U9495 ( .C1(n5324), .C2(n10440), .A(n8090), .B(n8089), .ZN(n8091)
         );
  AOI21_X1 U9496 ( .B1(n10915), .B2(n10533), .A(n8091), .ZN(n8092) );
  OAI21_X1 U9497 ( .B1(n10537), .B2(n10452), .A(n8092), .ZN(P1_U3276) );
  NAND2_X1 U9498 ( .A1(n8094), .A2(n8093), .ZN(n8095) );
  AOI21_X1 U9499 ( .B1(n8096), .B2(n11078), .A(n8095), .ZN(n8099) );
  MUX2_X1 U9500 ( .A(n8097), .B(n8099), .S(n11081), .Z(n8098) );
  OAI21_X1 U9501 ( .B1(n8102), .B2(n10532), .A(n8098), .ZN(P1_U3538) );
  INV_X1 U9502 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n8100) );
  MUX2_X1 U9503 ( .A(n8100), .B(n8099), .S(n11085), .Z(n8101) );
  OAI21_X1 U9504 ( .B1(n8102), .B2(n10579), .A(n8101), .ZN(P1_U3501) );
  INV_X1 U9505 ( .A(n8103), .ZN(n8107) );
  OAI222_X1 U9506 ( .A1(n8618), .A2(n8105), .B1(n9719), .B2(n8107), .C1(n8104), 
        .C2(P2_U3151), .ZN(P2_U3269) );
  OAI222_X1 U9507 ( .A1(n8108), .A2(P1_U3086), .B1(n8657), .B2(n8107), .C1(
        n8106), .C2(n10595), .ZN(P1_U3329) );
  NAND2_X1 U9508 ( .A1(n8128), .A2(n8938), .ZN(n8110) );
  NAND2_X1 U9509 ( .A1(n8976), .A2(n10161), .ZN(n8109) );
  NAND2_X1 U9510 ( .A1(n8110), .A2(n8109), .ZN(n8163) );
  INV_X1 U9511 ( .A(n8111), .ZN(n8112) );
  NAND2_X1 U9512 ( .A1(n8113), .A2(n8112), .ZN(n8119) );
  NAND2_X1 U9513 ( .A1(n8122), .A2(n8119), .ZN(n8118) );
  NAND2_X1 U9514 ( .A1(n8128), .A2(n9000), .ZN(n8115) );
  NAND2_X1 U9515 ( .A1(n8961), .A2(n10161), .ZN(n8114) );
  NAND2_X1 U9516 ( .A1(n8115), .A2(n8114), .ZN(n8116) );
  XNOR2_X1 U9517 ( .A(n8116), .B(n8974), .ZN(n8120) );
  INV_X1 U9518 ( .A(n8120), .ZN(n8117) );
  NAND2_X1 U9519 ( .A1(n8118), .A2(n8117), .ZN(n8165) );
  AND2_X1 U9520 ( .A1(n8120), .A2(n8119), .ZN(n8121) );
  NAND2_X1 U9521 ( .A1(n8165), .A2(n8164), .ZN(n8123) );
  XOR2_X1 U9522 ( .A(n8163), .B(n8123), .Z(n8130) );
  NAND2_X1 U9523 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n10731) );
  OAI21_X1 U9524 ( .B1(n9874), .B2(n8124), .A(n10731), .ZN(n8127) );
  OAI22_X1 U9525 ( .A1(n8125), .A2(n9876), .B1(n9877), .B2(n9787), .ZN(n8126)
         );
  AOI211_X1 U9526 ( .C1(n8128), .C2(n9863), .A(n8127), .B(n8126), .ZN(n8129)
         );
  OAI21_X1 U9527 ( .B1(n8130), .B2(n9866), .A(n8129), .ZN(P1_U3215) );
  NAND2_X1 U9528 ( .A1(n8134), .A2(n5180), .ZN(n8132) );
  OAI211_X1 U9529 ( .C1(n8618), .C2(n8133), .A(n8132), .B(n8131), .ZN(P2_U3268) );
  INV_X1 U9530 ( .A(n8134), .ZN(n8135) );
  OAI222_X1 U9531 ( .A1(n10660), .A2(P1_U3086), .B1(n8657), .B2(n8135), .C1(
        n8290), .C2(n10595), .ZN(P1_U3328) );
  INV_X1 U9532 ( .A(n8136), .ZN(n8138) );
  OAI21_X1 U9533 ( .B1(n8139), .B2(n8138), .A(n8137), .ZN(n8140) );
  XNOR2_X1 U9534 ( .A(n8140), .B(n8144), .ZN(n8142) );
  OAI22_X1 U9535 ( .A1(n9860), .A2(n10900), .B1(n10448), .B2(n10902), .ZN(
        n8141) );
  AOI21_X1 U9536 ( .B1(n8142), .B2(n10402), .A(n8141), .ZN(n10526) );
  OAI21_X1 U9537 ( .B1(n8145), .B2(n8144), .A(n8143), .ZN(n10528) );
  NAND2_X1 U9538 ( .A1(n10528), .A2(n10458), .ZN(n8151) );
  INV_X1 U9539 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n10261) );
  INV_X1 U9540 ( .A(n8146), .ZN(n9859) );
  OAI22_X1 U9541 ( .A1(n10915), .A2(n10261), .B1(n9859), .B2(n11050), .ZN(
        n8149) );
  INV_X1 U9542 ( .A(n8147), .ZN(n8154) );
  OAI211_X1 U9543 ( .C1(n10580), .C2(n5166), .A(n8154), .B(n11035), .ZN(n10525) );
  NOR2_X1 U9544 ( .A1(n10525), .A2(n10335), .ZN(n8148) );
  AOI211_X1 U9545 ( .C1(n11056), .C2(n9864), .A(n8149), .B(n8148), .ZN(n8150)
         );
  OAI211_X1 U9546 ( .C1(n11051), .C2(n10526), .A(n8151), .B(n8150), .ZN(
        P1_U3275) );
  XNOR2_X1 U9547 ( .A(n8152), .B(n10093), .ZN(n10524) );
  INV_X1 U9548 ( .A(n10439), .ZN(n8153) );
  AOI211_X1 U9549 ( .C1(n10522), .C2(n8154), .A(n10438), .B(n8153), .ZN(n10521) );
  NOR2_X1 U9550 ( .A1(n8155), .A2(n10440), .ZN(n8158) );
  OAI22_X1 U9551 ( .A1(n10915), .A2(n8156), .B1(n9752), .B2(n11050), .ZN(n8157) );
  AOI211_X1 U9552 ( .C1(n10521), .C2(n11045), .A(n8158), .B(n8157), .ZN(n8162)
         );
  XOR2_X1 U9553 ( .A(n8159), .B(n10093), .Z(n8160) );
  OAI222_X1 U9554 ( .A1(n10902), .A2(n10426), .B1(n10900), .B2(n9799), .C1(
        n11030), .C2(n8160), .ZN(n10520) );
  NAND2_X1 U9555 ( .A1(n10520), .A2(n10915), .ZN(n8161) );
  OAI211_X1 U9556 ( .C1(n10524), .C2(n10452), .A(n8162), .B(n8161), .ZN(
        P1_U3274) );
  NAND2_X1 U9557 ( .A1(n8164), .A2(n8163), .ZN(n8166) );
  NAND2_X1 U9558 ( .A1(n10540), .A2(n9000), .ZN(n8168) );
  OR2_X1 U9559 ( .A1(n9787), .A2(n7115), .ZN(n8167) );
  NAND2_X1 U9560 ( .A1(n8168), .A2(n8167), .ZN(n8169) );
  XNOR2_X1 U9561 ( .A(n8169), .B(n9002), .ZN(n8171) );
  NAND2_X1 U9562 ( .A1(n5121), .A2(n8902), .ZN(n8174) );
  NOR2_X1 U9563 ( .A1(n9787), .A2(n9001), .ZN(n8173) );
  AOI21_X1 U9564 ( .B1(n10540), .B2(n8938), .A(n8173), .ZN(n8901) );
  XNOR2_X1 U9565 ( .A(n8174), .B(n8901), .ZN(n8180) );
  INV_X1 U9566 ( .A(n8175), .ZN(n8627) );
  NAND2_X1 U9567 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10742) );
  INV_X1 U9568 ( .A(n10742), .ZN(n8177) );
  OAI22_X1 U9569 ( .A1(n8622), .A2(n9876), .B1(n9877), .B2(n9798), .ZN(n8176)
         );
  AOI211_X1 U9570 ( .C1(n9803), .C2(n8627), .A(n8177), .B(n8176), .ZN(n8179)
         );
  NAND2_X1 U9571 ( .A1(n10540), .A2(n9863), .ZN(n8178) );
  OAI211_X1 U9572 ( .C1(n8180), .C2(n9866), .A(n8179), .B(n8178), .ZN(P1_U3241) );
  INV_X1 U9573 ( .A(n8609), .ZN(n8182) );
  OAI222_X1 U9574 ( .A1(P1_U3086), .A2(n6210), .B1(n8657), .B2(n8182), .C1(
        n8181), .C2(n10595), .ZN(P1_U3327) );
  XNOR2_X1 U9575 ( .A(SI_31_), .B(keyinput_129), .ZN(n8185) );
  XNOR2_X1 U9576 ( .A(SI_30_), .B(keyinput_130), .ZN(n8184) );
  XNOR2_X1 U9577 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_128), .ZN(n8183) );
  NOR3_X1 U9578 ( .A1(n8185), .A2(n8184), .A3(n8183), .ZN(n8188) );
  XNOR2_X1 U9579 ( .A(SI_28_), .B(keyinput_132), .ZN(n8187) );
  XNOR2_X1 U9580 ( .A(SI_29_), .B(keyinput_131), .ZN(n8186) );
  NOR3_X1 U9581 ( .A1(n8188), .A2(n8187), .A3(n8186), .ZN(n8196) );
  XNOR2_X1 U9582 ( .A(n8388), .B(keyinput_136), .ZN(n8192) );
  XNOR2_X1 U9583 ( .A(SI_26_), .B(keyinput_134), .ZN(n8191) );
  XNOR2_X1 U9584 ( .A(SI_27_), .B(keyinput_133), .ZN(n8190) );
  XNOR2_X1 U9585 ( .A(SI_25_), .B(keyinput_135), .ZN(n8189) );
  NAND4_X1 U9586 ( .A1(n8192), .A2(n8191), .A3(n8190), .A4(n8189), .ZN(n8195)
         );
  XNOR2_X1 U9587 ( .A(n8401), .B(keyinput_137), .ZN(n8194) );
  XNOR2_X1 U9588 ( .A(n8400), .B(keyinput_138), .ZN(n8193) );
  OAI211_X1 U9589 ( .C1(n8196), .C2(n8195), .A(n8194), .B(n8193), .ZN(n8205)
         );
  XNOR2_X1 U9590 ( .A(n8197), .B(keyinput_139), .ZN(n8204) );
  XNOR2_X1 U9591 ( .A(n8407), .B(keyinput_141), .ZN(n8201) );
  XNOR2_X1 U9592 ( .A(n8198), .B(keyinput_143), .ZN(n8200) );
  XNOR2_X1 U9593 ( .A(SI_20_), .B(keyinput_140), .ZN(n8199) );
  NOR3_X1 U9594 ( .A1(n8201), .A2(n8200), .A3(n8199), .ZN(n8203) );
  XNOR2_X1 U9595 ( .A(SI_18_), .B(keyinput_142), .ZN(n8202) );
  NAND4_X1 U9596 ( .A1(n8205), .A2(n8204), .A3(n8203), .A4(n8202), .ZN(n8211)
         );
  XNOR2_X1 U9597 ( .A(n8206), .B(keyinput_144), .ZN(n8210) );
  XNOR2_X1 U9598 ( .A(n8418), .B(keyinput_145), .ZN(n8209) );
  XOR2_X1 U9599 ( .A(SI_13_), .B(keyinput_147), .Z(n8208) );
  XNOR2_X1 U9600 ( .A(SI_12_), .B(keyinput_148), .ZN(n8207) );
  NAND2_X1 U9601 ( .A1(n8208), .A2(n8207), .ZN(n8214) );
  AOI211_X1 U9602 ( .C1(n8211), .C2(n8210), .A(n8209), .B(n8214), .ZN(n8217)
         );
  XNOR2_X1 U9603 ( .A(n8422), .B(keyinput_146), .ZN(n8213) );
  XNOR2_X1 U9604 ( .A(SI_11_), .B(keyinput_149), .ZN(n8212) );
  OAI21_X1 U9605 ( .B1(n8214), .B2(n8213), .A(n8212), .ZN(n8216) );
  XNOR2_X1 U9606 ( .A(SI_10_), .B(keyinput_150), .ZN(n8215) );
  OAI21_X1 U9607 ( .B1(n8217), .B2(n8216), .A(n8215), .ZN(n8233) );
  XOR2_X1 U9608 ( .A(SI_7_), .B(keyinput_153), .Z(n8228) );
  XNOR2_X1 U9609 ( .A(n8218), .B(keyinput_157), .ZN(n8223) );
  XNOR2_X1 U9610 ( .A(n8219), .B(keyinput_151), .ZN(n8222) );
  XNOR2_X1 U9611 ( .A(SI_4_), .B(keyinput_156), .ZN(n8221) );
  XNOR2_X1 U9612 ( .A(SI_5_), .B(keyinput_155), .ZN(n8220) );
  NAND4_X1 U9613 ( .A1(n8223), .A2(n8222), .A3(n8221), .A4(n8220), .ZN(n8227)
         );
  XNOR2_X1 U9614 ( .A(n8224), .B(keyinput_152), .ZN(n8226) );
  XNOR2_X1 U9615 ( .A(SI_6_), .B(keyinput_154), .ZN(n8225) );
  NOR4_X1 U9616 ( .A1(n8228), .A2(n8227), .A3(n8226), .A4(n8225), .ZN(n8232)
         );
  XNOR2_X1 U9617 ( .A(n8229), .B(keyinput_158), .ZN(n8231) );
  XNOR2_X1 U9618 ( .A(n8441), .B(keyinput_159), .ZN(n8230) );
  AOI211_X1 U9619 ( .C1(n8233), .C2(n8232), .A(n8231), .B(n8230), .ZN(n8239)
         );
  XNOR2_X1 U9620 ( .A(SI_0_), .B(keyinput_160), .ZN(n8238) );
  XNOR2_X1 U9621 ( .A(P2_U3151), .B(keyinput_162), .ZN(n8236) );
  XNOR2_X1 U9622 ( .A(n8447), .B(keyinput_163), .ZN(n8235) );
  XNOR2_X1 U9623 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_161), .ZN(n8234) );
  NOR3_X1 U9624 ( .A1(n8236), .A2(n8235), .A3(n8234), .ZN(n8237) );
  OAI21_X1 U9625 ( .B1(n8239), .B2(n8238), .A(n8237), .ZN(n8243) );
  XOR2_X1 U9626 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput_165), .Z(n8242) );
  XNOR2_X1 U9627 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput_166), .ZN(n8241)
         );
  XNOR2_X1 U9628 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_164), .ZN(n8240)
         );
  NAND4_X1 U9629 ( .A1(n8243), .A2(n8242), .A3(n8241), .A4(n8240), .ZN(n8246)
         );
  XOR2_X1 U9630 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_167), .Z(n8245) );
  XNOR2_X1 U9631 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_168), .ZN(n8244) );
  AOI21_X1 U9632 ( .B1(n8246), .B2(n8245), .A(n8244), .ZN(n8251) );
  XNOR2_X1 U9633 ( .A(n8247), .B(keyinput_169), .ZN(n8250) );
  XOR2_X1 U9634 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput_171), .Z(n8249) );
  XNOR2_X1 U9635 ( .A(P2_REG3_REG_28__SCAN_IN), .B(keyinput_170), .ZN(n8248)
         );
  OAI211_X1 U9636 ( .C1(n8251), .C2(n8250), .A(n8249), .B(n8248), .ZN(n8254)
         );
  XNOR2_X1 U9637 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_172), .ZN(n8253) );
  XNOR2_X1 U9638 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput_173), .ZN(n8252)
         );
  AOI21_X1 U9639 ( .B1(n8254), .B2(n8253), .A(n8252), .ZN(n8258) );
  XNOR2_X1 U9640 ( .A(n8255), .B(keyinput_174), .ZN(n8257) );
  XNOR2_X1 U9641 ( .A(P2_REG3_REG_25__SCAN_IN), .B(keyinput_175), .ZN(n8256)
         );
  NOR3_X1 U9642 ( .A1(n8258), .A2(n8257), .A3(n8256), .ZN(n8262) );
  XOR2_X1 U9643 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_176), .Z(n8261) );
  XNOR2_X1 U9644 ( .A(n8259), .B(keyinput_177), .ZN(n8260) );
  NOR3_X1 U9645 ( .A1(n8262), .A2(n8261), .A3(n8260), .ZN(n8266) );
  XNOR2_X1 U9646 ( .A(n8476), .B(keyinput_178), .ZN(n8265) );
  XNOR2_X1 U9647 ( .A(n8263), .B(keyinput_179), .ZN(n8264) );
  NOR3_X1 U9648 ( .A1(n8266), .A2(n8265), .A3(n8264), .ZN(n8269) );
  XNOR2_X1 U9649 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_180), .ZN(n8268) );
  XNOR2_X1 U9650 ( .A(n8480), .B(keyinput_181), .ZN(n8267) );
  OAI21_X1 U9651 ( .B1(n8269), .B2(n8268), .A(n8267), .ZN(n8272) );
  XOR2_X1 U9652 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_182), .Z(n8271) );
  XNOR2_X1 U9653 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput_183), .ZN(n8270)
         );
  AOI21_X1 U9654 ( .B1(n8272), .B2(n8271), .A(n8270), .ZN(n8275) );
  XNOR2_X1 U9655 ( .A(P2_REG3_REG_13__SCAN_IN), .B(keyinput_184), .ZN(n8274)
         );
  XNOR2_X1 U9656 ( .A(P2_REG3_REG_22__SCAN_IN), .B(keyinput_185), .ZN(n8273)
         );
  NOR3_X1 U9657 ( .A1(n8275), .A2(n8274), .A3(n8273), .ZN(n8278) );
  XOR2_X1 U9658 ( .A(P2_REG3_REG_11__SCAN_IN), .B(keyinput_186), .Z(n8277) );
  XNOR2_X1 U9659 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_187), .ZN(n8276) );
  OAI21_X1 U9660 ( .B1(n8278), .B2(n8277), .A(n8276), .ZN(n8282) );
  XNOR2_X1 U9661 ( .A(P2_REG3_REG_26__SCAN_IN), .B(keyinput_190), .ZN(n8281)
         );
  XNOR2_X1 U9662 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput_189), .ZN(n8280) );
  XNOR2_X1 U9663 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput_188), .ZN(n8279)
         );
  NAND4_X1 U9664 ( .A1(n8282), .A2(n8281), .A3(n8280), .A4(n8279), .ZN(n8285)
         );
  XNOR2_X1 U9665 ( .A(P2_B_REG_SCAN_IN), .B(keyinput_192), .ZN(n8284) );
  XNOR2_X1 U9666 ( .A(P2_REG3_REG_15__SCAN_IN), .B(keyinput_191), .ZN(n8283)
         );
  NAND3_X1 U9667 ( .A1(n8285), .A2(n8284), .A3(n8283), .ZN(n8289) );
  INV_X1 U9668 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9894) );
  XNOR2_X1 U9669 ( .A(n9894), .B(keyinput_194), .ZN(n8288) );
  XNOR2_X1 U9670 ( .A(n10596), .B(keyinput_195), .ZN(n8287) );
  XNOR2_X1 U9671 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(keyinput_193), .ZN(n8286)
         );
  NAND4_X1 U9672 ( .A1(n8289), .A2(n8288), .A3(n8287), .A4(n8286), .ZN(n8300)
         );
  XOR2_X1 U9673 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput_196), .Z(n8299) );
  XNOR2_X1 U9674 ( .A(n8508), .B(keyinput_200), .ZN(n8293) );
  XNOR2_X1 U9675 ( .A(n8290), .B(keyinput_197), .ZN(n8292) );
  XNOR2_X1 U9676 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(keyinput_198), .ZN(n8291)
         );
  NOR3_X1 U9677 ( .A1(n8293), .A2(n8292), .A3(n8291), .ZN(n8297) );
  XNOR2_X1 U9678 ( .A(n8294), .B(keyinput_201), .ZN(n8296) );
  XNOR2_X1 U9679 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput_199), .ZN(n8295)
         );
  NAND3_X1 U9680 ( .A1(n8297), .A2(n8296), .A3(n8295), .ZN(n8298) );
  AOI21_X1 U9681 ( .B1(n8300), .B2(n8299), .A(n8298), .ZN(n8303) );
  XOR2_X1 U9682 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_203), .Z(n8302) );
  XNOR2_X1 U9683 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_202), .ZN(n8301)
         );
  NOR3_X1 U9684 ( .A1(n8303), .A2(n8302), .A3(n8301), .ZN(n8308) );
  XNOR2_X1 U9685 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(keyinput_204), .ZN(n8307)
         );
  XNOR2_X1 U9686 ( .A(n8304), .B(keyinput_205), .ZN(n8306) );
  XOR2_X1 U9687 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_206), .Z(n8305) );
  OAI211_X1 U9688 ( .C1(n8308), .C2(n8307), .A(n8306), .B(n8305), .ZN(n8312)
         );
  XNOR2_X1 U9689 ( .A(n8309), .B(keyinput_207), .ZN(n8311) );
  XNOR2_X1 U9690 ( .A(n8525), .B(keyinput_208), .ZN(n8310) );
  NAND3_X1 U9691 ( .A1(n8312), .A2(n8311), .A3(n8310), .ZN(n8315) );
  XNOR2_X1 U9692 ( .A(n8529), .B(keyinput_210), .ZN(n8314) );
  XNOR2_X1 U9693 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput_209), .ZN(n8313)
         );
  NAND3_X1 U9694 ( .A1(n8315), .A2(n8314), .A3(n8313), .ZN(n8318) );
  XNOR2_X1 U9695 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput_211), .ZN(n8317)
         );
  XOR2_X1 U9696 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput_212), .Z(n8316) );
  AOI21_X1 U9697 ( .B1(n8318), .B2(n8317), .A(n8316), .ZN(n8321) );
  XNOR2_X1 U9698 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput_213), .ZN(n8320)
         );
  XNOR2_X1 U9699 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput_214), .ZN(n8319)
         );
  NOR3_X1 U9700 ( .A1(n8321), .A2(n8320), .A3(n8319), .ZN(n8325) );
  XNOR2_X1 U9701 ( .A(n8539), .B(keyinput_215), .ZN(n8324) );
  XNOR2_X1 U9702 ( .A(n8322), .B(keyinput_216), .ZN(n8323) );
  NOR3_X1 U9703 ( .A1(n8325), .A2(n8324), .A3(n8323), .ZN(n8331) );
  XOR2_X1 U9704 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_217), .Z(n8330) );
  XOR2_X1 U9705 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_218), .Z(n8328) );
  XNOR2_X1 U9706 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_220), .ZN(n8327) );
  XNOR2_X1 U9707 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_219), .ZN(n8326) );
  NOR3_X1 U9708 ( .A1(n8328), .A2(n8327), .A3(n8326), .ZN(n8329) );
  OAI21_X1 U9709 ( .B1(n8331), .B2(n8330), .A(n8329), .ZN(n8335) );
  XNOR2_X1 U9710 ( .A(n8332), .B(keyinput_221), .ZN(n8334) );
  XNOR2_X1 U9711 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_222), .ZN(n8333) );
  AOI21_X1 U9712 ( .B1(n8335), .B2(n8334), .A(n8333), .ZN(n8341) );
  XOR2_X1 U9713 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_223), .Z(n8340) );
  XOR2_X1 U9714 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_225), .Z(n8338) );
  XNOR2_X1 U9715 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_226), .ZN(n8337) );
  XNOR2_X1 U9716 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_224), .ZN(n8336) );
  NOR3_X1 U9717 ( .A1(n8338), .A2(n8337), .A3(n8336), .ZN(n8339) );
  OAI21_X1 U9718 ( .B1(n8341), .B2(n8340), .A(n8339), .ZN(n8346) );
  XNOR2_X1 U9719 ( .A(n8558), .B(keyinput_228), .ZN(n8345) );
  XNOR2_X1 U9720 ( .A(n8559), .B(keyinput_229), .ZN(n8344) );
  XNOR2_X1 U9721 ( .A(n8342), .B(keyinput_227), .ZN(n8343) );
  NAND4_X1 U9722 ( .A1(n8346), .A2(n8345), .A3(n8344), .A4(n8343), .ZN(n8349)
         );
  XOR2_X1 U9723 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_230), .Z(n8348) );
  XNOR2_X1 U9724 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_231), .ZN(n8347) );
  AOI21_X1 U9725 ( .B1(n8349), .B2(n8348), .A(n8347), .ZN(n8355) );
  XOR2_X1 U9726 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_232), .Z(n8354) );
  XNOR2_X1 U9727 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_233), .ZN(n8352) );
  XNOR2_X1 U9728 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_235), .ZN(n8351) );
  XNOR2_X1 U9729 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_234), .ZN(n8350) );
  NOR3_X1 U9730 ( .A1(n8352), .A2(n8351), .A3(n8350), .ZN(n8353) );
  OAI21_X1 U9731 ( .B1(n8355), .B2(n8354), .A(n8353), .ZN(n8358) );
  XNOR2_X1 U9732 ( .A(n8573), .B(keyinput_236), .ZN(n8357) );
  XNOR2_X1 U9733 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_237), .ZN(n8356) );
  AOI21_X1 U9734 ( .B1(n8358), .B2(n8357), .A(n8356), .ZN(n8362) );
  XNOR2_X1 U9735 ( .A(n8577), .B(keyinput_238), .ZN(n8361) );
  XNOR2_X1 U9736 ( .A(n8359), .B(keyinput_239), .ZN(n8360) );
  OAI21_X1 U9737 ( .B1(n8362), .B2(n8361), .A(n8360), .ZN(n8368) );
  XNOR2_X1 U9738 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_240), .ZN(n8367) );
  XNOR2_X1 U9739 ( .A(n8582), .B(keyinput_242), .ZN(n8365) );
  XNOR2_X1 U9740 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_243), .ZN(n8364) );
  XNOR2_X1 U9741 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput_241), .ZN(n8363) );
  NAND3_X1 U9742 ( .A1(n8365), .A2(n8364), .A3(n8363), .ZN(n8366) );
  AOI21_X1 U9743 ( .B1(n8368), .B2(n8367), .A(n8366), .ZN(n8375) );
  XOR2_X1 U9744 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_244), .Z(n8374) );
  XNOR2_X1 U9745 ( .A(n8369), .B(keyinput_247), .ZN(n8372) );
  XNOR2_X1 U9746 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_246), .ZN(n8371) );
  XNOR2_X1 U9747 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_245), .ZN(n8370) );
  NOR3_X1 U9748 ( .A1(n8372), .A2(n8371), .A3(n8370), .ZN(n8373) );
  OAI21_X1 U9749 ( .B1(n8375), .B2(n8374), .A(n8373), .ZN(n8378) );
  XNOR2_X1 U9750 ( .A(n10588), .B(keyinput_248), .ZN(n8377) );
  XOR2_X1 U9751 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_249), .Z(n8376) );
  AOI21_X1 U9752 ( .B1(n8378), .B2(n8377), .A(n8376), .ZN(n8385) );
  XNOR2_X1 U9753 ( .A(P1_D_REG_2__SCAN_IN), .B(keyinput_252), .ZN(n8384) );
  XNOR2_X1 U9754 ( .A(P1_D_REG_1__SCAN_IN), .B(keyinput_251), .ZN(n8383) );
  XOR2_X1 U9755 ( .A(P1_D_REG_0__SCAN_IN), .B(keyinput_250), .Z(n8381) );
  XOR2_X1 U9756 ( .A(P1_D_REG_3__SCAN_IN), .B(keyinput_253), .Z(n8380) );
  XNOR2_X1 U9757 ( .A(keyinput_254), .B(P1_D_REG_4__SCAN_IN), .ZN(n8379) );
  NAND3_X1 U9758 ( .A1(n8381), .A2(n8380), .A3(n8379), .ZN(n8382) );
  NOR4_X1 U9759 ( .A1(n8385), .A2(n8384), .A3(n8383), .A4(n8382), .ZN(n8608)
         );
  XOR2_X1 U9760 ( .A(keyinput_127), .B(keyinput_255), .Z(n8607) );
  XNOR2_X1 U9761 ( .A(n8386), .B(keyinput_6), .ZN(n8392) );
  XNOR2_X1 U9762 ( .A(n8387), .B(keyinput_5), .ZN(n8391) );
  XNOR2_X1 U9763 ( .A(n8388), .B(keyinput_8), .ZN(n8390) );
  XNOR2_X1 U9764 ( .A(SI_25_), .B(keyinput_7), .ZN(n8389) );
  NOR4_X1 U9765 ( .A1(n8392), .A2(n8391), .A3(n8390), .A4(n8389), .ZN(n8405)
         );
  XOR2_X1 U9766 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_0), .Z(n8395) );
  INV_X1 U9767 ( .A(SI_31_), .ZN(n8663) );
  XNOR2_X1 U9768 ( .A(n8663), .B(keyinput_1), .ZN(n8394) );
  XNOR2_X1 U9769 ( .A(SI_30_), .B(keyinput_2), .ZN(n8393) );
  NAND3_X1 U9770 ( .A1(n8395), .A2(n8394), .A3(n8393), .ZN(n8399) );
  XNOR2_X1 U9771 ( .A(n8396), .B(keyinput_4), .ZN(n8398) );
  XNOR2_X1 U9772 ( .A(SI_29_), .B(keyinput_3), .ZN(n8397) );
  NAND3_X1 U9773 ( .A1(n8399), .A2(n8398), .A3(n8397), .ZN(n8404) );
  XNOR2_X1 U9774 ( .A(n8400), .B(keyinput_10), .ZN(n8403) );
  XNOR2_X1 U9775 ( .A(n8401), .B(keyinput_9), .ZN(n8402) );
  AOI211_X1 U9776 ( .C1(n8405), .C2(n8404), .A(n8403), .B(n8402), .ZN(n8414)
         );
  XNOR2_X1 U9777 ( .A(SI_18_), .B(keyinput_14), .ZN(n8413) );
  XNOR2_X1 U9778 ( .A(SI_21_), .B(keyinput_11), .ZN(n8412) );
  XNOR2_X1 U9779 ( .A(n8406), .B(keyinput_12), .ZN(n8410) );
  XNOR2_X1 U9780 ( .A(n8407), .B(keyinput_13), .ZN(n8409) );
  XNOR2_X1 U9781 ( .A(SI_17_), .B(keyinput_15), .ZN(n8408) );
  NAND3_X1 U9782 ( .A1(n8410), .A2(n8409), .A3(n8408), .ZN(n8411) );
  NOR4_X1 U9783 ( .A1(n8414), .A2(n8413), .A3(n8412), .A4(n8411), .ZN(n8421)
         );
  XNOR2_X1 U9784 ( .A(SI_16_), .B(keyinput_16), .ZN(n8420) );
  XOR2_X1 U9785 ( .A(SI_13_), .B(keyinput_19), .Z(n8417) );
  XNOR2_X1 U9786 ( .A(n8415), .B(keyinput_20), .ZN(n8416) );
  NOR2_X1 U9787 ( .A1(n8417), .A2(n8416), .ZN(n8426) );
  XNOR2_X1 U9788 ( .A(n8418), .B(keyinput_17), .ZN(n8419) );
  OAI211_X1 U9789 ( .C1(n8421), .C2(n8420), .A(n8426), .B(n8419), .ZN(n8430)
         );
  XNOR2_X1 U9790 ( .A(n8422), .B(keyinput_18), .ZN(n8425) );
  XNOR2_X1 U9791 ( .A(n8423), .B(keyinput_21), .ZN(n8424) );
  AOI21_X1 U9792 ( .B1(n8426), .B2(n8425), .A(n8424), .ZN(n8429) );
  XNOR2_X1 U9793 ( .A(n8427), .B(keyinput_22), .ZN(n8428) );
  AOI21_X1 U9794 ( .B1(n8430), .B2(n8429), .A(n8428), .ZN(n8445) );
  XNOR2_X1 U9795 ( .A(n8431), .B(keyinput_27), .ZN(n8435) );
  XNOR2_X1 U9796 ( .A(SI_4_), .B(keyinput_28), .ZN(n8434) );
  XNOR2_X1 U9797 ( .A(SI_3_), .B(keyinput_29), .ZN(n8433) );
  XNOR2_X1 U9798 ( .A(SI_7_), .B(keyinput_25), .ZN(n8432) );
  NOR4_X1 U9799 ( .A1(n8435), .A2(n8434), .A3(n8433), .A4(n8432), .ZN(n8440)
         );
  XNOR2_X1 U9800 ( .A(n8436), .B(keyinput_26), .ZN(n8439) );
  XNOR2_X1 U9801 ( .A(SI_9_), .B(keyinput_23), .ZN(n8438) );
  XNOR2_X1 U9802 ( .A(SI_8_), .B(keyinput_24), .ZN(n8437) );
  NAND4_X1 U9803 ( .A1(n8440), .A2(n8439), .A3(n8438), .A4(n8437), .ZN(n8444)
         );
  XNOR2_X1 U9804 ( .A(n8441), .B(keyinput_31), .ZN(n8443) );
  XNOR2_X1 U9805 ( .A(SI_2_), .B(keyinput_30), .ZN(n8442) );
  OAI211_X1 U9806 ( .C1(n8445), .C2(n8444), .A(n8443), .B(n8442), .ZN(n8453)
         );
  XOR2_X1 U9807 ( .A(SI_0_), .B(keyinput_32), .Z(n8452) );
  XNOR2_X1 U9808 ( .A(P2_U3151), .B(keyinput_34), .ZN(n8450) );
  XNOR2_X1 U9809 ( .A(n8447), .B(keyinput_35), .ZN(n8449) );
  XNOR2_X1 U9810 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_33), .ZN(n8448) );
  NAND3_X1 U9811 ( .A1(n8450), .A2(n8449), .A3(n8448), .ZN(n8451) );
  AOI21_X1 U9812 ( .B1(n8453), .B2(n8452), .A(n8451), .ZN(n8458) );
  XOR2_X1 U9813 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput_38), .Z(n8457) );
  XNOR2_X1 U9814 ( .A(n8454), .B(keyinput_36), .ZN(n8456) );
  XNOR2_X1 U9815 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput_37), .ZN(n8455) );
  NOR4_X1 U9816 ( .A1(n8458), .A2(n8457), .A3(n8456), .A4(n8455), .ZN(n8461)
         );
  XOR2_X1 U9817 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_39), .Z(n8460) );
  XNOR2_X1 U9818 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_40), .ZN(n8459) );
  OAI21_X1 U9819 ( .B1(n8461), .B2(n8460), .A(n8459), .ZN(n8465) );
  XNOR2_X1 U9820 ( .A(P2_REG3_REG_19__SCAN_IN), .B(keyinput_41), .ZN(n8464) );
  XNOR2_X1 U9821 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput_43), .ZN(n8463) );
  XNOR2_X1 U9822 ( .A(P2_REG3_REG_28__SCAN_IN), .B(keyinput_42), .ZN(n8462) );
  AOI211_X1 U9823 ( .C1(n8465), .C2(n8464), .A(n8463), .B(n8462), .ZN(n8468)
         );
  XOR2_X1 U9824 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_44), .Z(n8467) );
  XNOR2_X1 U9825 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput_45), .ZN(n8466) );
  OAI21_X1 U9826 ( .B1(n8468), .B2(n8467), .A(n8466), .ZN(n8472) );
  XNOR2_X1 U9827 ( .A(n8469), .B(keyinput_47), .ZN(n8471) );
  XNOR2_X1 U9828 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput_46), .ZN(n8470) );
  NAND3_X1 U9829 ( .A1(n8472), .A2(n8471), .A3(n8470), .ZN(n8475) );
  XNOR2_X1 U9830 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_48), .ZN(n8474) );
  XNOR2_X1 U9831 ( .A(P2_REG3_REG_5__SCAN_IN), .B(keyinput_49), .ZN(n8473) );
  NAND3_X1 U9832 ( .A1(n8475), .A2(n8474), .A3(n8473), .ZN(n8479) );
  XNOR2_X1 U9833 ( .A(n8476), .B(keyinput_50), .ZN(n8478) );
  XNOR2_X1 U9834 ( .A(P2_REG3_REG_24__SCAN_IN), .B(keyinput_51), .ZN(n8477) );
  NAND3_X1 U9835 ( .A1(n8479), .A2(n8478), .A3(n8477), .ZN(n8483) );
  XNOR2_X1 U9836 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_52), .ZN(n8482) );
  XNOR2_X1 U9837 ( .A(n8480), .B(keyinput_53), .ZN(n8481) );
  AOI21_X1 U9838 ( .B1(n8483), .B2(n8482), .A(n8481), .ZN(n8487) );
  XNOR2_X1 U9839 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_54), .ZN(n8486) );
  XNOR2_X1 U9840 ( .A(n8484), .B(keyinput_55), .ZN(n8485) );
  OAI21_X1 U9841 ( .B1(n8487), .B2(n8486), .A(n8485), .ZN(n8491) );
  XNOR2_X1 U9842 ( .A(n8488), .B(keyinput_56), .ZN(n8490) );
  XOR2_X1 U9843 ( .A(P2_REG3_REG_22__SCAN_IN), .B(keyinput_57), .Z(n8489) );
  NAND3_X1 U9844 ( .A1(n8491), .A2(n8490), .A3(n8489), .ZN(n8494) );
  XNOR2_X1 U9845 ( .A(P2_REG3_REG_11__SCAN_IN), .B(keyinput_58), .ZN(n8493) );
  XNOR2_X1 U9846 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_59), .ZN(n8492) );
  AOI21_X1 U9847 ( .B1(n8494), .B2(n8493), .A(n8492), .ZN(n8499) );
  XNOR2_X1 U9848 ( .A(n8495), .B(keyinput_61), .ZN(n8498) );
  XNOR2_X1 U9849 ( .A(P2_REG3_REG_26__SCAN_IN), .B(keyinput_62), .ZN(n8497) );
  XNOR2_X1 U9850 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput_60), .ZN(n8496) );
  NOR4_X1 U9851 ( .A1(n8499), .A2(n8498), .A3(n8497), .A4(n8496), .ZN(n8503)
         );
  XNOR2_X1 U9852 ( .A(n8500), .B(keyinput_63), .ZN(n8502) );
  XNOR2_X1 U9853 ( .A(P2_B_REG_SCAN_IN), .B(keyinput_64), .ZN(n8501) );
  NOR3_X1 U9854 ( .A1(n8503), .A2(n8502), .A3(n8501), .ZN(n8507) );
  XNOR2_X1 U9855 ( .A(n9894), .B(keyinput_66), .ZN(n8506) );
  XOR2_X1 U9856 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(keyinput_65), .Z(n8505) );
  XNOR2_X1 U9857 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(keyinput_67), .ZN(n8504)
         );
  NOR4_X1 U9858 ( .A1(n8507), .A2(n8506), .A3(n8505), .A4(n8504), .ZN(n8517)
         );
  XNOR2_X1 U9859 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput_68), .ZN(n8516)
         );
  XNOR2_X1 U9860 ( .A(n8508), .B(keyinput_72), .ZN(n8511) );
  XNOR2_X1 U9861 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(keyinput_73), .ZN(n8510)
         );
  XNOR2_X1 U9862 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(keyinput_70), .ZN(n8509)
         );
  NAND3_X1 U9863 ( .A1(n8511), .A2(n8510), .A3(n8509), .ZN(n8514) );
  XNOR2_X1 U9864 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput_71), .ZN(n8513)
         );
  XNOR2_X1 U9865 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(keyinput_69), .ZN(n8512)
         );
  NOR3_X1 U9866 ( .A1(n8514), .A2(n8513), .A3(n8512), .ZN(n8515) );
  OAI21_X1 U9867 ( .B1(n8517), .B2(n8516), .A(n8515), .ZN(n8520) );
  XOR2_X1 U9868 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_75), .Z(n8519) );
  XNOR2_X1 U9869 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_74), .ZN(n8518)
         );
  NAND3_X1 U9870 ( .A1(n8520), .A2(n8519), .A3(n8518), .ZN(n8524) );
  XNOR2_X1 U9871 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(keyinput_76), .ZN(n8523)
         );
  XOR2_X1 U9872 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_78), .Z(n8522) );
  XNOR2_X1 U9873 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput_77), .ZN(n8521)
         );
  AOI211_X1 U9874 ( .C1(n8524), .C2(n8523), .A(n8522), .B(n8521), .ZN(n8528)
         );
  XNOR2_X1 U9875 ( .A(n8525), .B(keyinput_80), .ZN(n8527) );
  XNOR2_X1 U9876 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput_79), .ZN(n8526)
         );
  NOR3_X1 U9877 ( .A1(n8528), .A2(n8527), .A3(n8526), .ZN(n8532) );
  XNOR2_X1 U9878 ( .A(n8529), .B(keyinput_82), .ZN(n8531) );
  XNOR2_X1 U9879 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput_81), .ZN(n8530)
         );
  NOR3_X1 U9880 ( .A1(n8532), .A2(n8531), .A3(n8530), .ZN(n8535) );
  XOR2_X1 U9881 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput_83), .Z(n8534) );
  XOR2_X1 U9882 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput_84), .Z(n8533) );
  OAI21_X1 U9883 ( .B1(n8535), .B2(n8534), .A(n8533), .ZN(n8538) );
  XNOR2_X1 U9884 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput_85), .ZN(n8537)
         );
  XNOR2_X1 U9885 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput_86), .ZN(n8536)
         );
  NAND3_X1 U9886 ( .A1(n8538), .A2(n8537), .A3(n8536), .ZN(n8542) );
  XNOR2_X1 U9887 ( .A(n8539), .B(keyinput_87), .ZN(n8541) );
  XNOR2_X1 U9888 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput_88), .ZN(n8540) );
  NAND3_X1 U9889 ( .A1(n8542), .A2(n8541), .A3(n8540), .ZN(n8548) );
  XNOR2_X1 U9890 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_89), .ZN(n8547) );
  XOR2_X1 U9891 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_90), .Z(n8545) );
  XNOR2_X1 U9892 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_91), .ZN(n8544) );
  XNOR2_X1 U9893 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_92), .ZN(n8543) );
  NAND3_X1 U9894 ( .A1(n8545), .A2(n8544), .A3(n8543), .ZN(n8546) );
  AOI21_X1 U9895 ( .B1(n8548), .B2(n8547), .A(n8546), .ZN(n8551) );
  XNOR2_X1 U9896 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_93), .ZN(n8550) );
  XNOR2_X1 U9897 ( .A(n5679), .B(keyinput_94), .ZN(n8549) );
  OAI21_X1 U9898 ( .B1(n8551), .B2(n8550), .A(n8549), .ZN(n8557) );
  XNOR2_X1 U9899 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_95), .ZN(n8556) );
  XOR2_X1 U9900 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_98), .Z(n8554) );
  XNOR2_X1 U9901 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_97), .ZN(n8553) );
  XNOR2_X1 U9902 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_96), .ZN(n8552) );
  NAND3_X1 U9903 ( .A1(n8554), .A2(n8553), .A3(n8552), .ZN(n8555) );
  AOI21_X1 U9904 ( .B1(n8557), .B2(n8556), .A(n8555), .ZN(n8563) );
  XNOR2_X1 U9905 ( .A(n8558), .B(keyinput_100), .ZN(n8562) );
  XNOR2_X1 U9906 ( .A(n8559), .B(keyinput_101), .ZN(n8561) );
  XNOR2_X1 U9907 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_99), .ZN(n8560) );
  NOR4_X1 U9908 ( .A1(n8563), .A2(n8562), .A3(n8561), .A4(n8560), .ZN(n8566)
         );
  XOR2_X1 U9909 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_102), .Z(n8565) );
  XNOR2_X1 U9910 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_103), .ZN(n8564) );
  OAI21_X1 U9911 ( .B1(n8566), .B2(n8565), .A(n8564), .ZN(n8572) );
  XNOR2_X1 U9912 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_104), .ZN(n8571) );
  XNOR2_X1 U9913 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_106), .ZN(n8569) );
  XNOR2_X1 U9914 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_105), .ZN(n8568) );
  XNOR2_X1 U9915 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_107), .ZN(n8567) );
  NAND3_X1 U9916 ( .A1(n8569), .A2(n8568), .A3(n8567), .ZN(n8570) );
  AOI21_X1 U9917 ( .B1(n8572), .B2(n8571), .A(n8570), .ZN(n8576) );
  XNOR2_X1 U9918 ( .A(n8573), .B(keyinput_108), .ZN(n8575) );
  XNOR2_X1 U9919 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_109), .ZN(n8574) );
  OAI21_X1 U9920 ( .B1(n8576), .B2(n8575), .A(n8574), .ZN(n8580) );
  XNOR2_X1 U9921 ( .A(n8577), .B(keyinput_110), .ZN(n8579) );
  XNOR2_X1 U9922 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput_111), .ZN(n8578) );
  AOI21_X1 U9923 ( .B1(n8580), .B2(n8579), .A(n8578), .ZN(n8588) );
  XNOR2_X1 U9924 ( .A(n8581), .B(keyinput_112), .ZN(n8587) );
  XNOR2_X1 U9925 ( .A(n8582), .B(keyinput_114), .ZN(n8585) );
  XNOR2_X1 U9926 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_115), .ZN(n8584) );
  XNOR2_X1 U9927 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput_113), .ZN(n8583) );
  NOR3_X1 U9928 ( .A1(n8585), .A2(n8584), .A3(n8583), .ZN(n8586) );
  OAI21_X1 U9929 ( .B1(n8588), .B2(n8587), .A(n8586), .ZN(n8594) );
  XNOR2_X1 U9930 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_116), .ZN(n8593) );
  XNOR2_X1 U9931 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_119), .ZN(n8591) );
  XNOR2_X1 U9932 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_118), .ZN(n8590) );
  XNOR2_X1 U9933 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_117), .ZN(n8589) );
  NAND3_X1 U9934 ( .A1(n8591), .A2(n8590), .A3(n8589), .ZN(n8592) );
  AOI21_X1 U9935 ( .B1(n8594), .B2(n8593), .A(n8592), .ZN(n8597) );
  XNOR2_X1 U9936 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_120), .ZN(n8596) );
  XNOR2_X1 U9937 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_121), .ZN(n8595) );
  OAI21_X1 U9938 ( .B1(n8597), .B2(n8596), .A(n8595), .ZN(n8604) );
  INV_X1 U9939 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10600) );
  OAI22_X1 U9940 ( .A1(n10600), .A2(keyinput_124), .B1(P1_D_REG_4__SCAN_IN), 
        .B2(keyinput_126), .ZN(n8598) );
  AOI221_X1 U9941 ( .B1(n10600), .B2(keyinput_124), .C1(keyinput_126), .C2(
        P1_D_REG_4__SCAN_IN), .A(n8598), .ZN(n8603) );
  XOR2_X1 U9942 ( .A(P1_D_REG_1__SCAN_IN), .B(keyinput_123), .Z(n8602) );
  INV_X1 U9943 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n8600) );
  OAI22_X1 U9944 ( .A1(n8600), .A2(keyinput_122), .B1(keyinput_125), .B2(
        P1_D_REG_3__SCAN_IN), .ZN(n8599) );
  AOI221_X1 U9945 ( .B1(n8600), .B2(keyinput_122), .C1(P1_D_REG_3__SCAN_IN), 
        .C2(keyinput_125), .A(n8599), .ZN(n8601) );
  NAND4_X1 U9946 ( .A1(n8604), .A2(n8603), .A3(n8602), .A4(n8601), .ZN(n8606)
         );
  XNOR2_X1 U9947 ( .A(keyinput_127), .B(P1_D_REG_5__SCAN_IN), .ZN(n8605) );
  OAI211_X1 U9948 ( .C1(n8608), .C2(n8607), .A(n8606), .B(n8605), .ZN(n8614)
         );
  NAND2_X1 U9949 ( .A1(n8609), .A2(n5180), .ZN(n8611) );
  OAI211_X1 U9950 ( .C1(n8618), .C2(n8612), .A(n8611), .B(n8610), .ZN(n8613)
         );
  XNOR2_X1 U9951 ( .A(n8614), .B(n8613), .ZN(P2_U3267) );
  OAI222_X1 U9952 ( .A1(n8618), .A2(n8617), .B1(n9719), .B2(n8616), .C1(n8615), 
        .C2(P2_U3151), .ZN(P2_U3270) );
  XOR2_X1 U9953 ( .A(n10088), .B(n8619), .Z(n10544) );
  XNOR2_X1 U9954 ( .A(n8620), .B(n10088), .ZN(n8621) );
  OAI222_X1 U9955 ( .A1(n10902), .A2(n9798), .B1(n10900), .B2(n8622), .C1(
        n11030), .C2(n8621), .ZN(n10538) );
  INV_X1 U9956 ( .A(n8623), .ZN(n8626) );
  INV_X1 U9957 ( .A(n8624), .ZN(n8625) );
  AOI211_X1 U9958 ( .C1(n10540), .C2(n8626), .A(n10438), .B(n8625), .ZN(n10539) );
  NAND2_X1 U9959 ( .A1(n10539), .A2(n11045), .ZN(n8629) );
  AOI22_X1 U9960 ( .A1(n11051), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8627), .B2(
        n10393), .ZN(n8628) );
  OAI211_X1 U9961 ( .C1(n8630), .C2(n10440), .A(n8629), .B(n8628), .ZN(n8631)
         );
  AOI21_X1 U9962 ( .B1(n10915), .B2(n10538), .A(n8631), .ZN(n8632) );
  OAI21_X1 U9963 ( .B1(n10544), .B2(n10452), .A(n8632), .ZN(P1_U3278) );
  XNOR2_X1 U9964 ( .A(n8633), .B(n9199), .ZN(n8641) );
  OAI21_X1 U9965 ( .B1(n9173), .B2(n8635), .A(n8634), .ZN(n8636) );
  AOI21_X1 U9966 ( .B1(n9152), .B2(n9200), .A(n8636), .ZN(n8637) );
  OAI21_X1 U9967 ( .B1(n8638), .B2(n9183), .A(n8637), .ZN(n8639) );
  AOI21_X1 U9968 ( .B1(n11010), .B2(n9190), .A(n8639), .ZN(n8640) );
  OAI21_X1 U9969 ( .B1(n8641), .B2(n9185), .A(n8640), .ZN(P2_U3157) );
  INV_X1 U9970 ( .A(n8642), .ZN(n8643) );
  NAND2_X1 U9971 ( .A1(n8643), .A2(SI_29_), .ZN(n8647) );
  NAND2_X1 U9972 ( .A1(n8647), .A2(n8646), .ZN(n8655) );
  INV_X1 U9973 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9030) );
  INV_X1 U9974 ( .A(SI_30_), .ZN(n8648) );
  NAND2_X1 U9975 ( .A1(n8649), .A2(n8648), .ZN(n8660) );
  INV_X1 U9976 ( .A(n8649), .ZN(n8650) );
  NAND2_X1 U9977 ( .A1(n8650), .A2(SI_30_), .ZN(n8651) );
  NAND2_X1 U9978 ( .A1(n8660), .A2(n8651), .ZN(n8654) );
  INV_X1 U9979 ( .A(n8654), .ZN(n8652) );
  NAND2_X1 U9980 ( .A1(n8655), .A2(n8654), .ZN(n8656) );
  INV_X1 U9981 ( .A(n8658), .ZN(n9029) );
  OAI222_X1 U9982 ( .A1(n5707), .A2(P1_U3086), .B1(n8657), .B2(n9029), .C1(
        n9894), .C2(n10595), .ZN(P1_U3325) );
  OR2_X1 U9983 ( .A1(n6360), .A2(n9030), .ZN(n8659) );
  MUX2_X1 U9984 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n8662), .Z(n8664) );
  XNOR2_X1 U9985 ( .A(n8664), .B(n8663), .ZN(n8665) );
  NAND2_X1 U9986 ( .A1(n10593), .A2(n6416), .ZN(n8668) );
  INV_X1 U9987 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9712) );
  OR2_X1 U9988 ( .A1(n6360), .A2(n9712), .ZN(n8667) );
  INV_X1 U9989 ( .A(n9380), .ZN(n9080) );
  NAND2_X1 U9990 ( .A1(n9072), .A2(n9080), .ZN(n8669) );
  NAND2_X1 U9991 ( .A1(n8670), .A2(n8669), .ZN(n8672) );
  OR2_X1 U9992 ( .A1(n9072), .A2(n9080), .ZN(n8671) );
  INV_X1 U9993 ( .A(n9018), .ZN(n8677) );
  NAND2_X1 U9994 ( .A1(n9716), .A2(n6416), .ZN(n8674) );
  OR2_X1 U9995 ( .A1(n6360), .A2(n9717), .ZN(n8673) );
  NAND2_X1 U9996 ( .A1(n9596), .A2(n8675), .ZN(n8842) );
  INV_X1 U9997 ( .A(n8842), .ZN(n8848) );
  OR2_X1 U9998 ( .A1(n8885), .A2(n9365), .ZN(n8688) );
  INV_X1 U9999 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8683) );
  NAND2_X1 U10000 ( .A1(n8678), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8682) );
  INV_X1 U10001 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8679) );
  OR2_X1 U10002 ( .A1(n6338), .A2(n8679), .ZN(n8681) );
  OAI211_X1 U10003 ( .C1(n8683), .C2(n5110), .A(n8682), .B(n8681), .ZN(n8684)
         );
  INV_X1 U10004 ( .A(n8684), .ZN(n8685) );
  NAND2_X1 U10005 ( .A1(n8686), .A2(n8685), .ZN(n9192) );
  INV_X1 U10006 ( .A(n9192), .ZN(n8690) );
  NAND2_X1 U10007 ( .A1(n8691), .A2(n8690), .ZN(n8687) );
  OAI211_X1 U10008 ( .C1(n9661), .C2(n8885), .A(n8689), .B(n8854), .ZN(n8891)
         );
  NAND3_X1 U10009 ( .A1(n8883), .A2(n8836), .A3(n8843), .ZN(n8851) );
  NOR2_X1 U10010 ( .A1(n9072), .A2(n8847), .ZN(n8692) );
  NOR2_X1 U10011 ( .A1(n9072), .A2(n9380), .ZN(n9014) );
  MUX2_X1 U10012 ( .A(n8694), .B(n8693), .S(n8836), .Z(n8835) );
  OR2_X1 U10013 ( .A1(n8830), .A2(n5605), .ZN(n9409) );
  INV_X1 U10014 ( .A(n9409), .ZN(n9412) );
  INV_X1 U10015 ( .A(n9429), .ZN(n8825) );
  MUX2_X1 U10016 ( .A(n8825), .B(n8826), .S(n8836), .Z(n8698) );
  NAND2_X1 U10017 ( .A1(n9421), .A2(n9437), .ZN(n8695) );
  MUX2_X1 U10018 ( .A(n8696), .B(n8695), .S(n8836), .Z(n8697) );
  OAI21_X1 U10019 ( .B1(n9422), .B2(n8698), .A(n8697), .ZN(n8829) );
  NAND2_X1 U10020 ( .A1(n8699), .A2(n8879), .ZN(n8701) );
  NAND3_X1 U10021 ( .A1(n8706), .A2(n8701), .A3(n8700), .ZN(n8702) );
  NAND2_X1 U10022 ( .A1(n8702), .A2(n6683), .ZN(n8703) );
  NAND2_X1 U10023 ( .A1(n8703), .A2(n8859), .ZN(n8704) );
  NAND3_X1 U10024 ( .A1(n8704), .A2(n8721), .A3(n10929), .ZN(n8713) );
  NAND2_X1 U10025 ( .A1(n6683), .A2(n8705), .ZN(n8707) );
  NAND2_X1 U10026 ( .A1(n8707), .A2(n8706), .ZN(n8708) );
  NAND2_X1 U10027 ( .A1(n8859), .A2(n8708), .ZN(n8709) );
  OAI211_X1 U10028 ( .C1(n8711), .C2(n8710), .A(n8709), .B(n8716), .ZN(n8712)
         );
  MUX2_X1 U10029 ( .A(n8713), .B(n8712), .S(n8836), .Z(n8715) );
  NAND2_X1 U10030 ( .A1(n8715), .A2(n8714), .ZN(n8724) );
  INV_X1 U10031 ( .A(n8716), .ZN(n8718) );
  OAI211_X1 U10032 ( .C1(n8724), .C2(n8718), .A(n8725), .B(n8717), .ZN(n8720)
         );
  NAND3_X1 U10033 ( .A1(n8720), .A2(n8719), .A3(n8726), .ZN(n8731) );
  INV_X1 U10034 ( .A(n8721), .ZN(n8723) );
  OAI21_X1 U10035 ( .B1(n8724), .B2(n8723), .A(n8722), .ZN(n8729) );
  AND2_X1 U10036 ( .A1(n8725), .A2(n8745), .ZN(n8728) );
  INV_X1 U10037 ( .A(n8726), .ZN(n8727) );
  AOI21_X1 U10038 ( .B1(n8729), .B2(n8728), .A(n8727), .ZN(n8730) );
  MUX2_X1 U10039 ( .A(n8731), .B(n8730), .S(n8836), .Z(n8738) );
  NAND2_X1 U10040 ( .A1(n8733), .A2(n8732), .ZN(n8735) );
  INV_X1 U10041 ( .A(n8740), .ZN(n8734) );
  MUX2_X1 U10042 ( .A(n8735), .B(n8734), .S(n8847), .Z(n8743) );
  INV_X1 U10043 ( .A(n8741), .ZN(n8736) );
  NOR2_X1 U10044 ( .A1(n8743), .A2(n8736), .ZN(n8749) );
  NAND3_X1 U10045 ( .A1(n8738), .A2(n8737), .A3(n8749), .ZN(n8748) );
  AND2_X1 U10046 ( .A1(n8740), .A2(n8739), .ZN(n8742) );
  OAI211_X1 U10047 ( .C1(n8743), .C2(n8742), .A(n8741), .B(n8753), .ZN(n8744)
         );
  NAND2_X1 U10048 ( .A1(n8744), .A2(n8836), .ZN(n8747) );
  NOR2_X1 U10049 ( .A1(n8745), .A2(n8836), .ZN(n8746) );
  AOI21_X1 U10050 ( .B1(n8748), .B2(n8747), .A(n8746), .ZN(n8756) );
  INV_X1 U10051 ( .A(n8749), .ZN(n8752) );
  OAI21_X1 U10052 ( .B1(n8752), .B2(n8751), .A(n8750), .ZN(n8754) );
  OAI211_X1 U10053 ( .C1(n8756), .C2(n8754), .A(n8753), .B(n8759), .ZN(n8755)
         );
  NAND2_X1 U10054 ( .A1(n8755), .A2(n8758), .ZN(n8763) );
  INV_X1 U10055 ( .A(n8756), .ZN(n8761) );
  NAND2_X1 U10056 ( .A1(n8758), .A2(n8757), .ZN(n8760) );
  OAI21_X1 U10057 ( .B1(n8761), .B2(n8760), .A(n8759), .ZN(n8762) );
  MUX2_X1 U10058 ( .A(n8763), .B(n8762), .S(n8836), .Z(n8764) );
  NAND2_X1 U10059 ( .A1(n8764), .A2(n8868), .ZN(n8768) );
  MUX2_X1 U10060 ( .A(n8766), .B(n8765), .S(n8836), .Z(n8767) );
  NAND3_X1 U10061 ( .A1(n8768), .A2(n9585), .A3(n8767), .ZN(n8772) );
  MUX2_X1 U10062 ( .A(n8770), .B(n8769), .S(n8847), .Z(n8771) );
  NAND2_X1 U10063 ( .A1(n8772), .A2(n8771), .ZN(n8783) );
  NAND2_X1 U10064 ( .A1(n8783), .A2(n6699), .ZN(n8780) );
  INV_X1 U10065 ( .A(n8773), .ZN(n11094) );
  AND2_X1 U10066 ( .A1(n8777), .A2(n11094), .ZN(n8775) );
  INV_X1 U10067 ( .A(n8776), .ZN(n8774) );
  AOI21_X1 U10068 ( .B1(n8780), .B2(n8775), .A(n8774), .ZN(n8782) );
  AND2_X1 U10069 ( .A1(n8776), .A2(n9179), .ZN(n8779) );
  INV_X1 U10070 ( .A(n8777), .ZN(n8778) );
  AOI21_X1 U10071 ( .B1(n8780), .B2(n8779), .A(n8778), .ZN(n8781) );
  MUX2_X1 U10072 ( .A(n8782), .B(n8781), .S(n8836), .Z(n8792) );
  INV_X1 U10073 ( .A(n8783), .ZN(n8786) );
  NOR2_X1 U10074 ( .A1(n9551), .A2(n8784), .ZN(n8785) );
  AOI21_X1 U10075 ( .B1(n8786), .B2(n8785), .A(n9536), .ZN(n8791) );
  MUX2_X1 U10076 ( .A(n8788), .B(n8787), .S(n8836), .Z(n8789) );
  INV_X1 U10077 ( .A(n8789), .ZN(n8790) );
  AOI21_X1 U10078 ( .B1(n8792), .B2(n8791), .A(n8790), .ZN(n8796) );
  MUX2_X1 U10079 ( .A(n9530), .B(n9521), .S(n8836), .Z(n8797) );
  NAND2_X1 U10080 ( .A1(n8801), .A2(n9530), .ZN(n8794) );
  NAND2_X1 U10081 ( .A1(n8800), .A2(n9521), .ZN(n8793) );
  MUX2_X1 U10082 ( .A(n8794), .B(n8793), .S(n8847), .Z(n8795) );
  AOI21_X1 U10083 ( .B1(n8796), .B2(n8797), .A(n8795), .ZN(n8808) );
  INV_X1 U10084 ( .A(n8796), .ZN(n8799) );
  INV_X1 U10085 ( .A(n8797), .ZN(n8798) );
  NAND3_X1 U10086 ( .A1(n8799), .A2(n9501), .A3(n8798), .ZN(n8803) );
  MUX2_X1 U10087 ( .A(n8801), .B(n8800), .S(n8836), .Z(n8802) );
  NAND3_X1 U10088 ( .A1(n8803), .A2(n9041), .A3(n8802), .ZN(n8807) );
  NAND2_X1 U10089 ( .A1(n9092), .A2(n9504), .ZN(n8804) );
  MUX2_X1 U10090 ( .A(n8805), .B(n8804), .S(n8836), .Z(n8806) );
  OAI211_X1 U10091 ( .C1(n8808), .C2(n8807), .A(n8806), .B(n9469), .ZN(n8814)
         );
  INV_X1 U10092 ( .A(n9105), .ZN(n9684) );
  MUX2_X1 U10093 ( .A(n9471), .B(n9684), .S(n8836), .Z(n8815) );
  NAND2_X1 U10094 ( .A1(n9195), .A2(n8836), .ZN(n8810) );
  NAND3_X1 U10095 ( .A1(n9474), .A2(n9488), .A3(n8847), .ZN(n8809) );
  OAI21_X1 U10096 ( .B1(n8810), .B2(n9474), .A(n8809), .ZN(n8811) );
  AOI21_X1 U10097 ( .B1(n8815), .B2(n8812), .A(n8811), .ZN(n8813) );
  NAND2_X1 U10098 ( .A1(n8814), .A2(n8813), .ZN(n8820) );
  INV_X1 U10099 ( .A(n9451), .ZN(n8819) );
  INV_X1 U10100 ( .A(n8815), .ZN(n8817) );
  NAND2_X1 U10101 ( .A1(n9105), .A2(n9447), .ZN(n8816) );
  NAND2_X1 U10102 ( .A1(n8817), .A2(n8816), .ZN(n8818) );
  NAND3_X1 U10103 ( .A1(n8820), .A2(n8819), .A3(n8818), .ZN(n8824) );
  MUX2_X1 U10104 ( .A(n8822), .B(n8821), .S(n8847), .Z(n8823) );
  NAND2_X1 U10105 ( .A1(n8824), .A2(n8823), .ZN(n8827) );
  OR2_X1 U10106 ( .A1(n8826), .A2(n8825), .ZN(n9438) );
  INV_X1 U10107 ( .A(n9438), .ZN(n9434) );
  NAND3_X1 U10108 ( .A1(n8827), .A2(n6708), .A3(n9434), .ZN(n8828) );
  NAND3_X1 U10109 ( .A1(n9412), .A2(n8829), .A3(n8828), .ZN(n8833) );
  MUX2_X1 U10110 ( .A(n8830), .B(n5605), .S(n8836), .Z(n8831) );
  INV_X1 U10111 ( .A(n8831), .ZN(n8832) );
  NAND3_X1 U10112 ( .A1(n8833), .A2(n9395), .A3(n8832), .ZN(n8834) );
  NAND3_X1 U10113 ( .A1(n9387), .A2(n8835), .A3(n8834), .ZN(n8840) );
  NAND2_X1 U10114 ( .A1(n9601), .A2(n9174), .ZN(n8837) );
  MUX2_X1 U10115 ( .A(n8838), .B(n8837), .S(n8836), .Z(n8839) );
  NAND2_X1 U10116 ( .A1(n8840), .A2(n8839), .ZN(n8841) );
  OAI21_X1 U10117 ( .B1(n8844), .B2(n9014), .A(n8841), .ZN(n8846) );
  NAND2_X1 U10118 ( .A1(n9072), .A2(n9380), .ZN(n9013) );
  AOI21_X1 U10119 ( .B1(n8844), .B2(n9013), .A(n9016), .ZN(n8845) );
  OAI211_X1 U10120 ( .C1(n8852), .C2(n8848), .A(n8847), .B(n8883), .ZN(n8850)
         );
  INV_X1 U10121 ( .A(n8854), .ZN(n8881) );
  INV_X1 U10122 ( .A(n9387), .ZN(n8877) );
  INV_X1 U10123 ( .A(n9041), .ZN(n9489) );
  NOR4_X1 U10124 ( .A1(n8858), .A2(n8855), .A3(n8857), .A4(n8856), .ZN(n8862)
         );
  NAND4_X1 U10125 ( .A1(n8862), .A2(n8861), .A3(n8860), .A4(n8859), .ZN(n8866)
         );
  NOR4_X1 U10126 ( .A1(n8866), .A2(n8865), .A3(n8864), .A4(n8863), .ZN(n8870)
         );
  NAND4_X1 U10127 ( .A1(n8870), .A2(n8869), .A3(n8868), .A4(n8867), .ZN(n8871)
         );
  NOR4_X1 U10128 ( .A1(n9551), .A2(n9570), .A3(n6483), .A4(n8871), .ZN(n8873)
         );
  NAND4_X1 U10129 ( .A1(n9501), .A2(n6701), .A3(n8873), .A4(n8872), .ZN(n8874)
         );
  NOR4_X1 U10130 ( .A1(n9451), .A2(n9489), .A3(n9473), .A4(n8874), .ZN(n8875)
         );
  NAND4_X1 U10131 ( .A1(n9412), .A2(n9434), .A3(n8875), .A4(n9457), .ZN(n8876)
         );
  NOR4_X1 U10132 ( .A1(n8877), .A2(n9422), .A3(n8876), .A4(n5343), .ZN(n8878)
         );
  NAND4_X1 U10133 ( .A1(n8883), .A2(n9017), .A3(n8878), .A4(n9067), .ZN(n8880)
         );
  OAI21_X1 U10134 ( .B1(n8881), .B2(n8880), .A(n8879), .ZN(n8882) );
  INV_X1 U10135 ( .A(n8883), .ZN(n8884) );
  NOR2_X1 U10136 ( .A1(n8884), .A2(n9365), .ZN(n8886) );
  XNOR2_X1 U10137 ( .A(n8893), .B(n8892), .ZN(n8900) );
  NAND3_X1 U10138 ( .A1(n8895), .A2(n8894), .A3(n9327), .ZN(n8896) );
  OAI211_X1 U10139 ( .C1(n8897), .C2(n8899), .A(n8896), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8898) );
  OAI21_X1 U10140 ( .B1(n8900), .B2(n8899), .A(n8898), .ZN(P2_U3296) );
  NAND2_X1 U10141 ( .A1(n9789), .A2(n9000), .ZN(n8904) );
  OR2_X1 U10142 ( .A1(n9798), .A2(n7115), .ZN(n8903) );
  NAND2_X1 U10143 ( .A1(n8904), .A2(n8903), .ZN(n8905) );
  XNOR2_X1 U10144 ( .A(n8905), .B(n8974), .ZN(n8908) );
  NOR2_X1 U10145 ( .A1(n9798), .A2(n9001), .ZN(n8906) );
  AOI21_X1 U10146 ( .B1(n9789), .B2(n8938), .A(n8906), .ZN(n8907) );
  NAND2_X1 U10147 ( .A1(n8908), .A2(n8907), .ZN(n8910) );
  OR2_X1 U10148 ( .A1(n8908), .A2(n8907), .ZN(n8909) );
  AND2_X1 U10149 ( .A1(n8910), .A2(n8909), .ZN(n9782) );
  NAND2_X1 U10150 ( .A1(n9780), .A2(n8910), .ZN(n9797) );
  NAND2_X1 U10151 ( .A1(n10535), .A2(n9000), .ZN(n8912) );
  OR2_X1 U10152 ( .A1(n9860), .A2(n7115), .ZN(n8911) );
  NAND2_X1 U10153 ( .A1(n8912), .A2(n8911), .ZN(n8913) );
  XNOR2_X1 U10154 ( .A(n8913), .B(n9002), .ZN(n8916) );
  NAND2_X1 U10155 ( .A1(n10535), .A2(n8961), .ZN(n8915) );
  OR2_X1 U10156 ( .A1(n9860), .A2(n9001), .ZN(n8914) );
  NAND2_X1 U10157 ( .A1(n8915), .A2(n8914), .ZN(n8917) );
  NAND2_X1 U10158 ( .A1(n8916), .A2(n8917), .ZN(n9795) );
  NAND2_X1 U10159 ( .A1(n9797), .A2(n9795), .ZN(n8920) );
  INV_X1 U10160 ( .A(n8916), .ZN(n8919) );
  INV_X1 U10161 ( .A(n8917), .ZN(n8918) );
  NAND2_X1 U10162 ( .A1(n8919), .A2(n8918), .ZN(n9794) );
  NOR2_X1 U10163 ( .A1(n9799), .A2(n7115), .ZN(n8921) );
  AOI21_X1 U10164 ( .B1(n9864), .B2(n9000), .A(n8921), .ZN(n8922) );
  XNOR2_X1 U10165 ( .A(n8922), .B(n9002), .ZN(n8942) );
  NAND2_X1 U10166 ( .A1(n10522), .A2(n9000), .ZN(n8924) );
  NAND2_X1 U10167 ( .A1(n8961), .A2(n10157), .ZN(n8923) );
  NAND2_X1 U10168 ( .A1(n8924), .A2(n8923), .ZN(n8925) );
  XNOR2_X1 U10169 ( .A(n8925), .B(n9002), .ZN(n8945) );
  INV_X1 U10170 ( .A(n8945), .ZN(n8927) );
  AND2_X1 U10171 ( .A1(n8976), .A2(n10157), .ZN(n8926) );
  AOI21_X1 U10172 ( .B1(n10522), .B2(n8961), .A(n8926), .ZN(n8944) );
  NAND2_X1 U10173 ( .A1(n8927), .A2(n8944), .ZN(n9759) );
  NAND2_X1 U10174 ( .A1(n10432), .A2(n9000), .ZN(n8929) );
  OR2_X1 U10175 ( .A1(n10449), .A2(n7115), .ZN(n8928) );
  NAND2_X1 U10176 ( .A1(n8929), .A2(n8928), .ZN(n8930) );
  XNOR2_X1 U10177 ( .A(n8930), .B(n8974), .ZN(n8933) );
  NOR2_X1 U10178 ( .A1(n10449), .A2(n9001), .ZN(n8931) );
  AOI21_X1 U10179 ( .B1(n10432), .B2(n8961), .A(n8931), .ZN(n8932) );
  OR2_X1 U10180 ( .A1(n8933), .A2(n8932), .ZN(n8949) );
  INV_X1 U10181 ( .A(n8949), .ZN(n8941) );
  XNOR2_X1 U10182 ( .A(n8933), .B(n8932), .ZN(n9762) );
  INV_X1 U10183 ( .A(n9762), .ZN(n8940) );
  NAND2_X1 U10184 ( .A1(n10517), .A2(n9000), .ZN(n8935) );
  OR2_X1 U10185 ( .A1(n10426), .A2(n7115), .ZN(n8934) );
  NAND2_X1 U10186 ( .A1(n8935), .A2(n8934), .ZN(n8936) );
  XNOR2_X1 U10187 ( .A(n8936), .B(n9002), .ZN(n8948) );
  INV_X1 U10188 ( .A(n8948), .ZN(n8939) );
  NOR2_X1 U10189 ( .A1(n10426), .A2(n9001), .ZN(n8937) );
  AOI21_X1 U10190 ( .B1(n10517), .B2(n8938), .A(n8937), .ZN(n8947) );
  NAND2_X1 U10191 ( .A1(n8939), .A2(n8947), .ZN(n9761) );
  AND2_X1 U10192 ( .A1(n8940), .A2(n9761), .ZN(n9764) );
  NOR2_X1 U10193 ( .A1(n9799), .A2(n9001), .ZN(n8943) );
  AOI21_X1 U10194 ( .B1(n9864), .B2(n8961), .A(n8943), .ZN(n9857) );
  XNOR2_X1 U10195 ( .A(n8945), .B(n8944), .ZN(n9757) );
  INV_X1 U10196 ( .A(n8946), .ZN(n8951) );
  XNOR2_X1 U10197 ( .A(n8948), .B(n8947), .ZN(n9827) );
  AND2_X1 U10198 ( .A1(n9827), .A2(n8949), .ZN(n8950) );
  INV_X1 U10199 ( .A(n9732), .ZN(n8971) );
  AOI22_X1 U10200 ( .A1(n10501), .A2(n9000), .B1(n8961), .B2(n10376), .ZN(
        n8954) );
  XOR2_X1 U10201 ( .A(n9002), .B(n8954), .Z(n9734) );
  NAND2_X1 U10202 ( .A1(n10501), .A2(n8961), .ZN(n8956) );
  NAND2_X1 U10203 ( .A1(n8976), .A2(n10376), .ZN(n8955) );
  NAND2_X1 U10204 ( .A1(n8956), .A2(n8955), .ZN(n8965) );
  NAND2_X1 U10205 ( .A1(n10507), .A2(n9000), .ZN(n8958) );
  OR2_X1 U10206 ( .A1(n10425), .A2(n7115), .ZN(n8957) );
  NAND2_X1 U10207 ( .A1(n8958), .A2(n8957), .ZN(n8959) );
  XNOR2_X1 U10208 ( .A(n8959), .B(n8974), .ZN(n9730) );
  NOR2_X1 U10209 ( .A1(n10425), .A2(n9001), .ZN(n8960) );
  AOI21_X1 U10210 ( .B1(n10507), .B2(n8961), .A(n8960), .ZN(n9838) );
  NOR2_X1 U10211 ( .A1(n9730), .A2(n9838), .ZN(n8962) );
  NAND2_X1 U10212 ( .A1(n9730), .A2(n9838), .ZN(n8964) );
  AOI21_X1 U10213 ( .B1(n8965), .B2(n8964), .A(n9734), .ZN(n8963) );
  INV_X1 U10214 ( .A(n8963), .ZN(n8968) );
  INV_X1 U10215 ( .A(n8964), .ZN(n8966) );
  INV_X1 U10216 ( .A(n8965), .ZN(n9733) );
  NAND2_X1 U10217 ( .A1(n10382), .A2(n9000), .ZN(n8973) );
  NAND2_X1 U10218 ( .A1(n8938), .A2(n10400), .ZN(n8972) );
  NAND2_X1 U10219 ( .A1(n8973), .A2(n8972), .ZN(n8975) );
  XNOR2_X1 U10220 ( .A(n8975), .B(n8974), .ZN(n8979) );
  AND2_X1 U10221 ( .A1(n8976), .A2(n10400), .ZN(n8977) );
  AOI21_X1 U10222 ( .B1(n10382), .B2(n8938), .A(n8977), .ZN(n8978) );
  NOR2_X1 U10223 ( .A1(n8979), .A2(n8978), .ZN(n9808) );
  NAND2_X1 U10224 ( .A1(n8979), .A2(n8978), .ZN(n9807) );
  OAI22_X1 U10225 ( .A1(n10365), .A2(n7115), .B1(n9875), .B2(n9001), .ZN(n8988) );
  NAND2_X1 U10226 ( .A1(n10491), .A2(n9000), .ZN(n8981) );
  NAND2_X1 U10227 ( .A1(n8938), .A2(n10375), .ZN(n8980) );
  NAND2_X1 U10228 ( .A1(n8981), .A2(n8980), .ZN(n8982) );
  XNOR2_X1 U10229 ( .A(n8982), .B(n9002), .ZN(n8987) );
  XOR2_X1 U10230 ( .A(n8988), .B(n8987), .Z(n9773) );
  NAND2_X1 U10231 ( .A1(n10350), .A2(n9000), .ZN(n8984) );
  OR2_X1 U10232 ( .A1(n10325), .A2(n7115), .ZN(n8983) );
  NAND2_X1 U10233 ( .A1(n8984), .A2(n8983), .ZN(n8985) );
  XNOR2_X1 U10234 ( .A(n8985), .B(n9002), .ZN(n8997) );
  NOR2_X1 U10235 ( .A1(n10325), .A2(n9001), .ZN(n8986) );
  AOI21_X1 U10236 ( .B1(n10350), .B2(n8961), .A(n8986), .ZN(n8995) );
  XNOR2_X1 U10237 ( .A(n8997), .B(n8995), .ZN(n9872) );
  INV_X1 U10238 ( .A(n8987), .ZN(n8990) );
  INV_X1 U10239 ( .A(n8988), .ZN(n8989) );
  NAND2_X1 U10240 ( .A1(n8990), .A2(n8989), .ZN(n9868) );
  OAI22_X1 U10241 ( .A1(n10484), .A2(n8991), .B1(n10309), .B2(n7115), .ZN(
        n8992) );
  XNOR2_X1 U10242 ( .A(n8992), .B(n9002), .ZN(n8994) );
  OAI22_X1 U10243 ( .A1(n10484), .A2(n7115), .B1(n10309), .B2(n9001), .ZN(
        n8993) );
  NOR2_X1 U10244 ( .A1(n8994), .A2(n8993), .ZN(n8998) );
  AOI21_X1 U10245 ( .B1(n8994), .B2(n8993), .A(n8998), .ZN(n9722) );
  INV_X1 U10246 ( .A(n8995), .ZN(n8996) );
  NAND2_X1 U10247 ( .A1(n8997), .A2(n8996), .ZN(n9723) );
  NAND3_X1 U10248 ( .A1(n9870), .A2(n9722), .A3(n9723), .ZN(n9721) );
  INV_X1 U10249 ( .A(n8998), .ZN(n8999) );
  NAND2_X1 U10250 ( .A1(n9721), .A2(n8999), .ZN(n9007) );
  AOI22_X1 U10251 ( .A1(n10553), .A2(n9000), .B1(n8938), .B2(n6159), .ZN(n9005) );
  OAI22_X1 U10252 ( .A1(n10477), .A2(n7115), .B1(n10326), .B2(n9001), .ZN(
        n9003) );
  XNOR2_X1 U10253 ( .A(n9003), .B(n9002), .ZN(n9004) );
  XOR2_X1 U10254 ( .A(n9005), .B(n9004), .Z(n9006) );
  XNOR2_X1 U10255 ( .A(n9007), .B(n9006), .ZN(n9012) );
  OAI22_X1 U10256 ( .A1(n9874), .A2(n10317), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9008), .ZN(n9010) );
  OAI22_X1 U10257 ( .A1(n10310), .A2(n9877), .B1(n9876), .B2(n10309), .ZN(
        n9009) );
  AOI211_X1 U10258 ( .C1(n10553), .C2(n9863), .A(n9010), .B(n9009), .ZN(n9011)
         );
  OAI21_X1 U10259 ( .B1(n9012), .B2(n9866), .A(n9011), .ZN(P1_U3220) );
  NAND2_X1 U10260 ( .A1(n6313), .A2(P2_B_REG_SCAN_IN), .ZN(n9019) );
  AND2_X1 U10261 ( .A1(n10926), .A2(n9019), .ZN(n9363) );
  AOI22_X1 U10262 ( .A1(n6677), .A2(n9380), .B1(n9192), .B2(n9363), .ZN(n9020)
         );
  OAI21_X1 U10263 ( .B1(n9593), .B2(n9021), .A(n9020), .ZN(n9022) );
  NAND2_X1 U10264 ( .A1(n9023), .A2(n9550), .ZN(n9366) );
  OAI21_X1 U10265 ( .B1(n10944), .B2(n9024), .A(n9366), .ZN(n9027) );
  NOR2_X1 U10266 ( .A1(n9593), .A2(n9025), .ZN(n9026) );
  AOI211_X1 U10267 ( .C1(n9509), .C2(n9596), .A(n9027), .B(n9026), .ZN(n9028)
         );
  OAI21_X1 U10268 ( .B1(n9600), .B2(n10946), .A(n9028), .ZN(P2_U3204) );
  OAI222_X1 U10269 ( .A1(n8618), .A2(n9030), .B1(n9719), .B2(n9029), .C1(n6293), .C2(P2_U3151), .ZN(P2_U3265) );
  XNOR2_X1 U10270 ( .A(n9553), .B(n9050), .ZN(n9035) );
  INV_X1 U10271 ( .A(n9035), .ZN(n9036) );
  INV_X1 U10272 ( .A(n9031), .ZN(n9032) );
  XOR2_X1 U10273 ( .A(n9529), .B(n9035), .Z(n9187) );
  NOR2_X1 U10274 ( .A1(n9186), .A2(n9187), .ZN(n9184) );
  XOR2_X1 U10275 ( .A(n9050), .B(n9537), .Z(n9115) );
  XNOR2_X1 U10276 ( .A(n9521), .B(n9050), .ZN(n9124) );
  NOR2_X1 U10277 ( .A1(n9124), .A2(n9503), .ZN(n9039) );
  INV_X1 U10278 ( .A(n9124), .ZN(n9038) );
  XNOR2_X1 U10279 ( .A(n9510), .B(n9050), .ZN(n9040) );
  XOR2_X1 U10280 ( .A(n9516), .B(n9040), .Z(n9158) );
  OR2_X1 U10281 ( .A1(n9094), .A2(n9504), .ZN(n9042) );
  XNOR2_X1 U10282 ( .A(n9474), .B(n9050), .ZN(n9043) );
  XOR2_X1 U10283 ( .A(n9195), .B(n9043), .Z(n9142) );
  NAND2_X1 U10284 ( .A1(n9043), .A2(n9488), .ZN(n9044) );
  XNOR2_X1 U10285 ( .A(n9105), .B(n9050), .ZN(n9045) );
  XNOR2_X1 U10286 ( .A(n9045), .B(n9447), .ZN(n9101) );
  XOR2_X1 U10287 ( .A(n9460), .B(n9046), .Z(n9150) );
  XNOR2_X1 U10288 ( .A(n9440), .B(n9050), .ZN(n9052) );
  NAND2_X1 U10289 ( .A1(n9085), .A2(n9426), .ZN(n9055) );
  INV_X1 U10290 ( .A(n9051), .ZN(n9053) );
  NAND2_X1 U10291 ( .A1(n9055), .A2(n9054), .ZN(n9132) );
  XNOR2_X1 U10292 ( .A(n9421), .B(n9050), .ZN(n9056) );
  NAND2_X1 U10293 ( .A1(n9132), .A2(n9133), .ZN(n9058) );
  NAND2_X1 U10294 ( .A1(n9056), .A2(n9437), .ZN(n9057) );
  NAND2_X1 U10295 ( .A1(n9058), .A2(n9057), .ZN(n9108) );
  XNOR2_X1 U10296 ( .A(n9411), .B(n9050), .ZN(n9059) );
  XNOR2_X1 U10297 ( .A(n9059), .B(n9398), .ZN(n9109) );
  NAND2_X1 U10298 ( .A1(n9108), .A2(n9109), .ZN(n9061) );
  NAND2_X1 U10299 ( .A1(n9059), .A2(n9425), .ZN(n9060) );
  NAND2_X1 U10300 ( .A1(n9061), .A2(n9060), .ZN(n9167) );
  XNOR2_X1 U10301 ( .A(n9406), .B(n9050), .ZN(n9062) );
  XNOR2_X1 U10302 ( .A(n9062), .B(n9381), .ZN(n9168) );
  NAND2_X1 U10303 ( .A1(n9167), .A2(n9168), .ZN(n9064) );
  NAND2_X1 U10304 ( .A1(n9062), .A2(n9415), .ZN(n9063) );
  XNOR2_X1 U10305 ( .A(n9601), .B(n7079), .ZN(n9065) );
  NAND2_X1 U10306 ( .A1(n9065), .A2(n9399), .ZN(n9066) );
  OAI21_X1 U10307 ( .B1(n9065), .B2(n9399), .A(n9066), .ZN(n9076) );
  XNOR2_X1 U10308 ( .A(n9067), .B(n9050), .ZN(n9068) );
  NAND2_X1 U10309 ( .A1(n9193), .A2(n9181), .ZN(n9070) );
  AOI22_X1 U10310 ( .A1(n9372), .A2(n9171), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n9069) );
  OAI211_X1 U10311 ( .C1(n9174), .C2(n9178), .A(n9070), .B(n9069), .ZN(n9071)
         );
  AOI21_X1 U10312 ( .B1(n9072), .B2(n9190), .A(n9071), .ZN(n9073) );
  OAI21_X1 U10313 ( .B1(n9074), .B2(n9185), .A(n9073), .ZN(P2_U3160) );
  INV_X1 U10314 ( .A(n9601), .ZN(n9084) );
  AOI21_X1 U10315 ( .B1(n9075), .B2(n9076), .A(n9185), .ZN(n9078) );
  NAND2_X1 U10316 ( .A1(n9078), .A2(n9077), .ZN(n9083) );
  AOI22_X1 U10317 ( .A1(n9389), .A2(n9171), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n9079) );
  OAI21_X1 U10318 ( .B1(n9080), .B2(n9173), .A(n9079), .ZN(n9081) );
  AOI21_X1 U10319 ( .B1(n9152), .B2(n9381), .A(n9081), .ZN(n9082) );
  OAI211_X1 U10320 ( .C1(n9084), .C2(n9166), .A(n9083), .B(n9082), .ZN(
        P2_U3154) );
  XNOR2_X1 U10321 ( .A(n9085), .B(n9448), .ZN(n9091) );
  INV_X1 U10322 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9086) );
  OAI22_X1 U10323 ( .A1(n9460), .A2(n9178), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9086), .ZN(n9088) );
  NOR2_X1 U10324 ( .A1(n9437), .A2(n9173), .ZN(n9087) );
  AOI211_X1 U10325 ( .C1(n9441), .C2(n9171), .A(n9088), .B(n9087), .ZN(n9090)
         );
  NAND2_X1 U10326 ( .A1(n9440), .A2(n9190), .ZN(n9089) );
  OAI211_X1 U10327 ( .C1(n9091), .C2(n9185), .A(n9090), .B(n9089), .ZN(
        P2_U3156) );
  INV_X1 U10328 ( .A(n9092), .ZN(n9692) );
  OAI211_X1 U10329 ( .C1(n9095), .C2(n9094), .A(n9093), .B(n9148), .ZN(n9099)
         );
  NAND2_X1 U10330 ( .A1(n9195), .A2(n9181), .ZN(n9096) );
  NAND2_X1 U10331 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n9355) );
  OAI211_X1 U10332 ( .C1(n9487), .C2(n9178), .A(n9096), .B(n9355), .ZN(n9097)
         );
  AOI21_X1 U10333 ( .B1(n9491), .B2(n9171), .A(n9097), .ZN(n9098) );
  OAI211_X1 U10334 ( .C1(n9692), .C2(n9166), .A(n9099), .B(n9098), .ZN(
        P2_U3159) );
  XOR2_X1 U10335 ( .A(n9100), .B(n9101), .Z(n9107) );
  AOI22_X1 U10336 ( .A1(n9047), .A2(n9181), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n9103) );
  NAND2_X1 U10337 ( .A1(n9171), .A2(n9463), .ZN(n9102) );
  OAI211_X1 U10338 ( .C1(n9488), .C2(n9178), .A(n9103), .B(n9102), .ZN(n9104)
         );
  AOI21_X1 U10339 ( .B1(n9105), .B2(n9190), .A(n9104), .ZN(n9106) );
  OAI21_X1 U10340 ( .B1(n9107), .B2(n9185), .A(n9106), .ZN(P2_U3163) );
  XOR2_X1 U10341 ( .A(n9109), .B(n9108), .Z(n9114) );
  AOI22_X1 U10342 ( .A1(n9194), .A2(n9152), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n9111) );
  NAND2_X1 U10343 ( .A1(n9418), .A2(n9171), .ZN(n9110) );
  OAI211_X1 U10344 ( .C1(n9415), .C2(n9173), .A(n9111), .B(n9110), .ZN(n9112)
         );
  AOI21_X1 U10345 ( .B1(n9411), .B2(n9190), .A(n9112), .ZN(n9113) );
  OAI21_X1 U10346 ( .B1(n9114), .B2(n9185), .A(n9113), .ZN(P2_U3165) );
  XNOR2_X1 U10347 ( .A(n9115), .B(n9546), .ZN(n9116) );
  XNOR2_X1 U10348 ( .A(n9117), .B(n9116), .ZN(n9123) );
  INV_X1 U10349 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9118) );
  NOR2_X1 U10350 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9118), .ZN(n9284) );
  NOR2_X1 U10351 ( .A1(n9563), .A2(n9178), .ZN(n9119) );
  AOI211_X1 U10352 ( .C1(n9181), .C2(n9530), .A(n9284), .B(n9119), .ZN(n9120)
         );
  OAI21_X1 U10353 ( .B1(n9538), .B2(n9183), .A(n9120), .ZN(n9121) );
  AOI21_X1 U10354 ( .B1(n9537), .B2(n9190), .A(n9121), .ZN(n9122) );
  OAI21_X1 U10355 ( .B1(n9123), .B2(n9185), .A(n9122), .ZN(P2_U3166) );
  XNOR2_X1 U10356 ( .A(n9124), .B(n9530), .ZN(n9125) );
  XNOR2_X1 U10357 ( .A(n9126), .B(n9125), .ZN(n9131) );
  NAND2_X1 U10358 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9308) );
  OAI21_X1 U10359 ( .B1(n9173), .B2(n9487), .A(n9308), .ZN(n9127) );
  AOI21_X1 U10360 ( .B1(n9152), .B2(n9546), .A(n9127), .ZN(n9128) );
  OAI21_X1 U10361 ( .B1(n9522), .B2(n9183), .A(n9128), .ZN(n9129) );
  AOI21_X1 U10362 ( .B1(n9521), .B2(n9190), .A(n9129), .ZN(n9130) );
  OAI21_X1 U10363 ( .B1(n9131), .B2(n9185), .A(n9130), .ZN(P2_U3168) );
  XOR2_X1 U10364 ( .A(n9133), .B(n9132), .Z(n9138) );
  AOI22_X1 U10365 ( .A1(n9448), .A2(n9152), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n9135) );
  NAND2_X1 U10366 ( .A1(n9428), .A2(n9171), .ZN(n9134) );
  OAI211_X1 U10367 ( .C1(n9425), .C2(n9173), .A(n9135), .B(n9134), .ZN(n9136)
         );
  AOI21_X1 U10368 ( .B1(n9421), .B2(n9190), .A(n9136), .ZN(n9137) );
  OAI21_X1 U10369 ( .B1(n9138), .B2(n9185), .A(n9137), .ZN(P2_U3169) );
  INV_X1 U10370 ( .A(n9139), .ZN(n9140) );
  AOI21_X1 U10371 ( .B1(n9142), .B2(n9141), .A(n9140), .ZN(n9147) );
  AOI22_X1 U10372 ( .A1(n9447), .A2(n9181), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n9144) );
  NAND2_X1 U10373 ( .A1(n9171), .A2(n9475), .ZN(n9143) );
  OAI211_X1 U10374 ( .C1(n9504), .C2(n9178), .A(n9144), .B(n9143), .ZN(n9145)
         );
  AOI21_X1 U10375 ( .B1(n9474), .B2(n9190), .A(n9145), .ZN(n9146) );
  OAI21_X1 U10376 ( .B1(n9147), .B2(n9185), .A(n9146), .ZN(P2_U3173) );
  INV_X1 U10377 ( .A(n9622), .ZN(n9157) );
  OAI211_X1 U10378 ( .C1(n9151), .C2(n9150), .A(n9149), .B(n9148), .ZN(n9156)
         );
  AOI22_X1 U10379 ( .A1(n9447), .A2(n9152), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n9153) );
  OAI21_X1 U10380 ( .B1(n9426), .B2(n9173), .A(n9153), .ZN(n9154) );
  AOI21_X1 U10381 ( .B1(n9452), .B2(n9171), .A(n9154), .ZN(n9155) );
  OAI211_X1 U10382 ( .C1(n9157), .C2(n9166), .A(n9156), .B(n9155), .ZN(
        P2_U3175) );
  INV_X1 U10383 ( .A(n9510), .ZN(n9696) );
  AOI21_X1 U10384 ( .B1(n9159), .B2(n9158), .A(n9185), .ZN(n9161) );
  NAND2_X1 U10385 ( .A1(n9161), .A2(n9160), .ZN(n9165) );
  NAND2_X1 U10386 ( .A1(n9196), .A2(n9181), .ZN(n9162) );
  NAND2_X1 U10387 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9333) );
  OAI211_X1 U10388 ( .C1(n9503), .C2(n9178), .A(n9162), .B(n9333), .ZN(n9163)
         );
  AOI21_X1 U10389 ( .B1(n9505), .B2(n9171), .A(n9163), .ZN(n9164) );
  OAI211_X1 U10390 ( .C1(n9696), .C2(n9166), .A(n9165), .B(n9164), .ZN(
        P2_U3178) );
  XOR2_X1 U10391 ( .A(n9168), .B(n9167), .Z(n9177) );
  OAI22_X1 U10392 ( .A1(n9425), .A2(n9178), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9169), .ZN(n9170) );
  AOI21_X1 U10393 ( .B1(n9402), .B2(n9171), .A(n9170), .ZN(n9172) );
  OAI21_X1 U10394 ( .B1(n9174), .B2(n9173), .A(n9172), .ZN(n9175) );
  AOI21_X1 U10395 ( .B1(n9406), .B2(n9190), .A(n9175), .ZN(n9176) );
  OAI21_X1 U10396 ( .B1(n9177), .B2(n9185), .A(n9176), .ZN(P2_U3180) );
  NAND2_X1 U10397 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9259) );
  OAI21_X1 U10398 ( .B1(n9179), .B2(n9178), .A(n9259), .ZN(n9180) );
  AOI21_X1 U10399 ( .B1(n9181), .B2(n9546), .A(n9180), .ZN(n9182) );
  OAI21_X1 U10400 ( .B1(n9544), .B2(n9183), .A(n9182), .ZN(n9189) );
  AOI211_X1 U10401 ( .C1(n9187), .C2(n9186), .A(n9185), .B(n9184), .ZN(n9188)
         );
  AOI211_X1 U10402 ( .C1(n9553), .C2(n9190), .A(n9189), .B(n9188), .ZN(n9191)
         );
  INV_X1 U10403 ( .A(n9191), .ZN(P2_U3181) );
  MUX2_X1 U10404 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n9192), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10405 ( .A(n9193), .B(P2_DATAO_REG_29__SCAN_IN), .S(n9331), .Z(
        P2_U3520) );
  MUX2_X1 U10406 ( .A(n9380), .B(P2_DATAO_REG_28__SCAN_IN), .S(n9331), .Z(
        P2_U3519) );
  MUX2_X1 U10407 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n9399), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10408 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n9381), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10409 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n9398), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10410 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n9194), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10411 ( .A(n9448), .B(P2_DATAO_REG_23__SCAN_IN), .S(n9331), .Z(
        P2_U3514) );
  MUX2_X1 U10412 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9047), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10413 ( .A(n9447), .B(P2_DATAO_REG_21__SCAN_IN), .S(n9331), .Z(
        P2_U3512) );
  MUX2_X1 U10414 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n9195), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10415 ( .A(n9196), .B(P2_DATAO_REG_19__SCAN_IN), .S(n9331), .Z(
        P2_U3510) );
  MUX2_X1 U10416 ( .A(n9516), .B(P2_DATAO_REG_18__SCAN_IN), .S(n9331), .Z(
        P2_U3509) );
  MUX2_X1 U10417 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9530), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10418 ( .A(n9546), .B(P2_DATAO_REG_16__SCAN_IN), .S(n9331), .Z(
        P2_U3507) );
  MUX2_X1 U10419 ( .A(n9529), .B(P2_DATAO_REG_15__SCAN_IN), .S(n9331), .Z(
        P2_U3506) );
  MUX2_X1 U10420 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n9577), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U10421 ( .A(n9197), .B(P2_DATAO_REG_13__SCAN_IN), .S(n9331), .Z(
        P2_U3504) );
  MUX2_X1 U10422 ( .A(n9578), .B(P2_DATAO_REG_12__SCAN_IN), .S(n9331), .Z(
        P2_U3503) );
  MUX2_X1 U10423 ( .A(n9198), .B(P2_DATAO_REG_11__SCAN_IN), .S(n9331), .Z(
        P2_U3502) );
  MUX2_X1 U10424 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n9199), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U10425 ( .A(n9200), .B(P2_DATAO_REG_9__SCAN_IN), .S(n9331), .Z(
        P2_U3500) );
  MUX2_X1 U10426 ( .A(n9201), .B(P2_DATAO_REG_8__SCAN_IN), .S(n9331), .Z(
        P2_U3499) );
  MUX2_X1 U10427 ( .A(n9202), .B(P2_DATAO_REG_7__SCAN_IN), .S(n9331), .Z(
        P2_U3498) );
  MUX2_X1 U10428 ( .A(n9203), .B(P2_DATAO_REG_6__SCAN_IN), .S(n9331), .Z(
        P2_U3497) );
  MUX2_X1 U10429 ( .A(n7171), .B(P2_DATAO_REG_5__SCAN_IN), .S(n9331), .Z(
        P2_U3496) );
  MUX2_X1 U10430 ( .A(n9204), .B(P2_DATAO_REG_3__SCAN_IN), .S(n9331), .Z(
        P2_U3494) );
  MUX2_X1 U10431 ( .A(n10925), .B(P2_DATAO_REG_2__SCAN_IN), .S(n9331), .Z(
        P2_U3493) );
  MUX2_X1 U10432 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n6953), .S(P2_U3893), .Z(
        P2_U3492) );
  MUX2_X1 U10433 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n6912), .S(P2_U3893), .Z(
        P2_U3491) );
  NAND2_X1 U10434 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n9207), .ZN(n9243) );
  OAI21_X1 U10435 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n9207), .A(n9243), .ZN(
        n9223) );
  AOI21_X1 U10436 ( .B1(n9209), .B2(n6477), .A(n9228), .ZN(n9211) );
  OAI21_X1 U10437 ( .B1(n10854), .B2(n9211), .A(n9210), .ZN(n9212) );
  AOI21_X1 U10438 ( .B1(n10858), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n9212), .ZN(
        n9221) );
  MUX2_X1 U10439 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n9327), .Z(n9231) );
  XNOR2_X1 U10440 ( .A(n9231), .B(n9226), .ZN(n9218) );
  OR2_X1 U10441 ( .A1(n9214), .A2(n9213), .ZN(n9216) );
  NAND2_X1 U10442 ( .A1(n9218), .A2(n9217), .ZN(n9232) );
  OAI21_X1 U10443 ( .B1(n9218), .B2(n9217), .A(n9232), .ZN(n9219) );
  NAND2_X1 U10444 ( .A1(n9219), .A2(n10859), .ZN(n9220) );
  OAI211_X1 U10445 ( .C1(n9330), .C2(n9242), .A(n9221), .B(n9220), .ZN(n9222)
         );
  AOI21_X1 U10446 ( .B1(n9223), .B2(n10849), .A(n9222), .ZN(n9224) );
  INV_X1 U10447 ( .A(n9224), .ZN(P2_U3195) );
  NOR2_X1 U10448 ( .A1(n9226), .A2(n9225), .ZN(n9227) );
  NAND2_X1 U10449 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n9264), .ZN(n9229) );
  OAI21_X1 U10450 ( .B1(n9264), .B2(P2_REG2_REG_14__SCAN_IN), .A(n9229), .ZN(
        n9230) );
  AOI21_X1 U10451 ( .B1(n5173), .B2(n9230), .A(n9255), .ZN(n9250) );
  MUX2_X1 U10452 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n9327), .Z(n9265) );
  XNOR2_X1 U10453 ( .A(n9265), .B(n9240), .ZN(n9235) );
  OR2_X1 U10454 ( .A1(n9231), .A2(n9242), .ZN(n9233) );
  NAND2_X1 U10455 ( .A1(n9233), .A2(n9232), .ZN(n9234) );
  OAI21_X1 U10456 ( .B1(n9235), .B2(n9234), .A(n9266), .ZN(n9239) );
  NAND2_X1 U10457 ( .A1(n10858), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n9237) );
  OAI211_X1 U10458 ( .C1(n9330), .C2(n9264), .A(n9237), .B(n9236), .ZN(n9238)
         );
  AOI21_X1 U10459 ( .B1(n10859), .B2(n9239), .A(n9238), .ZN(n9249) );
  AOI22_X1 U10460 ( .A1(n9240), .A2(n6491), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n9264), .ZN(n9246) );
  NAND2_X1 U10461 ( .A1(n9242), .A2(n9241), .ZN(n9244) );
  NAND2_X1 U10462 ( .A1(n9244), .A2(n9243), .ZN(n9245) );
  NAND2_X1 U10463 ( .A1(n9246), .A2(n9245), .ZN(n9251) );
  OAI21_X1 U10464 ( .B1(n9246), .B2(n9245), .A(n9251), .ZN(n9247) );
  NAND2_X1 U10465 ( .A1(n9247), .A2(n10849), .ZN(n9248) );
  OAI211_X1 U10466 ( .C1(n9250), .C2(n10854), .A(n9249), .B(n9248), .ZN(
        P2_U3196) );
  NAND2_X1 U10467 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n9264), .ZN(n9252) );
  NAND2_X1 U10468 ( .A1(n9252), .A2(n9251), .ZN(n9278) );
  XNOR2_X1 U10469 ( .A(n9278), .B(n9263), .ZN(n9253) );
  NAND2_X1 U10470 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n9253), .ZN(n9279) );
  OAI21_X1 U10471 ( .B1(n9253), .B2(P2_REG1_REG_15__SCAN_IN), .A(n9279), .ZN(
        n9254) );
  NAND2_X1 U10472 ( .A1(n9254), .A2(n10849), .ZN(n9273) );
  NAND2_X1 U10473 ( .A1(n9256), .A2(n9263), .ZN(n9257) );
  AOI21_X1 U10474 ( .B1(n9258), .B2(n9554), .A(n9275), .ZN(n9261) );
  NAND2_X1 U10475 ( .A1(n10858), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n9260) );
  OAI211_X1 U10476 ( .C1(n9261), .C2(n10854), .A(n9260), .B(n9259), .ZN(n9262)
         );
  AOI21_X1 U10477 ( .B1(n9263), .B2(n10848), .A(n9262), .ZN(n9272) );
  MUX2_X1 U10478 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n9327), .Z(n9286) );
  XNOR2_X1 U10479 ( .A(n9286), .B(n9263), .ZN(n9269) );
  OR2_X1 U10480 ( .A1(n9265), .A2(n9264), .ZN(n9267) );
  OAI21_X1 U10481 ( .B1(n9269), .B2(n9268), .A(n9287), .ZN(n9270) );
  NAND2_X1 U10482 ( .A1(n9270), .A2(n10859), .ZN(n9271) );
  NAND3_X1 U10483 ( .A1(n9273), .A2(n9272), .A3(n9271), .ZN(P2_U3197) );
  AOI22_X1 U10484 ( .A1(n9313), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n9539), .B2(
        n9301), .ZN(n9277) );
  AOI21_X1 U10485 ( .B1(n5169), .B2(n9277), .A(n9298), .ZN(n9297) );
  AOI22_X1 U10486 ( .A1(n9313), .A2(n9649), .B1(P2_REG1_REG_16__SCAN_IN), .B2(
        n9301), .ZN(n9282) );
  NAND2_X1 U10487 ( .A1(n9278), .A2(n9285), .ZN(n9280) );
  NAND2_X1 U10488 ( .A1(n9280), .A2(n9279), .ZN(n9281) );
  OAI21_X1 U10489 ( .B1(n9282), .B2(n9281), .A(n9312), .ZN(n9295) );
  NOR2_X1 U10490 ( .A1(n9330), .A2(n9301), .ZN(n9283) );
  AOI211_X1 U10491 ( .C1(n10858), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n9284), .B(
        n9283), .ZN(n9293) );
  MUX2_X1 U10492 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n9327), .Z(n9302) );
  XNOR2_X1 U10493 ( .A(n9302), .B(n9313), .ZN(n9290) );
  OR2_X1 U10494 ( .A1(n9286), .A2(n9285), .ZN(n9288) );
  NAND2_X1 U10495 ( .A1(n9290), .A2(n9289), .ZN(n9303) );
  OAI21_X1 U10496 ( .B1(n9290), .B2(n9289), .A(n9303), .ZN(n9291) );
  NAND2_X1 U10497 ( .A1(n9291), .A2(n10859), .ZN(n9292) );
  NAND2_X1 U10498 ( .A1(n9293), .A2(n9292), .ZN(n9294) );
  AOI21_X1 U10499 ( .B1(n9295), .B2(n10849), .A(n9294), .ZN(n9296) );
  OAI21_X1 U10500 ( .B1(n9297), .B2(n10854), .A(n9296), .ZN(P2_U3198) );
  INV_X1 U10501 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9300) );
  AOI21_X1 U10502 ( .B1(n9300), .B2(n9299), .A(n9322), .ZN(n9318) );
  MUX2_X1 U10503 ( .A(n9300), .B(n9645), .S(n9327), .Z(n9326) );
  XNOR2_X1 U10504 ( .A(n9326), .B(n9337), .ZN(n9306) );
  OR2_X1 U10505 ( .A1(n9302), .A2(n9301), .ZN(n9304) );
  NAND2_X1 U10506 ( .A1(n9304), .A2(n9303), .ZN(n9305) );
  NAND2_X1 U10507 ( .A1(n9306), .A2(n9305), .ZN(n9324) );
  OAI21_X1 U10508 ( .B1(n9306), .B2(n9305), .A(n9324), .ZN(n9311) );
  INV_X1 U10509 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n9309) );
  OR2_X1 U10510 ( .A1(n9330), .A2(n9337), .ZN(n9307) );
  OAI211_X1 U10511 ( .C1(n10843), .C2(n9309), .A(n9308), .B(n9307), .ZN(n9310)
         );
  AOI21_X1 U10512 ( .B1(n10859), .B2(n9311), .A(n9310), .ZN(n9317) );
  OAI21_X1 U10513 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n9314), .A(n9338), .ZN(
        n9315) );
  NAND2_X1 U10514 ( .A1(n9315), .A2(n10849), .ZN(n9316) );
  OAI211_X1 U10515 ( .C1(n9318), .C2(n10854), .A(n9317), .B(n9316), .ZN(
        P2_U3199) );
  NOR2_X1 U10516 ( .A1(n9356), .A2(n9507), .ZN(n9319) );
  AOI21_X1 U10517 ( .B1(n9356), .B2(n9507), .A(n9319), .ZN(n9323) );
  NOR2_X1 U10518 ( .A1(n9325), .A2(n9320), .ZN(n9321) );
  AOI21_X1 U10519 ( .B1(n9323), .B2(n5138), .A(n9346), .ZN(n9345) );
  MUX2_X1 U10520 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n9327), .Z(n9328) );
  NAND2_X1 U10521 ( .A1(n9329), .A2(n9328), .ZN(n9348) );
  OAI21_X1 U10522 ( .B1(n9332), .B2(n9331), .A(n9330), .ZN(n9343) );
  INV_X1 U10523 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n9335) );
  NAND3_X1 U10524 ( .A1(n9332), .A2(n10859), .A3(n9356), .ZN(n9334) );
  OAI211_X1 U10525 ( .C1(n10843), .C2(n9335), .A(n9334), .B(n9333), .ZN(n9342)
         );
  XNOR2_X1 U10526 ( .A(n9349), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n9357) );
  NAND2_X1 U10527 ( .A1(n9337), .A2(n9336), .ZN(n9339) );
  NAND2_X1 U10528 ( .A1(n9339), .A2(n9338), .ZN(n9358) );
  XOR2_X1 U10529 ( .A(n9357), .B(n9358), .Z(n9340) );
  NOR2_X1 U10530 ( .A1(n9340), .A2(n10833), .ZN(n9341) );
  AOI211_X1 U10531 ( .C1(n9349), .C2(n9343), .A(n9342), .B(n9341), .ZN(n9344)
         );
  OAI21_X1 U10532 ( .B1(n9345), .B2(n10854), .A(n9344), .ZN(P2_U3200) );
  MUX2_X1 U10533 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n6560), .S(n6711), .Z(n9351) );
  AOI21_X1 U10534 ( .B1(n9349), .B2(n9348), .A(n9347), .ZN(n9353) );
  XNOR2_X1 U10535 ( .A(n6711), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n9359) );
  INV_X1 U10536 ( .A(n9359), .ZN(n9350) );
  MUX2_X1 U10537 ( .A(n9351), .B(n9350), .S(n9327), .Z(n9352) );
  XNOR2_X1 U10538 ( .A(n9353), .B(n9352), .ZN(n9362) );
  NAND2_X1 U10539 ( .A1(n10848), .A2(n6711), .ZN(n9354) );
  OAI211_X1 U10540 ( .C1(n10843), .C2(n5371), .A(n9355), .B(n9354), .ZN(n9361)
         );
  AOI22_X1 U10541 ( .A1(n9358), .A2(n9357), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n9356), .ZN(n9360) );
  INV_X1 U10542 ( .A(n9363), .ZN(n9364) );
  NOR2_X1 U10543 ( .A1(n9365), .A2(n9364), .ZN(n9656) );
  INV_X1 U10544 ( .A(n9656), .ZN(n9367) );
  NAND3_X1 U10545 ( .A1(n9367), .A2(n10944), .A3(n9366), .ZN(n9369) );
  OAI21_X1 U10546 ( .B1(P2_REG2_REG_31__SCAN_IN), .B2(n10944), .A(n9369), .ZN(
        n9368) );
  OAI21_X1 U10547 ( .B1(n9658), .B2(n10939), .A(n9368), .ZN(P2_U3202) );
  OAI21_X1 U10548 ( .B1(P2_REG2_REG_30__SCAN_IN), .B2(n10944), .A(n9369), .ZN(
        n9370) );
  OAI21_X1 U10549 ( .B1(n9661), .B2(n10939), .A(n9370), .ZN(P2_U3203) );
  INV_X1 U10550 ( .A(n9371), .ZN(n9378) );
  AOI22_X1 U10551 ( .A1(n9372), .A2(n9550), .B1(n10946), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n9373) );
  OAI21_X1 U10552 ( .B1(n9374), .B2(n10939), .A(n9373), .ZN(n9375) );
  AOI21_X1 U10553 ( .B1(n9376), .B2(n10941), .A(n9375), .ZN(n9377) );
  OAI21_X1 U10554 ( .B1(n9378), .B2(n10946), .A(n9377), .ZN(P2_U3205) );
  XNOR2_X1 U10555 ( .A(n9379), .B(n9387), .ZN(n9385) );
  OAI21_X1 U10556 ( .B1(n9388), .B2(n9387), .A(n9386), .ZN(n9604) );
  AOI22_X1 U10557 ( .A1(n9389), .A2(n9550), .B1(n10946), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n9391) );
  NAND2_X1 U10558 ( .A1(n9601), .A2(n9509), .ZN(n9390) );
  OAI211_X1 U10559 ( .C1(n9604), .C2(n9513), .A(n9391), .B(n9390), .ZN(n9392)
         );
  INV_X1 U10560 ( .A(n9392), .ZN(n9393) );
  OAI21_X1 U10561 ( .B1(n9603), .B2(n10946), .A(n9393), .ZN(P2_U3206) );
  OAI21_X1 U10562 ( .B1(n5164), .B2(n9395), .A(n9394), .ZN(n9605) );
  XNOR2_X1 U10563 ( .A(n9396), .B(n9395), .ZN(n9397) );
  NAND2_X1 U10564 ( .A1(n9397), .A2(n10928), .ZN(n9401) );
  AOI22_X1 U10565 ( .A1(n9399), .A2(n10926), .B1(n6677), .B2(n9398), .ZN(n9400) );
  NAND2_X1 U10566 ( .A1(n9401), .A2(n9400), .ZN(n9607) );
  NAND2_X1 U10567 ( .A1(n9607), .A2(n10944), .ZN(n9408) );
  INV_X1 U10568 ( .A(n9402), .ZN(n9404) );
  OAI22_X1 U10569 ( .A1(n9404), .A2(n10937), .B1(n9403), .B2(n10944), .ZN(
        n9405) );
  AOI21_X1 U10570 ( .B1(n9406), .B2(n9509), .A(n9405), .ZN(n9407) );
  OAI211_X1 U10571 ( .C1(n9513), .C2(n9605), .A(n9408), .B(n9407), .ZN(
        P2_U3207) );
  XNOR2_X1 U10572 ( .A(n9410), .B(n9409), .ZN(n9611) );
  INV_X1 U10573 ( .A(n9411), .ZN(n9671) );
  NOR2_X1 U10574 ( .A1(n9671), .A2(n9583), .ZN(n9416) );
  XNOR2_X1 U10575 ( .A(n9413), .B(n9412), .ZN(n9414) );
  OAI222_X1 U10576 ( .A1(n9562), .A2(n9437), .B1(n9564), .B2(n9415), .C1(n9559), .C2(n9414), .ZN(n9610) );
  AOI211_X1 U10577 ( .C1(n9417), .C2(n9611), .A(n9416), .B(n9610), .ZN(n9420)
         );
  AOI22_X1 U10578 ( .A1(n9418), .A2(n9550), .B1(n10946), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n9419) );
  OAI21_X1 U10579 ( .B1(n9420), .B2(n10946), .A(n9419), .ZN(P2_U3208) );
  INV_X1 U10580 ( .A(n9421), .ZN(n9675) );
  NOR2_X1 U10581 ( .A1(n9675), .A2(n9583), .ZN(n9427) );
  XNOR2_X1 U10582 ( .A(n9423), .B(n9422), .ZN(n9424) );
  OAI222_X1 U10583 ( .A1(n9562), .A2(n9426), .B1(n9564), .B2(n9425), .C1(n9559), .C2(n9424), .ZN(n9614) );
  AOI211_X1 U10584 ( .C1(n9550), .C2(n9428), .A(n9427), .B(n9614), .ZN(n9433)
         );
  NAND2_X1 U10585 ( .A1(n9430), .A2(n9429), .ZN(n9431) );
  XNOR2_X1 U10586 ( .A(n9431), .B(n6708), .ZN(n9615) );
  AOI22_X1 U10587 ( .A1(n9615), .A2(n10941), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n10946), .ZN(n9432) );
  OAI21_X1 U10588 ( .B1(n9433), .B2(n10946), .A(n9432), .ZN(P2_U3209) );
  XNOR2_X1 U10589 ( .A(n9435), .B(n9434), .ZN(n9436) );
  OAI222_X1 U10590 ( .A1(n9562), .A2(n9460), .B1(n9564), .B2(n9437), .C1(n9559), .C2(n9436), .ZN(n9618) );
  INV_X1 U10591 ( .A(n9618), .ZN(n9445) );
  XNOR2_X1 U10592 ( .A(n9439), .B(n9438), .ZN(n9619) );
  INV_X1 U10593 ( .A(n9440), .ZN(n9679) );
  AOI22_X1 U10594 ( .A1(n9441), .A2(n9550), .B1(n10946), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n9442) );
  OAI21_X1 U10595 ( .B1(n9679), .B2(n10939), .A(n9442), .ZN(n9443) );
  AOI21_X1 U10596 ( .B1(n9619), .B2(n10941), .A(n9443), .ZN(n9444) );
  OAI21_X1 U10597 ( .B1(n9445), .B2(n10946), .A(n9444), .ZN(P2_U3210) );
  XNOR2_X1 U10598 ( .A(n9446), .B(n9451), .ZN(n9449) );
  AOI222_X1 U10599 ( .A1(n10928), .A2(n9449), .B1(n9448), .B2(n10926), .C1(
        n9447), .C2(n6677), .ZN(n9625) );
  XNOR2_X1 U10600 ( .A(n9450), .B(n9451), .ZN(n9623) );
  NAND2_X1 U10601 ( .A1(n9622), .A2(n9509), .ZN(n9454) );
  AOI22_X1 U10602 ( .A1(n10946), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9452), 
        .B2(n9550), .ZN(n9453) );
  NAND2_X1 U10603 ( .A1(n9454), .A2(n9453), .ZN(n9455) );
  AOI21_X1 U10604 ( .B1(n9623), .B2(n10941), .A(n9455), .ZN(n9456) );
  OAI21_X1 U10605 ( .B1(n9625), .B2(n10946), .A(n9456), .ZN(P2_U3211) );
  XNOR2_X1 U10606 ( .A(n9458), .B(n9457), .ZN(n9459) );
  OAI222_X1 U10607 ( .A1(n9564), .A2(n9460), .B1(n9562), .B2(n9488), .C1(n9459), .C2(n9559), .ZN(n9626) );
  INV_X1 U10608 ( .A(n9626), .ZN(n9467) );
  XNOR2_X1 U10609 ( .A(n9461), .B(n9462), .ZN(n9627) );
  AOI22_X1 U10610 ( .A1(n10946), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n9550), 
        .B2(n9463), .ZN(n9464) );
  OAI21_X1 U10611 ( .B1(n9684), .B2(n10939), .A(n9464), .ZN(n9465) );
  AOI21_X1 U10612 ( .B1(n9627), .B2(n10941), .A(n9465), .ZN(n9466) );
  OAI21_X1 U10613 ( .B1(n9467), .B2(n10946), .A(n9466), .ZN(P2_U3212) );
  XNOR2_X1 U10614 ( .A(n9468), .B(n9469), .ZN(n9470) );
  OAI222_X1 U10615 ( .A1(n9562), .A2(n9504), .B1(n9564), .B2(n9471), .C1(n9470), .C2(n9559), .ZN(n9630) );
  INV_X1 U10616 ( .A(n9630), .ZN(n9479) );
  XNOR2_X1 U10617 ( .A(n9472), .B(n9473), .ZN(n9631) );
  INV_X1 U10618 ( .A(n9474), .ZN(n9688) );
  AOI22_X1 U10619 ( .A1(n10946), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9475), 
        .B2(n9550), .ZN(n9476) );
  OAI21_X1 U10620 ( .B1(n9688), .B2(n10939), .A(n9476), .ZN(n9477) );
  AOI21_X1 U10621 ( .B1(n9631), .B2(n10941), .A(n9477), .ZN(n9478) );
  OAI21_X1 U10622 ( .B1(n9479), .B2(n10946), .A(n9478), .ZN(P2_U3213) );
  NAND2_X1 U10623 ( .A1(n9528), .A2(n9482), .ZN(n9484) );
  NAND2_X1 U10624 ( .A1(n9484), .A2(n9483), .ZN(n9485) );
  XNOR2_X1 U10625 ( .A(n9485), .B(n9489), .ZN(n9486) );
  OAI222_X1 U10626 ( .A1(n9564), .A2(n9488), .B1(n9562), .B2(n9487), .C1(n9559), .C2(n9486), .ZN(n9634) );
  INV_X1 U10627 ( .A(n9634), .ZN(n9495) );
  XNOR2_X1 U10628 ( .A(n9490), .B(n9489), .ZN(n9635) );
  AOI22_X1 U10629 ( .A1(n10946), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n9550), 
        .B2(n9491), .ZN(n9492) );
  OAI21_X1 U10630 ( .B1(n9692), .B2(n10939), .A(n9492), .ZN(n9493) );
  AOI21_X1 U10631 ( .B1(n9635), .B2(n10941), .A(n9493), .ZN(n9494) );
  OAI21_X1 U10632 ( .B1(n9495), .B2(n10946), .A(n9494), .ZN(P2_U3214) );
  OAI21_X1 U10633 ( .B1(n9497), .B2(n9501), .A(n9496), .ZN(n9638) );
  NAND2_X1 U10634 ( .A1(n9528), .A2(n9536), .ZN(n9527) );
  NAND2_X1 U10635 ( .A1(n9527), .A2(n9498), .ZN(n9515) );
  NAND2_X1 U10636 ( .A1(n9515), .A2(n9519), .ZN(n9514) );
  NAND2_X1 U10637 ( .A1(n9514), .A2(n9499), .ZN(n9500) );
  XOR2_X1 U10638 ( .A(n9501), .B(n9500), .Z(n9502) );
  OAI222_X1 U10639 ( .A1(n9564), .A2(n9504), .B1(n9562), .B2(n9503), .C1(n9502), .C2(n9559), .ZN(n9639) );
  NAND2_X1 U10640 ( .A1(n9639), .A2(n10944), .ZN(n9512) );
  INV_X1 U10641 ( .A(n9505), .ZN(n9506) );
  OAI22_X1 U10642 ( .A1(n9589), .A2(n9507), .B1(n9506), .B2(n10937), .ZN(n9508) );
  AOI21_X1 U10643 ( .B1(n9510), .B2(n9509), .A(n9508), .ZN(n9511) );
  OAI211_X1 U10644 ( .C1(n9638), .C2(n9513), .A(n9512), .B(n9511), .ZN(
        P2_U3215) );
  OAI211_X1 U10645 ( .C1(n9515), .C2(n9519), .A(n9514), .B(n10928), .ZN(n9518)
         );
  AOI22_X1 U10646 ( .A1(n6677), .A2(n9546), .B1(n9516), .B2(n10926), .ZN(n9517) );
  NAND2_X1 U10647 ( .A1(n9518), .A2(n9517), .ZN(n9643) );
  INV_X1 U10648 ( .A(n9643), .ZN(n9526) );
  XNOR2_X1 U10649 ( .A(n9520), .B(n9519), .ZN(n9644) );
  INV_X1 U10650 ( .A(n9521), .ZN(n9700) );
  NOR2_X1 U10651 ( .A1(n9700), .A2(n10939), .ZN(n9524) );
  OAI22_X1 U10652 ( .A1(n9589), .A2(n9300), .B1(n9522), .B2(n10937), .ZN(n9523) );
  AOI211_X1 U10653 ( .C1(n9644), .C2(n10941), .A(n9524), .B(n9523), .ZN(n9525)
         );
  OAI21_X1 U10654 ( .B1(n9526), .B2(n10946), .A(n9525), .ZN(P2_U3216) );
  OAI211_X1 U10655 ( .C1(n9528), .C2(n9536), .A(n9527), .B(n10928), .ZN(n9532)
         );
  AOI22_X1 U10656 ( .A1(n9530), .A2(n10926), .B1(n6677), .B2(n9529), .ZN(n9531) );
  NAND2_X1 U10657 ( .A1(n9532), .A2(n9531), .ZN(n9647) );
  INV_X1 U10658 ( .A(n9647), .ZN(n9543) );
  INV_X1 U10659 ( .A(n9533), .ZN(n9534) );
  AOI21_X1 U10660 ( .B1(n9536), .B2(n9535), .A(n9534), .ZN(n9648) );
  INV_X1 U10661 ( .A(n9537), .ZN(n9704) );
  NOR2_X1 U10662 ( .A1(n9704), .A2(n10939), .ZN(n9541) );
  OAI22_X1 U10663 ( .A1(n9589), .A2(n9539), .B1(n9538), .B2(n10937), .ZN(n9540) );
  AOI211_X1 U10664 ( .C1(n9648), .C2(n10941), .A(n9541), .B(n9540), .ZN(n9542)
         );
  OAI21_X1 U10665 ( .B1(n9543), .B2(n10946), .A(n9542), .ZN(P2_U3217) );
  INV_X1 U10666 ( .A(n9544), .ZN(n9549) );
  OAI211_X1 U10667 ( .C1(n9545), .C2(n9551), .A(n9480), .B(n10928), .ZN(n9548)
         );
  AOI22_X1 U10668 ( .A1(n6677), .A2(n9577), .B1(n9546), .B2(n10926), .ZN(n9547) );
  NAND2_X1 U10669 ( .A1(n9548), .A2(n9547), .ZN(n9651) );
  AOI21_X1 U10670 ( .B1(n9550), .B2(n9549), .A(n9651), .ZN(n9557) );
  XNOR2_X1 U10671 ( .A(n9552), .B(n9551), .ZN(n9652) );
  INV_X1 U10672 ( .A(n9553), .ZN(n9709) );
  OAI22_X1 U10673 ( .A1(n9709), .A2(n10939), .B1(n9554), .B2(n9589), .ZN(n9555) );
  AOI21_X1 U10674 ( .B1(n9652), .B2(n10941), .A(n9555), .ZN(n9556) );
  OAI21_X1 U10675 ( .B1(n9557), .B2(n10946), .A(n9556), .ZN(P2_U3218) );
  XNOR2_X1 U10676 ( .A(n9558), .B(n6699), .ZN(n9560) );
  OAI222_X1 U10677 ( .A1(n9564), .A2(n9563), .B1(n9562), .B2(n9561), .C1(n9560), .C2(n9559), .ZN(n11095) );
  OAI22_X1 U10678 ( .A1(n11094), .A2(n9583), .B1(n9565), .B2(n10937), .ZN(
        n9566) );
  OAI21_X1 U10679 ( .B1(n11095), .B2(n9566), .A(n9589), .ZN(n9572) );
  INV_X1 U10680 ( .A(n9567), .ZN(n9568) );
  AOI21_X1 U10681 ( .B1(n9570), .B2(n9569), .A(n9568), .ZN(n11098) );
  NAND2_X1 U10682 ( .A1(n11098), .A2(n10941), .ZN(n9571) );
  OAI211_X1 U10683 ( .C1(n6494), .C2(n9589), .A(n9572), .B(n9571), .ZN(
        P2_U3219) );
  NAND2_X1 U10684 ( .A1(n9574), .A2(n9585), .ZN(n9575) );
  NAND2_X1 U10685 ( .A1(n9573), .A2(n9575), .ZN(n9576) );
  NAND2_X1 U10686 ( .A1(n9576), .A2(n10928), .ZN(n9580) );
  AOI22_X1 U10687 ( .A1(n6677), .A2(n9578), .B1(n9577), .B2(n10926), .ZN(n9579) );
  NAND2_X1 U10688 ( .A1(n9580), .A2(n9579), .ZN(n11090) );
  INV_X1 U10689 ( .A(n9581), .ZN(n11088) );
  OAI22_X1 U10690 ( .A1(n11088), .A2(n9583), .B1(n9582), .B2(n10937), .ZN(
        n9584) );
  OAI21_X1 U10691 ( .B1(n11090), .B2(n9584), .A(n9589), .ZN(n9588) );
  XNOR2_X1 U10692 ( .A(n9586), .B(n9585), .ZN(n11086) );
  NAND2_X1 U10693 ( .A1(n11086), .A2(n10941), .ZN(n9587) );
  OAI211_X1 U10694 ( .C1(n6477), .C2(n9589), .A(n9588), .B(n9587), .ZN(
        P2_U3220) );
  NAND2_X1 U10695 ( .A1(n9656), .A2(n11100), .ZN(n9591) );
  NAND2_X1 U10696 ( .A1(n11099), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n9590) );
  OAI211_X1 U10697 ( .C1(n9658), .C2(n9655), .A(n9591), .B(n9590), .ZN(
        P2_U3490) );
  NAND2_X1 U10698 ( .A1(n11099), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n9592) );
  OAI211_X1 U10699 ( .C1(n9661), .C2(n9655), .A(n9592), .B(n9591), .ZN(
        P2_U3489) );
  INV_X1 U10700 ( .A(n9593), .ZN(n9595) );
  NAND2_X1 U10701 ( .A1(n9595), .A2(n9594), .ZN(n9598) );
  NAND2_X1 U10702 ( .A1(n9600), .A2(n9599), .ZN(n9662) );
  MUX2_X1 U10703 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9662), .S(n11100), .Z(
        P2_U3488) );
  INV_X1 U10704 ( .A(n11097), .ZN(n11012) );
  NAND2_X1 U10705 ( .A1(n9601), .A2(n11017), .ZN(n9602) );
  OAI211_X1 U10706 ( .C1(n11012), .C2(n9604), .A(n9603), .B(n9602), .ZN(n9663)
         );
  MUX2_X1 U10707 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9663), .S(n11100), .Z(
        P2_U3486) );
  NOR2_X1 U10708 ( .A1(n9605), .A2(n11012), .ZN(n9606) );
  MUX2_X1 U10709 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9664), .S(n11100), .Z(
        n9608) );
  INV_X1 U10710 ( .A(n9608), .ZN(n9609) );
  OAI21_X1 U10711 ( .B1(n9667), .B2(n9655), .A(n9609), .ZN(P2_U3485) );
  INV_X1 U10712 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9612) );
  AOI21_X1 U10713 ( .B1(n11097), .B2(n9611), .A(n9610), .ZN(n9668) );
  MUX2_X1 U10714 ( .A(n9612), .B(n9668), .S(n11100), .Z(n9613) );
  OAI21_X1 U10715 ( .B1(n9671), .B2(n9655), .A(n9613), .ZN(P2_U3484) );
  INV_X1 U10716 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9616) );
  AOI21_X1 U10717 ( .B1(n11097), .B2(n9615), .A(n9614), .ZN(n9672) );
  MUX2_X1 U10718 ( .A(n9616), .B(n9672), .S(n11100), .Z(n9617) );
  OAI21_X1 U10719 ( .B1(n9675), .B2(n9655), .A(n9617), .ZN(P2_U3483) );
  INV_X1 U10720 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9620) );
  AOI21_X1 U10721 ( .B1(n11097), .B2(n9619), .A(n9618), .ZN(n9676) );
  MUX2_X1 U10722 ( .A(n9620), .B(n9676), .S(n11100), .Z(n9621) );
  OAI21_X1 U10723 ( .B1(n9679), .B2(n9655), .A(n9621), .ZN(P2_U3482) );
  AOI22_X1 U10724 ( .A1(n9623), .A2(n11097), .B1(n11017), .B2(n9622), .ZN(
        n9624) );
  NAND2_X1 U10725 ( .A1(n9625), .A2(n9624), .ZN(n9680) );
  MUX2_X1 U10726 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9680), .S(n11100), .Z(
        P2_U3481) );
  INV_X1 U10727 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9628) );
  AOI21_X1 U10728 ( .B1(n9627), .B2(n11097), .A(n9626), .ZN(n9681) );
  MUX2_X1 U10729 ( .A(n9628), .B(n9681), .S(n11100), .Z(n9629) );
  OAI21_X1 U10730 ( .B1(n9684), .B2(n9655), .A(n9629), .ZN(P2_U3480) );
  INV_X1 U10731 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9632) );
  AOI21_X1 U10732 ( .B1(n9631), .B2(n11097), .A(n9630), .ZN(n9685) );
  MUX2_X1 U10733 ( .A(n9632), .B(n9685), .S(n11100), .Z(n9633) );
  OAI21_X1 U10734 ( .B1(n9688), .B2(n9655), .A(n9633), .ZN(P2_U3479) );
  INV_X1 U10735 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9636) );
  AOI21_X1 U10736 ( .B1(n9635), .B2(n11097), .A(n9634), .ZN(n9689) );
  MUX2_X1 U10737 ( .A(n9636), .B(n9689), .S(n11100), .Z(n9637) );
  OAI21_X1 U10738 ( .B1(n9692), .B2(n9655), .A(n9637), .ZN(P2_U3478) );
  INV_X1 U10739 ( .A(n9638), .ZN(n9640) );
  AOI21_X1 U10740 ( .B1(n9640), .B2(n11097), .A(n9639), .ZN(n9693) );
  MUX2_X1 U10741 ( .A(n9641), .B(n9693), .S(n11100), .Z(n9642) );
  OAI21_X1 U10742 ( .B1(n9696), .B2(n9655), .A(n9642), .ZN(P2_U3477) );
  AOI21_X1 U10743 ( .B1(n9644), .B2(n11097), .A(n9643), .ZN(n9697) );
  MUX2_X1 U10744 ( .A(n9645), .B(n9697), .S(n11100), .Z(n9646) );
  OAI21_X1 U10745 ( .B1(n9700), .B2(n9655), .A(n9646), .ZN(P2_U3476) );
  AOI21_X1 U10746 ( .B1(n9648), .B2(n11097), .A(n9647), .ZN(n9701) );
  MUX2_X1 U10747 ( .A(n9649), .B(n9701), .S(n11100), .Z(n9650) );
  OAI21_X1 U10748 ( .B1(n9704), .B2(n9655), .A(n9650), .ZN(P2_U3475) );
  AOI21_X1 U10749 ( .B1(n11097), .B2(n9652), .A(n9651), .ZN(n9705) );
  MUX2_X1 U10750 ( .A(n9653), .B(n9705), .S(n11100), .Z(n9654) );
  OAI21_X1 U10751 ( .B1(n9709), .B2(n9655), .A(n9654), .ZN(P2_U3474) );
  NAND2_X1 U10752 ( .A1(n9656), .A2(n11104), .ZN(n9659) );
  NAND2_X1 U10753 ( .A1(n11101), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9657) );
  OAI211_X1 U10754 ( .C1(n9658), .C2(n9708), .A(n9659), .B(n9657), .ZN(
        P2_U3458) );
  NAND2_X1 U10755 ( .A1(n11101), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9660) );
  OAI211_X1 U10756 ( .C1(n9661), .C2(n9708), .A(n9660), .B(n9659), .ZN(
        P2_U3457) );
  MUX2_X1 U10757 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9662), .S(n11104), .Z(
        P2_U3456) );
  MUX2_X1 U10758 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9663), .S(n11104), .Z(
        P2_U3454) );
  MUX2_X1 U10759 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9664), .S(n11104), .Z(
        n9665) );
  INV_X1 U10760 ( .A(n9665), .ZN(n9666) );
  OAI21_X1 U10761 ( .B1(n9667), .B2(n9708), .A(n9666), .ZN(P2_U3453) );
  INV_X1 U10762 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9669) );
  MUX2_X1 U10763 ( .A(n9669), .B(n9668), .S(n11104), .Z(n9670) );
  OAI21_X1 U10764 ( .B1(n9671), .B2(n9708), .A(n9670), .ZN(P2_U3452) );
  INV_X1 U10765 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9673) );
  MUX2_X1 U10766 ( .A(n9673), .B(n9672), .S(n11104), .Z(n9674) );
  OAI21_X1 U10767 ( .B1(n9675), .B2(n9708), .A(n9674), .ZN(P2_U3451) );
  INV_X1 U10768 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9677) );
  MUX2_X1 U10769 ( .A(n9677), .B(n9676), .S(n11104), .Z(n9678) );
  OAI21_X1 U10770 ( .B1(n9679), .B2(n9708), .A(n9678), .ZN(P2_U3450) );
  MUX2_X1 U10771 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9680), .S(n11104), .Z(
        P2_U3449) );
  INV_X1 U10772 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9682) );
  MUX2_X1 U10773 ( .A(n9682), .B(n9681), .S(n11104), .Z(n9683) );
  OAI21_X1 U10774 ( .B1(n9684), .B2(n9708), .A(n9683), .ZN(P2_U3448) );
  INV_X1 U10775 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9686) );
  MUX2_X1 U10776 ( .A(n9686), .B(n9685), .S(n11104), .Z(n9687) );
  OAI21_X1 U10777 ( .B1(n9688), .B2(n9708), .A(n9687), .ZN(P2_U3447) );
  INV_X1 U10778 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9690) );
  MUX2_X1 U10779 ( .A(n9690), .B(n9689), .S(n11104), .Z(n9691) );
  OAI21_X1 U10780 ( .B1(n9692), .B2(n9708), .A(n9691), .ZN(P2_U3446) );
  MUX2_X1 U10781 ( .A(n9694), .B(n9693), .S(n11104), .Z(n9695) );
  OAI21_X1 U10782 ( .B1(n9696), .B2(n9708), .A(n9695), .ZN(P2_U3444) );
  INV_X1 U10783 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9698) );
  MUX2_X1 U10784 ( .A(n9698), .B(n9697), .S(n11104), .Z(n9699) );
  OAI21_X1 U10785 ( .B1(n9700), .B2(n9708), .A(n9699), .ZN(P2_U3441) );
  INV_X1 U10786 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9702) );
  MUX2_X1 U10787 ( .A(n9702), .B(n9701), .S(n11104), .Z(n9703) );
  OAI21_X1 U10788 ( .B1(n9704), .B2(n9708), .A(n9703), .ZN(P2_U3438) );
  INV_X1 U10789 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9706) );
  MUX2_X1 U10790 ( .A(n9706), .B(n9705), .S(n11104), .Z(n9707) );
  OAI21_X1 U10791 ( .B1(n9709), .B2(n9708), .A(n9707), .ZN(P2_U3435) );
  NAND3_X1 U10792 ( .A1(n9711), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n9713) );
  OAI22_X1 U10793 ( .A1(n9710), .A2(n9713), .B1(n9712), .B2(n8618), .ZN(n9714)
         );
  AOI21_X1 U10794 ( .B1(n10593), .B2(n5180), .A(n9714), .ZN(n9715) );
  INV_X1 U10795 ( .A(n9715), .ZN(P2_U3264) );
  INV_X1 U10796 ( .A(n9716), .ZN(n10597) );
  MUX2_X1 U10797 ( .A(n9720), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U10798 ( .A(n9721), .ZN(n9725) );
  AOI21_X1 U10799 ( .B1(n9870), .B2(n9723), .A(n9722), .ZN(n9724) );
  OAI21_X1 U10800 ( .B1(n9725), .B2(n9724), .A(n9871), .ZN(n9729) );
  NOR2_X1 U10801 ( .A1(n9874), .A2(n10332), .ZN(n9727) );
  OAI22_X1 U10802 ( .A1(n10326), .A2(n9877), .B1(n9876), .B2(n10325), .ZN(
        n9726) );
  AOI211_X1 U10803 ( .C1(P1_REG3_REG_27__SCAN_IN), .C2(P1_U3086), .A(n9727), 
        .B(n9726), .ZN(n9728) );
  OAI211_X1 U10804 ( .C1(n10484), .C2(n9882), .A(n9729), .B(n9728), .ZN(
        P1_U3214) );
  INV_X1 U10805 ( .A(n9730), .ZN(n9731) );
  NOR2_X1 U10806 ( .A1(n9732), .A2(n9731), .ZN(n9836) );
  OR2_X1 U10807 ( .A1(n9836), .A2(n9838), .ZN(n9835) );
  NAND2_X1 U10808 ( .A1(n9732), .A2(n9731), .ZN(n9833) );
  NAND2_X1 U10809 ( .A1(n9835), .A2(n9833), .ZN(n9837) );
  XNOR2_X1 U10810 ( .A(n9734), .B(n9733), .ZN(n9735) );
  XNOR2_X1 U10811 ( .A(n9837), .B(n9735), .ZN(n9740) );
  OAI22_X1 U10812 ( .A1(n9874), .A2(n10392), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9736), .ZN(n9738) );
  OAI22_X1 U10813 ( .A1(n10425), .A2(n9876), .B1(n9877), .B2(n9775), .ZN(n9737) );
  AOI211_X1 U10814 ( .C1(n10501), .C2(n9863), .A(n9738), .B(n9737), .ZN(n9739)
         );
  OAI21_X1 U10815 ( .B1(n9740), .B2(n9866), .A(n9739), .ZN(P1_U3216) );
  OAI21_X1 U10816 ( .B1(n9743), .B2(n9742), .A(n9741), .ZN(n9744) );
  NAND2_X1 U10817 ( .A1(n9744), .A2(n9871), .ZN(n9750) );
  AOI22_X1 U10818 ( .A1(n9845), .A2(n9745), .B1(n10917), .B2(n9863), .ZN(n9749) );
  NAND2_X1 U10819 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n10210) );
  INV_X1 U10820 ( .A(n10210), .ZN(n9747) );
  NOR2_X1 U10821 ( .A1(n9874), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9746) );
  AOI211_X1 U10822 ( .C1(n9846), .C2(n10170), .A(n9747), .B(n9746), .ZN(n9748)
         );
  NAND3_X1 U10823 ( .A1(n9750), .A2(n9749), .A3(n9748), .ZN(P1_U3218) );
  NAND2_X1 U10824 ( .A1(n9751), .A2(n5117), .ZN(n9758) );
  XOR2_X1 U10825 ( .A(n9757), .B(n9758), .Z(n9756) );
  NAND2_X1 U10826 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n10266)
         );
  OAI21_X1 U10827 ( .B1(n9874), .B2(n9752), .A(n10266), .ZN(n9754) );
  OAI22_X1 U10828 ( .A1(n9799), .A2(n9876), .B1(n9877), .B2(n10426), .ZN(n9753) );
  AOI211_X1 U10829 ( .C1(n10522), .C2(n9863), .A(n9754), .B(n9753), .ZN(n9755)
         );
  OAI21_X1 U10830 ( .B1(n9756), .B2(n9866), .A(n9755), .ZN(P1_U3219) );
  NAND2_X1 U10831 ( .A1(n9758), .A2(n9757), .ZN(n9760) );
  NAND2_X1 U10832 ( .A1(n9760), .A2(n9759), .ZN(n9826) );
  NAND2_X1 U10833 ( .A1(n9826), .A2(n9827), .ZN(n9765) );
  NAND2_X1 U10834 ( .A1(n9765), .A2(n9761), .ZN(n9763) );
  AOI21_X1 U10835 ( .B1(n9763), .B2(n9762), .A(n9866), .ZN(n9767) );
  NAND2_X1 U10836 ( .A1(n9765), .A2(n9764), .ZN(n9766) );
  NAND2_X1 U10837 ( .A1(n9767), .A2(n9766), .ZN(n9771) );
  NOR2_X1 U10838 ( .A1(n9874), .A2(n10429), .ZN(n9769) );
  OAI22_X1 U10839 ( .A1(n10425), .A2(n9877), .B1(n9876), .B2(n10426), .ZN(
        n9768) );
  AOI211_X1 U10840 ( .C1(P1_REG3_REG_21__SCAN_IN), .C2(P1_U3086), .A(n9769), 
        .B(n9768), .ZN(n9770) );
  OAI211_X1 U10841 ( .C1(n10573), .C2(n9882), .A(n9771), .B(n9770), .ZN(
        P1_U3223) );
  OAI21_X1 U10842 ( .B1(n9773), .B2(n9772), .A(n9869), .ZN(n9774) );
  NAND2_X1 U10843 ( .A1(n9774), .A2(n9871), .ZN(n9779) );
  NOR2_X1 U10844 ( .A1(n9874), .A2(n10362), .ZN(n9777) );
  OAI22_X1 U10845 ( .A1(n9775), .A2(n9876), .B1(n9877), .B2(n10325), .ZN(n9776) );
  AOI211_X1 U10846 ( .C1(P1_REG3_REG_25__SCAN_IN), .C2(P1_U3086), .A(n9777), 
        .B(n9776), .ZN(n9778) );
  OAI211_X1 U10847 ( .C1(n10365), .C2(n9882), .A(n9779), .B(n9778), .ZN(
        P1_U3225) );
  OAI21_X1 U10848 ( .B1(n9782), .B2(n9781), .A(n9780), .ZN(n9783) );
  NAND2_X1 U10849 ( .A1(n9783), .A2(n9871), .ZN(n9793) );
  INV_X1 U10850 ( .A(n9784), .ZN(n9786) );
  AOI21_X1 U10851 ( .B1(n9803), .B2(n9786), .A(n9785), .ZN(n9792) );
  OAI22_X1 U10852 ( .A1(n9787), .A2(n9876), .B1(n9877), .B2(n9860), .ZN(n9788)
         );
  INV_X1 U10853 ( .A(n9788), .ZN(n9791) );
  NAND2_X1 U10854 ( .A1(n9789), .A2(n9863), .ZN(n9790) );
  NAND4_X1 U10855 ( .A1(n9793), .A2(n9792), .A3(n9791), .A4(n9790), .ZN(
        P1_U3226) );
  NAND2_X1 U10856 ( .A1(n9795), .A2(n9794), .ZN(n9796) );
  XNOR2_X1 U10857 ( .A(n9797), .B(n9796), .ZN(n9806) );
  OAI22_X1 U10858 ( .A1(n9799), .A2(n9877), .B1(n9876), .B2(n9798), .ZN(n9800)
         );
  AOI211_X1 U10859 ( .C1(n9803), .C2(n9802), .A(n9801), .B(n9800), .ZN(n9805)
         );
  NAND2_X1 U10860 ( .A1(n10535), .A2(n9863), .ZN(n9804) );
  OAI211_X1 U10861 ( .C1(n9806), .C2(n9866), .A(n9805), .B(n9804), .ZN(
        P1_U3228) );
  NOR2_X1 U10862 ( .A1(n9808), .A2(n5461), .ZN(n9809) );
  XNOR2_X1 U10863 ( .A(n9810), .B(n9809), .ZN(n9815) );
  OAI22_X1 U10864 ( .A1(n9874), .A2(n10383), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9811), .ZN(n9813) );
  OAI22_X1 U10865 ( .A1(n10417), .A2(n9876), .B1(n9877), .B2(n9875), .ZN(n9812) );
  AOI211_X1 U10866 ( .C1(n10382), .C2(n9863), .A(n9813), .B(n9812), .ZN(n9814)
         );
  OAI21_X1 U10867 ( .B1(n9815), .B2(n9866), .A(n9814), .ZN(P1_U3229) );
  AOI21_X1 U10868 ( .B1(n9817), .B2(n9816), .A(n9866), .ZN(n9819) );
  NAND2_X1 U10869 ( .A1(n9819), .A2(n9818), .ZN(n9825) );
  AOI22_X1 U10870 ( .A1(n9846), .A2(n10169), .B1(n9820), .B2(n9863), .ZN(n9824) );
  AND2_X1 U10871 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n10218) );
  NOR2_X1 U10872 ( .A1(n9874), .A2(n9821), .ZN(n9822) );
  AOI211_X1 U10873 ( .C1(n9845), .C2(n10168), .A(n10218), .B(n9822), .ZN(n9823) );
  NAND3_X1 U10874 ( .A1(n9825), .A2(n9824), .A3(n9823), .ZN(P1_U3230) );
  XOR2_X1 U10875 ( .A(n9827), .B(n9826), .Z(n9832) );
  INV_X1 U10876 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9828) );
  OAI22_X1 U10877 ( .A1(n9874), .A2(n10441), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9828), .ZN(n9830) );
  OAI22_X1 U10878 ( .A1(n10448), .A2(n9876), .B1(n9877), .B2(n10449), .ZN(
        n9829) );
  AOI211_X1 U10879 ( .C1(n10517), .C2(n9863), .A(n9830), .B(n9829), .ZN(n9831)
         );
  OAI21_X1 U10880 ( .B1(n9832), .B2(n9866), .A(n9831), .ZN(P1_U3233) );
  INV_X1 U10881 ( .A(n9833), .ZN(n9834) );
  NOR2_X1 U10882 ( .A1(n9835), .A2(n9834), .ZN(n9839) );
  OAI22_X1 U10883 ( .A1(n9839), .A2(n9838), .B1(n9837), .B2(n9836), .ZN(n9840)
         );
  NAND2_X1 U10884 ( .A1(n9840), .A2(n9871), .ZN(n9844) );
  NOR2_X1 U10885 ( .A1(n9874), .A2(n10410), .ZN(n9842) );
  OAI22_X1 U10886 ( .A1(n10449), .A2(n9876), .B1(n9877), .B2(n10417), .ZN(
        n9841) );
  AOI211_X1 U10887 ( .C1(P1_REG3_REG_22__SCAN_IN), .C2(P1_U3086), .A(n9842), 
        .B(n9841), .ZN(n9843) );
  OAI211_X1 U10888 ( .C1(n10409), .C2(n9882), .A(n9844), .B(n9843), .ZN(
        P1_U3235) );
  AOI22_X1 U10889 ( .A1(n9846), .A2(n10171), .B1(n9845), .B2(n10169), .ZN(
        n9855) );
  AOI22_X1 U10890 ( .A1(n9863), .A2(n9848), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n9847), .ZN(n9854) );
  OAI21_X1 U10891 ( .B1(n9851), .B2(n9850), .A(n9849), .ZN(n9852) );
  NAND2_X1 U10892 ( .A1(n9852), .A2(n9871), .ZN(n9853) );
  NAND3_X1 U10893 ( .A1(n9855), .A2(n9854), .A3(n9853), .ZN(P1_U3237) );
  NAND2_X1 U10894 ( .A1(n9856), .A2(n5117), .ZN(n9858) );
  XNOR2_X1 U10895 ( .A(n9858), .B(n9857), .ZN(n9867) );
  NAND2_X1 U10896 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10756)
         );
  OAI21_X1 U10897 ( .B1(n9874), .B2(n9859), .A(n10756), .ZN(n9862) );
  OAI22_X1 U10898 ( .A1(n9860), .A2(n9876), .B1(n9877), .B2(n10448), .ZN(n9861) );
  AOI211_X1 U10899 ( .C1(n9864), .C2(n9863), .A(n9862), .B(n9861), .ZN(n9865)
         );
  OAI21_X1 U10900 ( .B1(n9867), .B2(n9866), .A(n9865), .ZN(P1_U3238) );
  AND2_X1 U10901 ( .A1(n9869), .A2(n9868), .ZN(n9873) );
  OAI211_X1 U10902 ( .C1(n9873), .C2(n9872), .A(n9871), .B(n9870), .ZN(n9881)
         );
  NOR2_X1 U10903 ( .A1(n9874), .A2(n10351), .ZN(n9879) );
  OAI22_X1 U10904 ( .A1(n10309), .A2(n9877), .B1(n9876), .B2(n9875), .ZN(n9878) );
  AOI211_X1 U10905 ( .C1(P1_REG3_REG_26__SCAN_IN), .C2(P1_U3086), .A(n9879), 
        .B(n9878), .ZN(n9880) );
  OAI211_X1 U10906 ( .C1(n10562), .C2(n9882), .A(n9881), .B(n9880), .ZN(
        P1_U3240) );
  NAND2_X1 U10907 ( .A1(n10593), .A2(n9893), .ZN(n9884) );
  INV_X1 U10908 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10589) );
  OR2_X1 U10909 ( .A1(n9895), .A2(n10589), .ZN(n9883) );
  NAND2_X1 U10910 ( .A1(n9885), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n9892) );
  INV_X1 U10911 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9886) );
  OR2_X1 U10912 ( .A1(n9887), .A2(n9886), .ZN(n9891) );
  INV_X1 U10913 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9888) );
  OR2_X1 U10914 ( .A1(n9889), .A2(n9888), .ZN(n9890) );
  AND3_X1 U10915 ( .A1(n9892), .A2(n9891), .A3(n9890), .ZN(n9940) );
  NAND2_X1 U10916 ( .A1(n10283), .A2(n9940), .ZN(n10139) );
  NAND2_X1 U10917 ( .A1(n8658), .A2(n9893), .ZN(n9897) );
  OR2_X1 U10918 ( .A1(n9895), .A2(n9894), .ZN(n9896) );
  INV_X1 U10919 ( .A(n10155), .ZN(n9935) );
  OR2_X1 U10920 ( .A1(n10291), .A2(n9935), .ZN(n10101) );
  NAND2_X1 U10921 ( .A1(n10061), .A2(n10056), .ZN(n10134) );
  NAND2_X1 U10922 ( .A1(n10057), .A2(n10052), .ZN(n10131) );
  NAND2_X1 U10923 ( .A1(n10044), .A2(n9898), .ZN(n10127) );
  NAND2_X1 U10924 ( .A1(n10036), .A2(n9899), .ZN(n9942) );
  NAND2_X1 U10925 ( .A1(n9942), .A2(n10037), .ZN(n9900) );
  NAND2_X1 U10926 ( .A1(n10048), .A2(n9900), .ZN(n9901) );
  NAND2_X1 U10927 ( .A1(n9901), .A2(n10040), .ZN(n9902) );
  AND2_X1 U10928 ( .A1(n9902), .A2(n10042), .ZN(n9903) );
  OAI211_X1 U10929 ( .C1(n10127), .C2(n9903), .A(n10053), .B(n10049), .ZN(
        n10129) );
  NAND2_X1 U10930 ( .A1(n10040), .A2(n10037), .ZN(n10125) );
  NAND2_X1 U10931 ( .A1(n10091), .A2(n10024), .ZN(n9904) );
  OAI21_X1 U10932 ( .B1(n10016), .B2(n10010), .A(n9904), .ZN(n9927) );
  INV_X1 U10933 ( .A(n10006), .ZN(n10009) );
  NAND2_X1 U10934 ( .A1(n10005), .A2(n9999), .ZN(n9991) );
  INV_X1 U10935 ( .A(n9991), .ZN(n9924) );
  NAND2_X1 U10936 ( .A1(n9989), .A2(n9980), .ZN(n9995) );
  NAND2_X1 U10937 ( .A1(n10171), .A2(n5729), .ZN(n9908) );
  NAND2_X1 U10938 ( .A1(n9906), .A2(n9905), .ZN(n9907) );
  NAND3_X1 U10939 ( .A1(n9908), .A2(n9907), .A3(n10107), .ZN(n9909) );
  NAND2_X1 U10940 ( .A1(n9909), .A2(n10904), .ZN(n9910) );
  OAI21_X1 U10941 ( .B1(n9949), .B2(n9910), .A(n9948), .ZN(n9911) );
  NAND2_X1 U10942 ( .A1(n9947), .A2(n9953), .ZN(n9943) );
  AOI21_X1 U10943 ( .B1(n9911), .B2(n9951), .A(n9943), .ZN(n9913) );
  NAND2_X1 U10944 ( .A1(n9912), .A2(n9950), .ZN(n9944) );
  OAI21_X1 U10945 ( .B1(n9913), .B2(n9944), .A(n9955), .ZN(n9914) );
  NAND2_X1 U10946 ( .A1(n9914), .A2(n10070), .ZN(n9915) );
  NAND2_X1 U10947 ( .A1(n9915), .A2(n10078), .ZN(n9917) );
  NAND3_X1 U10948 ( .A1(n9917), .A2(n9916), .A3(n11021), .ZN(n9919) );
  INV_X1 U10949 ( .A(n9983), .ZN(n9918) );
  AOI21_X1 U10950 ( .B1(n9919), .B2(n9975), .A(n9918), .ZN(n9920) );
  NAND2_X1 U10951 ( .A1(n9988), .A2(n9976), .ZN(n9986) );
  NOR2_X1 U10952 ( .A1(n9920), .A2(n9986), .ZN(n9921) );
  OAI211_X1 U10953 ( .C1(n9995), .C2(n9921), .A(n9994), .B(n9997), .ZN(n9923)
         );
  INV_X1 U10954 ( .A(n10003), .ZN(n9922) );
  AOI21_X1 U10955 ( .B1(n9924), .B2(n9923), .A(n9922), .ZN(n9925) );
  OR3_X1 U10956 ( .A1(n10091), .A2(n10009), .A3(n9925), .ZN(n9926) );
  NAND3_X1 U10957 ( .A1(n9927), .A2(n10019), .A3(n9926), .ZN(n9928) );
  NAND2_X1 U10958 ( .A1(n9928), .A2(n10027), .ZN(n9929) );
  NAND2_X1 U10959 ( .A1(n9930), .A2(n9929), .ZN(n9931) );
  NAND3_X1 U10960 ( .A1(n9932), .A2(n9931), .A3(n10124), .ZN(n9933) );
  NOR2_X1 U10961 ( .A1(n10129), .A2(n5607), .ZN(n9934) );
  NOR2_X1 U10962 ( .A1(n10131), .A2(n9934), .ZN(n9936) );
  NAND2_X1 U10963 ( .A1(n10291), .A2(n9935), .ZN(n10100) );
  OAI211_X1 U10964 ( .C1(n10134), .C2(n9936), .A(n10100), .B(n10132), .ZN(
        n9937) );
  NAND3_X1 U10965 ( .A1(n10139), .A2(n10101), .A3(n9937), .ZN(n9938) );
  OR2_X1 U10966 ( .A1(n10283), .A2(n9940), .ZN(n10119) );
  NAND2_X1 U10967 ( .A1(n9938), .A2(n10119), .ZN(n9939) );
  XNOR2_X1 U10968 ( .A(n9939), .B(n10274), .ZN(n10146) );
  INV_X1 U10969 ( .A(n9940), .ZN(n10287) );
  NAND2_X1 U10970 ( .A1(n10287), .A2(n10155), .ZN(n10062) );
  OR2_X1 U10971 ( .A1(n10291), .A2(n10062), .ZN(n10136) );
  NAND3_X1 U10972 ( .A1(n10139), .A2(n10138), .A3(n10136), .ZN(n10105) );
  INV_X1 U10973 ( .A(n10127), .ZN(n10041) );
  NAND2_X1 U10974 ( .A1(n10037), .A2(n10124), .ZN(n9941) );
  MUX2_X1 U10975 ( .A(n9942), .B(n9941), .S(n10060), .Z(n10039) );
  NAND3_X1 U10976 ( .A1(n10905), .A2(n9951), .A3(n10904), .ZN(n9946) );
  NOR2_X1 U10977 ( .A1(n10072), .A2(n9943), .ZN(n9945) );
  AOI22_X1 U10978 ( .A1(n9946), .A2(n9945), .B1(n9955), .B2(n9944), .ZN(n9960)
         );
  OAI211_X1 U10979 ( .C1(n9949), .C2(n10065), .A(n9948), .B(n9947), .ZN(n9952)
         );
  NAND3_X1 U10980 ( .A1(n9952), .A2(n9951), .A3(n9950), .ZN(n9954) );
  NAND2_X1 U10981 ( .A1(n9954), .A2(n9953), .ZN(n9958) );
  INV_X1 U10982 ( .A(n9955), .ZN(n9956) );
  AOI21_X1 U10983 ( .B1(n9958), .B2(n9957), .A(n9956), .ZN(n9959) );
  INV_X1 U10984 ( .A(n10060), .ZN(n10055) );
  MUX2_X1 U10985 ( .A(n9960), .B(n9959), .S(n10055), .Z(n9965) );
  MUX2_X1 U10986 ( .A(n9962), .B(n10070), .S(n10060), .Z(n9963) );
  OAI211_X1 U10987 ( .C1(n9965), .C2(n9964), .A(n5534), .B(n9963), .ZN(n9970)
         );
  MUX2_X1 U10988 ( .A(n9967), .B(n9966), .S(n10055), .Z(n9969) );
  NAND2_X1 U10989 ( .A1(n11021), .A2(n9971), .ZN(n9972) );
  MUX2_X1 U10990 ( .A(n9973), .B(n9972), .S(n10055), .Z(n9974) );
  INV_X1 U10991 ( .A(n9975), .ZN(n9984) );
  OAI211_X1 U10992 ( .C1(n9978), .C2(n9977), .A(n9976), .B(n9975), .ZN(n9979)
         );
  INV_X1 U10993 ( .A(n9979), .ZN(n9982) );
  NAND2_X1 U10994 ( .A1(n9980), .A2(n9983), .ZN(n9981) );
  OAI211_X1 U10995 ( .C1(n9984), .C2(n10075), .A(n9983), .B(n11021), .ZN(n9985) );
  INV_X1 U10996 ( .A(n9985), .ZN(n9987) );
  NAND2_X1 U10997 ( .A1(n9994), .A2(n9988), .ZN(n9990) );
  OAI21_X1 U10998 ( .B1(n9996), .B2(n9990), .A(n9989), .ZN(n9993) );
  AOI21_X1 U10999 ( .B1(n9993), .B2(n9992), .A(n9991), .ZN(n10002) );
  OAI21_X1 U11000 ( .B1(n9996), .B2(n9995), .A(n9994), .ZN(n10000) );
  NAND2_X1 U11001 ( .A1(n10003), .A2(n9997), .ZN(n9998) );
  AOI21_X1 U11002 ( .B1(n10000), .B2(n9999), .A(n9998), .ZN(n10001) );
  MUX2_X1 U11003 ( .A(n10002), .B(n10001), .S(n10060), .Z(n10015) );
  NAND2_X1 U11004 ( .A1(n10004), .A2(n10003), .ZN(n10008) );
  NAND2_X1 U11005 ( .A1(n10006), .A2(n10005), .ZN(n10007) );
  MUX2_X1 U11006 ( .A(n10008), .B(n10007), .S(n10060), .Z(n10014) );
  MUX2_X1 U11007 ( .A(n10010), .B(n10009), .S(n10055), .Z(n10011) );
  NOR2_X1 U11008 ( .A1(n10012), .A2(n10011), .ZN(n10013) );
  OAI21_X1 U11009 ( .B1(n10015), .B2(n10014), .A(n10013), .ZN(n10023) );
  INV_X1 U11010 ( .A(n10016), .ZN(n10094) );
  NAND2_X1 U11011 ( .A1(n10023), .A2(n10094), .ZN(n10018) );
  NAND3_X1 U11012 ( .A1(n10018), .A2(n10027), .A3(n10017), .ZN(n10020) );
  NAND3_X1 U11013 ( .A1(n10020), .A2(n10029), .A3(n10019), .ZN(n10021) );
  NAND2_X1 U11014 ( .A1(n10021), .A2(n10026), .ZN(n10032) );
  INV_X1 U11015 ( .A(n10091), .ZN(n10022) );
  NAND2_X1 U11016 ( .A1(n10023), .A2(n10022), .ZN(n10025) );
  NAND3_X1 U11017 ( .A1(n10093), .A2(n10025), .A3(n10024), .ZN(n10028) );
  NAND3_X1 U11018 ( .A1(n10028), .A2(n10027), .A3(n10026), .ZN(n10030) );
  NAND2_X1 U11019 ( .A1(n10030), .A2(n10029), .ZN(n10031) );
  MUX2_X1 U11020 ( .A(n10034), .B(n10033), .S(n10060), .Z(n10035) );
  MUX2_X1 U11021 ( .A(n10037), .B(n10036), .S(n10060), .Z(n10038) );
  NAND3_X1 U11022 ( .A1(n10041), .A2(n10040), .A3(n10047), .ZN(n10046) );
  INV_X1 U11023 ( .A(n10042), .ZN(n10043) );
  NAND2_X1 U11024 ( .A1(n10044), .A2(n10043), .ZN(n10045) );
  INV_X1 U11025 ( .A(n10358), .ZN(n10367) );
  NAND4_X1 U11026 ( .A1(n10346), .A2(n10367), .A3(n10048), .A4(n10047), .ZN(
        n10051) );
  NAND2_X1 U11027 ( .A1(n10127), .A2(n10049), .ZN(n10050) );
  MUX2_X1 U11028 ( .A(n10053), .B(n10052), .S(n10055), .Z(n10054) );
  MUX2_X1 U11029 ( .A(n10057), .B(n10056), .S(n10055), .Z(n10058) );
  NAND2_X1 U11030 ( .A1(n10059), .A2(n10058), .ZN(n10064) );
  MUX2_X1 U11031 ( .A(n10132), .B(n10061), .S(n10060), .Z(n10063) );
  AND2_X1 U11032 ( .A1(n10291), .A2(n10062), .ZN(n10135) );
  INV_X1 U11033 ( .A(n10135), .ZN(n10113) );
  OAI211_X1 U11034 ( .C1(n10102), .C2(n10064), .A(n10063), .B(n10113), .ZN(
        n10115) );
  INV_X1 U11035 ( .A(n11023), .ZN(n10082) );
  NOR2_X1 U11036 ( .A1(n10065), .A2(n10107), .ZN(n10068) );
  NAND4_X1 U11037 ( .A1(n10069), .A2(n10068), .A3(n10067), .A4(n10066), .ZN(
        n10074) );
  INV_X1 U11038 ( .A(n10070), .ZN(n10073) );
  NOR4_X1 U11039 ( .A1(n10074), .A2(n10073), .A3(n10072), .A4(n10071), .ZN(
        n10076) );
  NAND4_X1 U11040 ( .A1(n10078), .A2(n10077), .A3(n10076), .A4(n10075), .ZN(
        n10080) );
  NOR2_X1 U11041 ( .A1(n10080), .A2(n10079), .ZN(n10081) );
  NAND3_X1 U11042 ( .A1(n10083), .A2(n10082), .A3(n10081), .ZN(n10084) );
  NOR3_X1 U11043 ( .A1(n10086), .A2(n10085), .A3(n10084), .ZN(n10087) );
  NAND3_X1 U11044 ( .A1(n10089), .A2(n10088), .A3(n10087), .ZN(n10090) );
  NOR2_X1 U11045 ( .A1(n10091), .A2(n10090), .ZN(n10092) );
  AND4_X1 U11046 ( .A1(n10446), .A2(n10094), .A3(n10093), .A4(n10092), .ZN(
        n10095) );
  NAND4_X1 U11047 ( .A1(n10398), .A2(n5528), .A3(n10415), .A4(n10095), .ZN(
        n10096) );
  NOR2_X1 U11048 ( .A1(n10358), .A2(n10096), .ZN(n10097) );
  NAND4_X1 U11049 ( .A1(n10329), .A2(n10346), .A3(n10379), .A4(n10097), .ZN(
        n10098) );
  NOR2_X1 U11050 ( .A1(n10314), .A2(n10098), .ZN(n10099) );
  NAND3_X1 U11051 ( .A1(n10101), .A2(n10100), .A3(n10099), .ZN(n10103) );
  NOR2_X1 U11052 ( .A1(n10103), .A2(n10102), .ZN(n10104) );
  NAND3_X1 U11053 ( .A1(n10119), .A2(n10104), .A3(n10139), .ZN(n10140) );
  NOR2_X1 U11054 ( .A1(n10113), .A2(n10106), .ZN(n10110) );
  NAND2_X1 U11055 ( .A1(n10287), .A2(n10138), .ZN(n10108) );
  OAI22_X1 U11056 ( .A1(n10113), .A2(n10108), .B1(n10107), .B2(n10280), .ZN(
        n10109) );
  AOI21_X1 U11057 ( .B1(n10547), .B2(n10110), .A(n10109), .ZN(n10123) );
  OAI21_X1 U11058 ( .B1(n10111), .B2(n10117), .A(n10280), .ZN(n10112) );
  OAI211_X1 U11059 ( .C1(n10113), .C2(n10280), .A(n10112), .B(n10136), .ZN(
        n10114) );
  INV_X1 U11060 ( .A(n10114), .ZN(n10116) );
  NAND4_X1 U11061 ( .A1(n10116), .A2(n10119), .A3(n10115), .A4(n10139), .ZN(
        n10122) );
  OR2_X1 U11062 ( .A1(n10117), .A2(n10274), .ZN(n10118) );
  AOI21_X1 U11063 ( .B1(n10136), .B2(n10287), .A(n10280), .ZN(n10120) );
  NAND2_X1 U11064 ( .A1(n10120), .A2(n10283), .ZN(n10121) );
  OR3_X1 U11065 ( .A1(n10125), .A2(n5229), .A3(n10414), .ZN(n10126) );
  NOR2_X1 U11066 ( .A1(n10127), .A2(n10126), .ZN(n10128) );
  NOR2_X1 U11067 ( .A1(n10129), .A2(n10128), .ZN(n10130) );
  NOR2_X1 U11068 ( .A1(n10131), .A2(n10130), .ZN(n10133) );
  OAI21_X1 U11069 ( .B1(n10134), .B2(n10133), .A(n10132), .ZN(n10137) );
  AOI21_X1 U11070 ( .B1(n10137), .B2(n10136), .A(n10135), .ZN(n10142) );
  NAND2_X1 U11071 ( .A1(n10139), .A2(n10138), .ZN(n10141) );
  OAI21_X1 U11072 ( .B1(n10142), .B2(n10141), .A(n10140), .ZN(n10143) );
  NAND2_X1 U11073 ( .A1(n10143), .A2(n10274), .ZN(n10144) );
  NOR3_X1 U11074 ( .A1(n10148), .A2(n10147), .A3(n10663), .ZN(n10149) );
  AOI211_X1 U11075 ( .C1(n10153), .C2(n10151), .A(n10150), .B(n10149), .ZN(
        n10152) );
  INV_X1 U11076 ( .A(n10154), .ZN(P1_U3242) );
  MUX2_X1 U11077 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n10287), .S(P1_U3973), .Z(
        P1_U3585) );
  MUX2_X1 U11078 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n10155), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U11079 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n6159), .S(P1_U3973), .Z(
        P1_U3582) );
  INV_X1 U11080 ( .A(n10309), .ZN(n10343) );
  MUX2_X1 U11081 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n10343), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U11082 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n10368), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U11083 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n10375), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U11084 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n10400), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U11085 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n10399), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U11086 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n10156), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U11087 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n10157), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U11088 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n10158), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U11089 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n10159), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U11090 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n10160), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U11091 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n10161), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U11092 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n10162), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U11093 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n11025), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U11094 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n10163), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U11095 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n11028), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U11096 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n10164), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U11097 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n10165), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U11098 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n10166), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U11099 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n10167), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U11100 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n10168), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U11101 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n10169), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U11102 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n10170), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U11103 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n10171), .S(P1_U3973), .Z(
        P1_U3555) );
  OAI211_X1 U11104 ( .C1(n10174), .C2(n10173), .A(n10776), .B(n10172), .ZN(
        n10184) );
  OAI211_X1 U11105 ( .C1(n10177), .C2(n10176), .A(n10782), .B(n10175), .ZN(
        n10183) );
  INV_X1 U11106 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10179) );
  OAI22_X1 U11107 ( .A1(n10808), .A2(n10179), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10178), .ZN(n10180) );
  AOI21_X1 U11108 ( .B1(n10799), .B2(n10181), .A(n10180), .ZN(n10182) );
  NAND3_X1 U11109 ( .A1(n10184), .A2(n10183), .A3(n10182), .ZN(P1_U3244) );
  INV_X1 U11110 ( .A(n10660), .ZN(n10185) );
  OR2_X1 U11111 ( .A1(n10185), .A2(n6210), .ZN(n10189) );
  NOR2_X1 U11112 ( .A1(n6210), .A2(n10662), .ZN(n10186) );
  XNOR2_X1 U11113 ( .A(n10186), .B(P1_IR_REG_0__SCAN_IN), .ZN(n10187) );
  NAND2_X1 U11114 ( .A1(n10187), .A2(n10189), .ZN(n10188) );
  OAI211_X1 U11115 ( .C1(n10190), .C2(n10189), .A(P1_U3973), .B(n10188), .ZN(
        n10232) );
  INV_X1 U11116 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10192) );
  OAI22_X1 U11117 ( .A1(n10808), .A2(n10192), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10191), .ZN(n10193) );
  AOI21_X1 U11118 ( .B1(n10799), .B2(n10194), .A(n10193), .ZN(n10203) );
  OAI211_X1 U11119 ( .C1(n10197), .C2(n10196), .A(n10782), .B(n10195), .ZN(
        n10202) );
  OAI211_X1 U11120 ( .C1(n10200), .C2(n10199), .A(n10776), .B(n10198), .ZN(
        n10201) );
  NAND4_X1 U11121 ( .A1(n10232), .A2(n10203), .A3(n10202), .A4(n10201), .ZN(
        P1_U3245) );
  OAI211_X1 U11122 ( .C1(n10206), .C2(n10205), .A(n10776), .B(n10204), .ZN(
        n10216) );
  OAI211_X1 U11123 ( .C1(n10209), .C2(n10208), .A(n10782), .B(n10207), .ZN(
        n10215) );
  INV_X1 U11124 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10211) );
  OAI21_X1 U11125 ( .B1(n10808), .B2(n10211), .A(n10210), .ZN(n10212) );
  AOI21_X1 U11126 ( .B1(n10799), .B2(n10213), .A(n10212), .ZN(n10214) );
  NAND3_X1 U11127 ( .A1(n10216), .A2(n10215), .A3(n10214), .ZN(P1_U3246) );
  INV_X1 U11128 ( .A(n10217), .ZN(n10222) );
  INV_X1 U11129 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10220) );
  INV_X1 U11130 ( .A(n10218), .ZN(n10219) );
  OAI21_X1 U11131 ( .B1(n10808), .B2(n10220), .A(n10219), .ZN(n10221) );
  AOI21_X1 U11132 ( .B1(n10799), .B2(n10222), .A(n10221), .ZN(n10231) );
  OAI211_X1 U11133 ( .C1(n10225), .C2(n10224), .A(n10776), .B(n10223), .ZN(
        n10230) );
  OAI211_X1 U11134 ( .C1(n10228), .C2(n10227), .A(n10782), .B(n10226), .ZN(
        n10229) );
  NAND4_X1 U11135 ( .A1(n10232), .A2(n10231), .A3(n10230), .A4(n10229), .ZN(
        P1_U3247) );
  OAI211_X1 U11136 ( .C1(n10235), .C2(n10234), .A(n10776), .B(n10233), .ZN(
        n10245) );
  OAI211_X1 U11137 ( .C1(n10238), .C2(n10237), .A(n10782), .B(n10236), .ZN(
        n10244) );
  INV_X1 U11138 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10240) );
  OAI21_X1 U11139 ( .B1(n10808), .B2(n10240), .A(n10239), .ZN(n10241) );
  AOI21_X1 U11140 ( .B1(n10799), .B2(n10242), .A(n10241), .ZN(n10243) );
  NAND3_X1 U11141 ( .A1(n10245), .A2(n10244), .A3(n10243), .ZN(P1_U3248) );
  OAI211_X1 U11142 ( .C1(n10248), .C2(n10247), .A(n10776), .B(n10246), .ZN(
        n10257) );
  OAI211_X1 U11143 ( .C1(n10251), .C2(n10250), .A(n10782), .B(n10249), .ZN(
        n10256) );
  AOI21_X1 U11144 ( .B1(n10666), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n10252), .ZN(
        n10255) );
  NAND2_X1 U11145 ( .A1(n10799), .A2(n10253), .ZN(n10254) );
  NAND4_X1 U11146 ( .A1(n10257), .A2(n10256), .A3(n10255), .A4(n10254), .ZN(
        P1_U3249) );
  MUX2_X1 U11147 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n8156), .S(n10274), .Z(
        n10265) );
  AOI22_X1 U11148 ( .A1(n10260), .A2(n10259), .B1(n10258), .B2(n10267), .ZN(
        n10747) );
  AND2_X1 U11149 ( .A1(n10271), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n10262) );
  AOI21_X1 U11150 ( .B1(n10261), .B2(n10753), .A(n10262), .ZN(n10746) );
  NAND2_X1 U11151 ( .A1(n10747), .A2(n10746), .ZN(n10745) );
  INV_X1 U11152 ( .A(n10262), .ZN(n10263) );
  NAND2_X1 U11153 ( .A1(n10745), .A2(n10263), .ZN(n10264) );
  XOR2_X1 U11154 ( .A(n10265), .B(n10264), .Z(n10282) );
  OAI21_X1 U11155 ( .B1(n10808), .B2(n7276), .A(n10266), .ZN(n10279) );
  AOI22_X1 U11156 ( .A1(n10270), .A2(n10269), .B1(n10268), .B2(n10267), .ZN(
        n10750) );
  INV_X1 U11157 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n10530) );
  AND2_X1 U11158 ( .A1(n10271), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n10272) );
  AOI21_X1 U11159 ( .B1(n10530), .B2(n10753), .A(n10272), .ZN(n10749) );
  NAND2_X1 U11160 ( .A1(n10750), .A2(n10749), .ZN(n10748) );
  INV_X1 U11161 ( .A(n10272), .ZN(n10273) );
  NAND2_X1 U11162 ( .A1(n10748), .A2(n10273), .ZN(n10276) );
  XNOR2_X1 U11163 ( .A(n10274), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n10275) );
  XNOR2_X1 U11164 ( .A(n10276), .B(n10275), .ZN(n10277) );
  NOR2_X1 U11165 ( .A1(n10277), .A2(n10803), .ZN(n10278) );
  AOI211_X1 U11166 ( .C1(n10280), .C2(n10799), .A(n10279), .B(n10278), .ZN(
        n10281) );
  OAI21_X1 U11167 ( .B1(n10797), .B2(n10282), .A(n10281), .ZN(P1_U3262) );
  NOR2_X1 U11168 ( .A1(n10291), .A2(n10290), .ZN(n10284) );
  XNOR2_X1 U11169 ( .A(n10284), .B(n10283), .ZN(n10466) );
  NAND2_X1 U11170 ( .A1(n10466), .A2(n10285), .ZN(n10289) );
  AND2_X1 U11171 ( .A1(n10287), .A2(n10286), .ZN(n10465) );
  INV_X1 U11172 ( .A(n10465), .ZN(n10469) );
  NOR2_X1 U11173 ( .A1(n11051), .A2(n10469), .ZN(n10293) );
  AOI21_X1 U11174 ( .B1(n11051), .B2(P1_REG2_REG_31__SCAN_IN), .A(n10293), 
        .ZN(n10288) );
  OAI211_X1 U11175 ( .C1(n10547), .C2(n10440), .A(n10289), .B(n10288), .ZN(
        P1_U3263) );
  INV_X1 U11176 ( .A(n10291), .ZN(n10551) );
  NOR2_X1 U11177 ( .A1(n10551), .A2(n10440), .ZN(n10292) );
  AOI211_X1 U11178 ( .C1(n11051), .C2(P1_REG2_REG_30__SCAN_IN), .A(n10293), 
        .B(n10292), .ZN(n10294) );
  OAI21_X1 U11179 ( .B1(n10470), .B2(n10335), .A(n10294), .ZN(P1_U3264) );
  INV_X1 U11180 ( .A(n10295), .ZN(n10303) );
  NAND2_X1 U11181 ( .A1(n11051), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n10296) );
  OAI21_X1 U11182 ( .B1(n11050), .B2(n10297), .A(n10296), .ZN(n10298) );
  AOI21_X1 U11183 ( .B1(n10299), .B2(n11056), .A(n10298), .ZN(n10300) );
  OAI21_X1 U11184 ( .B1(n10301), .B2(n10335), .A(n10300), .ZN(n10302) );
  AOI21_X1 U11185 ( .B1(n10303), .B2(n10458), .A(n10302), .ZN(n10304) );
  OAI21_X1 U11186 ( .B1(n10305), .B2(n11051), .A(n10304), .ZN(P1_U3356) );
  OAI21_X1 U11187 ( .B1(n10308), .B2(n10307), .A(n10306), .ZN(n10312) );
  OAI22_X1 U11188 ( .A1(n10310), .A2(n10902), .B1(n10309), .B2(n10900), .ZN(
        n10311) );
  AOI21_X1 U11189 ( .B1(n10312), .B2(n10402), .A(n10311), .ZN(n10472) );
  OAI21_X1 U11190 ( .B1(n10315), .B2(n10314), .A(n10313), .ZN(n10473) );
  INV_X1 U11191 ( .A(n10473), .ZN(n10316) );
  NAND2_X1 U11192 ( .A1(n10316), .A2(n10458), .ZN(n10323) );
  OAI22_X1 U11193 ( .A1(n10915), .A2(n10318), .B1(n10317), .B2(n11050), .ZN(
        n10321) );
  INV_X1 U11194 ( .A(n10334), .ZN(n10319) );
  OAI211_X1 U11195 ( .C1(n10477), .C2(n10319), .A(n11035), .B(n5135), .ZN(
        n10471) );
  NOR2_X1 U11196 ( .A1(n10471), .A2(n10335), .ZN(n10320) );
  AOI211_X1 U11197 ( .C1(n11056), .C2(n10553), .A(n10321), .B(n10320), .ZN(
        n10322) );
  OAI211_X1 U11198 ( .C1(n11051), .C2(n10472), .A(n10323), .B(n10322), .ZN(
        P1_U3265) );
  XNOR2_X1 U11199 ( .A(n10324), .B(n10329), .ZN(n10328) );
  OAI22_X1 U11200 ( .A1(n10326), .A2(n10902), .B1(n10325), .B2(n10900), .ZN(
        n10327) );
  AOI21_X1 U11201 ( .B1(n10328), .B2(n10402), .A(n10327), .ZN(n10479) );
  XNOR2_X1 U11202 ( .A(n10330), .B(n10329), .ZN(n10480) );
  INV_X1 U11203 ( .A(n10480), .ZN(n10331) );
  NAND2_X1 U11204 ( .A1(n10331), .A2(n10458), .ZN(n10339) );
  OAI22_X1 U11205 ( .A1(n10915), .A2(n10333), .B1(n10332), .B2(n11050), .ZN(
        n10337) );
  OAI211_X1 U11206 ( .C1(n10484), .C2(n10348), .A(n11035), .B(n10334), .ZN(
        n10478) );
  NOR2_X1 U11207 ( .A1(n10478), .A2(n10335), .ZN(n10336) );
  AOI211_X1 U11208 ( .C1(n11056), .C2(n10556), .A(n10337), .B(n10336), .ZN(
        n10338) );
  OAI211_X1 U11209 ( .C1(n11051), .C2(n10479), .A(n10339), .B(n10338), .ZN(
        P1_U3266) );
  OAI21_X1 U11210 ( .B1(n10346), .B2(n10341), .A(n10340), .ZN(n10342) );
  NAND2_X1 U11211 ( .A1(n10342), .A2(n10402), .ZN(n10345) );
  AOI22_X1 U11212 ( .A1(n10343), .A2(n11026), .B1(n11027), .B2(n10375), .ZN(
        n10344) );
  NAND2_X1 U11213 ( .A1(n10345), .A2(n10344), .ZN(n10485) );
  INV_X1 U11214 ( .A(n10485), .ZN(n10357) );
  XNOR2_X1 U11215 ( .A(n10347), .B(n10346), .ZN(n10487) );
  NAND2_X1 U11216 ( .A1(n10487), .A2(n10458), .ZN(n10356) );
  INV_X1 U11217 ( .A(n10360), .ZN(n10349) );
  AOI211_X1 U11218 ( .C1(n10350), .C2(n10349), .A(n10438), .B(n10348), .ZN(
        n10486) );
  NOR2_X1 U11219 ( .A1(n10562), .A2(n10440), .ZN(n10354) );
  OAI22_X1 U11220 ( .A1(n10915), .A2(n10352), .B1(n10351), .B2(n11050), .ZN(
        n10353) );
  AOI211_X1 U11221 ( .C1(n10486), .C2(n11045), .A(n10354), .B(n10353), .ZN(
        n10355) );
  OAI211_X1 U11222 ( .C1(n11051), .C2(n10357), .A(n10356), .B(n10355), .ZN(
        P1_U3267) );
  XNOR2_X1 U11223 ( .A(n10359), .B(n10358), .ZN(n10494) );
  INV_X1 U11224 ( .A(n10381), .ZN(n10361) );
  AOI211_X1 U11225 ( .C1(n10491), .C2(n10361), .A(n10438), .B(n10360), .ZN(
        n10490) );
  INV_X1 U11226 ( .A(n10362), .ZN(n10363) );
  AOI22_X1 U11227 ( .A1(n11051), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n10363), 
        .B2(n10393), .ZN(n10364) );
  OAI21_X1 U11228 ( .B1(n10365), .B2(n10440), .A(n10364), .ZN(n10371) );
  OAI21_X1 U11229 ( .B1(n5140), .B2(n10367), .A(n10366), .ZN(n10369) );
  AOI222_X1 U11230 ( .A1(n10402), .A2(n10369), .B1(n10368), .B2(n11026), .C1(
        n10400), .C2(n11027), .ZN(n10493) );
  NOR2_X1 U11231 ( .A1(n10493), .A2(n11051), .ZN(n10370) );
  AOI211_X1 U11232 ( .C1(n10490), .C2(n11045), .A(n10371), .B(n10370), .ZN(
        n10372) );
  OAI21_X1 U11233 ( .B1(n10494), .B2(n10452), .A(n10372), .ZN(P1_U3268) );
  OAI211_X1 U11234 ( .C1(n10379), .C2(n10374), .A(n10373), .B(n10402), .ZN(
        n10378) );
  AOI22_X1 U11235 ( .A1(n11027), .A2(n10376), .B1(n10375), .B2(n11026), .ZN(
        n10377) );
  NAND2_X1 U11236 ( .A1(n10378), .A2(n10377), .ZN(n10495) );
  INV_X1 U11237 ( .A(n10495), .ZN(n10389) );
  XNOR2_X1 U11238 ( .A(n10380), .B(n10379), .ZN(n10497) );
  NAND2_X1 U11239 ( .A1(n10497), .A2(n10458), .ZN(n10388) );
  AOI211_X1 U11240 ( .C1(n10382), .C2(n10391), .A(n10438), .B(n10381), .ZN(
        n10496) );
  NOR2_X1 U11241 ( .A1(n10567), .A2(n10440), .ZN(n10386) );
  OAI22_X1 U11242 ( .A1(n10915), .A2(n10384), .B1(n10383), .B2(n11050), .ZN(
        n10385) );
  AOI211_X1 U11243 ( .C1(n10496), .C2(n11045), .A(n10386), .B(n10385), .ZN(
        n10387) );
  OAI211_X1 U11244 ( .C1(n11051), .C2(n10389), .A(n10388), .B(n10387), .ZN(
        P1_U3269) );
  XNOR2_X1 U11245 ( .A(n10390), .B(n10398), .ZN(n10504) );
  AOI211_X1 U11246 ( .C1(n10501), .C2(n10407), .A(n10438), .B(n6213), .ZN(
        n10500) );
  INV_X1 U11247 ( .A(n10392), .ZN(n10394) );
  AOI22_X1 U11248 ( .A1(n11051), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n10394), 
        .B2(n10393), .ZN(n10395) );
  OAI21_X1 U11249 ( .B1(n10396), .B2(n10440), .A(n10395), .ZN(n10404) );
  XNOR2_X1 U11250 ( .A(n10398), .B(n10397), .ZN(n10401) );
  AOI222_X1 U11251 ( .A1(n10402), .A2(n10401), .B1(n10400), .B2(n11026), .C1(
        n10399), .C2(n11027), .ZN(n10503) );
  NOR2_X1 U11252 ( .A1(n10503), .A2(n11051), .ZN(n10403) );
  AOI211_X1 U11253 ( .C1(n10500), .C2(n11045), .A(n10404), .B(n10403), .ZN(
        n10405) );
  OAI21_X1 U11254 ( .B1(n10504), .B2(n10452), .A(n10405), .ZN(P1_U3270) );
  XOR2_X1 U11255 ( .A(n10406), .B(n10415), .Z(n10509) );
  INV_X1 U11256 ( .A(n10420), .ZN(n10408) );
  AOI211_X1 U11257 ( .C1(n10507), .C2(n10408), .A(n10438), .B(n5315), .ZN(
        n10506) );
  NOR2_X1 U11258 ( .A1(n10409), .A2(n10440), .ZN(n10413) );
  OAI22_X1 U11259 ( .A1(n10915), .A2(n10411), .B1(n10410), .B2(n11050), .ZN(
        n10412) );
  AOI211_X1 U11260 ( .C1(n10506), .C2(n11045), .A(n10413), .B(n10412), .ZN(
        n10419) );
  XOR2_X1 U11261 ( .A(n10415), .B(n10414), .Z(n10416) );
  OAI222_X1 U11262 ( .A1(n10902), .A2(n10417), .B1(n10900), .B2(n10449), .C1(
        n10416), .C2(n11030), .ZN(n10505) );
  NAND2_X1 U11263 ( .A1(n10505), .A2(n10915), .ZN(n10418) );
  OAI211_X1 U11264 ( .C1(n10509), .C2(n10452), .A(n10419), .B(n10418), .ZN(
        P1_U3271) );
  INV_X1 U11265 ( .A(n10437), .ZN(n10421) );
  AOI211_X1 U11266 ( .C1(n10432), .C2(n10421), .A(n10438), .B(n10420), .ZN(
        n10511) );
  AOI21_X1 U11267 ( .B1(n10446), .B2(n10445), .A(n10422), .ZN(n10423) );
  XNOR2_X1 U11268 ( .A(n5528), .B(n10423), .ZN(n10424) );
  OAI222_X1 U11269 ( .A1(n10900), .A2(n10426), .B1(n10902), .B2(n10425), .C1(
        n10424), .C2(n11030), .ZN(n10510) );
  AOI21_X1 U11270 ( .B1(n10511), .B2(n10274), .A(n10510), .ZN(n10435) );
  XNOR2_X1 U11271 ( .A(n10427), .B(n10428), .ZN(n10512) );
  NAND2_X1 U11272 ( .A1(n10512), .A2(n10458), .ZN(n10434) );
  OAI22_X1 U11273 ( .A1(n10915), .A2(n10430), .B1(n10429), .B2(n11050), .ZN(
        n10431) );
  AOI21_X1 U11274 ( .B1(n10432), .B2(n11056), .A(n10431), .ZN(n10433) );
  OAI211_X1 U11275 ( .C1(n11051), .C2(n10435), .A(n10434), .B(n10433), .ZN(
        P1_U3272) );
  XOR2_X1 U11276 ( .A(n10446), .B(n10436), .Z(n10519) );
  AOI211_X1 U11277 ( .C1(n10517), .C2(n10439), .A(n10438), .B(n10437), .ZN(
        n10516) );
  NOR2_X1 U11278 ( .A1(n5318), .A2(n10440), .ZN(n10444) );
  OAI22_X1 U11279 ( .A1(n10915), .A2(n10442), .B1(n10441), .B2(n11050), .ZN(
        n10443) );
  AOI211_X1 U11280 ( .C1(n10516), .C2(n11045), .A(n10444), .B(n10443), .ZN(
        n10451) );
  XOR2_X1 U11281 ( .A(n10446), .B(n10445), .Z(n10447) );
  OAI222_X1 U11282 ( .A1(n10902), .A2(n10449), .B1(n10900), .B2(n10448), .C1(
        n10447), .C2(n11030), .ZN(n10515) );
  NAND2_X1 U11283 ( .A1(n10515), .A2(n10915), .ZN(n10450) );
  OAI211_X1 U11284 ( .C1(n10519), .C2(n10452), .A(n10451), .B(n10450), .ZN(
        P1_U3273) );
  NAND2_X1 U11285 ( .A1(n10453), .A2(n10915), .ZN(n10464) );
  NAND2_X1 U11286 ( .A1(n11051), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10454) );
  OAI21_X1 U11287 ( .B1(n11050), .B2(n10455), .A(n10454), .ZN(n10456) );
  AOI21_X1 U11288 ( .B1(n11056), .B2(n10457), .A(n10456), .ZN(n10463) );
  NAND2_X1 U11289 ( .A1(n10459), .A2(n10458), .ZN(n10462) );
  NAND2_X1 U11290 ( .A1(n10460), .A2(n11045), .ZN(n10461) );
  NAND4_X1 U11291 ( .A1(n10464), .A2(n10463), .A3(n10462), .A4(n10461), .ZN(
        P1_U3284) );
  INV_X1 U11292 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n10467) );
  AOI21_X1 U11293 ( .B1(n10466), .B2(n11035), .A(n10465), .ZN(n10545) );
  MUX2_X1 U11294 ( .A(n10467), .B(n10545), .S(n11081), .Z(n10468) );
  OAI21_X1 U11295 ( .B1(n10547), .B2(n10532), .A(n10468), .ZN(P1_U3553) );
  INV_X1 U11296 ( .A(n10552), .ZN(n10474) );
  OAI21_X1 U11297 ( .B1(n10477), .B2(n10532), .A(n10476), .ZN(P1_U3550) );
  OAI211_X1 U11298 ( .C1(n10480), .C2(n10543), .A(n10479), .B(n10478), .ZN(
        n10554) );
  INV_X1 U11299 ( .A(n10554), .ZN(n10481) );
  MUX2_X1 U11300 ( .A(n10482), .B(n10481), .S(n10529), .Z(n10483) );
  OAI21_X1 U11301 ( .B1(n10484), .B2(n10532), .A(n10483), .ZN(P1_U3549) );
  AOI211_X1 U11302 ( .C1(n10487), .C2(n11078), .A(n10486), .B(n10485), .ZN(
        n10559) );
  MUX2_X1 U11303 ( .A(n10488), .B(n10559), .S(n10529), .Z(n10489) );
  OAI21_X1 U11304 ( .B1(n10562), .B2(n10532), .A(n10489), .ZN(P1_U3548) );
  AOI21_X1 U11305 ( .B1(n10541), .B2(n10491), .A(n10490), .ZN(n10492) );
  OAI211_X1 U11306 ( .C1(n10494), .C2(n10543), .A(n10493), .B(n10492), .ZN(
        n10563) );
  MUX2_X1 U11307 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10563), .S(n11081), .Z(
        P1_U3547) );
  AOI211_X1 U11308 ( .C1(n10497), .C2(n11078), .A(n10496), .B(n10495), .ZN(
        n10564) );
  MUX2_X1 U11309 ( .A(n10498), .B(n10564), .S(n10529), .Z(n10499) );
  OAI21_X1 U11310 ( .B1(n10567), .B2(n10532), .A(n10499), .ZN(P1_U3546) );
  AOI21_X1 U11311 ( .B1(n10541), .B2(n10501), .A(n10500), .ZN(n10502) );
  OAI211_X1 U11312 ( .C1(n10504), .C2(n10543), .A(n10503), .B(n10502), .ZN(
        n10568) );
  MUX2_X1 U11313 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10568), .S(n10529), .Z(
        P1_U3545) );
  AOI211_X1 U11314 ( .C1(n10541), .C2(n10507), .A(n10506), .B(n10505), .ZN(
        n10508) );
  OAI21_X1 U11315 ( .B1(n10509), .B2(n10543), .A(n10508), .ZN(n10569) );
  MUX2_X1 U11316 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10569), .S(n10529), .Z(
        P1_U3544) );
  AOI211_X1 U11317 ( .C1(n10512), .C2(n11078), .A(n10511), .B(n10510), .ZN(
        n10570) );
  MUX2_X1 U11318 ( .A(n10513), .B(n10570), .S(n10529), .Z(n10514) );
  OAI21_X1 U11319 ( .B1(n10573), .B2(n10532), .A(n10514), .ZN(P1_U3543) );
  AOI211_X1 U11320 ( .C1(n10541), .C2(n10517), .A(n10516), .B(n10515), .ZN(
        n10518) );
  OAI21_X1 U11321 ( .B1(n10519), .B2(n10543), .A(n10518), .ZN(n10574) );
  MUX2_X1 U11322 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10574), .S(n11081), .Z(
        P1_U3542) );
  AOI211_X1 U11323 ( .C1(n10541), .C2(n10522), .A(n10521), .B(n10520), .ZN(
        n10523) );
  OAI21_X1 U11324 ( .B1(n10524), .B2(n10543), .A(n10523), .ZN(n10575) );
  MUX2_X1 U11325 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10575), .S(n11081), .Z(
        P1_U3541) );
  NAND2_X1 U11326 ( .A1(n10526), .A2(n10525), .ZN(n10527) );
  AOI21_X1 U11327 ( .B1(n10528), .B2(n11078), .A(n10527), .ZN(n10576) );
  MUX2_X1 U11328 ( .A(n10530), .B(n10576), .S(n10529), .Z(n10531) );
  OAI21_X1 U11329 ( .B1(n10580), .B2(n10532), .A(n10531), .ZN(P1_U3540) );
  AOI211_X1 U11330 ( .C1(n10541), .C2(n10535), .A(n10534), .B(n10533), .ZN(
        n10536) );
  OAI21_X1 U11331 ( .B1(n10537), .B2(n10543), .A(n10536), .ZN(n10581) );
  MUX2_X1 U11332 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10581), .S(n11081), .Z(
        P1_U3539) );
  AOI211_X1 U11333 ( .C1(n10541), .C2(n10540), .A(n10539), .B(n10538), .ZN(
        n10542) );
  OAI21_X1 U11334 ( .B1(n10544), .B2(n10543), .A(n10542), .ZN(n10582) );
  MUX2_X1 U11335 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n10582), .S(n11081), .Z(
        P1_U3537) );
  MUX2_X1 U11336 ( .A(n9888), .B(n10545), .S(n11085), .Z(n10546) );
  OAI21_X1 U11337 ( .B1(n10547), .B2(n10579), .A(n10546), .ZN(P1_U3521) );
  INV_X1 U11338 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10548) );
  MUX2_X1 U11339 ( .A(n10549), .B(n10548), .S(n11082), .Z(n10550) );
  OAI21_X1 U11340 ( .B1(n10551), .B2(n10579), .A(n10550), .ZN(P1_U3520) );
  MUX2_X1 U11341 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10554), .S(n11085), .Z(
        n10555) );
  AOI21_X1 U11342 ( .B1(n10557), .B2(n10556), .A(n10555), .ZN(n10558) );
  INV_X1 U11343 ( .A(n10558), .ZN(P1_U3517) );
  INV_X1 U11344 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n10560) );
  MUX2_X1 U11345 ( .A(n10560), .B(n10559), .S(n11085), .Z(n10561) );
  OAI21_X1 U11346 ( .B1(n10562), .B2(n10579), .A(n10561), .ZN(P1_U3516) );
  MUX2_X1 U11347 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10563), .S(n11085), .Z(
        P1_U3515) );
  INV_X1 U11348 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n10565) );
  MUX2_X1 U11349 ( .A(n10565), .B(n10564), .S(n11085), .Z(n10566) );
  OAI21_X1 U11350 ( .B1(n10567), .B2(n10579), .A(n10566), .ZN(P1_U3514) );
  MUX2_X1 U11351 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10568), .S(n11085), .Z(
        P1_U3513) );
  MUX2_X1 U11352 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10569), .S(n11085), .Z(
        P1_U3512) );
  INV_X1 U11353 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n10571) );
  MUX2_X1 U11354 ( .A(n10571), .B(n10570), .S(n11085), .Z(n10572) );
  OAI21_X1 U11355 ( .B1(n10573), .B2(n10579), .A(n10572), .ZN(P1_U3511) );
  MUX2_X1 U11356 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10574), .S(n11085), .Z(
        P1_U3510) );
  MUX2_X1 U11357 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10575), .S(n11085), .Z(
        P1_U3509) );
  INV_X1 U11358 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10577) );
  MUX2_X1 U11359 ( .A(n10577), .B(n10576), .S(n11085), .Z(n10578) );
  OAI21_X1 U11360 ( .B1(n10580), .B2(n10579), .A(n10578), .ZN(P1_U3507) );
  MUX2_X1 U11361 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10581), .S(n11085), .Z(
        P1_U3504) );
  MUX2_X1 U11362 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n10582), .S(n11085), .Z(
        P1_U3498) );
  AND2_X1 U11363 ( .A1(n10584), .A2(n10583), .ZN(n10602) );
  MUX2_X1 U11364 ( .A(P1_D_REG_1__SCAN_IN), .B(n10585), .S(n10602), .Z(
        P1_U3440) );
  MUX2_X1 U11365 ( .A(P1_D_REG_0__SCAN_IN), .B(n10586), .S(n10602), .Z(
        P1_U3439) );
  NAND3_X1 U11366 ( .A1(n10588), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n10590) );
  OAI22_X1 U11367 ( .A1(n10587), .A2(n10590), .B1(n10589), .B2(n10595), .ZN(
        n10591) );
  AOI21_X1 U11368 ( .B1(n10593), .B2(n10592), .A(n10591), .ZN(n10594) );
  INV_X1 U11369 ( .A(n10594), .ZN(P1_U3324) );
  OAI222_X1 U11370 ( .A1(P1_U3086), .A2(n10598), .B1(n8657), .B2(n10597), .C1(
        n10596), .C2(n10595), .ZN(P1_U3326) );
  MUX2_X1 U11371 ( .A(n10599), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  NOR2_X1 U11372 ( .A1(n10602), .A2(n10600), .ZN(P1_U3323) );
  AND2_X1 U11373 ( .A1(n10603), .A2(P1_D_REG_3__SCAN_IN), .ZN(P1_U3322) );
  INV_X1 U11374 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10601) );
  NOR2_X1 U11375 ( .A1(n10602), .A2(n10601), .ZN(P1_U3321) );
  AND2_X1 U11376 ( .A1(n10603), .A2(P1_D_REG_5__SCAN_IN), .ZN(P1_U3320) );
  AND2_X1 U11377 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10603), .ZN(P1_U3319) );
  AND2_X1 U11378 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10603), .ZN(P1_U3318) );
  AND2_X1 U11379 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10603), .ZN(P1_U3317) );
  AND2_X1 U11380 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10603), .ZN(P1_U3316) );
  AND2_X1 U11381 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10603), .ZN(P1_U3315) );
  AND2_X1 U11382 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10603), .ZN(P1_U3314) );
  AND2_X1 U11383 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10603), .ZN(P1_U3313) );
  AND2_X1 U11384 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10603), .ZN(P1_U3312) );
  AND2_X1 U11385 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10603), .ZN(P1_U3311) );
  AND2_X1 U11386 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10603), .ZN(P1_U3310) );
  AND2_X1 U11387 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10603), .ZN(P1_U3309) );
  AND2_X1 U11388 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10603), .ZN(P1_U3308) );
  AND2_X1 U11389 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10603), .ZN(P1_U3307) );
  AND2_X1 U11390 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10603), .ZN(P1_U3306) );
  AND2_X1 U11391 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10603), .ZN(P1_U3305) );
  AND2_X1 U11392 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10603), .ZN(P1_U3304) );
  AND2_X1 U11393 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10603), .ZN(P1_U3303) );
  AND2_X1 U11394 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10603), .ZN(P1_U3302) );
  AND2_X1 U11395 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10603), .ZN(P1_U3301) );
  AND2_X1 U11396 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10603), .ZN(P1_U3300) );
  AND2_X1 U11397 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10603), .ZN(P1_U3299) );
  AND2_X1 U11398 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10603), .ZN(P1_U3298) );
  AND2_X1 U11399 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10603), .ZN(P1_U3297) );
  AND2_X1 U11400 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10603), .ZN(P1_U3296) );
  AND2_X1 U11401 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10603), .ZN(P1_U3295) );
  AND2_X1 U11402 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10603), .ZN(P1_U3294) );
  XOR2_X1 U11403 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  OAI222_X1 U11404 ( .A1(n10608), .A2(n10607), .B1(n10608), .B2(n10606), .C1(
        n10605), .C2(n10604), .ZN(ADD_1068_U5) );
  AOI21_X1 U11405 ( .B1(n10611), .B2(n10610), .A(n10609), .ZN(ADD_1068_U54) );
  AOI21_X1 U11406 ( .B1(n10614), .B2(n10613), .A(n10612), .ZN(ADD_1068_U53) );
  OAI21_X1 U11407 ( .B1(n10617), .B2(n10616), .A(n10615), .ZN(ADD_1068_U52) );
  OAI21_X1 U11408 ( .B1(n10620), .B2(n10619), .A(n10618), .ZN(ADD_1068_U51) );
  OAI21_X1 U11409 ( .B1(n10623), .B2(n10622), .A(n10621), .ZN(ADD_1068_U50) );
  OAI21_X1 U11410 ( .B1(n10626), .B2(n10625), .A(n10624), .ZN(ADD_1068_U49) );
  OAI21_X1 U11411 ( .B1(n10629), .B2(n10628), .A(n10627), .ZN(ADD_1068_U48) );
  OAI21_X1 U11412 ( .B1(n10632), .B2(n10631), .A(n10630), .ZN(ADD_1068_U47) );
  OAI21_X1 U11413 ( .B1(n10635), .B2(n10634), .A(n10633), .ZN(ADD_1068_U63) );
  OAI21_X1 U11414 ( .B1(n10638), .B2(n10637), .A(n10636), .ZN(ADD_1068_U62) );
  OAI21_X1 U11415 ( .B1(n10641), .B2(n10640), .A(n10639), .ZN(ADD_1068_U61) );
  OAI21_X1 U11416 ( .B1(n10644), .B2(n10643), .A(n10642), .ZN(ADD_1068_U60) );
  OAI21_X1 U11417 ( .B1(n10647), .B2(n10646), .A(n10645), .ZN(ADD_1068_U59) );
  OAI21_X1 U11418 ( .B1(n10650), .B2(n10649), .A(n10648), .ZN(ADD_1068_U58) );
  OAI21_X1 U11419 ( .B1(n10653), .B2(n10652), .A(n10651), .ZN(ADD_1068_U57) );
  OAI21_X1 U11420 ( .B1(n10656), .B2(n10655), .A(n10654), .ZN(ADD_1068_U56) );
  OAI21_X1 U11421 ( .B1(n10659), .B2(n10658), .A(n10657), .ZN(ADD_1068_U55) );
  NAND2_X1 U11422 ( .A1(n10660), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10661) );
  OAI21_X1 U11423 ( .B1(n10663), .B2(n10662), .A(n10661), .ZN(n10664) );
  XNOR2_X1 U11424 ( .A(n10664), .B(P1_IR_REG_0__SCAN_IN), .ZN(n10668) );
  AOI22_X1 U11425 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n10666), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n10667) );
  OAI21_X1 U11426 ( .B1(n10669), .B2(n10668), .A(n10667), .ZN(P1_U3243) );
  INV_X1 U11427 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10685) );
  OAI21_X1 U11428 ( .B1(n10672), .B2(n10671), .A(n10670), .ZN(n10681) );
  NOR2_X1 U11429 ( .A1(n10674), .A2(n10673), .ZN(n10675) );
  OR2_X1 U11430 ( .A1(n10676), .A2(n10675), .ZN(n10677) );
  OR2_X1 U11431 ( .A1(n10797), .A2(n10677), .ZN(n10680) );
  NAND2_X1 U11432 ( .A1(n10799), .A2(n10678), .ZN(n10679) );
  OAI211_X1 U11433 ( .C1(n10803), .C2(n10681), .A(n10680), .B(n10679), .ZN(
        n10682) );
  INV_X1 U11434 ( .A(n10682), .ZN(n10684) );
  OAI211_X1 U11435 ( .C1(n10808), .C2(n10685), .A(n10684), .B(n10683), .ZN(
        P1_U3250) );
  INV_X1 U11436 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10699) );
  OAI21_X1 U11437 ( .B1(n10688), .B2(n10687), .A(n10686), .ZN(n10695) );
  OAI211_X1 U11438 ( .C1(n10691), .C2(n10690), .A(n10782), .B(n10689), .ZN(
        n10694) );
  NAND2_X1 U11439 ( .A1(n10799), .A2(n10692), .ZN(n10693) );
  OAI211_X1 U11440 ( .C1(n10797), .C2(n10695), .A(n10694), .B(n10693), .ZN(
        n10696) );
  INV_X1 U11441 ( .A(n10696), .ZN(n10698) );
  OAI211_X1 U11442 ( .C1(n10808), .C2(n10699), .A(n10698), .B(n10697), .ZN(
        P1_U3251) );
  INV_X1 U11443 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10716) );
  NAND2_X1 U11444 ( .A1(n10701), .A2(n10700), .ZN(n10704) );
  INV_X1 U11445 ( .A(n10702), .ZN(n10703) );
  NAND2_X1 U11446 ( .A1(n10704), .A2(n10703), .ZN(n10712) );
  AOI21_X1 U11447 ( .B1(n10707), .B2(n10706), .A(n10705), .ZN(n10708) );
  NAND2_X1 U11448 ( .A1(n10782), .A2(n10708), .ZN(n10711) );
  NAND2_X1 U11449 ( .A1(n10799), .A2(n10709), .ZN(n10710) );
  OAI211_X1 U11450 ( .C1(n10712), .C2(n10797), .A(n10711), .B(n10710), .ZN(
        n10713) );
  INV_X1 U11451 ( .A(n10713), .ZN(n10715) );
  OAI211_X1 U11452 ( .C1(n10808), .C2(n10716), .A(n10715), .B(n10714), .ZN(
        P1_U3254) );
  INV_X1 U11453 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10733) );
  NAND2_X1 U11454 ( .A1(n10718), .A2(n10717), .ZN(n10721) );
  INV_X1 U11455 ( .A(n10719), .ZN(n10720) );
  NAND2_X1 U11456 ( .A1(n10721), .A2(n10720), .ZN(n10729) );
  AOI21_X1 U11457 ( .B1(n10724), .B2(n10723), .A(n10722), .ZN(n10725) );
  NAND2_X1 U11458 ( .A1(n10782), .A2(n10725), .ZN(n10728) );
  NAND2_X1 U11459 ( .A1(n10799), .A2(n10726), .ZN(n10727) );
  OAI211_X1 U11460 ( .C1(n10729), .C2(n10797), .A(n10728), .B(n10727), .ZN(
        n10730) );
  INV_X1 U11461 ( .A(n10730), .ZN(n10732) );
  OAI211_X1 U11462 ( .C1(n10808), .C2(n10733), .A(n10732), .B(n10731), .ZN(
        P1_U3257) );
  INV_X1 U11463 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10744) );
  AOI211_X1 U11464 ( .C1(n10736), .C2(n10735), .A(n10734), .B(n10803), .ZN(
        n10740) );
  AOI211_X1 U11465 ( .C1(n10738), .C2(n5943), .A(n10737), .B(n10797), .ZN(
        n10739) );
  AOI211_X1 U11466 ( .C1(n10799), .C2(n10741), .A(n10740), .B(n10739), .ZN(
        n10743) );
  OAI211_X1 U11467 ( .C1(n10808), .C2(n10744), .A(n10743), .B(n10742), .ZN(
        P1_U3258) );
  INV_X1 U11468 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10758) );
  OAI211_X1 U11469 ( .C1(n10747), .C2(n10746), .A(n10745), .B(n10776), .ZN(
        n10752) );
  OAI211_X1 U11470 ( .C1(n10750), .C2(n10749), .A(n10748), .B(n10782), .ZN(
        n10751) );
  OAI211_X1 U11471 ( .C1(n10754), .C2(n10753), .A(n10752), .B(n10751), .ZN(
        n10755) );
  INV_X1 U11472 ( .A(n10755), .ZN(n10757) );
  OAI211_X1 U11473 ( .C1(n10808), .C2(n10758), .A(n10757), .B(n10756), .ZN(
        P1_U3261) );
  INV_X1 U11474 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10770) );
  AOI211_X1 U11475 ( .C1(n10761), .C2(n10760), .A(n10759), .B(n10803), .ZN(
        n10766) );
  AOI211_X1 U11476 ( .C1(n10764), .C2(n10763), .A(n10762), .B(n10797), .ZN(
        n10765) );
  AOI211_X1 U11477 ( .C1(n10799), .C2(n10767), .A(n10766), .B(n10765), .ZN(
        n10769) );
  OAI211_X1 U11478 ( .C1(n10808), .C2(n10770), .A(n10769), .B(n10768), .ZN(
        P1_U3256) );
  INV_X1 U11479 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10787) );
  AOI21_X1 U11480 ( .B1(n10773), .B2(n10772), .A(n10771), .ZN(n10775) );
  AOI22_X1 U11481 ( .A1(n10776), .A2(n10775), .B1(n10774), .B2(n10799), .ZN(
        n10784) );
  NAND2_X1 U11482 ( .A1(n10778), .A2(n10777), .ZN(n10781) );
  INV_X1 U11483 ( .A(n10779), .ZN(n10780) );
  NAND3_X1 U11484 ( .A1(n10782), .A2(n10781), .A3(n10780), .ZN(n10783) );
  AND2_X1 U11485 ( .A1(n10784), .A2(n10783), .ZN(n10786) );
  OAI211_X1 U11486 ( .C1(n10808), .C2(n10787), .A(n10786), .B(n10785), .ZN(
        P1_U3253) );
  INV_X1 U11487 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10807) );
  NAND2_X1 U11488 ( .A1(n10789), .A2(n10788), .ZN(n10790) );
  AND2_X1 U11489 ( .A1(n10791), .A2(n10790), .ZN(n10802) );
  OR2_X1 U11490 ( .A1(n10793), .A2(n10792), .ZN(n10795) );
  AND2_X1 U11491 ( .A1(n10795), .A2(n10794), .ZN(n10796) );
  OR2_X1 U11492 ( .A1(n10797), .A2(n10796), .ZN(n10801) );
  NAND2_X1 U11493 ( .A1(n10799), .A2(n10798), .ZN(n10800) );
  OAI211_X1 U11494 ( .C1(n10803), .C2(n10802), .A(n10801), .B(n10800), .ZN(
        n10804) );
  INV_X1 U11495 ( .A(n10804), .ZN(n10806) );
  OAI211_X1 U11496 ( .C1(n10808), .C2(n10807), .A(n10806), .B(n10805), .ZN(
        P1_U3252) );
  INV_X1 U11497 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10827) );
  AOI21_X1 U11498 ( .B1(n10810), .B2(n6326), .A(n10809), .ZN(n10818) );
  OAI21_X1 U11499 ( .B1(P2_REG1_REG_3__SCAN_IN), .B2(n10812), .A(n10811), .ZN(
        n10814) );
  AOI21_X1 U11500 ( .B1(n10849), .B2(n10814), .A(n10813), .ZN(n10817) );
  NAND2_X1 U11501 ( .A1(n10848), .A2(n10815), .ZN(n10816) );
  OAI211_X1 U11502 ( .C1(n10818), .C2(n10854), .A(n10817), .B(n10816), .ZN(
        n10819) );
  INV_X1 U11503 ( .A(n10819), .ZN(n10826) );
  AOI21_X1 U11504 ( .B1(n10822), .B2(n10821), .A(n10820), .ZN(n10824) );
  OR2_X1 U11505 ( .A1(n10824), .A2(n10823), .ZN(n10825) );
  OAI211_X1 U11506 ( .C1(n10827), .C2(n10843), .A(n10826), .B(n10825), .ZN(
        P2_U3185) );
  INV_X1 U11507 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10844) );
  XOR2_X1 U11508 ( .A(n10829), .B(n10828), .Z(n10834) );
  AOI21_X1 U11509 ( .B1(n5126), .B2(n10831), .A(n10830), .ZN(n10832) );
  OAI22_X1 U11510 ( .A1(n10834), .A2(n10833), .B1(n10854), .B2(n10832), .ZN(
        n10835) );
  AOI211_X1 U11511 ( .C1(n10837), .C2(n10848), .A(n10836), .B(n10835), .ZN(
        n10842) );
  OAI211_X1 U11512 ( .C1(n10840), .C2(n10839), .A(n10838), .B(n10859), .ZN(
        n10841) );
  OAI211_X1 U11513 ( .C1(n10844), .C2(n10843), .A(n10842), .B(n10841), .ZN(
        P2_U3186) );
  OAI21_X1 U11514 ( .B1(P2_REG1_REG_5__SCAN_IN), .B2(n10846), .A(n10845), .ZN(
        n10850) );
  AOI22_X1 U11515 ( .A1(n10850), .A2(n10849), .B1(n10848), .B2(n10847), .ZN(
        n10865) );
  INV_X1 U11516 ( .A(n10851), .ZN(n10857) );
  AOI21_X1 U11517 ( .B1(n10853), .B2(n7513), .A(n10852), .ZN(n10855) );
  NOR2_X1 U11518 ( .A1(n10855), .A2(n10854), .ZN(n10856) );
  AOI211_X1 U11519 ( .C1(n10858), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n10857), .B(
        n10856), .ZN(n10864) );
  OAI211_X1 U11520 ( .C1(n10862), .C2(n10861), .A(n10860), .B(n10859), .ZN(
        n10863) );
  NAND3_X1 U11521 ( .A1(n10865), .A2(n10864), .A3(n10863), .ZN(P2_U3187) );
  XNOR2_X1 U11522 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U11523 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10866) );
  AOI22_X1 U11524 ( .A1(n11085), .A2(n10867), .B1(n10866), .B2(n11082), .ZN(
        P1_U3453) );
  INV_X1 U11525 ( .A(n10868), .ZN(n10872) );
  OAI22_X1 U11526 ( .A1(n10870), .A2(n11012), .B1(n10869), .B2(n11093), .ZN(
        n10871) );
  NOR2_X1 U11527 ( .A1(n10872), .A2(n10871), .ZN(n10874) );
  AOI22_X1 U11528 ( .A1(n11100), .A2(n10874), .B1(n6853), .B2(n11099), .ZN(
        P2_U3460) );
  INV_X1 U11529 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10873) );
  AOI22_X1 U11530 ( .A1(n11104), .A2(n10874), .B1(n10873), .B2(n11101), .ZN(
        P2_U3393) );
  INV_X1 U11531 ( .A(n10875), .ZN(n10880) );
  OAI21_X1 U11532 ( .B1(n5729), .B2(n11074), .A(n10876), .ZN(n10879) );
  INV_X1 U11533 ( .A(n10877), .ZN(n10878) );
  AOI211_X1 U11534 ( .C1(n11039), .C2(n10880), .A(n10879), .B(n10878), .ZN(
        n10882) );
  AOI22_X1 U11535 ( .A1(n11081), .A2(n10882), .B1(n10881), .B2(n11080), .ZN(
        P1_U3523) );
  AOI22_X1 U11536 ( .A1(n11085), .A2(n10882), .B1(n5713), .B2(n11082), .ZN(
        P1_U3456) );
  OAI21_X1 U11537 ( .B1(n10884), .B2(n11074), .A(n10883), .ZN(n10887) );
  INV_X1 U11538 ( .A(n10885), .ZN(n10886) );
  AOI211_X1 U11539 ( .C1(n11039), .C2(n10888), .A(n10887), .B(n10886), .ZN(
        n10890) );
  AOI22_X1 U11540 ( .A1(n11081), .A2(n10890), .B1(n10889), .B2(n11080), .ZN(
        P1_U3524) );
  AOI22_X1 U11541 ( .A1(n11085), .A2(n10890), .B1(n5732), .B2(n11082), .ZN(
        P1_U3459) );
  AOI211_X1 U11542 ( .C1(n11097), .C2(n10893), .A(n10892), .B(n10891), .ZN(
        n10895) );
  AOI22_X1 U11543 ( .A1(n11100), .A2(n10895), .B1(n7341), .B2(n11099), .ZN(
        P2_U3461) );
  INV_X1 U11544 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10894) );
  AOI22_X1 U11545 ( .A1(n11104), .A2(n10895), .B1(n10894), .B2(n11101), .ZN(
        P2_U3396) );
  XNOR2_X1 U11546 ( .A(n10896), .B(n10903), .ZN(n10920) );
  OAI211_X1 U11547 ( .C1(n10898), .C2(n10899), .A(n11035), .B(n10897), .ZN(
        n10918) );
  OAI21_X1 U11548 ( .B1(n10899), .B2(n11074), .A(n10918), .ZN(n10911) );
  OAI22_X1 U11549 ( .A1(n5245), .A2(n10902), .B1(n10901), .B2(n10900), .ZN(
        n10909) );
  NAND3_X1 U11550 ( .A1(n10905), .A2(n10904), .A3(n10903), .ZN(n10906) );
  AOI21_X1 U11551 ( .B1(n10907), .B2(n10906), .A(n11030), .ZN(n10908) );
  AOI211_X1 U11552 ( .C1(n11033), .C2(n10920), .A(n10909), .B(n10908), .ZN(
        n10923) );
  INV_X1 U11553 ( .A(n10923), .ZN(n10910) );
  AOI211_X1 U11554 ( .C1(n11039), .C2(n10920), .A(n10911), .B(n10910), .ZN(
        n10913) );
  INV_X1 U11555 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10912) );
  AOI22_X1 U11556 ( .A1(n11081), .A2(n10913), .B1(n10912), .B2(n11080), .ZN(
        P1_U3525) );
  AOI22_X1 U11557 ( .A1(n11085), .A2(n10913), .B1(n5746), .B2(n11082), .ZN(
        P1_U3462) );
  OAI22_X1 U11558 ( .A1(n10915), .A2(n10914), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n11050), .ZN(n10916) );
  AOI21_X1 U11559 ( .B1(n11056), .B2(n10917), .A(n10916), .ZN(n10922) );
  INV_X1 U11560 ( .A(n10918), .ZN(n10919) );
  AOI22_X1 U11561 ( .A1(n11046), .A2(n10920), .B1(n11045), .B2(n10919), .ZN(
        n10921) );
  OAI211_X1 U11562 ( .C1(n11051), .C2(n10923), .A(n10922), .B(n10921), .ZN(
        P1_U3290) );
  XNOR2_X1 U11563 ( .A(n10924), .B(n8855), .ZN(n10927) );
  AOI222_X1 U11564 ( .A1(n10928), .A2(n10927), .B1(n7154), .B2(n10926), .C1(
        n10925), .C2(n6677), .ZN(n10945) );
  NAND2_X1 U11565 ( .A1(n10930), .A2(n10929), .ZN(n10931) );
  XNOR2_X1 U11566 ( .A(n10932), .B(n10931), .ZN(n10942) );
  AOI22_X1 U11567 ( .A1(n10942), .A2(n11097), .B1(n11017), .B2(n10933), .ZN(
        n10934) );
  AND2_X1 U11568 ( .A1(n10945), .A2(n10934), .ZN(n10936) );
  AOI22_X1 U11569 ( .A1(n11100), .A2(n10936), .B1(n6327), .B2(n11099), .ZN(
        P2_U3462) );
  INV_X1 U11570 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10935) );
  AOI22_X1 U11571 ( .A1(n11104), .A2(n10936), .B1(n10935), .B2(n11101), .ZN(
        P2_U3399) );
  OAI22_X1 U11572 ( .A1(n10939), .A2(n10938), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n10937), .ZN(n10940) );
  AOI21_X1 U11573 ( .B1(n10942), .B2(n10941), .A(n10940), .ZN(n10943) );
  OAI221_X1 U11574 ( .B1(n10946), .B2(n10945), .C1(n10944), .C2(n6326), .A(
        n10943), .ZN(P2_U3230) );
  NOR2_X1 U11575 ( .A1(n10947), .A2(n11012), .ZN(n10950) );
  INV_X1 U11576 ( .A(n10948), .ZN(n10949) );
  AOI211_X1 U11577 ( .C1(n11017), .C2(n10951), .A(n10950), .B(n10949), .ZN(
        n10953) );
  AOI22_X1 U11578 ( .A1(n11100), .A2(n10953), .B1(n6337), .B2(n11099), .ZN(
        P2_U3463) );
  INV_X1 U11579 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10952) );
  AOI22_X1 U11580 ( .A1(n11104), .A2(n10953), .B1(n10952), .B2(n11101), .ZN(
        P2_U3402) );
  OAI21_X1 U11581 ( .B1(n10955), .B2(n11074), .A(n10954), .ZN(n10957) );
  AOI211_X1 U11582 ( .C1(n11078), .C2(n10958), .A(n10957), .B(n10956), .ZN(
        n10959) );
  AOI22_X1 U11583 ( .A1(n11081), .A2(n10959), .B1(n6995), .B2(n11080), .ZN(
        P1_U3526) );
  AOI22_X1 U11584 ( .A1(n11085), .A2(n10959), .B1(n5762), .B2(n11082), .ZN(
        P1_U3465) );
  INV_X1 U11585 ( .A(n10960), .ZN(n10964) );
  OAI22_X1 U11586 ( .A1(n10962), .A2(n11012), .B1(n10961), .B2(n11093), .ZN(
        n10963) );
  NOR2_X1 U11587 ( .A1(n10964), .A2(n10963), .ZN(n10966) );
  AOI22_X1 U11588 ( .A1(n11100), .A2(n10966), .B1(n6349), .B2(n11099), .ZN(
        P2_U3464) );
  INV_X1 U11589 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10965) );
  AOI22_X1 U11590 ( .A1(n11104), .A2(n10966), .B1(n10965), .B2(n11101), .ZN(
        P2_U3405) );
  AND2_X1 U11591 ( .A1(n10967), .A2(n11078), .ZN(n10972) );
  OAI21_X1 U11592 ( .B1(n10969), .B2(n11074), .A(n10968), .ZN(n10970) );
  NOR3_X1 U11593 ( .A1(n10972), .A2(n10971), .A3(n10970), .ZN(n10973) );
  AOI22_X1 U11594 ( .A1(n11081), .A2(n10973), .B1(n6997), .B2(n11080), .ZN(
        P1_U3527) );
  AOI22_X1 U11595 ( .A1(n11085), .A2(n10973), .B1(n5777), .B2(n11082), .ZN(
        P1_U3468) );
  NOR2_X1 U11596 ( .A1(n10974), .A2(n11093), .ZN(n10976) );
  AOI211_X1 U11597 ( .C1(n11097), .C2(n10977), .A(n10976), .B(n10975), .ZN(
        n10979) );
  AOI22_X1 U11598 ( .A1(n11100), .A2(n10979), .B1(n7348), .B2(n11099), .ZN(
        P2_U3465) );
  INV_X1 U11599 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10978) );
  AOI22_X1 U11600 ( .A1(n11104), .A2(n10979), .B1(n10978), .B2(n11101), .ZN(
        P2_U3408) );
  NAND2_X1 U11601 ( .A1(n10980), .A2(n11039), .ZN(n10982) );
  OAI211_X1 U11602 ( .C1(n10983), .C2(n11074), .A(n10982), .B(n10981), .ZN(
        n10984) );
  NOR2_X1 U11603 ( .A1(n10985), .A2(n10984), .ZN(n10987) );
  AOI22_X1 U11604 ( .A1(n11081), .A2(n10987), .B1(n5812), .B2(n11080), .ZN(
        P1_U3529) );
  INV_X1 U11605 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10986) );
  AOI22_X1 U11606 ( .A1(n11085), .A2(n10987), .B1(n10986), .B2(n11082), .ZN(
        P1_U3474) );
  OAI22_X1 U11607 ( .A1(n10989), .A2(n11012), .B1(n10988), .B2(n11093), .ZN(
        n10990) );
  NOR2_X1 U11608 ( .A1(n10991), .A2(n10990), .ZN(n10993) );
  AOI22_X1 U11609 ( .A1(n11100), .A2(n10993), .B1(n6395), .B2(n11099), .ZN(
        P2_U3466) );
  INV_X1 U11610 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10992) );
  AOI22_X1 U11611 ( .A1(n11104), .A2(n10993), .B1(n10992), .B2(n11101), .ZN(
        P2_U3411) );
  NOR2_X1 U11612 ( .A1(n10994), .A2(n11012), .ZN(n10996) );
  AOI211_X1 U11613 ( .C1(n11017), .C2(n10997), .A(n10996), .B(n10995), .ZN(
        n10999) );
  AOI22_X1 U11614 ( .A1(n11100), .A2(n10999), .B1(n7698), .B2(n11099), .ZN(
        P2_U3467) );
  INV_X1 U11615 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10998) );
  AOI22_X1 U11616 ( .A1(n11104), .A2(n10999), .B1(n10998), .B2(n11101), .ZN(
        P2_U3414) );
  NOR2_X1 U11617 ( .A1(n11000), .A2(n11093), .ZN(n11002) );
  AOI211_X1 U11618 ( .C1(n11003), .C2(n11097), .A(n11002), .B(n11001), .ZN(
        n11005) );
  AOI22_X1 U11619 ( .A1(n11100), .A2(n11005), .B1(n6421), .B2(n11099), .ZN(
        P2_U3468) );
  INV_X1 U11620 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n11004) );
  AOI22_X1 U11621 ( .A1(n11104), .A2(n11005), .B1(n11004), .B2(n11101), .ZN(
        P2_U3417) );
  NOR2_X1 U11622 ( .A1(n11007), .A2(n11006), .ZN(n11009) );
  AOI211_X1 U11623 ( .C1(n11017), .C2(n11010), .A(n11009), .B(n11008), .ZN(
        n11011) );
  AOI22_X1 U11624 ( .A1(n11100), .A2(n11011), .B1(n7792), .B2(n11099), .ZN(
        P2_U3469) );
  AOI22_X1 U11625 ( .A1(n11104), .A2(n11011), .B1(n6434), .B2(n11101), .ZN(
        P2_U3420) );
  NOR2_X1 U11626 ( .A1(n11013), .A2(n11012), .ZN(n11015) );
  AOI211_X1 U11627 ( .C1(n11017), .C2(n11016), .A(n11015), .B(n11014), .ZN(
        n11019) );
  AOI22_X1 U11628 ( .A1(n11100), .A2(n11019), .B1(n6450), .B2(n11099), .ZN(
        P2_U3470) );
  INV_X1 U11629 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n11018) );
  AOI22_X1 U11630 ( .A1(n11104), .A2(n11019), .B1(n11018), .B2(n11101), .ZN(
        P2_U3423) );
  XNOR2_X1 U11631 ( .A(n11020), .B(n11023), .ZN(n11047) );
  NAND2_X1 U11632 ( .A1(n11022), .A2(n11021), .ZN(n11024) );
  XNOR2_X1 U11633 ( .A(n11024), .B(n11023), .ZN(n11031) );
  AOI22_X1 U11634 ( .A1(n11028), .A2(n11027), .B1(n11026), .B2(n11025), .ZN(
        n11029) );
  OAI21_X1 U11635 ( .B1(n11031), .B2(n11030), .A(n11029), .ZN(n11032) );
  AOI21_X1 U11636 ( .B1(n11047), .B2(n11033), .A(n11032), .ZN(n11052) );
  OAI211_X1 U11637 ( .C1(n11036), .C2(n11037), .A(n11035), .B(n11034), .ZN(
        n11043) );
  OAI21_X1 U11638 ( .B1(n11037), .B2(n11074), .A(n11043), .ZN(n11038) );
  AOI21_X1 U11639 ( .B1(n11047), .B2(n11039), .A(n11038), .ZN(n11040) );
  AND2_X1 U11640 ( .A1(n11052), .A2(n11040), .ZN(n11042) );
  AOI22_X1 U11641 ( .A1(n11081), .A2(n11042), .B1(n7006), .B2(n11080), .ZN(
        P1_U3533) );
  INV_X1 U11642 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n11041) );
  AOI22_X1 U11643 ( .A1(n11085), .A2(n11042), .B1(n11041), .B2(n11082), .ZN(
        P1_U3486) );
  INV_X1 U11644 ( .A(n11043), .ZN(n11044) );
  AOI22_X1 U11645 ( .A1(n11047), .A2(n11046), .B1(n11045), .B2(n11044), .ZN(
        n11058) );
  NAND2_X1 U11646 ( .A1(n11051), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n11048) );
  OAI21_X1 U11647 ( .B1(n11050), .B2(n11049), .A(n11048), .ZN(n11054) );
  NOR2_X1 U11648 ( .A1(n11052), .A2(n11051), .ZN(n11053) );
  AOI211_X1 U11649 ( .C1(n11056), .C2(n11055), .A(n11054), .B(n11053), .ZN(
        n11057) );
  NAND2_X1 U11650 ( .A1(n11058), .A2(n11057), .ZN(P1_U3282) );
  NAND2_X1 U11651 ( .A1(n11059), .A2(n11097), .ZN(n11060) );
  OAI21_X1 U11652 ( .B1(n11061), .B2(n11093), .A(n11060), .ZN(n11062) );
  NOR2_X1 U11653 ( .A1(n11063), .A2(n11062), .ZN(n11065) );
  AOI22_X1 U11654 ( .A1(n11100), .A2(n11065), .B1(n6461), .B2(n11099), .ZN(
        P2_U3471) );
  INV_X1 U11655 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n11064) );
  AOI22_X1 U11656 ( .A1(n11104), .A2(n11065), .B1(n11064), .B2(n11101), .ZN(
        P2_U3426) );
  OAI21_X1 U11657 ( .B1(n11067), .B2(n11074), .A(n11066), .ZN(n11068) );
  AOI211_X1 U11658 ( .C1(n11070), .C2(n11078), .A(n11069), .B(n11068), .ZN(
        n11072) );
  AOI22_X1 U11659 ( .A1(n11081), .A2(n11072), .B1(n5893), .B2(n11080), .ZN(
        P1_U3534) );
  INV_X1 U11660 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n11071) );
  AOI22_X1 U11661 ( .A1(n11085), .A2(n11072), .B1(n11071), .B2(n11082), .ZN(
        P1_U3489) );
  OAI21_X1 U11662 ( .B1(n11075), .B2(n11074), .A(n11073), .ZN(n11076) );
  AOI211_X1 U11663 ( .C1(n11079), .C2(n11078), .A(n11077), .B(n11076), .ZN(
        n11084) );
  AOI22_X1 U11664 ( .A1(n11081), .A2(n11084), .B1(n7823), .B2(n11080), .ZN(
        P1_U3535) );
  INV_X1 U11665 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n11083) );
  AOI22_X1 U11666 ( .A1(n11085), .A2(n11084), .B1(n11083), .B2(n11082), .ZN(
        P1_U3492) );
  NAND2_X1 U11667 ( .A1(n11086), .A2(n11097), .ZN(n11087) );
  OAI21_X1 U11668 ( .B1(n11088), .B2(n11093), .A(n11087), .ZN(n11089) );
  NOR2_X1 U11669 ( .A1(n11090), .A2(n11089), .ZN(n11092) );
  AOI22_X1 U11670 ( .A1(n11100), .A2(n11092), .B1(n6474), .B2(n11099), .ZN(
        P2_U3472) );
  INV_X1 U11671 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n11091) );
  AOI22_X1 U11672 ( .A1(n11104), .A2(n11092), .B1(n11091), .B2(n11101), .ZN(
        P2_U3429) );
  NOR2_X1 U11673 ( .A1(n11094), .A2(n11093), .ZN(n11096) );
  AOI211_X1 U11674 ( .C1(n11098), .C2(n11097), .A(n11096), .B(n11095), .ZN(
        n11103) );
  AOI22_X1 U11675 ( .A1(n11100), .A2(n11103), .B1(n6491), .B2(n11099), .ZN(
        P2_U3473) );
  INV_X1 U11676 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n11102) );
  AOI22_X1 U11677 ( .A1(n11104), .A2(n11103), .B1(n11102), .B2(n11101), .ZN(
        P2_U3432) );
  XNOR2_X1 U11678 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  NAND3_X1 U6290 ( .A1(n5249), .A2(n5248), .A3(n5714), .ZN(n10171) );
  CLKBUF_X1 U5185 ( .A(n6307), .Z(n8678) );
  CLKBUF_X1 U5200 ( .A(n5791), .Z(n6167) );
  NAND2_X1 U5347 ( .A1(n8145), .A2(n8144), .ZN(n8143) );
endmodule

