

module b17_C_SARLock_k_128_5 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127, U355, U356, U357, U358, U359, U360, U361, 
        U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, U373, U374, 
        U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, U376, U247, 
        U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, 
        U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223, 
        U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254, U255, 
        U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, U266, U267, 
        U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, U278, U279, 
        U280, U281, U282, U212, U215, U213, U214, P3_U3274, P3_U3275, P3_U3276, 
        P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, P3_U3057, P3_U3056, 
        P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, P3_U3050, P3_U3049, 
        P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, P3_U3043, P3_U3042, 
        P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, P3_U3036, P3_U3035, 
        P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, P3_U3029, P3_U3280, 
        P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, P3_U3024, P3_U3023, 
        P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, P3_U3017, P3_U3016, 
        P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, P3_U3010, P3_U3009, 
        P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, P3_U3003, P3_U3002, 
        P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, P3_U2997, P3_U2996, 
        P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, P3_U2990, P3_U2989, 
        P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, P3_U2983, P3_U2982, 
        P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, P3_U2976, P3_U2975, 
        P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, P3_U2969, P3_U2968, 
        P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, P3_U2962, P3_U2961, 
        P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, P3_U2955, P3_U2954, 
        P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, P3_U2948, P3_U2947, 
        P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, P3_U2941, P3_U2940, 
        P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, P3_U2934, P3_U2933, 
        P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, P3_U2927, P3_U2926, 
        P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, P3_U2920, P3_U2919, 
        P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, P3_U2913, P3_U2912, 
        P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, P3_U2906, P3_U2905, 
        P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, P3_U2899, P3_U2898, 
        P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, P3_U2892, P3_U2891, 
        P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, P3_U2885, P3_U2884, 
        P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, P3_U2878, P3_U2877, 
        P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, P3_U2871, P3_U2870, 
        P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, P3_U3289, P3_U3290, 
        P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, P3_U2862, P3_U2861, 
        P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, P3_U2855, P3_U2854, 
        P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, P3_U2848, P3_U2847, 
        P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, P3_U2841, P3_U2840, 
        P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, P3_U2834, P3_U2833, 
        P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, P3_U2827, P3_U2826, 
        P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, P3_U2820, P3_U2819, 
        P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, P3_U2813, P3_U2812, 
        P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, P3_U2806, P3_U2805, 
        P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, P3_U2799, P3_U2798, 
        P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, P3_U2792, P3_U2791, 
        P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, P3_U2785, P3_U2784, 
        P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, P3_U2778, P3_U2777, 
        P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, P3_U2771, P3_U2770, 
        P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, P3_U2764, P3_U2763, 
        P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, P3_U2757, P3_U2756, 
        P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, P3_U2750, P3_U2749, 
        P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, P3_U2743, P3_U2742, 
        P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, P3_U2736, P3_U2735, 
        P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, P3_U2729, P3_U2728, 
        P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, P3_U2722, P3_U2721, 
        P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, P3_U2715, P3_U2714, 
        P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, P3_U2708, P3_U2707, 
        P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, P3_U2701, P3_U2700, 
        P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, P3_U2694, P3_U2693, 
        P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, P3_U2687, P3_U2686, 
        P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, P3_U2680, P3_U2679, 
        P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, P3_U2673, P3_U2672, 
        P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, P3_U2666, P3_U2665, 
        P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, P3_U2659, P3_U2658, 
        P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, P3_U2652, P3_U2651, 
        P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, P3_U2645, P3_U2644, 
        P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, P3_U3292, P3_U2638, 
        P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, P3_U3296, P3_U2635, 
        P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, P2_U3585, P2_U3586, 
        P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, 
        P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, P2_U3178, P2_U3177, 
        P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, 
        P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, 
        P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, 
        P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, P2_U3150, P2_U3149, 
        P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, P2_U3143, P2_U3142, 
        P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, P2_U3136, P2_U3135, 
        P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, P2_U3129, P2_U3128, 
        P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, P2_U3122, P2_U3121, 
        P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, P2_U3115, P2_U3114, 
        P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, P2_U3108, P2_U3107, 
        P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, P2_U3101, P2_U3100, 
        P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, P2_U3094, P2_U3093, 
        P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, P2_U3087, P2_U3086, 
        P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, P2_U3080, P2_U3079, 
        P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, P2_U3073, P2_U3072, 
        P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, P2_U3066, P2_U3065, 
        P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, P2_U3059, P2_U3058, 
        P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, P2_U3052, P2_U3051, 
        P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, P2_U3599, P2_U3600, 
        P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, P2_U3605, P2_U3046, 
        P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, P2_U3040, P2_U3039, 
        P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, P2_U3033, P2_U3032, 
        P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, P2_U3026, P2_U3025, 
        P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, P2_U3019, P2_U3018, 
        P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, P2_U3012, P2_U3011, 
        P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, P2_U3005, P2_U3004, 
        P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, P2_U2998, P2_U2997, 
        P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, P2_U2991, P2_U2990, 
        P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, P2_U2984, P2_U2983, 
        P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, P2_U2977, P2_U2976, 
        P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, P2_U2970, P2_U2969, 
        P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, P2_U2963, P2_U2962, 
        P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, P2_U2956, P2_U2955, 
        P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, P2_U2949, P2_U2948, 
        P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, P2_U2942, P2_U2941, 
        P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, P2_U2935, P2_U2934, 
        P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, P2_U2928, P2_U2927, 
        P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, P2_U2921, P2_U2920, 
        P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, P2_U2914, P2_U2913, 
        P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, P2_U2907, P2_U2906, 
        P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, P2_U2900, P2_U2899, 
        P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, P2_U2893, P2_U2892, 
        P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, P2_U2886, P2_U2885, 
        P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, P2_U2879, P2_U2878, 
        P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, P2_U2872, P2_U2871, 
        P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, P2_U2865, P2_U2864, 
        P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, P2_U2858, P2_U2857, 
        P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, P2_U2851, P2_U2850, 
        P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, P2_U2844, P2_U2843, 
        P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, P2_U2837, P2_U2836, 
        P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, P2_U2830, P2_U2829, 
        P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, P2_U2823, P2_U2822, 
        P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, P2_U2818, P2_U3610, 
        P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, P2_U2814, P1_U3458, 
        P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3210, P1_U3209, 
        P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, P1_U3203, P1_U3202, 
        P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, P1_U3196, P1_U3195, 
        P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, P1_U3191, P1_U3190, 
        P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, P1_U3184, P1_U3183, 
        P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, P1_U3177, P1_U3176, 
        P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, P1_U3170, P1_U3169, 
        P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, P1_U3466, P1_U3163, 
        P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, P1_U3157, P1_U3156, 
        P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, P1_U3150, P1_U3149, 
        P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, P1_U3143, P1_U3142, 
        P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, P1_U3136, P1_U3135, 
        P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, P1_U3129, P1_U3128, 
        P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, P1_U3122, P1_U3121, 
        P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, P1_U3115, P1_U3114, 
        P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, P1_U3108, P1_U3107, 
        P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, P1_U3101, P1_U3100, 
        P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, P1_U3094, P1_U3093, 
        P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, P1_U3087, P1_U3086, 
        P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, P1_U3080, P1_U3079, 
        P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, P1_U3073, P1_U3072, 
        P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, P1_U3066, P1_U3065, 
        P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, P1_U3059, P1_U3058, 
        P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, P1_U3052, P1_U3051, 
        P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, P1_U3045, P1_U3044, 
        P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, P1_U3038, P1_U3037, 
        P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, P1_U3469, P1_U3472, 
        P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, P1_U3477, P1_U3478, 
        P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, P1_U3026, P1_U3025, 
        P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, P1_U3019, P1_U3018, 
        P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, P1_U3012, P1_U3011, 
        P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, P1_U3005, P1_U3004, 
        P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, P1_U2998, P1_U2997, 
        P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, P1_U2991, P1_U2990, 
        P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, P1_U2984, P1_U2983, 
        P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, P1_U2977, P1_U2976, 
        P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, P1_U2970, P1_U2969, 
        P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, P1_U2963, P1_U2962, 
        P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, P1_U2956, P1_U2955, 
        P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, P1_U2949, P1_U2948, 
        P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, P1_U2942, P1_U2941, 
        P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, P1_U2935, P1_U2934, 
        P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, P1_U2928, P1_U2927, 
        P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, P1_U2921, P1_U2920, 
        P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, P1_U2914, P1_U2913, 
        P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, P1_U2907, P1_U2906, 
        P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, P1_U2900, P1_U2899, 
        P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, P1_U2893, P1_U2892, 
        P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, P1_U2886, P1_U2885, 
        P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, P1_U2879, P1_U2878, 
        P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, P1_U2872, P1_U2871, 
        P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, P1_U2865, P1_U2864, 
        P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, P1_U2858, P1_U2857, 
        P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, P1_U2851, P1_U2850, 
        P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, P1_U2844, P1_U2843, 
        P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, P1_U2837, P1_U2836, 
        P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, P1_U2830, P1_U2829, 
        P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, P1_U2823, P1_U2822, 
        P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, P1_U2816, P1_U2815, 
        P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, P1_U2809, P1_U2808, 
        P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, P1_U3484, P1_U2805, 
        P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, P1_U3487, P1_U2801
 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
         n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
         n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
         n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
         n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
         n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
         n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
         n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
         n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
         n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
         n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
         n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
         n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
         n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
         n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
         n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
         n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
         n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
         n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
         n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
         n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
         n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
         n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133,
         n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
         n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
         n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
         n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
         n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
         n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
         n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
         n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
         n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
         n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
         n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
         n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
         n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
         n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
         n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
         n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
         n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
         n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
         n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
         n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
         n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
         n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
         n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
         n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
         n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325,
         n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333,
         n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
         n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
         n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
         n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
         n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
         n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
         n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
         n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
         n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
         n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429,
         n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
         n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
         n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
         n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
         n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
         n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477,
         n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
         n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
         n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501,
         n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
         n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
         n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
         n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533,
         n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
         n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549,
         n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
         n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565,
         n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573,
         n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
         n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
         n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
         n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621,
         n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
         n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
         n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
         n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
         n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
         n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
         n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
         n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374,
         n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
         n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
         n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
         n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406,
         n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,
         n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422,
         n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430,
         n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438,
         n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446,
         n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454,
         n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462,
         n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470,
         n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478,
         n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486,
         n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494,
         n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502,
         n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510,
         n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518,
         n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526,
         n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534,
         n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542,
         n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550,
         n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558,
         n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566,
         n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574,
         n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582,
         n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590,
         n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598,
         n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606,
         n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614,
         n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622,
         n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630,
         n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638,
         n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646,
         n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654,
         n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662,
         n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670,
         n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678,
         n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686,
         n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694,
         n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702,
         n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710,
         n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718,
         n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726,
         n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734,
         n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742,
         n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750,
         n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758,
         n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766,
         n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774,
         n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782,
         n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790,
         n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798,
         n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806,
         n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814,
         n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822,
         n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830,
         n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838,
         n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846,
         n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854,
         n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862,
         n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870,
         n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878,
         n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886,
         n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894,
         n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902,
         n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910,
         n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918,
         n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926,
         n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934,
         n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942,
         n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950,
         n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958,
         n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966,
         n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974,
         n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982,
         n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990,
         n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998,
         n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006,
         n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014,
         n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022,
         n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030,
         n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038,
         n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046,
         n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054,
         n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062,
         n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070,
         n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078,
         n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086,
         n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094,
         n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102,
         n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110,
         n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118,
         n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126,
         n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134,
         n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142,
         n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150,
         n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158,
         n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166,
         n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174,
         n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182,
         n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190,
         n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198,
         n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206,
         n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214,
         n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222,
         n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230,
         n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238,
         n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246,
         n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254,
         n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262,
         n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270,
         n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278,
         n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286,
         n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294,
         n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302,
         n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310,
         n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318,
         n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326,
         n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334,
         n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342,
         n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350,
         n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358,
         n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366,
         n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374,
         n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382,
         n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390,
         n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398,
         n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406,
         n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414,
         n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422,
         n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430,
         n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438,
         n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446,
         n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454,
         n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462,
         n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470,
         n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478,
         n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486,
         n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494,
         n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502,
         n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510,
         n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518,
         n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526,
         n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534,
         n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542,
         n16543, n16544, n16546, n16547, n16548, n16549, n16550, n16551,
         n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559,
         n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567,
         n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575,
         n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583,
         n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591,
         n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599,
         n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607,
         n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615,
         n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623,
         n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631,
         n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639,
         n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647,
         n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655,
         n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663,
         n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671,
         n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679,
         n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687,
         n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695,
         n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703,
         n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711,
         n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719,
         n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
         n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735,
         n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743,
         n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751,
         n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759,
         n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767,
         n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775,
         n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783,
         n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791,
         n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799,
         n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807,
         n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815,
         n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823,
         n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831,
         n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839,
         n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847,
         n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855,
         n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863,
         n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871,
         n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879,
         n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887,
         n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895,
         n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903,
         n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911,
         n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919,
         n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927,
         n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935,
         n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943,
         n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951,
         n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959,
         n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967,
         n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975,
         n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983,
         n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991,
         n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999,
         n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007,
         n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015,
         n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023,
         n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031,
         n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039,
         n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047,
         n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055,
         n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063,
         n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071,
         n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079,
         n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087,
         n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095,
         n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103,
         n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111,
         n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119,
         n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127,
         n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135,
         n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143,
         n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151,
         n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159,
         n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167,
         n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175,
         n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183,
         n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191,
         n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199,
         n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207,
         n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215,
         n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223,
         n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231,
         n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239,
         n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247,
         n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255,
         n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263,
         n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271,
         n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279,
         n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287,
         n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295,
         n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303,
         n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311,
         n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319,
         n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327,
         n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335,
         n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343,
         n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351,
         n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359,
         n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367,
         n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375,
         n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383,
         n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391,
         n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399,
         n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407,
         n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415,
         n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423,
         n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431,
         n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439,
         n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447,
         n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455,
         n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463,
         n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471,
         n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479,
         n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487,
         n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495,
         n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503,
         n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511,
         n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519,
         n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527,
         n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535,
         n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543,
         n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551,
         n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559,
         n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567,
         n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575,
         n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583,
         n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591,
         n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599,
         n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607,
         n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615,
         n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623,
         n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631,
         n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639,
         n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647,
         n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655,
         n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663,
         n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671,
         n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679,
         n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687,
         n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695,
         n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703,
         n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711,
         n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719,
         n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727,
         n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735,
         n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743,
         n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751,
         n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759,
         n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767,
         n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775,
         n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783,
         n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791,
         n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799,
         n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807,
         n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815,
         n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823,
         n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831,
         n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839,
         n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847,
         n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855,
         n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863,
         n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871,
         n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879,
         n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887,
         n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895,
         n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903,
         n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911,
         n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919,
         n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927,
         n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935,
         n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943,
         n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951,
         n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959,
         n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967,
         n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975,
         n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983,
         n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991,
         n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999,
         n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007,
         n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015,
         n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023,
         n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031,
         n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039,
         n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047,
         n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055,
         n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063,
         n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071,
         n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079,
         n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087,
         n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095,
         n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103,
         n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111,
         n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119,
         n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127,
         n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135,
         n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143,
         n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151,
         n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159,
         n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167,
         n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175,
         n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183,
         n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191,
         n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199,
         n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207,
         n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215,
         n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223,
         n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231,
         n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239,
         n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247,
         n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255,
         n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263,
         n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271,
         n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279,
         n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287,
         n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295,
         n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303,
         n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311,
         n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319,
         n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327,
         n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335,
         n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343,
         n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351,
         n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359,
         n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367,
         n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375,
         n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383,
         n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391,
         n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399,
         n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407,
         n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415,
         n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423,
         n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431,
         n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439,
         n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447,
         n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455,
         n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463,
         n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471,
         n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479,
         n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487,
         n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495,
         n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503,
         n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511,
         n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519,
         n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527,
         n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535,
         n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543,
         n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551,
         n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559,
         n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567,
         n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575,
         n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583,
         n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591,
         n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599,
         n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607,
         n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615,
         n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623,
         n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631,
         n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639,
         n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647,
         n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655,
         n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663,
         n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671,
         n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679,
         n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687,
         n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695,
         n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703,
         n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711,
         n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719,
         n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727,
         n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735,
         n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743,
         n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751,
         n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759,
         n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767,
         n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775,
         n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783,
         n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791,
         n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799,
         n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807,
         n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815,
         n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823,
         n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831,
         n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839,
         n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847,
         n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855,
         n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863,
         n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871,
         n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879,
         n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887,
         n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895,
         n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903,
         n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911,
         n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919,
         n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927,
         n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935,
         n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943,
         n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951,
         n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959,
         n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967,
         n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975,
         n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983,
         n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991,
         n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999,
         n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007,
         n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015,
         n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023,
         n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031,
         n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039,
         n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047,
         n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055,
         n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063,
         n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071,
         n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079,
         n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087,
         n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095,
         n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103,
         n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111,
         n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119,
         n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127,
         n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135,
         n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143,
         n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151,
         n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159,
         n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167,
         n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175,
         n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183,
         n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191,
         n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199,
         n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207,
         n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215,
         n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223,
         n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231,
         n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239,
         n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247,
         n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255,
         n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263,
         n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271,
         n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279,
         n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287,
         n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295,
         n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303,
         n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311,
         n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319,
         n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327,
         n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335,
         n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343,
         n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351,
         n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359,
         n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367,
         n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375,
         n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383,
         n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391,
         n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399,
         n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407,
         n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415,
         n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423,
         n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431,
         n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439,
         n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447,
         n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455,
         n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463,
         n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471,
         n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479,
         n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487,
         n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495,
         n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503,
         n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511,
         n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519,
         n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527,
         n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535,
         n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543,
         n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551,
         n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559,
         n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567,
         n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575,
         n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583,
         n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591,
         n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599,
         n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607,
         n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615,
         n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623,
         n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631,
         n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639,
         n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647,
         n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655,
         n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663,
         n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671,
         n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679,
         n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687,
         n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695,
         n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703,
         n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711,
         n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719,
         n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727,
         n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735,
         n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743,
         n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751,
         n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759,
         n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767,
         n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775,
         n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783,
         n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791,
         n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799,
         n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807,
         n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815,
         n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823,
         n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831,
         n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839,
         n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847,
         n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855,
         n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863,
         n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871,
         n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879,
         n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887,
         n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895,
         n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903,
         n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911,
         n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919,
         n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927,
         n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935,
         n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943,
         n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951,
         n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959,
         n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967,
         n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975,
         n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983,
         n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991,
         n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999,
         n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007,
         n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015,
         n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023,
         n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031,
         n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039,
         n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047,
         n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055,
         n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063,
         n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071,
         n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079,
         n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087,
         n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095,
         n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103,
         n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111,
         n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119,
         n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127,
         n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135,
         n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143,
         n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151,
         n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159,
         n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167,
         n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175,
         n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183,
         n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191,
         n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199,
         n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207,
         n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215,
         n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223,
         n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231,
         n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239,
         n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247,
         n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255,
         n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263,
         n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271,
         n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279,
         n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287,
         n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295,
         n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303,
         n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311,
         n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319,
         n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327,
         n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335,
         n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343,
         n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351,
         n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359,
         n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367,
         n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375,
         n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383,
         n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391,
         n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399,
         n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407,
         n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415,
         n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423,
         n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431,
         n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439,
         n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447,
         n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455,
         n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463,
         n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471,
         n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479,
         n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487,
         n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495,
         n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503,
         n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511,
         n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519,
         n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527,
         n20528, n20529, n20530, n20531, n20532, n20533, n20534, n20535,
         n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543,
         n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551,
         n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559,
         n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567,
         n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575,
         n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583,
         n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591,
         n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599,
         n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607,
         n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615,
         n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623,
         n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631,
         n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639,
         n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647,
         n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655,
         n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663,
         n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671,
         n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679,
         n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687,
         n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695,
         n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703,
         n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711,
         n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719,
         n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727,
         n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735,
         n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743,
         n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751,
         n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759,
         n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767,
         n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775,
         n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783,
         n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791,
         n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799,
         n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807,
         n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815,
         n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823,
         n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831,
         n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839,
         n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847,
         n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855,
         n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863,
         n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871,
         n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879,
         n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887,
         n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895,
         n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903,
         n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911,
         n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919,
         n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927,
         n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935,
         n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943,
         n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951,
         n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959,
         n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967,
         n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975,
         n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983,
         n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991,
         n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999,
         n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007,
         n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015,
         n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023,
         n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031,
         n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039,
         n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047,
         n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055,
         n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063,
         n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071,
         n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079,
         n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087,
         n21088, n21089, n21090, n21091, n21092, n21093, n21094, n21095,
         n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103,
         n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111,
         n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119,
         n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127,
         n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135,
         n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143,
         n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151,
         n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159,
         n21160, n21161, n21162, n21163, n21164, n21165, n21166, n21167;

  NOR2_X1 U11191 ( .A1(n13643), .A2(n13644), .ZN(n19275) );
  NOR2_X1 U11192 ( .A1(n13645), .A2(n13644), .ZN(n19274) );
  INV_X2 U11193 ( .A(n19030), .ZN(n18957) );
  AND2_X1 U11194 ( .A1(n12912), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20116)
         );
  INV_X1 U11197 ( .A(n15594), .ZN(n17123) );
  AND2_X1 U11198 ( .A1(n9753), .A2(n15408), .ZN(n12695) );
  CLKBUF_X2 U11199 ( .A(n10339), .Z(n10343) );
  INV_X1 U11200 ( .A(n11202), .ZN(n12705) );
  BUF_X1 U11201 ( .A(n12374), .Z(n12452) );
  AND2_X1 U11202 ( .A1(n9750), .A2(n15408), .ZN(n10395) );
  BUF_X1 U11203 ( .A(n10243), .Z(n9759) );
  INV_X2 U11204 ( .A(n14175), .ZN(n13459) );
  NAND2_X1 U11205 ( .A1(n9795), .A2(n15408), .ZN(n12689) );
  AND2_X1 U11206 ( .A1(n10331), .A2(n9902), .ZN(n10340) );
  CLKBUF_X2 U11207 ( .A(n10826), .Z(n9782) );
  NAND2_X1 U11208 ( .A1(n12838), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12654) );
  NAND2_X1 U11209 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n10380), .ZN(
        n12699) );
  INV_X2 U11210 ( .A(n15474), .ZN(n17215) );
  CLKBUF_X2 U11211 ( .A(n15463), .Z(n17207) );
  INV_X1 U11212 ( .A(n15562), .ZN(n9758) );
  INV_X1 U11213 ( .A(n17175), .ZN(n17212) );
  INV_X1 U11214 ( .A(n17175), .ZN(n15550) );
  CLKBUF_X1 U11215 ( .A(n15463), .Z(n17173) );
  NOR2_X1 U11216 ( .A1(n12924), .A2(n12921), .ZN(n15538) );
  AND2_X2 U11217 ( .A1(n10312), .A2(n15502), .ZN(n11253) );
  CLKBUF_X1 U11218 ( .A(n11380), .Z(n12208) );
  CLKBUF_X2 U11219 ( .A(n11528), .Z(n12327) );
  CLKBUF_X2 U11220 ( .A(n9747), .Z(n12317) );
  CLKBUF_X1 U11221 ( .A(n11371), .Z(n12116) );
  AND2_X2 U11222 ( .A1(n10953), .A2(n10304), .ZN(n10826) );
  CLKBUF_X2 U11223 ( .A(n11438), .Z(n12326) );
  CLKBUF_X2 U11224 ( .A(n12243), .Z(n12323) );
  CLKBUF_X2 U11225 ( .A(n10267), .Z(n9755) );
  BUF_X1 U11226 ( .A(n11451), .Z(n20136) );
  CLKBUF_X1 U11227 ( .A(n11455), .Z(n20152) );
  INV_X1 U11228 ( .A(n11455), .ZN(n13244) );
  AND4_X2 U11229 ( .A1(n11347), .A2(n11346), .A3(n11345), .A4(n11344), .ZN(
        n12350) );
  AND4_X1 U11230 ( .A1(n11315), .A2(n11316), .A3(n11317), .A4(n11314), .ZN(
        n11327) );
  AND2_X1 U11231 ( .A1(n13411), .A2(n13392), .ZN(n9785) );
  AND2_X2 U11232 ( .A1(n11321), .A2(n11320), .ZN(n12243) );
  AND2_X1 U11233 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13388) );
  CLKBUF_X1 U11234 ( .A(n18730), .Z(n9746) );
  NOR2_X1 U11235 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18824), .ZN(n18730) );
  INV_X4 U11236 ( .A(n15697), .ZN(n9760) );
  CLKBUF_X2 U11238 ( .A(n11417), .Z(n12144) );
  INV_X2 U11239 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9780) );
  AND2_X1 U11240 ( .A1(n12350), .A2(n20160), .ZN(n11481) );
  OR2_X1 U11241 ( .A1(n11545), .A2(n11544), .ZN(n11558) );
  NAND2_X1 U11242 ( .A1(n9776), .A2(n10101), .ZN(n10185) );
  AND3_X1 U11243 ( .A1(n10257), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n10999), 
        .ZN(n9801) );
  INV_X1 U11244 ( .A(n13265), .ZN(n10353) );
  NOR2_X1 U11245 ( .A1(n9771), .A2(n14487), .ZN(n11759) );
  BUF_X2 U11246 ( .A(n10158), .Z(n9752) );
  NAND2_X1 U11247 ( .A1(n12861), .A2(n15408), .ZN(n15402) );
  OR2_X1 U11248 ( .A1(n12916), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12919) );
  AND2_X1 U11249 ( .A1(n12448), .A2(n10135), .ZN(n12441) );
  NAND2_X1 U11251 ( .A1(n11520), .A2(n11519), .ZN(n11664) );
  NAND2_X1 U11253 ( .A1(n11557), .A2(n11556), .ZN(n11840) );
  NOR2_X1 U11254 ( .A1(n13144), .A2(n14087), .ZN(n13175) );
  OAI21_X1 U11255 ( .B1(n10182), .B2(n10181), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10183) );
  AND2_X1 U11256 ( .A1(n9752), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10401) );
  AOI21_X1 U11257 ( .B1(n15048), .B2(n11301), .A(n11300), .ZN(n15038) );
  INV_X1 U11258 ( .A(n10539), .ZN(n10258) );
  INV_X2 U11259 ( .A(n12917), .ZN(n17224) );
  OR2_X1 U11260 ( .A1(n15693), .A2(n10128), .ZN(n15694) );
  NAND2_X1 U11261 ( .A1(n12811), .A2(n12810), .ZN(n14848) );
  OR2_X1 U11262 ( .A1(n12882), .A2(n11017), .ZN(n11249) );
  NAND2_X1 U11263 ( .A1(n18848), .A2(n12916), .ZN(n13030) );
  INV_X1 U11264 ( .A(n18874), .ZN(n18221) );
  AND2_X1 U11265 ( .A1(n14372), .A2(n14361), .ZN(n14284) );
  INV_X1 U11267 ( .A(n15648), .ZN(n17398) );
  NOR2_X1 U11269 ( .A1(n17781), .A2(n17779), .ZN(n17780) );
  INV_X1 U11270 ( .A(n19949), .ZN(n19926) );
  INV_X1 U11271 ( .A(n15861), .ZN(n19983) );
  OAI21_X1 U11272 ( .B1(n13605), .B2(n13603), .A(n13604), .ZN(n19854) );
  INV_X1 U11273 ( .A(n15600), .ZN(n12993) );
  INV_X2 U11274 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11311) );
  AND2_X2 U11275 ( .A1(n13393), .A2(n9883), .ZN(n9747) );
  AND2_X2 U11276 ( .A1(n11485), .A2(n11475), .ZN(n11820) );
  NAND2_X2 U11277 ( .A1(n16275), .A2(n10637), .ZN(n10119) );
  NOR2_X2 U11278 ( .A1(n20089), .A2(n13985), .ZN(n20052) );
  NAND2_X2 U11279 ( .A1(n10019), .A2(n10811), .ZN(n15098) );
  AND2_X1 U11280 ( .A1(n13617), .A2(n10361), .ZN(n13718) );
  NOR2_X2 U11281 ( .A1(n14808), .A2(n14810), .ZN(n14809) );
  NAND2_X4 U11282 ( .A1(n10223), .A2(n10222), .ZN(n10274) );
  BUF_X4 U11283 ( .A(n10171), .Z(n9748) );
  BUF_X4 U11284 ( .A(n10171), .Z(n9749) );
  BUF_X4 U11285 ( .A(n10171), .Z(n9750) );
  AOI21_X2 U11286 ( .B1(n13966), .B2(n14603), .A(n14606), .ZN(n14459) );
  NAND2_X2 U11287 ( .A1(n13965), .A2(n14505), .ZN(n13966) );
  NOR3_X2 U11288 ( .A1(n17573), .A2(n17584), .A3(n17925), .ZN(n17567) );
  NAND2_X2 U11289 ( .A1(n10199), .A2(n10198), .ZN(n10252) );
  INV_X2 U11290 ( .A(n10279), .ZN(n10257) );
  AND2_X4 U11291 ( .A1(n13411), .A2(n9883), .ZN(n11380) );
  AND2_X4 U11292 ( .A1(n11318), .A2(n13411), .ZN(n11371) );
  AND2_X2 U11293 ( .A1(n14006), .A2(n10080), .ZN(n14334) );
  NAND2_X2 U11294 ( .A1(n14002), .A2(n11949), .ZN(n14006) );
  NAND2_X2 U11295 ( .A1(n13621), .A2(n10785), .ZN(n13757) );
  NAND2_X2 U11296 ( .A1(n10783), .A2(n10782), .ZN(n13621) );
  NAND2_X2 U11297 ( .A1(n13246), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11669) );
  BUF_X4 U11298 ( .A(n10158), .Z(n9751) );
  BUF_X4 U11299 ( .A(n10158), .Z(n9753) );
  NAND2_X1 U11300 ( .A1(n10184), .A2(n10183), .ZN(n10267) );
  NOR3_X1 U11303 ( .A1(n18227), .A2(n18221), .A3(n15770), .ZN(n17256) );
  XNOR2_X2 U11304 ( .A(n11680), .B(n20069), .ZN(n13560) );
  NAND2_X2 U11305 ( .A1(n13425), .A2(n11674), .ZN(n11680) );
  AND2_X2 U11306 ( .A1(n11313), .A2(n13388), .ZN(n9757) );
  NOR2_X4 U11307 ( .A1(n12920), .A2(n12919), .ZN(n15559) );
  AND2_X4 U11308 ( .A1(n11319), .A2(n13392), .ZN(n12266) );
  NOR2_X4 U11309 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13392) );
  NOR3_X2 U11310 ( .A1(n13930), .A2(n18673), .A3(n13929), .ZN(n15642) );
  NAND2_X1 U11311 ( .A1(n14208), .A2(n14197), .ZN(n14199) );
  AND2_X1 U11312 ( .A1(n9777), .A2(n9778), .ZN(n10018) );
  AND2_X1 U11313 ( .A1(n13803), .A2(n13838), .ZN(n13839) );
  NOR2_X1 U11314 ( .A1(n14897), .A2(n14887), .ZN(n14886) );
  NAND2_X1 U11315 ( .A1(n17668), .A2(n18007), .ZN(n17667) );
  OR3_X1 U11316 ( .A1(n13709), .A2(n9841), .A3(n9959), .ZN(n9958) );
  AND3_X1 U11317 ( .A1(n15688), .A2(n15686), .A3(n15687), .ZN(n17668) );
  NAND2_X1 U11318 ( .A1(n13830), .A2(n13831), .ZN(n13709) );
  NAND2_X1 U11319 ( .A1(n11840), .A2(n11839), .ZN(n20214) );
  OR2_X1 U11320 ( .A1(n10369), .A2(n10370), .ZN(n10484) );
  OR2_X1 U11321 ( .A1(n10371), .A2(n10368), .ZN(n13815) );
  INV_X1 U11322 ( .A(n12528), .ZN(n13313) );
  INV_X1 U11323 ( .A(n17993), .ZN(n18086) );
  BUF_X1 U11324 ( .A(n12528), .Z(n9791) );
  INV_X1 U11325 ( .A(n10337), .ZN(n10348) );
  NAND2_X1 U11326 ( .A1(n17796), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17795) );
  NAND2_X1 U11327 ( .A1(n11819), .A2(n11818), .ZN(n13232) );
  AND2_X1 U11328 ( .A1(n10345), .A2(n10346), .ZN(n10322) );
  NOR2_X2 U11329 ( .A1(n18098), .A2(n18692), .ZN(n17930) );
  AOI21_X1 U11330 ( .B1(n15645), .B2(n9819), .A(n15644), .ZN(n18671) );
  NOR2_X1 U11331 ( .A1(n11031), .A2(n11030), .ZN(n11037) );
  OAI211_X1 U11332 ( .C1(n10333), .C2(n13758), .A(n10335), .B(n10334), .ZN(
        n10819) );
  AND2_X1 U11333 ( .A1(n13208), .A2(n13209), .ZN(n11028) );
  AND2_X1 U11334 ( .A1(n10295), .A2(n10999), .ZN(n10993) );
  OR2_X1 U11335 ( .A1(n10294), .A2(n10293), .ZN(n15502) );
  CLKBUF_X2 U11336 ( .A(n10258), .Z(n19265) );
  NAND2_X1 U11337 ( .A1(n10258), .A2(n10251), .ZN(n10283) );
  INV_X2 U11338 ( .A(n16394), .ZN(n18227) );
  INV_X2 U11339 ( .A(n9789), .ZN(n11013) );
  INV_X2 U11340 ( .A(n10274), .ZN(n14666) );
  INV_X4 U11342 ( .A(n10265), .ZN(n19259) );
  OR2_X1 U11344 ( .A1(n11378), .A2(n11377), .ZN(n11451) );
  NAND2_X2 U11345 ( .A1(n11327), .A2(n11326), .ZN(n20160) );
  OR2_X2 U11346 ( .A1(n11403), .A2(n11402), .ZN(n11456) );
  AND4_X1 U11347 ( .A1(n11343), .A2(n11342), .A3(n11341), .A4(n11340), .ZN(
        n11344) );
  AND4_X1 U11348 ( .A1(n11359), .A2(n11358), .A3(n11357), .A4(n11356), .ZN(
        n11365) );
  AND4_X1 U11349 ( .A1(n11325), .A2(n11324), .A3(n11323), .A4(n11322), .ZN(
        n11326) );
  AND4_X1 U11350 ( .A1(n11433), .A2(n11432), .A3(n11431), .A4(n11430), .ZN(
        n11445) );
  BUF_X2 U11351 ( .A(n11533), .Z(n12316) );
  BUF_X2 U11352 ( .A(n11372), .Z(n12299) );
  BUF_X2 U11353 ( .A(n11412), .Z(n12139) );
  BUF_X2 U11354 ( .A(n11496), .Z(n12325) );
  CLKBUF_X2 U11355 ( .A(n12266), .Z(n12324) );
  CLKBUF_X2 U11356 ( .A(n17176), .Z(n17194) );
  BUF_X2 U11357 ( .A(n12096), .Z(n12328) );
  AND2_X1 U11358 ( .A1(n11311), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11321) );
  AND2_X2 U11359 ( .A1(n13392), .A2(n13393), .ZN(n12096) );
  AND2_X1 U11360 ( .A1(n11311), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11312) );
  AND2_X1 U11361 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9883) );
  NOR2_X1 U11362 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11313) );
  INV_X1 U11363 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10328) );
  XNOR2_X1 U11364 ( .A(n13971), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14001) );
  AND2_X1 U11365 ( .A1(n9997), .A2(n9996), .ZN(n14095) );
  OAI21_X1 U11366 ( .B1(n10945), .B2(n10944), .A(n10137), .ZN(n10952) );
  AND2_X1 U11367 ( .A1(n15019), .A2(n11287), .ZN(n12506) );
  NAND2_X1 U11368 ( .A1(n11286), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15019) );
  AND2_X1 U11369 ( .A1(n10031), .A2(n14850), .ZN(n10032) );
  AOI21_X1 U11370 ( .B1(n9834), .B2(n10113), .A(n9802), .ZN(n12468) );
  NAND2_X1 U11371 ( .A1(n15016), .A2(n10108), .ZN(n10113) );
  AND2_X1 U11372 ( .A1(n15247), .A2(n11285), .ZN(n15225) );
  AND2_X1 U11373 ( .A1(n9915), .A2(n16230), .ZN(n15072) );
  NAND2_X1 U11374 ( .A1(n14221), .A2(n14222), .ZN(n14211) );
  OAI21_X1 U11375 ( .B1(n12811), .B2(n12810), .A(n14848), .ZN(n14857) );
  AND2_X1 U11376 ( .A1(n11284), .A2(n15241), .ZN(n15247) );
  INV_X1 U11377 ( .A(n11296), .ZN(n15077) );
  NAND2_X1 U11378 ( .A1(n9920), .A2(n9855), .ZN(n11296) );
  NAND2_X1 U11379 ( .A1(n10075), .A2(n10074), .ZN(n14331) );
  NAND2_X1 U11380 ( .A1(n10119), .A2(n9921), .ZN(n9920) );
  OAI22_X1 U11381 ( .A1(n12463), .A2(n19986), .B1(n20000), .B2(n14112), .ZN(
        n12464) );
  NAND2_X1 U11382 ( .A1(n14869), .A2(n12765), .ZN(n12785) );
  XNOR2_X1 U11383 ( .A(n9889), .B(n14177), .ZN(n14566) );
  OAI21_X1 U11384 ( .B1(n19503), .B2(n19481), .A(n19683), .ZN(n19506) );
  OAI21_X1 U11385 ( .B1(n17520), .B2(n16453), .A(n16452), .ZN(n16454) );
  OAI211_X1 U11386 ( .C1(n14840), .C2(n16299), .A(n11280), .B(n11279), .ZN(
        n11281) );
  NAND2_X1 U11387 ( .A1(n10917), .A2(n11009), .ZN(n14168) );
  NAND2_X1 U11388 ( .A1(n14544), .A2(n11738), .ZN(n14532) );
  OR2_X1 U11389 ( .A1(n14062), .A2(n14061), .ZN(n14063) );
  NAND2_X1 U11390 ( .A1(n10582), .A2(n10581), .ZN(n13853) );
  NAND2_X1 U11391 ( .A1(n19689), .A2(n19688), .ZN(n19714) );
  AND2_X1 U11392 ( .A1(n14892), .A2(n12713), .ZN(n12714) );
  XOR2_X1 U11393 ( .A(n11009), .B(n11008), .Z(n14840) );
  OR2_X1 U11394 ( .A1(n10913), .A2(n14843), .ZN(n16124) );
  AND2_X1 U11395 ( .A1(n9833), .A2(n11874), .ZN(n9803) );
  XNOR2_X1 U11396 ( .A(n12712), .B(n12737), .ZN(n14884) );
  NAND2_X1 U11397 ( .A1(n20040), .A2(n11689), .ZN(n15943) );
  NAND2_X1 U11398 ( .A1(n14842), .A2(n9957), .ZN(n11009) );
  AND2_X1 U11399 ( .A1(n11873), .A2(n10073), .ZN(n9833) );
  AND2_X1 U11400 ( .A1(n12879), .A2(n14915), .ZN(n16122) );
  XNOR2_X1 U11401 ( .A(n10807), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16274) );
  AND2_X1 U11402 ( .A1(n11709), .A2(n11708), .ZN(n15937) );
  AND2_X1 U11403 ( .A1(n14460), .A2(n11728), .ZN(n13845) );
  NOR2_X2 U11404 ( .A1(n9815), .A2(n12475), .ZN(n14842) );
  INV_X1 U11405 ( .A(n13594), .ZN(n11873) );
  OR2_X1 U11406 ( .A1(n9773), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n9778) );
  OR2_X1 U11407 ( .A1(n10810), .A2(n11055), .ZN(n10807) );
  OR2_X1 U11408 ( .A1(n10790), .A2(n13867), .ZN(n13855) );
  OAI21_X1 U11409 ( .B1(n10791), .B2(n10808), .A(n19027), .ZN(n10622) );
  NOR2_X1 U11410 ( .A1(n10745), .A2(n10744), .ZN(n10947) );
  INV_X1 U11411 ( .A(n19756), .ZN(n19743) );
  NAND2_X1 U11412 ( .A1(n19607), .A2(n19850), .ZN(n19598) );
  NOR2_X1 U11413 ( .A1(n17551), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17550) );
  NOR2_X2 U11414 ( .A1(n19419), .A2(n19650), .ZN(n19409) );
  OR2_X1 U11415 ( .A1(n10736), .A2(n10735), .ZN(n10745) );
  NOR2_X1 U11416 ( .A1(n19651), .A2(n19650), .ZN(n19713) );
  OR2_X1 U11417 ( .A1(n10739), .A2(n10896), .ZN(n14994) );
  AND2_X1 U11418 ( .A1(n13464), .A2(n13465), .ZN(n13574) );
  OR2_X2 U11419 ( .A1(n11703), .A2(n11702), .ZN(n11716) );
  NAND2_X1 U11420 ( .A1(n14950), .A2(n9865), .ZN(n14928) );
  AND2_X1 U11421 ( .A1(n11703), .A2(n11692), .ZN(n11872) );
  AND2_X1 U11422 ( .A1(n19854), .A2(n19881), .ZN(n19316) );
  OAI21_X1 U11423 ( .B1(n11858), .B2(n11770), .A(n11687), .ZN(n11688) );
  OR2_X1 U11424 ( .A1(n10690), .A2(n9938), .ZN(n10107) );
  NAND2_X1 U11425 ( .A1(n13609), .A2(n9859), .ZN(n13581) );
  OAI21_X1 U11426 ( .B1(n20107), .B2(n12062), .A(n11829), .ZN(n13464) );
  AND2_X1 U11427 ( .A1(n10512), .A2(n10511), .ZN(n10515) );
  AND2_X1 U11428 ( .A1(n10720), .A2(n10716), .ZN(n16144) );
  NAND2_X1 U11429 ( .A1(n10619), .A2(n10618), .ZN(n10800) );
  OR3_X1 U11430 ( .A1(n10600), .A2(n10599), .A3(n10598), .ZN(n10619) );
  NAND2_X1 U11431 ( .A1(n13259), .A2(n13264), .ZN(n19864) );
  NAND2_X1 U11432 ( .A1(n17995), .A2(n9754), .ZN(n17685) );
  AOI21_X1 U11433 ( .B1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n10490), .A(
        n10356), .ZN(n10379) );
  NAND2_X1 U11434 ( .A1(n13259), .A2(n12534), .ZN(n13605) );
  AND4_X1 U11435 ( .A1(n10429), .A2(n10428), .A3(n10427), .A4(n10426), .ZN(
        n10435) );
  OR2_X1 U11436 ( .A1(n10695), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15036) );
  NOR2_X1 U11437 ( .A1(n10711), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10726) );
  NOR2_X1 U11438 ( .A1(n17037), .A2(n17038), .ZN(n17010) );
  OR2_X1 U11439 ( .A1(n10710), .A2(n10709), .ZN(n10711) );
  AND2_X1 U11440 ( .A1(n10697), .A2(n12500), .ZN(n15026) );
  NOR2_X2 U11441 ( .A1(n14380), .A2(n12413), .ZN(n14372) );
  NAND2_X1 U11442 ( .A1(n17721), .A2(n17995), .ZN(n15685) );
  NAND2_X1 U11443 ( .A1(n19214), .A2(n19213), .ZN(n16294) );
  OR2_X1 U11444 ( .A1(n10683), .A2(n10701), .ZN(n14748) );
  AND2_X1 U11445 ( .A1(n18946), .A2(n10808), .ZN(n10696) );
  AND2_X1 U11446 ( .A1(n13626), .A2(n10361), .ZN(n19640) );
  AND2_X1 U11447 ( .A1(n13626), .A2(n10362), .ZN(n19573) );
  AND2_X1 U11448 ( .A1(n10668), .A2(n10669), .ZN(n18946) );
  OR2_X1 U11449 ( .A1(n10371), .A2(n10370), .ZN(n10485) );
  CLKBUF_X1 U11450 ( .A(n14089), .Z(n14441) );
  NAND4_X1 U11451 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(P3_EBX_REG_17__SCAN_IN), 
        .A3(P3_EBX_REG_16__SCAN_IN), .A4(n17101), .ZN(n17065) );
  AND2_X1 U11452 ( .A1(n13262), .A2(n13261), .ZN(n12530) );
  NAND2_X1 U11453 ( .A1(n11609), .A2(n11608), .ZN(n13471) );
  NAND2_X1 U11454 ( .A1(n11558), .A2(n11546), .ZN(n11838) );
  NAND2_X1 U11455 ( .A1(n10674), .A2(n10673), .ZN(n10676) );
  INV_X1 U11456 ( .A(n17078), .ZN(n17101) );
  NAND2_X1 U11457 ( .A1(n13171), .A2(n13170), .ZN(n13262) );
  AND2_X1 U11458 ( .A1(n10674), .A2(n9941), .ZN(n10682) );
  INV_X2 U11459 ( .A(n13356), .ZN(n9761) );
  AND2_X1 U11460 ( .A1(n13216), .A2(n10349), .ZN(n10359) );
  NAND2_X1 U11461 ( .A1(n11575), .A2(n11574), .ZN(n11590) );
  OR2_X1 U11462 ( .A1(n11575), .A2(n11574), .ZN(n10005) );
  NOR2_X2 U11463 ( .A1(n9788), .A2(n19278), .ZN(n19247) );
  AND2_X1 U11464 ( .A1(n9829), .A2(n17795), .ZN(n17754) );
  NAND2_X1 U11465 ( .A1(n11564), .A2(n11563), .ZN(n11575) );
  NOR2_X1 U11466 ( .A1(n13207), .A2(n13643), .ZN(n19078) );
  AND2_X1 U11467 ( .A1(n16074), .A2(n16073), .ZN(n16076) );
  OR2_X1 U11468 ( .A1(n13807), .A2(n9960), .ZN(n9959) );
  XNOR2_X1 U11469 ( .A(n10820), .B(n10819), .ZN(n10817) );
  OAI21_X1 U11470 ( .B1(n18672), .B2(n15646), .A(n18671), .ZN(n18692) );
  OR2_X1 U11471 ( .A1(n10640), .A2(n19265), .ZN(n10729) );
  CLKBUF_X1 U11472 ( .A(n13045), .Z(n13118) );
  INV_X1 U11473 ( .A(n10333), .ZN(n10907) );
  NOR2_X2 U11474 ( .A1(n21019), .A2(n17201), .ZN(n17202) );
  OR2_X1 U11475 ( .A1(n13003), .A2(n9974), .ZN(n15646) );
  NAND2_X1 U11476 ( .A1(n13133), .A2(n13142), .ZN(n13243) );
  NOR2_X1 U11477 ( .A1(n9937), .A2(n10576), .ZN(n10631) );
  NOR2_X1 U11478 ( .A1(n11471), .A2(n13198), .ZN(n11493) );
  NAND2_X1 U11479 ( .A1(n17852), .A2(n15616), .ZN(n17840) );
  XNOR2_X1 U11480 ( .A(n11028), .B(n11029), .ZN(n13446) );
  AND2_X1 U11481 ( .A1(n10288), .A2(n10287), .ZN(n11254) );
  NAND2_X1 U11482 ( .A1(n17853), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n17852) );
  NAND2_X2 U11483 ( .A1(n10288), .A2(n9770), .ZN(n10297) );
  NOR2_X1 U11484 ( .A1(n10094), .A2(n17824), .ZN(n10093) );
  OAI21_X1 U11485 ( .B1(n13221), .B2(n11195), .A(n11021), .ZN(n13209) );
  NOR2_X1 U11486 ( .A1(n12035), .A2(n14033), .ZN(n12020) );
  INV_X1 U11487 ( .A(n10905), .ZN(n10823) );
  NOR2_X1 U11488 ( .A1(n18232), .A2(n13014), .ZN(n13921) );
  INV_X1 U11489 ( .A(n10905), .ZN(n9762) );
  NAND2_X1 U11490 ( .A1(n17862), .A2(n15611), .ZN(n15614) );
  NAND2_X1 U11491 ( .A1(n14666), .A2(n11013), .ZN(n10926) );
  NOR2_X1 U11492 ( .A1(n17381), .A2(n15590), .ZN(n15618) );
  AND2_X2 U11494 ( .A1(n10273), .A2(n10013), .ZN(n10953) );
  INV_X1 U11495 ( .A(n10254), .ZN(n10992) );
  INV_X1 U11496 ( .A(n17267), .ZN(n18247) );
  NAND2_X2 U11497 ( .A1(n9789), .A2(n10274), .ZN(n10279) );
  NAND2_X1 U11498 ( .A1(n11777), .A2(n11597), .ZN(n11814) );
  BUF_X2 U11499 ( .A(n11014), .Z(n9789) );
  CLKBUF_X1 U11500 ( .A(n10539), .Z(n10742) );
  NAND3_X1 U11501 ( .A1(n13002), .A2(n13001), .A3(n13000), .ZN(n16394) );
  INV_X1 U11502 ( .A(n10268), .ZN(n10282) );
  CLKBUF_X3 U11503 ( .A(n11014), .Z(n9790) );
  INV_X1 U11504 ( .A(n20842), .ZN(n15742) );
  NAND3_X1 U11505 ( .A1(n12953), .A2(n12952), .A3(n12951), .ZN(n17267) );
  NAND3_X1 U11506 ( .A1(n12991), .A2(n12990), .A3(n12989), .ZN(n15635) );
  NAND2_X1 U11507 ( .A1(n13183), .A2(n12355), .ZN(n13685) );
  NAND2_X1 U11508 ( .A1(n13291), .A2(n11464), .ZN(n20842) );
  NOR2_X2 U11509 ( .A1(n12963), .A2(n12962), .ZN(n18232) );
  AOI211_X1 U11510 ( .C1(n17215), .C2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n12950), .B(n12949), .ZN(n12951) );
  AOI211_X1 U11511 ( .C1(n17213), .C2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A(
        n12999), .B(n12998), .ZN(n13000) );
  CLKBUF_X3 U11512 ( .A(n12460), .Z(n9787) );
  INV_X2 U11513 ( .A(U212), .ZN(n16509) );
  NAND2_X1 U11514 ( .A1(n10170), .A2(n10169), .ZN(n10265) );
  OR2_X1 U11515 ( .A1(n15606), .A2(n15607), .ZN(n15774) );
  AOI211_X1 U11516 ( .C1(n17224), .C2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n12930), .B(n12929), .ZN(n12931) );
  INV_X1 U11517 ( .A(n12355), .ZN(n13291) );
  NOR2_X1 U11518 ( .A1(n11464), .A2(n12355), .ZN(n13677) );
  OR2_X2 U11519 ( .A1(n16510), .A2(n16468), .ZN(n16512) );
  AND4_X1 U11520 ( .A1(n15549), .A2(n15544), .A3(n15548), .A4(n15547), .ZN(
        n15648) );
  OAI21_X1 U11521 ( .B1(n9918), .B2(n9917), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9919) );
  NAND2_X1 U11522 ( .A1(n9749), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11202) );
  AND4_X1 U11523 ( .A1(n11437), .A2(n11436), .A3(n11435), .A4(n11434), .ZN(
        n11444) );
  AND2_X2 U11524 ( .A1(n9759), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10467) );
  AND4_X1 U11525 ( .A1(n11339), .A2(n11338), .A3(n11337), .A4(n11336), .ZN(
        n11345) );
  AND4_X1 U11526 ( .A1(n11442), .A2(n11441), .A3(n11440), .A4(n11439), .ZN(
        n11443) );
  AND4_X1 U11527 ( .A1(n11363), .A2(n11362), .A3(n11361), .A4(n11360), .ZN(
        n11364) );
  AND4_X1 U11528 ( .A1(n11331), .A2(n11330), .A3(n11329), .A4(n11328), .ZN(
        n11347) );
  AND4_X1 U11529 ( .A1(n11335), .A2(n11334), .A3(n11333), .A4(n11332), .ZN(
        n11346) );
  AND4_X1 U11530 ( .A1(n11411), .A2(n11410), .A3(n11409), .A4(n11408), .ZN(
        n11424) );
  AND4_X1 U11531 ( .A1(n11429), .A2(n11428), .A3(n11427), .A4(n11426), .ZN(
        n11446) );
  AND4_X1 U11532 ( .A1(n11416), .A2(n11415), .A3(n11414), .A4(n11413), .ZN(
        n11423) );
  AND4_X1 U11533 ( .A1(n11421), .A2(n11420), .A3(n11419), .A4(n11418), .ZN(
        n11422) );
  AND4_X1 U11534 ( .A1(n11351), .A2(n11350), .A3(n11349), .A4(n11348), .ZN(
        n11366) );
  INV_X2 U11535 ( .A(n13645), .ZN(n13643) );
  AND4_X1 U11536 ( .A1(n11407), .A2(n11406), .A3(n11405), .A4(n11404), .ZN(
        n11425) );
  BUF_X2 U11537 ( .A(n11379), .Z(n12329) );
  BUF_X2 U11538 ( .A(n15560), .Z(n17117) );
  BUF_X4 U11539 ( .A(n15559), .Z(n17208) );
  INV_X2 U11540 ( .A(n16045), .ZN(n20099) );
  INV_X2 U11541 ( .A(n18749), .ZN(n18801) );
  NAND2_X2 U11542 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19891), .ZN(n19835) );
  NAND2_X2 U11543 ( .A1(n19891), .A2(n19792), .ZN(n19839) );
  BUF_X2 U11544 ( .A(n17176), .Z(n17206) );
  CLKBUF_X3 U11545 ( .A(n15538), .Z(n17217) );
  AND2_X2 U11546 ( .A1(n15382), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10171) );
  AND2_X1 U11547 ( .A1(n12862), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10205) );
  INV_X2 U11548 ( .A(n10185), .ZN(n12720) );
  OR2_X1 U11549 ( .A1(n12922), .A2(n16921), .ZN(n15562) );
  NOR2_X4 U11550 ( .A1(n13030), .A2(n12921), .ZN(n15600) );
  BUF_X4 U11551 ( .A(n15553), .Z(n9763) );
  INV_X2 U11552 ( .A(n18882), .ZN(n18864) );
  BUF_X4 U11553 ( .A(n15435), .Z(n9764) );
  INV_X2 U11554 ( .A(n16550), .ZN(n16552) );
  OR3_X2 U11555 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), 
        .A3(n18837), .ZN(n15697) );
  NAND2_X1 U11556 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18826), .ZN(
        n12922) );
  AND2_X2 U11557 ( .A1(n11313), .A2(n13388), .ZN(n11501) );
  AND2_X1 U11558 ( .A1(n10101), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10385) );
  NOR2_X1 U11559 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10144) );
  AND2_X2 U11560 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10388) );
  NOR2_X1 U11561 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12672) );
  NAND2_X1 U11562 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16921) );
  INV_X1 U11563 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18826) );
  AND2_X2 U11565 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13393) );
  NAND2_X1 U11566 ( .A1(n13560), .A2(n13559), .ZN(n9765) );
  INV_X1 U11567 ( .A(n10011), .ZN(n9766) );
  NAND2_X1 U11568 ( .A1(n9905), .A2(n9903), .ZN(n10331) );
  AND2_X1 U11569 ( .A1(n13471), .A2(n11652), .ZN(n9767) );
  NAND2_X1 U11570 ( .A1(n11589), .A2(n11652), .ZN(n9768) );
  OR2_X1 U11571 ( .A1(n11545), .A2(n11544), .ZN(n9769) );
  NAND2_X1 U11572 ( .A1(n12355), .A2(n20145), .ZN(n12460) );
  XNOR2_X1 U11573 ( .A(n11716), .B(n11715), .ZN(n11880) );
  AND2_X1 U11574 ( .A1(n10287), .A2(n10999), .ZN(n9770) );
  AND2_X1 U11575 ( .A1(n10986), .A2(n10280), .ZN(n10288) );
  NAND2_X1 U11576 ( .A1(n10926), .A2(n10279), .ZN(n10986) );
  AND2_X1 U11577 ( .A1(n14460), .A2(n14603), .ZN(n9771) );
  AND2_X2 U11578 ( .A1(n11313), .A2(n13388), .ZN(n9772) );
  AND2_X1 U11579 ( .A1(n10514), .A2(n10788), .ZN(n9773) );
  NAND2_X1 U11581 ( .A1(n10789), .A2(n13866), .ZN(n9775) );
  AND2_X1 U11582 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9776) );
  NAND2_X1 U11583 ( .A1(n11755), .A2(n11754), .ZN(n14511) );
  NOR2_X1 U11584 ( .A1(n14211), .A2(n10084), .ZN(n14186) );
  OR3_X2 U11585 ( .A1(n14211), .A2(n10084), .A3(n10083), .ZN(n9797) );
  NAND2_X1 U11586 ( .A1(n13621), .A2(n9779), .ZN(n9777) );
  AND2_X1 U11587 ( .A1(n10785), .A2(n13755), .ZN(n9779) );
  NOR2_X2 U11588 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n15695), .ZN(
        n16462) );
  OAI21_X2 U11589 ( .B1(n13622), .B2(n10808), .A(n14163), .ZN(n13614) );
  NAND2_X1 U11590 ( .A1(n11751), .A2(n11750), .ZN(n14526) );
  XNOR2_X1 U11591 ( .A(n11763), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14586) );
  INV_X1 U11592 ( .A(n9781), .ZN(n15089) );
  INV_X4 U11593 ( .A(n12350), .ZN(n11473) );
  AND2_X2 U11594 ( .A1(n15098), .A2(n11264), .ZN(n9781) );
  NAND2_X2 U11595 ( .A1(n10786), .A2(n10021), .ZN(n13622) );
  NOR2_X2 U11596 ( .A1(n15256), .A2(n15257), .ZN(n13886) );
  NOR2_X2 U11597 ( .A1(n14790), .A2(n14792), .ZN(n14791) );
  NAND2_X1 U11598 ( .A1(n10806), .A2(n10805), .ZN(n15106) );
  AND2_X2 U11599 ( .A1(n15384), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10387) );
  NOR4_X1 U11601 ( .A1(n18221), .A2(n13917), .A3(n17267), .A4(n15635), .ZN(
        n17463) );
  OAI21_X2 U11602 ( .B1(n14300), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11555), 
        .ZN(n11837) );
  AND2_X1 U11603 ( .A1(n13617), .A2(n10358), .ZN(n19287) );
  AND2_X1 U11604 ( .A1(n13617), .A2(n10362), .ZN(n19348) );
  NOR2_X1 U11606 ( .A1(n10369), .A2(n10374), .ZN(n19483) );
  INV_X1 U11607 ( .A(n12317), .ZN(n9784) );
  AND2_X1 U11608 ( .A1(n13411), .A2(n13392), .ZN(n11417) );
  AND2_X4 U11609 ( .A1(n10387), .A2(n9780), .ZN(n10243) );
  AND2_X2 U11610 ( .A1(n13626), .A2(n10363), .ZN(n10476) );
  OR2_X1 U11611 ( .A1(n10341), .A2(n10340), .ZN(n10342) );
  AND2_X4 U11612 ( .A1(n11312), .A2(n13388), .ZN(n11438) );
  NAND2_X2 U11613 ( .A1(n11253), .A2(n10313), .ZN(n11010) );
  NOR2_X2 U11614 ( .A1(n10328), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15382) );
  NAND2_X2 U11615 ( .A1(n10157), .A2(n10156), .ZN(n10539) );
  AOI21_X1 U11616 ( .B1(n10477), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A(n9788), .ZN(n10355) );
  AND2_X2 U11617 ( .A1(n10358), .A2(n10351), .ZN(n10477) );
  AND2_X2 U11618 ( .A1(n10363), .A2(n13617), .ZN(n10478) );
  AOI21_X1 U11619 ( .B1(n10822), .B2(n10818), .A(n10821), .ZN(n13760) );
  NOR2_X2 U11620 ( .A1(n10375), .A2(n13313), .ZN(n10490) );
  INV_X2 U11621 ( .A(n10252), .ZN(n10251) );
  NAND2_X2 U11622 ( .A1(n10953), .A2(n10274), .ZN(n10312) );
  NAND2_X2 U11623 ( .A1(n15007), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13951) );
  NOR2_X2 U11624 ( .A1(n15006), .A2(n15180), .ZN(n15007) );
  OAI211_X2 U11625 ( .C1(n9794), .C2(n13219), .A(n10310), .B(n10309), .ZN(
        n10338) );
  NAND3_X2 U11626 ( .A1(n16362), .A2(n10298), .A3(n10297), .ZN(n10299) );
  OAI21_X2 U11627 ( .B1(n15370), .B2(n9793), .A(n10319), .ZN(n10346) );
  AND2_X2 U11628 ( .A1(n15382), .A2(n10101), .ZN(n10158) );
  AND2_X2 U11629 ( .A1(n10979), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10981) );
  NOR2_X4 U11630 ( .A1(n14050), .A2(n14067), .ZN(n10979) );
  NAND2_X2 U11631 ( .A1(n13953), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14050) );
  NOR2_X4 U11632 ( .A1(n13951), .A2(n10896), .ZN(n13953) );
  OAI21_X1 U11633 ( .B1(n14126), .B2(n12523), .A(n12522), .ZN(n15355) );
  OAI21_X2 U11634 ( .B1(n10338), .B2(n10336), .A(n10348), .ZN(n14126) );
  NAND2_X1 U11635 ( .A1(n10299), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9793) );
  NAND2_X1 U11636 ( .A1(n10299), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9794) );
  NAND2_X4 U11637 ( .A1(n10299), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10333) );
  INV_X2 U11638 ( .A(n10185), .ZN(n9795) );
  NAND2_X1 U11639 ( .A1(n11622), .A2(n11682), .ZN(n11691) );
  INV_X1 U11640 ( .A(n12654), .ZN(n12706) );
  INV_X1 U11641 ( .A(n15402), .ZN(n12690) );
  INV_X1 U11642 ( .A(n10514), .ZN(n10513) );
  OAI21_X1 U11643 ( .B1(n14477), .B2(n13968), .A(n15893), .ZN(n14469) );
  AND2_X1 U11644 ( .A1(n11474), .A2(n11456), .ZN(n11485) );
  NAND2_X1 U11645 ( .A1(n11637), .A2(n11636), .ZN(n11703) );
  INV_X1 U11646 ( .A(n11690), .ZN(n11636) );
  AOI21_X1 U11647 ( .B1(n19861), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n10556), .ZN(n10754) );
  NOR2_X1 U11648 ( .A1(n10555), .A2(n10554), .ZN(n10556) );
  INV_X1 U11649 ( .A(n10553), .ZN(n10555) );
  NAND2_X1 U11650 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n12916), .ZN(
        n12924) );
  AND2_X1 U11651 ( .A1(n12072), .A2(n10082), .ZN(n10081) );
  INV_X1 U11652 ( .A(n14346), .ZN(n10082) );
  INV_X1 U11653 ( .A(n12340), .ZN(n12345) );
  OR2_X1 U11654 ( .A1(n11456), .A2(n20742), .ZN(n12343) );
  INV_X1 U11655 ( .A(n13671), .ZN(n12340) );
  NOR2_X2 U11656 ( .A1(n11473), .A2(n20742), .ZN(n12044) );
  NAND2_X1 U11657 ( .A1(n14553), .A2(n11734), .ZN(n14009) );
  OR2_X1 U11658 ( .A1(n20152), .A2(n11495), .ZN(n11777) );
  NAND2_X1 U11659 ( .A1(n10631), .A2(n10630), .ZN(n10640) );
  NAND2_X1 U11660 ( .A1(n14863), .A2(n10121), .ZN(n12811) );
  AND2_X1 U11661 ( .A1(n10043), .A2(n14891), .ZN(n10042) );
  OAI211_X1 U11662 ( .C1(n10300), .C2(n10991), .A(n10275), .B(n10312), .ZN(
        n10302) );
  AND2_X1 U11663 ( .A1(n10257), .A2(n10999), .ZN(n10277) );
  NAND2_X1 U11664 ( .A1(n9847), .A2(n10058), .ZN(n10057) );
  INV_X1 U11665 ( .A(n14754), .ZN(n10058) );
  INV_X1 U11666 ( .A(n11195), .ZN(n11223) );
  NAND2_X1 U11667 ( .A1(n10065), .A2(n13864), .ZN(n10064) );
  INV_X1 U11668 ( .A(n13606), .ZN(n10065) );
  NAND2_X1 U11669 ( .A1(n10517), .A2(n10799), .ZN(n10790) );
  AND4_X1 U11670 ( .A1(n10460), .A2(n10459), .A3(n10458), .A4(n10457), .ZN(
        n10475) );
  NAND2_X1 U11671 ( .A1(n9925), .A2(n10453), .ZN(n10562) );
  NAND2_X1 U11672 ( .A1(n9926), .A2(n10425), .ZN(n10561) );
  NAND2_X1 U11673 ( .A1(n12878), .A2(n10268), .ZN(n10286) );
  NOR2_X1 U11674 ( .A1(n10266), .A2(n10268), .ZN(n10999) );
  AOI221_X1 U11675 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n10754), 
        .C1(n15505), .C2(n10754), .A(n10753), .ZN(n10936) );
  NOR2_X1 U11676 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15769), .ZN(
        n10753) );
  INV_X1 U11677 ( .A(n15551), .ZN(n15594) );
  INV_X1 U11678 ( .A(n15537), .ZN(n17175) );
  NAND2_X1 U11679 ( .A1(n13018), .A2(n18826), .ZN(n12921) );
  NAND2_X1 U11680 ( .A1(n13429), .A2(n11857), .ZN(n13465) );
  AND2_X1 U11681 ( .A1(n15747), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13317) );
  AND2_X1 U11682 ( .A1(n20742), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14083) );
  INV_X1 U11683 ( .A(n14329), .ZN(n10074) );
  INV_X1 U11684 ( .A(n14328), .ZN(n10075) );
  NAND2_X1 U11685 ( .A1(n14460), .A2(n14588), .ZN(n9994) );
  AOI21_X1 U11686 ( .B1(n14511), .B2(n15893), .A(n10002), .ZN(n10001) );
  INV_X1 U11687 ( .A(n10003), .ZN(n10002) );
  AOI21_X1 U11688 ( .B1(n15893), .B2(n9813), .A(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n10003) );
  INV_X1 U11689 ( .A(n11249), .ZN(n11251) );
  INV_X1 U11690 ( .A(n14850), .ZN(n10030) );
  NAND2_X1 U11691 ( .A1(n10107), .A2(n9831), .ZN(n10104) );
  AND4_X1 U11692 ( .A1(n10522), .A2(n10521), .A3(n10520), .A4(n10519), .ZN(
        n10537) );
  AND4_X1 U11693 ( .A1(n10526), .A2(n10525), .A3(n10524), .A4(n10523), .ZN(
        n10536) );
  NAND2_X1 U11694 ( .A1(n9805), .A2(n9916), .ZN(n9911) );
  INV_X1 U11695 ( .A(n15070), .ZN(n9914) );
  AOI21_X1 U11696 ( .B1(n18684), .B2(n13931), .A(n9987), .ZN(n15771) );
  OR2_X1 U11697 ( .A1(n18660), .A2(n18870), .ZN(n9987) );
  NAND2_X1 U11698 ( .A1(n10089), .A2(n10092), .ZN(n10088) );
  NAND2_X1 U11699 ( .A1(n15617), .A2(n18145), .ZN(n10092) );
  INV_X1 U11700 ( .A(n10093), .ZN(n10089) );
  AND2_X1 U11701 ( .A1(n20001), .A2(n13325), .ZN(n14440) );
  OR2_X1 U11702 ( .A1(n13023), .A2(n13024), .ZN(n13019) );
  NAND2_X1 U11703 ( .A1(n11768), .A2(n11767), .ZN(n11772) );
  NAND2_X1 U11704 ( .A1(n11675), .A2(n11683), .ZN(n11684) );
  NAND2_X1 U11705 ( .A1(n11822), .A2(n12350), .ZN(n11475) );
  NOR2_X1 U11706 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20105), .ZN(
        n11811) );
  INV_X1 U11707 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11549) );
  NAND2_X1 U11708 ( .A1(n9822), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11560) );
  AND2_X1 U11709 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n9928) );
  NOR2_X1 U11710 ( .A1(n9873), .A2(n9934), .ZN(n12776) );
  AND2_X1 U11711 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n9934) );
  NAND2_X1 U11712 ( .A1(n10051), .A2(n14741), .ZN(n10050) );
  INV_X1 U11713 ( .A(n12498), .ZN(n10051) );
  NAND2_X1 U11714 ( .A1(n10254), .A2(n10282), .ZN(n10255) );
  AOI22_X1 U11715 ( .A1(n9753), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10243), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10240) );
  AOI22_X1 U11716 ( .A1(n9752), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10243), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10245) );
  XNOR2_X1 U11717 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10765) );
  NOR2_X1 U11718 ( .A1(n18874), .A2(n9796), .ZN(n13016) );
  OR2_X1 U11719 ( .A1(n13195), .A2(n12353), .ZN(n13147) );
  AND2_X1 U11720 ( .A1(n12070), .A2(n14358), .ZN(n14274) );
  OR2_X1 U11721 ( .A1(n11669), .A2(n11671), .ZN(n11672) );
  OR2_X1 U11722 ( .A1(n11607), .A2(n11606), .ZN(n11694) );
  NAND2_X1 U11723 ( .A1(n20258), .A2(n11552), .ZN(n11564) );
  OR2_X1 U11724 ( .A1(n11464), .A2(n11495), .ZN(n11597) );
  NOR2_X1 U11725 ( .A1(n11585), .A2(n11584), .ZN(n11677) );
  NAND3_X1 U11726 ( .A1(n20152), .A2(n11464), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11809) );
  NAND2_X1 U11727 ( .A1(n11596), .A2(n11595), .ZN(n20295) );
  INV_X1 U11728 ( .A(n10671), .ZN(n9944) );
  NAND2_X1 U11729 ( .A1(n10682), .A2(n14903), .ZN(n10703) );
  NAND2_X1 U11730 ( .A1(n10666), .A2(n10729), .ZN(n10674) );
  NAND2_X1 U11731 ( .A1(n9955), .A2(n9954), .ZN(n10666) );
  INV_X1 U11732 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n9954) );
  INV_X1 U11733 ( .A(n10664), .ZN(n9955) );
  NAND2_X1 U11734 ( .A1(n10651), .A2(n10654), .ZN(n10680) );
  NAND2_X1 U11735 ( .A1(n12764), .A2(n12759), .ZN(n12765) );
  INV_X1 U11736 ( .A(n14875), .ZN(n10038) );
  NAND2_X1 U11737 ( .A1(n10053), .A2(n14971), .ZN(n10052) );
  INV_X1 U11738 ( .A(n15234), .ZN(n10053) );
  INV_X1 U11739 ( .A(n13905), .ZN(n10044) );
  NOR2_X1 U11740 ( .A1(n21034), .A2(n10067), .ZN(n10066) );
  INV_X1 U11741 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10067) );
  NOR2_X1 U11742 ( .A1(n15100), .A2(n10061), .ZN(n10060) );
  INV_X1 U11743 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10061) );
  NOR2_X1 U11744 ( .A1(n19211), .A2(n10071), .ZN(n10070) );
  INV_X1 U11745 ( .A(n14131), .ZN(n10069) );
  AND2_X1 U11746 ( .A1(n13383), .A2(n13759), .ZN(n9968) );
  OAI21_X1 U11747 ( .B1(n10332), .B2(n9780), .A(n10330), .ZN(n9904) );
  AND2_X1 U11748 ( .A1(n15502), .A2(n10313), .ZN(n10298) );
  AND2_X1 U11749 ( .A1(n13945), .A2(n14878), .ZN(n9970) );
  NAND2_X1 U11750 ( .A1(n13577), .A2(n9962), .ZN(n13780) );
  AND2_X1 U11751 ( .A1(n9828), .A2(n13781), .ZN(n9962) );
  INV_X1 U11752 ( .A(n16238), .ZN(n9923) );
  NOR2_X1 U11753 ( .A1(n10115), .A2(n10120), .ZN(n10114) );
  INV_X1 U11754 ( .A(n9867), .ZN(n10120) );
  INV_X1 U11755 ( .A(n10117), .ZN(n10115) );
  INV_X1 U11756 ( .A(n10799), .ZN(n10802) );
  NOR2_X1 U11757 ( .A1(n16277), .A2(n10118), .ZN(n10117) );
  INV_X1 U11758 ( .A(n15304), .ZN(n10118) );
  NAND2_X1 U11759 ( .A1(n15324), .A2(n15323), .ZN(n14808) );
  NAND2_X1 U11760 ( .A1(n10045), .A2(n10798), .ZN(n10803) );
  AND4_X1 U11761 ( .A1(n10605), .A2(n10604), .A3(n10603), .A4(n10602), .ZN(
        n10616) );
  AND4_X1 U11762 ( .A1(n10612), .A2(n10611), .A3(n10610), .A4(n10609), .ZN(
        n10615) );
  AND2_X1 U11763 ( .A1(n10453), .A2(n11044), .ZN(n9924) );
  INV_X1 U11764 ( .A(n10562), .ZN(n10454) );
  INV_X1 U11765 ( .A(n10561), .ZN(n10455) );
  NOR2_X1 U11766 ( .A1(n12541), .A2(n12521), .ZN(n12533) );
  AND2_X1 U11767 ( .A1(n13265), .A2(n10359), .ZN(n10361) );
  OAI21_X1 U11768 ( .B1(n10192), .B2(n10191), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10199) );
  NOR2_X1 U11769 ( .A1(n19785), .A2(n14667), .ZN(n15359) );
  NAND2_X1 U11770 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19886), .ZN(
        n10755) );
  AND2_X1 U11771 ( .A1(n10766), .A2(n10752), .ZN(n10932) );
  OR2_X1 U11772 ( .A1(n15564), .A2(n15563), .ZN(n15565) );
  NAND2_X1 U11773 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12920) );
  NAND2_X1 U11774 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13018), .ZN(
        n12923) );
  NAND2_X1 U11775 ( .A1(n17811), .A2(n15620), .ZN(n15623) );
  OR2_X1 U11776 ( .A1(n13232), .A2(n13147), .ZN(n13190) );
  AND2_X1 U11777 ( .A1(n13389), .A2(n13178), .ZN(n13314) );
  INV_X1 U11778 ( .A(n13234), .ZN(n14088) );
  NOR3_X1 U11779 ( .A1(n13329), .A2(n13328), .A3(n13327), .ZN(n13331) );
  NAND2_X1 U11780 ( .A1(n12292), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13674) );
  AND2_X1 U11781 ( .A1(n12138), .A2(n12137), .ZN(n14335) );
  OR2_X1 U11782 ( .A1(n15797), .A2(n12340), .ZN(n12137) );
  AND2_X1 U11783 ( .A1(n10081), .A2(n14343), .ZN(n10080) );
  OR2_X1 U11784 ( .A1(n15892), .A2(n12340), .ZN(n12094) );
  NOR2_X1 U11785 ( .A1(n11918), .A2(n19921), .ZN(n11934) );
  AND3_X1 U11786 ( .A1(n11901), .A2(n11900), .A3(n11899), .ZN(n13789) );
  INV_X1 U11787 ( .A(n11875), .ZN(n11876) );
  NAND2_X1 U11788 ( .A1(n11876), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11881) );
  OR2_X1 U11789 ( .A1(n11836), .A2(n11835), .ZN(n13427) );
  AND2_X1 U11790 ( .A1(n13420), .A2(n12044), .ZN(n11836) );
  NAND2_X1 U11791 ( .A1(n13427), .A2(n11856), .ZN(n13429) );
  INV_X1 U11792 ( .A(n13431), .ZN(n11856) );
  NAND2_X1 U11793 ( .A1(n13232), .A2(n13317), .ZN(n13329) );
  NAND2_X1 U11794 ( .A1(n15893), .A2(n9881), .ZN(n9995) );
  INV_X1 U11795 ( .A(n14223), .ZN(n9884) );
  NAND2_X1 U11796 ( .A1(n14284), .A2(n14285), .ZN(n14353) );
  AND2_X1 U11797 ( .A1(n11650), .A2(n12351), .ZN(n11651) );
  INV_X1 U11798 ( .A(n13467), .ZN(n9886) );
  INV_X1 U11799 ( .A(n13468), .ZN(n9885) );
  NOR2_X1 U11800 ( .A1(n20214), .A2(n11846), .ZN(n20610) );
  AND2_X1 U11801 ( .A1(n20471), .A2(n20299), .ZN(n20649) );
  AND2_X1 U11802 ( .A1(n20214), .A2(n11846), .ZN(n20639) );
  AND2_X1 U11803 ( .A1(n13420), .A2(n13471), .ZN(n20679) );
  AND2_X1 U11804 ( .A1(n10985), .A2(n10984), .ZN(n15379) );
  INV_X1 U11805 ( .A(n10720), .ZN(n10949) );
  AOI21_X1 U11806 ( .B1(n14132), .B2(n18894), .A(n10049), .ZN(n14707) );
  AND2_X1 U11807 ( .A1(n10980), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10049) );
  OR2_X1 U11808 ( .A1(n13072), .A2(n13042), .ZN(n14137) );
  AND3_X1 U11809 ( .A1(n10136), .A2(n11151), .A3(n11150), .ZN(n13782) );
  NAND2_X1 U11810 ( .A1(n10023), .A2(n10025), .ZN(n10022) );
  AOI21_X1 U11811 ( .B1(n10029), .B2(n10034), .A(n10026), .ZN(n10025) );
  NAND2_X1 U11812 ( .A1(n12829), .A2(n10029), .ZN(n10023) );
  NAND2_X1 U11813 ( .A1(n14848), .A2(n14856), .ZN(n10031) );
  NAND2_X1 U11814 ( .A1(n14848), .A2(n14857), .ZN(n10033) );
  AOI21_X1 U11815 ( .B1(n9795), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A(n9930), 
        .ZN(n12816) );
  XNOR2_X1 U11816 ( .A(n12785), .B(n9875), .ZN(n14866) );
  NAND2_X1 U11817 ( .A1(n10258), .A2(n9755), .ZN(n12882) );
  INV_X1 U11818 ( .A(n13046), .ZN(n14143) );
  AND2_X1 U11819 ( .A1(n14681), .A2(n9878), .ZN(n14677) );
  NOR2_X1 U11820 ( .A1(n14708), .A2(n16155), .ZN(n14681) );
  NOR2_X1 U11821 ( .A1(n14697), .A2(n15084), .ZN(n14696) );
  NAND2_X1 U11822 ( .A1(n15105), .A2(n16326), .ZN(n10020) );
  AOI21_X1 U11823 ( .B1(n12472), .B2(n9880), .A(n9802), .ZN(n9946) );
  NOR2_X1 U11824 ( .A1(n12472), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9947) );
  NAND2_X1 U11825 ( .A1(n14950), .A2(n10072), .ZN(n14933) );
  INV_X1 U11826 ( .A(n11303), .ZN(n9940) );
  NAND2_X1 U11827 ( .A1(n11296), .A2(n10690), .ZN(n10106) );
  INV_X1 U11828 ( .A(n15035), .ZN(n11286) );
  AOI21_X1 U11829 ( .B1(n9911), .B2(n9913), .A(n9909), .ZN(n9908) );
  INV_X1 U11830 ( .A(n9911), .ZN(n9910) );
  INV_X1 U11831 ( .A(n15059), .ZN(n9909) );
  INV_X1 U11832 ( .A(n14781), .ZN(n10059) );
  AND3_X1 U11833 ( .A1(n11047), .A2(n11046), .A3(n11045), .ZN(n13606) );
  OR2_X1 U11834 ( .A1(n13601), .A2(n10064), .ZN(n13863) );
  AND2_X1 U11835 ( .A1(n11259), .A2(n10978), .ZN(n10982) );
  INV_X1 U11836 ( .A(n19871), .ZN(n19852) );
  AOI21_X1 U11837 ( .B1(n9791), .B2(n12527), .A(n12526), .ZN(n13170) );
  XNOR2_X1 U11838 ( .A(n15355), .B(n12529), .ZN(n13171) );
  NAND2_X1 U11839 ( .A1(n10972), .A2(n10937), .ZN(n13074) );
  AND2_X1 U11840 ( .A1(n19854), .A2(n13724), .ZN(n19448) );
  AND2_X1 U11841 ( .A1(n19864), .A2(n19871), .ZN(n19509) );
  AND2_X1 U11842 ( .A1(n19864), .A2(n19852), .ZN(n19850) );
  OAI21_X1 U11843 ( .B1(n10229), .B2(n10228), .A(n15408), .ZN(n10236) );
  NAND2_X1 U11844 ( .A1(n10234), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10235) );
  INV_X1 U11845 ( .A(n10484), .ZN(n19687) );
  OR2_X1 U11846 ( .A1(n19854), .A2(n19881), .ZN(n19651) );
  OR2_X1 U11847 ( .A1(n19854), .A2(n13724), .ZN(n19477) );
  NAND2_X1 U11848 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19683), .ZN(n19278) );
  AND3_X1 U11850 ( .A1(n9796), .A2(n18242), .A3(n15418), .ZN(n15419) );
  AOI22_X1 U11851 ( .A1(n17209), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13002) );
  AOI22_X1 U11852 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13001) );
  OAI21_X1 U11853 ( .B1(n17537), .B2(n10096), .A(n10095), .ZN(n17520) );
  NAND2_X1 U11854 ( .A1(n10099), .A2(n17674), .ZN(n10096) );
  INV_X1 U11855 ( .A(n17521), .ZN(n10099) );
  NAND2_X1 U11856 ( .A1(n16441), .A2(n16442), .ZN(n17537) );
  OR2_X1 U11857 ( .A1(n17537), .A2(n17781), .ZN(n10097) );
  NAND3_X1 U11858 ( .A1(n15516), .A2(n15515), .A3(n15514), .ZN(n16436) );
  INV_X1 U11859 ( .A(n17824), .ZN(n10091) );
  INV_X1 U11860 ( .A(n15617), .ZN(n10094) );
  XNOR2_X1 U11861 ( .A(n15614), .B(n15613), .ZN(n17853) );
  NAND2_X1 U11862 ( .A1(n18679), .A2(n15641), .ZN(n18684) );
  OR2_X1 U11863 ( .A1(n13329), .A2(n9766), .ZN(n19893) );
  AND2_X1 U11864 ( .A1(n15776), .A2(n13676), .ZN(n19949) );
  NOR2_X1 U11865 ( .A1(n14097), .A2(n20739), .ZN(n13676) );
  INV_X1 U11866 ( .A(n20642), .ZN(n20645) );
  AND2_X1 U11867 ( .A1(n14097), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13690) );
  INV_X1 U11868 ( .A(n11456), .ZN(n14087) );
  INV_X1 U11869 ( .A(n15902), .ZN(n14437) );
  INV_X1 U11870 ( .A(n20001), .ZN(n15884) );
  OR2_X1 U11871 ( .A1(n14440), .A2(n13326), .ZN(n15883) );
  AND2_X1 U11872 ( .A1(n14518), .A2(n12284), .ZN(n15919) );
  INV_X1 U11873 ( .A(n20045), .ZN(n20115) );
  OR2_X1 U11874 ( .A1(n13329), .A2(n15735), .ZN(n19904) );
  NAND2_X1 U11875 ( .A1(n14188), .A2(n14172), .ZN(n14173) );
  OAI21_X1 U11876 ( .B1(n14092), .B2(n9991), .A(n9989), .ZN(n9996) );
  AND2_X1 U11877 ( .A1(n13256), .A2(n13245), .ZN(n20079) );
  INV_X1 U11878 ( .A(n20079), .ZN(n20088) );
  CLKBUF_X1 U11879 ( .A(n11845), .Z(n11846) );
  INV_X1 U11880 ( .A(n20247), .ZN(n20217) );
  NAND2_X1 U11881 ( .A1(n20389), .A2(n20513), .ZN(n20433) );
  NAND2_X1 U11882 ( .A1(n10971), .A2(n10776), .ZN(n18899) );
  INV_X1 U11883 ( .A(n19881), .ZN(n13724) );
  AOI211_X1 U11884 ( .C1(n16247), .C2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n14070), .B(n10938), .ZN(n10941) );
  NAND2_X1 U11885 ( .A1(n16116), .A2(n19228), .ZN(n11280) );
  NAND2_X1 U11886 ( .A1(n14072), .A2(n14071), .ZN(n14073) );
  INV_X1 U11887 ( .A(n15346), .ZN(n19228) );
  AND2_X1 U11888 ( .A1(n10982), .A2(n9788), .ZN(n19233) );
  INV_X1 U11889 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19886) );
  INV_X1 U11890 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19877) );
  INV_X1 U11891 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19861) );
  NOR2_X2 U11892 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19856) );
  INV_X1 U11893 ( .A(n19864), .ZN(n15394) );
  AND2_X1 U11894 ( .A1(n13074), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16368) );
  NAND2_X1 U11895 ( .A1(n10204), .A2(n15408), .ZN(n10211) );
  INV_X1 U11896 ( .A(n17277), .ZN(n17273) );
  NAND2_X1 U11897 ( .A1(n17347), .A2(n9979), .ZN(n17301) );
  NOR3_X1 U11898 ( .A1(n9870), .A2(n9983), .A3(n9980), .ZN(n9979) );
  NAND2_X1 U11899 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_21__SCAN_IN), 
        .ZN(n9983) );
  INV_X1 U11900 ( .A(n9981), .ZN(n9980) );
  NAND2_X1 U11901 ( .A1(n17347), .A2(P3_EAX_REG_15__SCAN_IN), .ZN(n17342) );
  NOR2_X1 U11902 ( .A1(n9796), .A2(n15772), .ZN(n17348) );
  INV_X1 U11903 ( .A(n17260), .ZN(n15772) );
  NAND2_X1 U11904 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17260), .ZN(n17402) );
  NAND2_X1 U11905 ( .A1(n10011), .A2(n11449), .ZN(n10010) );
  INV_X1 U11906 ( .A(n13157), .ZN(n10011) );
  NAND2_X1 U11907 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12681) );
  OAI22_X1 U11908 ( .A1(n19608), .A2(n12774), .B1(n10484), .B2(n12600), .ZN(
        n10431) );
  AND2_X1 U11909 ( .A1(n12862), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n10186) );
  NAND2_X1 U11910 ( .A1(n10551), .A2(n10550), .ZN(n10553) );
  XNOR2_X1 U11911 ( .A(n15408), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10554) );
  OR2_X1 U11912 ( .A1(n11619), .A2(n11618), .ZN(n11693) );
  AND2_X1 U11913 ( .A1(n12351), .A2(n12350), .ZN(n13225) );
  OR2_X1 U11914 ( .A1(n11507), .A2(n11506), .ZN(n11720) );
  AND2_X1 U11915 ( .A1(n11455), .A2(n11456), .ZN(n12352) );
  AND2_X2 U11916 ( .A1(n11549), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11319) );
  AOI21_X1 U11917 ( .B1(n9795), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A(n9929), .ZN(n12796) );
  AND2_X1 U11918 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n9929) );
  NOR2_X1 U11919 ( .A1(n9874), .A2(n9935), .ZN(n12789) );
  AND2_X1 U11920 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n9935) );
  NOR2_X1 U11921 ( .A1(n9872), .A2(n9933), .ZN(n12752) );
  AND2_X1 U11922 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n9933) );
  NOR2_X1 U11923 ( .A1(n19235), .A2(n18894), .ZN(n9901) );
  NOR3_X1 U11924 ( .A1(n10640), .A2(n9948), .A3(P2_EBX_REG_10__SCAN_IN), .ZN(
        n10643) );
  AND2_X1 U11925 ( .A1(n10961), .A2(n9755), .ZN(n10253) );
  AND2_X1 U11926 ( .A1(n10265), .A2(n9755), .ZN(n10280) );
  AND2_X1 U11927 ( .A1(n12862), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n10150) );
  XNOR2_X1 U11928 ( .A(n9780), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10547) );
  NOR2_X1 U11929 ( .A1(n12922), .A2(n12924), .ZN(n15537) );
  AND2_X1 U11930 ( .A1(n13015), .A2(n18232), .ZN(n13004) );
  AND2_X1 U11931 ( .A1(n15774), .A2(n17398), .ZN(n15659) );
  AOI21_X1 U11932 ( .B1(n18699), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n13017), .ZN(n13024) );
  NAND2_X1 U11933 ( .A1(n12278), .A2(n10086), .ZN(n10085) );
  INV_X1 U11934 ( .A(n14212), .ZN(n10086) );
  OR2_X1 U11935 ( .A1(n14652), .A2(n11495), .ZN(n12310) );
  AND2_X1 U11936 ( .A1(n12069), .A2(n14366), .ZN(n14358) );
  NAND2_X1 U11937 ( .A1(n10079), .A2(n11902), .ZN(n10078) );
  INV_X1 U11938 ( .A(n13876), .ZN(n10079) );
  INV_X1 U11939 ( .A(n11720), .ZN(n11726) );
  INV_X1 U11940 ( .A(n13595), .ZN(n11874) );
  INV_X1 U11941 ( .A(n11466), .ZN(n11822) );
  AND2_X1 U11942 ( .A1(n11820), .A2(n11821), .ZN(n13185) );
  NOR2_X1 U11943 ( .A1(n14340), .A2(n14332), .ZN(n9891) );
  NOR2_X1 U11944 ( .A1(n11777), .A2(n11726), .ZN(n11650) );
  INV_X1 U11945 ( .A(n11701), .ZN(n10008) );
  INV_X1 U11946 ( .A(n11770), .ZN(n12351) );
  AND2_X1 U11947 ( .A1(n13685), .A2(n20842), .ZN(n13142) );
  OR2_X1 U11948 ( .A1(n11517), .A2(n11516), .ZN(n11666) );
  OAI211_X1 U11949 ( .C1(n11565), .C2(n11566), .A(n11573), .B(n11572), .ZN(
        n11574) );
  NOR2_X1 U11950 ( .A1(n11809), .A2(n11770), .ZN(n11817) );
  AOI21_X1 U11951 ( .B1(n11813), .B2(n11812), .A(n11811), .ZN(n13139) );
  CLKBUF_X1 U11952 ( .A(n13148), .Z(n13149) );
  INV_X1 U11953 ( .A(n20220), .ZN(n20260) );
  XNOR2_X1 U11954 ( .A(n10000), .B(n11560), .ZN(n20258) );
  INV_X1 U11955 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20555) );
  INV_X1 U11956 ( .A(n11846), .ZN(n20109) );
  NAND2_X1 U11957 ( .A1(n20416), .A2(n11495), .ZN(n11609) );
  NAND2_X1 U11958 ( .A1(n10539), .A2(n10252), .ZN(n10270) );
  AOI22_X1 U11959 ( .A1(n9753), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10243), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10219) );
  NOR2_X1 U11960 ( .A1(n10731), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n10722) );
  NOR2_X1 U11961 ( .A1(n9953), .A2(n10678), .ZN(n9952) );
  INV_X1 U11962 ( .A(n10654), .ZN(n9953) );
  NAND2_X1 U11963 ( .A1(n10643), .A2(n13704), .ZN(n10652) );
  NAND2_X1 U11964 ( .A1(n9949), .A2(n10845), .ZN(n9948) );
  INV_X1 U11965 ( .A(n10632), .ZN(n9949) );
  NOR2_X1 U11966 ( .A1(n10640), .A2(n10632), .ZN(n10639) );
  INV_X1 U11967 ( .A(n10558), .ZN(n10576) );
  NOR2_X1 U11968 ( .A1(n10577), .A2(n10576), .ZN(n10575) );
  INV_X1 U11969 ( .A(n14739), .ZN(n9966) );
  OAI22_X1 U11971 ( .A1(n10332), .A2(n15408), .B1(n16363), .B2(n19861), .ZN(
        n10820) );
  INV_X1 U11972 ( .A(n12852), .ZN(n10026) );
  AND2_X1 U11973 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n9930) );
  AOI21_X1 U11974 ( .B1(n9795), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A(n9931), .ZN(n12823) );
  AND2_X1 U11975 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n9931) );
  AOI21_X1 U11976 ( .B1(n9795), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A(n9928), 
        .ZN(n12769) );
  AND2_X1 U11977 ( .A1(n9863), .A2(n14902), .ZN(n10043) );
  INV_X1 U11978 ( .A(n13701), .ZN(n9963) );
  INV_X1 U11979 ( .A(n9904), .ZN(n9903) );
  INV_X1 U11980 ( .A(n9906), .ZN(n9905) );
  NOR2_X1 U11981 ( .A1(n10733), .A2(n10732), .ZN(n10734) );
  NOR2_X1 U11982 ( .A1(n12470), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10733) );
  NOR2_X1 U11983 ( .A1(n14996), .A2(n10112), .ZN(n10111) );
  INV_X1 U11984 ( .A(n15162), .ZN(n10112) );
  AND2_X1 U11985 ( .A1(n13947), .A2(n14934), .ZN(n10072) );
  OR2_X1 U11986 ( .A1(n16156), .A2(n11055), .ZN(n10739) );
  NOR2_X1 U11987 ( .A1(n10109), .A2(n10110), .ZN(n10108) );
  INV_X1 U11988 ( .A(n10708), .ZN(n10110) );
  INV_X1 U11989 ( .A(n9851), .ZN(n10109) );
  NAND2_X1 U11990 ( .A1(n15037), .A2(n15226), .ZN(n11303) );
  CLKBUF_X1 U11991 ( .A(n14742), .Z(n15194) );
  AND2_X1 U11992 ( .A1(n11230), .A2(n11229), .ZN(n15234) );
  INV_X1 U11993 ( .A(n13771), .ZN(n9961) );
  NOR2_X1 U11994 ( .A1(n10057), .A2(n10056), .ZN(n10055) );
  INV_X1 U11995 ( .A(n15267), .ZN(n10056) );
  NOR2_X1 U11996 ( .A1(n16233), .A2(n15279), .ZN(n10041) );
  OAI21_X1 U11997 ( .B1(n10247), .B2(n10248), .A(n15408), .ZN(n10249) );
  AND2_X1 U11998 ( .A1(n9978), .A2(n9977), .ZN(n13916) );
  INV_X1 U11999 ( .A(n15552), .ZN(n15474) );
  NOR2_X1 U12000 ( .A1(n12922), .A2(n12919), .ZN(n15554) );
  AND3_X1 U12001 ( .A1(n12916), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n18685), .ZN(n15595) );
  NOR2_X1 U12002 ( .A1(n12923), .A2(n16921), .ZN(n15551) );
  NOR2_X1 U12003 ( .A1(n17715), .A2(n17717), .ZN(n16776) );
  NAND2_X1 U12004 ( .A1(n15684), .A2(n17781), .ZN(n15688) );
  NOR2_X1 U12005 ( .A1(n17801), .A2(n15671), .ZN(n15672) );
  NAND2_X1 U12006 ( .A1(n13921), .A2(n9977), .ZN(n9976) );
  INV_X1 U12007 ( .A(n15646), .ZN(n18679) );
  NOR2_X1 U12008 ( .A1(n13014), .A2(n15644), .ZN(n15641) );
  AOI211_X1 U12009 ( .C1(n17213), .C2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n12988), .B(n12987), .ZN(n12989) );
  OAI221_X1 U12010 ( .B1(n18888), .B2(P3_STATE2_REG_1__SCAN_IN), .C1(
        P3_STATE2_REG_2__SCAN_IN), .C2(n18834), .A(n18836), .ZN(n18219) );
  OR2_X1 U12011 ( .A1(n20840), .A2(n13673), .ZN(n15776) );
  AND2_X1 U12012 ( .A1(n12445), .A2(n12444), .ZN(n14223) );
  AND2_X1 U12013 ( .A1(n12422), .A2(n12421), .ZN(n14352) );
  OR2_X1 U12014 ( .A1(n14187), .A2(n10085), .ZN(n10084) );
  OR2_X1 U12015 ( .A1(n11759), .A2(n11758), .ZN(n11760) );
  NAND2_X1 U12016 ( .A1(n12238), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12239) );
  INV_X1 U12017 ( .A(n12237), .ZN(n12238) );
  OR2_X1 U12018 ( .A1(n12239), .A2(n14214), .ZN(n12291) );
  OR2_X1 U12019 ( .A1(n12202), .A2(n21030), .ZN(n12237) );
  INV_X1 U12020 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n21030) );
  OR2_X1 U12021 ( .A1(n12158), .A2(n14265), .ZN(n12184) );
  AND2_X1 U12022 ( .A1(n12088), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12089) );
  AND2_X1 U12023 ( .A1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n12089), .ZN(
        n12132) );
  NOR2_X1 U12024 ( .A1(n11970), .A2(n11951), .ZN(n12088) );
  NAND2_X1 U12025 ( .A1(n12020), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12004) );
  INV_X1 U12026 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11950) );
  AND2_X1 U12027 ( .A1(n11934), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11935) );
  AND2_X1 U12028 ( .A1(n12044), .A2(n11948), .ZN(n15874) );
  AND3_X1 U12029 ( .A1(n11931), .A2(n11930), .A3(n11929), .ZN(n11932) );
  NAND2_X1 U12030 ( .A1(n11903), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11918) );
  INV_X1 U12031 ( .A(n13749), .ZN(n10077) );
  NOR2_X1 U12032 ( .A1(n21005), .A2(n11881), .ZN(n11903) );
  AOI21_X1 U12033 ( .B1(n11879), .B2(n12044), .A(n11878), .ZN(n13732) );
  NAND2_X1 U12034 ( .A1(n11868), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11875) );
  NAND2_X1 U12035 ( .A1(n11844), .A2(n11843), .ZN(n13296) );
  AOI21_X1 U12036 ( .B1(n9990), .B2(n9994), .A(n9860), .ZN(n9989) );
  INV_X1 U12037 ( .A(n9995), .ZN(n9990) );
  INV_X1 U12038 ( .A(n9994), .ZN(n9991) );
  NAND2_X1 U12039 ( .A1(n9993), .A2(n9998), .ZN(n9992) );
  INV_X1 U12040 ( .A(n14449), .ZN(n9993) );
  INV_X1 U12041 ( .A(n12440), .ZN(n14238) );
  NOR2_X1 U12042 ( .A1(n14327), .A2(n14260), .ZN(n14261) );
  OAI21_X2 U12043 ( .B1(n14511), .B2(n9813), .A(n15893), .ZN(n14505) );
  AND2_X1 U12044 ( .A1(n14525), .A2(n10127), .ZN(n10012) );
  NAND2_X1 U12045 ( .A1(n9891), .A2(n9890), .ZN(n14327) );
  INV_X1 U12046 ( .A(n14325), .ZN(n9890) );
  OR2_X1 U12047 ( .A1(n14353), .A2(n14352), .ZN(n14355) );
  NOR2_X2 U12048 ( .A1(n14355), .A2(n14348), .ZN(n14347) );
  OR3_X1 U12049 ( .A1(n16001), .A2(n15971), .A3(n13983), .ZN(n14641) );
  AND2_X1 U12050 ( .A1(n12399), .A2(n12398), .ZN(n13910) );
  OR2_X1 U12051 ( .A1(n16053), .A2(n13910), .ZN(n15867) );
  NAND2_X1 U12052 ( .A1(n11484), .A2(n11495), .ZN(n20835) );
  CLKBUF_X1 U12053 ( .A(n14009), .Z(n14554) );
  AND2_X1 U12054 ( .A1(n11732), .A2(n10123), .ZN(n10009) );
  NAND2_X1 U12055 ( .A1(n12395), .A2(n12394), .ZN(n16053) );
  INV_X1 U12056 ( .A(n16051), .ZN(n12394) );
  INV_X1 U12057 ( .A(n13790), .ZN(n12395) );
  INV_X1 U12058 ( .A(n16089), .ZN(n12381) );
  NAND2_X1 U12059 ( .A1(n15943), .A2(n15942), .ZN(n15941) );
  NAND2_X1 U12060 ( .A1(n12370), .A2(n12369), .ZN(n13468) );
  NOR2_X1 U12061 ( .A1(n13467), .A2(n13468), .ZN(n13570) );
  NAND2_X1 U12062 ( .A1(n13994), .A2(n20094), .ZN(n20054) );
  INV_X1 U12063 ( .A(n16024), .ZN(n20072) );
  NAND2_X1 U12064 ( .A1(n13240), .A2(n13239), .ZN(n13256) );
  OR2_X1 U12065 ( .A1(n13329), .A2(n13238), .ZN(n13239) );
  AND2_X1 U12066 ( .A1(n9787), .A2(n12452), .ZN(n13247) );
  NAND2_X1 U12067 ( .A1(n20188), .A2(n11564), .ZN(n14300) );
  NAND2_X1 U12068 ( .A1(n10004), .A2(n9853), .ZN(n11588) );
  INV_X1 U12069 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13387) );
  NOR2_X1 U12070 ( .A1(n13405), .A2(n9877), .ZN(n13397) );
  OAI21_X1 U12071 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n21100), .A(
        n20299), .ZN(n20261) );
  INV_X1 U12072 ( .A(n20522), .ZN(n20514) );
  OR2_X1 U12073 ( .A1(n20107), .A2(n13420), .ZN(n20522) );
  OR2_X2 U12074 ( .A1(n11390), .A2(n11389), .ZN(n20145) );
  AND3_X1 U12075 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n11495), .A3(n20119), 
        .ZN(n20177) );
  NOR2_X1 U12076 ( .A1(n20214), .A2(n20109), .ZN(n20548) );
  AND2_X1 U12077 ( .A1(n20214), .A2(n20109), .ZN(n20513) );
  INV_X1 U12078 ( .A(n20261), .ZN(n20684) );
  NOR2_X2 U12079 ( .A1(n20116), .A2(n20115), .ZN(n20173) );
  NOR2_X2 U12080 ( .A1(n20115), .A2(n20114), .ZN(n20172) );
  CLKBUF_X1 U12081 ( .A(n13175), .Z(n13176) );
  OR2_X1 U12082 ( .A1(n13141), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n13327) );
  NAND2_X1 U12083 ( .A1(n10949), .A2(n10721), .ZN(n10736) );
  NAND2_X1 U12084 ( .A1(n14681), .A2(n9811), .ZN(n14678) );
  NOR2_X1 U12085 ( .A1(n10722), .A2(n10715), .ZN(n10720) );
  INV_X1 U12086 ( .A(n10729), .ZN(n10715) );
  NOR2_X1 U12087 ( .A1(n9945), .A2(n9942), .ZN(n9941) );
  NAND2_X1 U12088 ( .A1(n9944), .A2(n9943), .ZN(n9942) );
  INV_X1 U12089 ( .A(n10673), .ZN(n9945) );
  AND2_X1 U12090 ( .A1(n14707), .A2(n10048), .ZN(n14733) );
  INV_X1 U12091 ( .A(n14732), .ZN(n10048) );
  NOR2_X1 U12092 ( .A1(n14698), .A2(n18975), .ZN(n14701) );
  NAND2_X1 U12093 ( .A1(n10651), .A2(n9950), .ZN(n10664) );
  NOR2_X1 U12094 ( .A1(n9951), .A2(n9956), .ZN(n9950) );
  INV_X1 U12095 ( .A(n10658), .ZN(n9956) );
  INV_X1 U12096 ( .A(n9952), .ZN(n9951) );
  AND2_X1 U12097 ( .A1(n9970), .A2(n14861), .ZN(n9969) );
  NAND2_X1 U12098 ( .A1(n11293), .A2(n9964), .ZN(n14897) );
  AND2_X1 U12099 ( .A1(n9848), .A2(n9965), .ZN(n9964) );
  INV_X1 U12100 ( .A(n14895), .ZN(n9965) );
  AND2_X1 U12101 ( .A1(n13707), .A2(n13705), .ZN(n13706) );
  AOI21_X1 U12102 ( .B1(n9748), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A(n9932), 
        .ZN(n12859) );
  AND2_X1 U12103 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n9932) );
  AOI21_X1 U12104 ( .B1(n9759), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A(n9936), .ZN(n12857) );
  AND2_X1 U12105 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n9936) );
  NOR2_X2 U12106 ( .A1(n14928), .A2(n12477), .ZN(n14914) );
  OAI21_X1 U12107 ( .B1(n14884), .B2(n10036), .A(n10035), .ZN(n14874) );
  NAND2_X1 U12108 ( .A1(n10038), .A2(n10037), .ZN(n10036) );
  INV_X1 U12109 ( .A(n14883), .ZN(n10037) );
  NOR2_X1 U12110 ( .A1(n14884), .A2(n14883), .ZN(n14882) );
  AND2_X1 U12111 ( .A1(n11233), .A2(n11232), .ZN(n12498) );
  AND4_X1 U12112 ( .A1(n12634), .A2(n12633), .A3(n12632), .A4(n12631), .ZN(
        n13905) );
  NAND2_X1 U12113 ( .A1(n13839), .A2(n14906), .ZN(n14905) );
  AND2_X1 U12114 ( .A1(n11227), .A2(n11226), .ZN(n15257) );
  INV_X1 U12115 ( .A(n10281), .ZN(n12878) );
  NAND2_X1 U12116 ( .A1(n19110), .A2(n12897), .ZN(n13207) );
  OAI21_X1 U12117 ( .B1(n11249), .B2(n18912), .A(n11016), .ZN(n13208) );
  INV_X1 U12118 ( .A(n10935), .ZN(n19140) );
  AND2_X1 U12119 ( .A1(n19139), .A2(n19778), .ZN(n19169) );
  INV_X1 U12120 ( .A(n12893), .ZN(n13645) );
  OAI21_X1 U12121 ( .B1(n12892), .B2(n12891), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12893) );
  AND2_X1 U12122 ( .A1(n14681), .A2(n9871), .ZN(n14042) );
  NOR2_X1 U12123 ( .A1(n14706), .A2(n15010), .ZN(n14709) );
  NAND2_X1 U12124 ( .A1(n14685), .A2(n9812), .ZN(n14684) );
  NOR2_X1 U12125 ( .A1(n14684), .A2(n15029), .ZN(n14705) );
  INV_X1 U12126 ( .A(n14700), .ZN(n14685) );
  NAND2_X1 U12127 ( .A1(n14685), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14703) );
  INV_X1 U12128 ( .A(n14686), .ZN(n14699) );
  NAND2_X1 U12129 ( .A1(n14692), .A2(n9808), .ZN(n14697) );
  NAND2_X1 U12130 ( .A1(n14692), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14695) );
  NOR2_X1 U12131 ( .A1(n16271), .A2(n14693), .ZN(n14692) );
  NOR2_X1 U12132 ( .A1(n14690), .A2(n16282), .ZN(n14687) );
  AND2_X1 U12133 ( .A1(n10636), .A2(n16327), .ZN(n16277) );
  AND2_X1 U12134 ( .A1(n10069), .A2(n9806), .ZN(n14691) );
  NAND2_X1 U12135 ( .A1(n14691), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14690) );
  INV_X1 U12136 ( .A(n13376), .ZN(n9967) );
  NAND2_X1 U12137 ( .A1(n10069), .A2(n10070), .ZN(n14688) );
  AND2_X1 U12138 ( .A1(n13760), .A2(n13759), .ZN(n13762) );
  NOR2_X1 U12139 ( .A1(n14131), .A2(n19211), .ZN(n14130) );
  NAND2_X1 U12140 ( .A1(n10341), .A2(n10340), .ZN(n10339) );
  AND2_X1 U12141 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13618) );
  OAI22_X1 U12142 ( .A1(n9762), .A2(n10278), .B1(n10311), .B2(n10277), .ZN(
        n10292) );
  NOR2_X1 U12143 ( .A1(n10394), .A2(n10393), .ZN(n13221) );
  AND2_X1 U12144 ( .A1(n14841), .A2(n10914), .ZN(n9957) );
  NOR2_X1 U12145 ( .A1(n16135), .A2(n11055), .ZN(n12470) );
  AND2_X1 U12146 ( .A1(n10814), .A2(n10041), .ZN(n10040) );
  NAND2_X1 U12147 ( .A1(n9939), .A2(n9864), .ZN(n15023) );
  INV_X1 U12148 ( .A(n14748), .ZN(n9939) );
  OR2_X1 U12149 ( .A1(n10697), .A2(n12500), .ZN(n15024) );
  AND2_X1 U12150 ( .A1(n10114), .A2(n9922), .ZN(n9921) );
  INV_X1 U12151 ( .A(n15095), .ZN(n9922) );
  AND2_X1 U12152 ( .A1(n10677), .A2(n16305), .ZN(n16239) );
  AND3_X1 U12153 ( .A1(n11154), .A2(n11153), .A3(n11152), .ZN(n14781) );
  AND2_X1 U12154 ( .A1(n11112), .A2(n11111), .ZN(n14792) );
  CLKBUF_X1 U12155 ( .A(n14790), .Z(n15309) );
  NAND2_X1 U12156 ( .A1(n13763), .A2(n11263), .ZN(n15289) );
  OR2_X1 U12157 ( .A1(n10810), .A2(n10809), .ZN(n10811) );
  INV_X1 U12158 ( .A(n16277), .ZN(n10116) );
  AND3_X1 U12159 ( .A1(n11073), .A2(n11072), .A3(n11071), .ZN(n14810) );
  NOR2_X1 U12160 ( .A1(n10063), .A2(n9856), .ZN(n10062) );
  NOR2_X1 U12161 ( .A1(n15331), .A2(n11052), .ZN(n10063) );
  INV_X1 U12162 ( .A(n10791), .ZN(n10792) );
  NAND2_X1 U12163 ( .A1(n10514), .A2(n10788), .ZN(n13755) );
  NAND2_X1 U12164 ( .A1(n10561), .A2(n10562), .ZN(n10021) );
  INV_X1 U12165 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13758) );
  AND2_X1 U12166 ( .A1(n11259), .A2(n15379), .ZN(n15245) );
  INV_X1 U12167 ( .A(n16361), .ZN(n15768) );
  NAND2_X1 U12168 ( .A1(n12535), .A2(n19680), .ZN(n12524) );
  INV_X1 U12169 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15370) );
  OAI21_X1 U12170 ( .B1(n13617), .B2(n12523), .A(n10015), .ZN(n10014) );
  NOR2_X1 U12171 ( .A1(n9852), .A2(n10016), .ZN(n10015) );
  AOI21_X1 U12172 ( .B1(n9749), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A(
        n10205), .ZN(n10210) );
  NAND2_X1 U12173 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10207) );
  NAND2_X1 U12174 ( .A1(n12861), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10206) );
  NAND2_X1 U12175 ( .A1(n10209), .A2(n10208), .ZN(n9918) );
  AND2_X1 U12176 ( .A1(n19346), .A2(n19856), .ZN(n19350) );
  INV_X1 U12177 ( .A(n19477), .ZN(n19607) );
  INV_X1 U12178 ( .A(n19644), .ZN(n19650) );
  INV_X1 U12179 ( .A(n19274), .ZN(n19276) );
  INV_X1 U12180 ( .A(n19275), .ZN(n19277) );
  INV_X1 U12181 ( .A(n9755), .ZN(n19279) );
  NOR2_X1 U12182 ( .A1(n15362), .A2(n15361), .ZN(n16354) );
  OR2_X1 U12183 ( .A1(n10936), .A2(n10757), .ZN(n13072) );
  OR2_X1 U12184 ( .A1(n13921), .A2(n9783), .ZN(n9978) );
  NOR2_X1 U12185 ( .A1(n16610), .A2(n9897), .ZN(n16601) );
  NOR2_X1 U12186 ( .A1(n16624), .A2(n9897), .ZN(n16611) );
  NOR2_X1 U12187 ( .A1(n16611), .A2(n16612), .ZN(n16610) );
  NOR2_X1 U12188 ( .A1(n16625), .A2(n17519), .ZN(n16624) );
  NOR2_X1 U12189 ( .A1(n16634), .A2(n16633), .ZN(n16632) );
  NOR2_X1 U12190 ( .A1(n16668), .A2(n9897), .ZN(n16654) );
  NOR2_X1 U12191 ( .A1(n16654), .A2(n16655), .ZN(n16653) );
  NOR2_X1 U12192 ( .A1(n16669), .A2(n17575), .ZN(n16668) );
  NOR2_X1 U12193 ( .A1(n16687), .A2(n9897), .ZN(n16676) );
  NOR2_X1 U12194 ( .A1(n17587), .A2(n16676), .ZN(n16675) );
  NOR2_X1 U12195 ( .A1(n16698), .A2(n9897), .ZN(n16688) );
  NOR2_X1 U12196 ( .A1(n16688), .A2(n16689), .ZN(n16687) );
  NAND2_X1 U12197 ( .A1(n17122), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n9973) );
  NAND2_X1 U12198 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n9972) );
  NAND2_X1 U12199 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17234), .ZN(n17201) );
  NOR2_X1 U12200 ( .A1(n17479), .A2(n9985), .ZN(n9984) );
  NOR2_X1 U12201 ( .A1(n17432), .A2(n9982), .ZN(n9981) );
  NOR2_X1 U12202 ( .A1(n15566), .A2(n15565), .ZN(n15567) );
  NOR2_X1 U12203 ( .A1(n17464), .A2(n17407), .ZN(n17433) );
  NOR2_X1 U12204 ( .A1(n18724), .A2(n18660), .ZN(n17462) );
  NOR2_X1 U12205 ( .A1(n16390), .A2(n17875), .ZN(n16412) );
  NAND2_X1 U12206 ( .A1(n16415), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16390) );
  NOR2_X1 U12207 ( .A1(n17530), .A2(n17531), .ZN(n16415) );
  NAND2_X1 U12208 ( .A1(n17627), .A2(n9893), .ZN(n17561) );
  AND2_X1 U12209 ( .A1(n9894), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9893) );
  AND2_X1 U12210 ( .A1(n16583), .A2(n9895), .ZN(n9894) );
  INV_X1 U12211 ( .A(n17604), .ZN(n9895) );
  OR2_X1 U12212 ( .A1(n17604), .A2(n16588), .ZN(n17560) );
  NAND2_X1 U12213 ( .A1(n17627), .A2(n16583), .ZN(n17603) );
  INV_X1 U12214 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17629) );
  NOR2_X1 U12215 ( .A1(n17677), .A2(n17678), .ZN(n17627) );
  NAND2_X1 U12216 ( .A1(n16776), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17677) );
  NAND2_X1 U12217 ( .A1(n16844), .A2(n17700), .ZN(n17715) );
  NOR2_X1 U12218 ( .A1(n16812), .A2(n9898), .ZN(n17700) );
  NAND2_X1 U12219 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n9898) );
  NOR2_X1 U12220 ( .A1(n17814), .A2(n17815), .ZN(n16844) );
  NOR2_X1 U12221 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18888), .ZN(n17713) );
  AOI21_X1 U12222 ( .B1(n16448), .B2(n16447), .A(n16446), .ZN(n16449) );
  AOI21_X1 U12223 ( .B1(n16451), .B2(n18062), .A(n16450), .ZN(n16452) );
  NOR2_X1 U12224 ( .A1(n17907), .A2(n17945), .ZN(n17921) );
  NOR2_X1 U12225 ( .A1(n17707), .A2(n18063), .ZN(n17706) );
  NOR2_X1 U12226 ( .A1(n17730), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17698) );
  NOR2_X1 U12227 ( .A1(n17765), .A2(n17761), .ZN(n17745) );
  NAND2_X1 U12228 ( .A1(n18694), .A2(n18665), .ZN(n18098) );
  NAND2_X1 U12229 ( .A1(n17795), .A2(n15624), .ZN(n15680) );
  INV_X1 U12230 ( .A(n18084), .ZN(n17994) );
  NOR2_X1 U12231 ( .A1(n17803), .A2(n17802), .ZN(n17801) );
  NAND2_X1 U12232 ( .A1(n15642), .A2(n18884), .ZN(n18665) );
  XNOR2_X1 U12233 ( .A(n15648), .B(n15608), .ZN(n17872) );
  OAI21_X1 U12234 ( .B1(n15633), .B2(n15632), .A(n15631), .ZN(n18661) );
  AND2_X1 U12235 ( .A1(n15774), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17880) );
  OR2_X1 U12236 ( .A1(n15774), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17873) );
  NOR2_X1 U12237 ( .A1(n15641), .A2(n15646), .ZN(n18694) );
  INV_X1 U12238 ( .A(n18665), .ZN(n18690) );
  NOR2_X1 U12239 ( .A1(n12981), .A2(n12980), .ZN(n18238) );
  INV_X1 U12240 ( .A(n15635), .ZN(n18242) );
  NOR2_X1 U12241 ( .A1(n12943), .A2(n12942), .ZN(n18253) );
  INV_X1 U12242 ( .A(n18515), .ZN(n18331) );
  NAND2_X1 U12243 ( .A1(n18727), .A2(n18219), .ZN(n18515) );
  NAND2_X1 U12244 ( .A1(n19893), .A2(n19895), .ZN(n20840) );
  AND2_X1 U12245 ( .A1(n19937), .A2(n15776), .ZN(n14281) );
  AND2_X1 U12246 ( .A1(n14331), .A2(n14330), .ZN(n15784) );
  INV_X1 U12247 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15839) );
  NAND2_X1 U12248 ( .A1(n19964), .A2(n13793), .ZN(n19954) );
  NAND2_X1 U12249 ( .A1(n13688), .A2(n13687), .ZN(n19937) );
  INV_X1 U12250 ( .A(n19937), .ZN(n19964) );
  INV_X1 U12251 ( .A(n19977), .ZN(n19942) );
  AND2_X1 U12252 ( .A1(n15776), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19960) );
  NOR2_X1 U12253 ( .A1(n13190), .A2(n19899), .ZN(n12357) );
  INV_X1 U12254 ( .A(n14410), .ZN(n14438) );
  OR2_X1 U12255 ( .A1(n14388), .A2(n14387), .ZN(n15881) );
  OR2_X1 U12256 ( .A1(n13574), .A2(n13466), .ZN(n13566) );
  NAND2_X1 U12257 ( .A1(n13320), .A2(n13319), .ZN(n20001) );
  AOI21_X1 U12258 ( .B1(n13318), .B2(n13317), .A(n13316), .ZN(n13319) );
  OR2_X1 U12259 ( .A1(n13329), .A2(n13314), .ZN(n13320) );
  NAND2_X1 U12260 ( .A1(n13517), .A2(n13332), .ZN(n20007) );
  NOR2_X1 U12261 ( .A1(n20007), .A2(n20006), .ZN(n20008) );
  INV_X1 U12262 ( .A(n20007), .ZN(n13556) );
  INV_X2 U12263 ( .A(n13334), .ZN(n20036) );
  AND2_X1 U12264 ( .A1(n20842), .A2(n20838), .ZN(n13290) );
  NOR2_X2 U12265 ( .A1(n9761), .A2(n13291), .ZN(n20022) );
  XNOR2_X1 U12266 ( .A(n13675), .B(n14179), .ZN(n14097) );
  INV_X1 U12267 ( .A(n15784), .ZN(n14509) );
  AND2_X1 U12268 ( .A1(n14328), .A2(n14336), .ZN(n15794) );
  NAND2_X1 U12269 ( .A1(n14006), .A2(n12072), .ZN(n14345) );
  AND2_X1 U12270 ( .A1(n14277), .A2(n14350), .ZN(n15902) );
  INV_X1 U12271 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13564) );
  INV_X1 U12272 ( .A(n14518), .ZN(n20039) );
  AND2_X2 U12273 ( .A1(n12279), .A2(n20613), .ZN(n20045) );
  NAND2_X1 U12274 ( .A1(n9988), .A2(n9994), .ZN(n14451) );
  NAND2_X1 U12275 ( .A1(n14092), .A2(n9995), .ZN(n9988) );
  AND2_X1 U12276 ( .A1(n14199), .A2(n14198), .ZN(n14589) );
  AND2_X1 U12277 ( .A1(n14630), .A2(n13984), .ZN(n14600) );
  OR2_X1 U12278 ( .A1(n20835), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16045) );
  CLKBUF_X1 U12279 ( .A(n11848), .Z(n11849) );
  INV_X1 U12280 ( .A(n20613), .ZN(n20836) );
  NAND2_X1 U12281 ( .A1(n10005), .A2(n11590), .ZN(n20552) );
  NAND2_X1 U12282 ( .A1(n13419), .A2(n20182), .ZN(n20104) );
  INV_X1 U12283 ( .A(n20213), .ZN(n20205) );
  OAI21_X1 U12284 ( .B1(n20225), .B2(n20222), .A(n20221), .ZN(n20250) );
  OR2_X1 U12285 ( .A1(n20257), .A2(n20187), .ZN(n20247) );
  INV_X1 U12286 ( .A(n20311), .ZN(n20318) );
  NAND2_X1 U12287 ( .A1(n20389), .A2(n20548), .ZN(n20348) );
  OAI21_X1 U12288 ( .B1(n20394), .B2(n20393), .A(n20684), .ZN(n20412) );
  OAI211_X1 U12289 ( .C1(n20439), .C2(n21100), .A(n20477), .B(n20422), .ZN(
        n20441) );
  INV_X1 U12290 ( .A(n20433), .ZN(n20440) );
  INV_X1 U12291 ( .A(n20482), .ZN(n20509) );
  NAND2_X1 U12292 ( .A1(n20514), .A2(n20639), .ZN(n20546) );
  OAI211_X1 U12293 ( .C1(n20563), .C2(n21100), .A(n20649), .B(n20562), .ZN(
        n20605) );
  OAI211_X1 U12294 ( .C1(n20669), .C2(n20650), .A(n20649), .B(n20648), .ZN(
        n20671) );
  INV_X1 U12295 ( .A(n20556), .ZN(n20678) );
  INV_X1 U12296 ( .A(n20567), .ZN(n20691) );
  INV_X1 U12297 ( .A(n20572), .ZN(n20697) );
  INV_X1 U12298 ( .A(n20579), .ZN(n20703) );
  INV_X1 U12299 ( .A(n20584), .ZN(n20709) );
  NAND2_X1 U12300 ( .A1(n20679), .A2(n20639), .ZN(n20720) );
  INV_X1 U12301 ( .A(n20591), .ZN(n20715) );
  INV_X1 U12302 ( .A(n20596), .ZN(n20723) );
  NAND2_X1 U12303 ( .A1(n20679), .A2(n20513), .ZN(n20737) );
  INV_X1 U12304 ( .A(n20720), .ZN(n20733) );
  INV_X1 U12305 ( .A(n20602), .ZN(n20731) );
  NOR2_X1 U12306 ( .A1(n20742), .A2(n20739), .ZN(n16110) );
  NOR2_X1 U12307 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20843) );
  INV_X1 U12308 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20739) );
  INV_X1 U12309 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n21100) );
  NAND2_X1 U12310 ( .A1(n20746), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20833) );
  INV_X1 U12311 ( .A(n14137), .ZN(n18895) );
  NOR2_X1 U12312 ( .A1(n14733), .A2(n10047), .ZN(n15712) );
  AND2_X1 U12313 ( .A1(n14707), .A2(n15032), .ZN(n10047) );
  CLKBUF_X1 U12314 ( .A(n19003), .Z(n19024) );
  INV_X1 U12315 ( .A(n19054), .ZN(n19028) );
  INV_X1 U12316 ( .A(n19003), .ZN(n19057) );
  OR2_X1 U12317 ( .A1(n19136), .A2(n14145), .ZN(n19063) );
  AND2_X1 U12318 ( .A1(n14146), .A2(n14145), .ZN(n19054) );
  INV_X1 U12319 ( .A(n19771), .ZN(n19050) );
  AND2_X1 U12320 ( .A1(n13828), .A2(n13827), .ZN(n13880) );
  NOR2_X1 U12321 ( .A1(n13659), .A2(n13658), .ZN(n13775) );
  INV_X1 U12322 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n20987) );
  NAND2_X1 U12323 ( .A1(n9755), .A2(n14901), .ZN(n14911) );
  NAND2_X1 U12324 ( .A1(n10024), .A2(n10022), .ZN(n12873) );
  NAND2_X1 U12325 ( .A1(n10032), .A2(n10033), .ZN(n14845) );
  NAND2_X1 U12326 ( .A1(n10031), .A2(n10029), .ZN(n10028) );
  INV_X1 U12327 ( .A(n10033), .ZN(n10027) );
  NOR2_X1 U12328 ( .A1(n14857), .A2(n14856), .ZN(n14855) );
  INV_X1 U12329 ( .A(n14863), .ZN(n14864) );
  NAND2_X1 U12330 ( .A1(n19110), .A2(n12883), .ZN(n14973) );
  AND2_X1 U12331 ( .A1(n12877), .A2(n19768), .ZN(n19110) );
  AND2_X1 U12332 ( .A1(n19084), .A2(n19112), .ZN(n19118) );
  NAND2_X1 U12333 ( .A1(n12878), .A2(n19110), .ZN(n19112) );
  NAND2_X1 U12334 ( .A1(n14973), .A2(n13207), .ZN(n19102) );
  AND2_X1 U12335 ( .A1(n19110), .A2(n19279), .ZN(n19127) );
  INV_X1 U12336 ( .A(n19112), .ZN(n19131) );
  NAND2_X1 U12337 ( .A1(n14143), .A2(n9788), .ZN(n19136) );
  XNOR2_X1 U12338 ( .A(n14058), .B(n14057), .ZN(n14132) );
  INV_X1 U12339 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15010) );
  INV_X1 U12340 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n21034) );
  INV_X1 U12341 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15084) );
  INV_X1 U12342 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n15100) );
  INV_X1 U12343 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19211) );
  NAND2_X1 U12344 ( .A1(n18899), .A2(n10816), .ZN(n19212) );
  INV_X1 U12345 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14833) );
  INV_X1 U12346 ( .A(n19212), .ZN(n16247) );
  INV_X1 U12347 ( .A(n19204), .ZN(n16265) );
  NOR2_X1 U12348 ( .A1(n16114), .A2(n11055), .ZN(n10950) );
  AND2_X1 U12349 ( .A1(n14950), .A2(n13947), .ZN(n14935) );
  NAND2_X1 U12350 ( .A1(n9907), .A2(n9911), .ZN(n15060) );
  NAND2_X1 U12351 ( .A1(n16232), .A2(n9912), .ZN(n9907) );
  NOR2_X1 U12352 ( .A1(n16233), .A2(n16292), .ZN(n15272) );
  NAND2_X1 U12353 ( .A1(n16232), .A2(n16229), .ZN(n9915) );
  NAND2_X1 U12354 ( .A1(n10054), .A2(n9847), .ZN(n14753) );
  INV_X1 U12355 ( .A(n19233), .ZN(n16318) );
  NOR2_X1 U12356 ( .A1(n13601), .A2(n13606), .ZN(n13865) );
  INV_X1 U12357 ( .A(n15245), .ZN(n19214) );
  NAND2_X1 U12358 ( .A1(n11259), .A2(n11257), .ZN(n15346) );
  INV_X1 U12359 ( .A(n19225), .ZN(n16323) );
  NAND2_X1 U12360 ( .A1(n13165), .A2(n13164), .ZN(n19881) );
  INV_X1 U12361 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19868) );
  NAND2_X1 U12362 ( .A1(n13260), .A2(n13263), .ZN(n13264) );
  AND2_X1 U12363 ( .A1(n13172), .A2(n13262), .ZN(n19871) );
  OR2_X1 U12364 ( .A1(n13171), .A2(n13170), .ZN(n13172) );
  CLKBUF_X1 U12365 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n16336) );
  INV_X1 U12366 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15505) );
  OAI21_X1 U12367 ( .B1(n13723), .B2(n13812), .A(n13717), .ZN(n19410) );
  OAI21_X1 U12368 ( .B1(n13723), .B2(n13722), .A(n13721), .ZN(n19407) );
  AND2_X1 U12369 ( .A1(n19448), .A2(n19447), .ZN(n19504) );
  OAI21_X1 U12370 ( .B1(n19519), .B2(n19518), .A(n19517), .ZN(n19536) );
  OAI21_X1 U12371 ( .B1(n19548), .B2(n19563), .A(n19683), .ZN(n19566) );
  NOR2_X2 U12372 ( .A1(n19651), .A2(n19511), .ZN(n19565) );
  INV_X1 U12373 ( .A(n19733), .ZN(n19592) );
  OAI22_X1 U12374 ( .A1(n19270), .A2(n19277), .B1(n19269), .B2(n19276), .ZN(
        n19595) );
  OAI22_X1 U12375 ( .A1(n21050), .A2(n19276), .B1(n19264), .B2(n19277), .ZN(
        n19628) );
  INV_X1 U12376 ( .A(n19720), .ZN(n19658) );
  INV_X1 U12377 ( .A(n19667), .ZN(n19671) );
  NOR2_X1 U12378 ( .A1(n19646), .A2(n19642), .ZN(n19670) );
  AND2_X1 U12379 ( .A1(n10266), .A2(n13651), .ZN(n19697) );
  OAI22_X1 U12380 ( .A1(n20139), .A2(n19277), .B1(n18233), .B2(n19276), .ZN(
        n19698) );
  OAI21_X1 U12381 ( .B1(n19712), .B2(n19684), .A(n19683), .ZN(n19715) );
  OAI22_X1 U12382 ( .A1(n20118), .A2(n19277), .B1(n18223), .B2(n19276), .ZN(
        n19677) );
  NOR2_X2 U12383 ( .A1(n19651), .A2(n19451), .ZN(n19740) );
  INV_X1 U12384 ( .A(n19631), .ZN(n19739) );
  INV_X1 U12385 ( .A(n19628), .ZN(n19744) );
  AND2_X1 U12386 ( .A1(n16371), .A2(n16370), .ZN(n19763) );
  INV_X1 U12387 ( .A(n17462), .ZN(n17464) );
  AOI21_X1 U12388 ( .B1(n9819), .B2(n18684), .A(n17464), .ZN(n18887) );
  NAND2_X1 U12389 ( .A1(n18868), .A2(n18714), .ZN(n16562) );
  NOR2_X1 U12390 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16660), .ZN(n16645) );
  NOR2_X1 U12391 ( .A1(n16653), .A2(n9897), .ZN(n16647) );
  NOR2_X1 U12392 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16680), .ZN(n16667) );
  NOR2_X1 U12393 ( .A1(n16699), .A2(n17615), .ZN(n16698) );
  NOR2_X1 U12394 ( .A1(n16858), .A2(n16590), .ZN(n16707) );
  NOR2_X1 U12395 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16746), .ZN(n16729) );
  NOR2_X1 U12396 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16818), .ZN(n16805) );
  INV_X1 U12397 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n20968) );
  INV_X1 U12398 ( .A(n16935), .ZN(n16909) );
  INV_X1 U12399 ( .A(n16946), .ZN(n16937) );
  INV_X1 U12400 ( .A(n16947), .ZN(n16911) );
  NAND4_X1 U12401 ( .A1(n15697), .A2(n18885), .A3(n16926), .A4(n18722), .ZN(
        n16945) );
  AND2_X1 U12402 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17131), .ZN(n17115) );
  NOR2_X1 U12403 ( .A1(n16796), .A2(n17156), .ZN(n17131) );
  NAND2_X1 U12404 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17172), .ZN(n17156) );
  NAND2_X1 U12405 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17202), .ZN(n17186) );
  NAND2_X1 U12406 ( .A1(n17256), .A2(n17236), .ZN(n17231) );
  NAND2_X1 U12407 ( .A1(n17289), .A2(n9814), .ZN(n17277) );
  NAND2_X1 U12408 ( .A1(n17289), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n17285) );
  NOR2_X1 U12409 ( .A1(n17416), .A2(n17295), .ZN(n17289) );
  OR2_X1 U12410 ( .A1(n17475), .A2(n17294), .ZN(n17295) );
  NOR2_X1 U12411 ( .A1(n17301), .A2(n17419), .ZN(n17300) );
  NOR2_X1 U12412 ( .A1(n17467), .A2(n17329), .ZN(n17330) );
  NOR3_X1 U12413 ( .A1(n17370), .A2(n17346), .A3(n17263), .ZN(n17347) );
  NOR3_X1 U12414 ( .A1(n17402), .A2(n17262), .A3(n17261), .ZN(n17371) );
  NOR2_X1 U12415 ( .A1(n15536), .A2(n15535), .ZN(n17388) );
  AND2_X1 U12416 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17391), .ZN(n17396) );
  NAND2_X1 U12417 ( .A1(n9986), .A2(n9823), .ZN(n17260) );
  NAND2_X1 U12418 ( .A1(n15771), .A2(n18868), .ZN(n9986) );
  INV_X1 U12419 ( .A(n17397), .ZN(n17400) );
  CLKBUF_X1 U12420 ( .A(n17505), .Z(n17501) );
  NOR2_X1 U12421 ( .A1(n17464), .A2(n18717), .ZN(n17505) );
  CLKBUF_X1 U12422 ( .A(n17504), .Z(n17511) );
  NOR2_X1 U12423 ( .A1(n17511), .A2(n18227), .ZN(n17512) );
  INV_X1 U12424 ( .A(n16858), .ZN(n16907) );
  NOR2_X1 U12425 ( .A1(n18834), .A2(n17877), .ZN(n17538) );
  OR2_X1 U12426 ( .A1(n17526), .A2(n17525), .ZN(n17527) );
  NOR2_X1 U12427 ( .A1(n17561), .A2(n17562), .ZN(n17548) );
  NOR2_X1 U12428 ( .A1(n16436), .A2(n17885), .ZN(n17711) );
  INV_X1 U12429 ( .A(n17538), .ZN(n17740) );
  INV_X1 U12430 ( .A(n17794), .ZN(n17748) );
  OAI22_X1 U12431 ( .A1(n17994), .A2(n17886), .B1(n17993), .B2(n17789), .ZN(
        n17775) );
  AND2_X1 U12432 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17782) );
  INV_X1 U12433 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17785) );
  INV_X1 U12434 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17798) );
  INV_X1 U12435 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17815) );
  NOR2_X1 U12436 ( .A1(n18227), .A2(n16562), .ZN(n17832) );
  NAND2_X1 U12437 ( .A1(n17515), .A2(n17882), .ZN(n17877) );
  NOR2_X1 U12438 ( .A1(n16394), .A2(n16562), .ZN(n17874) );
  INV_X1 U12439 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18834) );
  OAI21_X1 U12440 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18867), .A(n16562), 
        .ZN(n17882) );
  INV_X1 U12441 ( .A(n17874), .ZN(n17886) );
  OR2_X1 U12442 ( .A1(n18199), .A2(n17781), .ZN(n10098) );
  INV_X1 U12443 ( .A(n10097), .ZN(n17536) );
  NOR2_X1 U12444 ( .A1(n17993), .A2(n17672), .ZN(n18025) );
  AND2_X1 U12445 ( .A1(n10090), .A2(n9804), .ZN(n17813) );
  NAND2_X1 U12446 ( .A1(n17839), .A2(n15617), .ZN(n17823) );
  INV_X1 U12447 ( .A(n18185), .ZN(n18190) );
  NOR2_X1 U12448 ( .A1(n9760), .A2(n18184), .ZN(n18185) );
  INV_X1 U12449 ( .A(n18694), .ZN(n18206) );
  NOR2_X1 U12450 ( .A1(n18205), .A2(n18664), .ZN(n18204) );
  NOR2_X1 U12451 ( .A1(n10087), .A2(n17880), .ZN(n18201) );
  INV_X1 U12452 ( .A(n17873), .ZN(n10087) );
  INV_X1 U12453 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18217) );
  NOR2_X1 U12454 ( .A1(n18873), .A2(n16556), .ZN(n18470) );
  INV_X1 U12455 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18704) );
  INV_X1 U12456 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18708) );
  INV_X1 U12457 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18848) );
  INV_X1 U12458 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18230) );
  NAND2_X1 U12459 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18834), .ZN(n18729) );
  NAND2_X1 U12460 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n18875) );
  CLKBUF_X1 U12461 ( .A(n16546), .Z(n16544) );
  OAI21_X1 U12462 ( .B1(n14396), .B2(n20115), .A(n12286), .ZN(n12287) );
  OAI21_X1 U12463 ( .B1(n14566), .B2(n20102), .A(n9888), .ZN(n9887) );
  AOI211_X1 U12464 ( .C1(n14078), .C2(n19233), .A(n14077), .B(n14076), .ZN(
        n14079) );
  NAND2_X1 U12465 ( .A1(n14075), .A2(n14074), .ZN(n14076) );
  INV_X1 U12466 ( .A(n9927), .ZN(n12508) );
  NOR2_X1 U12467 ( .A1(n10369), .A2(n9800), .ZN(n10491) );
  INV_X2 U12468 ( .A(n14460), .ZN(n15893) );
  NOR2_X2 U12469 ( .A1(n12971), .A2(n9971), .ZN(n9796) );
  AND2_X1 U12470 ( .A1(n13839), .A2(n9863), .ZN(n13904) );
  OR2_X1 U12471 ( .A1(n13888), .A2(n10052), .ZN(n9798) );
  OR2_X1 U12472 ( .A1(n13709), .A2(n9841), .ZN(n9799) );
  NAND2_X1 U12473 ( .A1(n10119), .A2(n10117), .ZN(n15303) );
  AND2_X1 U12474 ( .A1(n14006), .A2(n10081), .ZN(n14341) );
  NAND2_X1 U12475 ( .A1(n11293), .A2(n9848), .ZN(n14738) );
  OR2_X1 U12476 ( .A1(n13313), .A2(n13265), .ZN(n9800) );
  INV_X1 U12477 ( .A(n14707), .ZN(n14704) );
  OR2_X1 U12478 ( .A1(n14211), .A2(n10085), .ZN(n12313) );
  INV_X1 U12479 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17741) );
  NAND2_X1 U12480 ( .A1(n14994), .A2(n10740), .ZN(n9802) );
  NAND2_X1 U12481 ( .A1(n10091), .A2(n18145), .ZN(n9804) );
  OR2_X1 U12482 ( .A1(n11299), .A2(n9914), .ZN(n9805) );
  AND2_X1 U12483 ( .A1(n10070), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9806) );
  OR4_X1 U12484 ( .A1(n19030), .A2(n19050), .A3(n18895), .A4(n16359), .ZN(
        n9807) );
  NAND2_X1 U12485 ( .A1(n13577), .A2(n9820), .ZN(n13663) );
  INV_X1 U12486 ( .A(n12515), .ZN(n10016) );
  AND2_X1 U12487 ( .A1(n10060), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9808) );
  OR2_X1 U12488 ( .A1(n10078), .A2(n9876), .ZN(n9809) );
  AND2_X1 U12489 ( .A1(n13608), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n9810) );
  AND2_X1 U12490 ( .A1(n9871), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9811) );
  AND2_X1 U12491 ( .A1(n10066), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9812) );
  NAND2_X1 U12492 ( .A1(n11756), .A2(n14521), .ZN(n9813) );
  AND2_X1 U12493 ( .A1(n9984), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n9814) );
  NOR2_X1 U12494 ( .A1(n12920), .A2(n16921), .ZN(n15601) );
  INV_X1 U12495 ( .A(n15601), .ZN(n12917) );
  OR2_X1 U12496 ( .A1(n14045), .A2(n14046), .ZN(n9815) );
  AND2_X2 U12497 ( .A1(n12863), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10456) );
  INV_X1 U12498 ( .A(n15559), .ZN(n17012) );
  NAND2_X1 U12499 ( .A1(n10250), .A2(n10249), .ZN(n10268) );
  NAND2_X1 U12500 ( .A1(n14526), .A2(n14525), .ZN(n14510) );
  INV_X2 U12501 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n11495) );
  INV_X2 U12502 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15408) );
  INV_X1 U12503 ( .A(n9938), .ZN(n10699) );
  NAND2_X1 U12504 ( .A1(n10113), .A2(n15162), .ZN(n13941) );
  AND2_X1 U12505 ( .A1(n10651), .A2(n9952), .ZN(n9816) );
  AND2_X1 U12506 ( .A1(n17347), .A2(n9981), .ZN(n9817) );
  OAI21_X1 U12507 ( .B1(n16232), .B2(n9910), .A(n9908), .ZN(n15048) );
  NAND2_X1 U12508 ( .A1(n10339), .A2(n10331), .ZN(n10818) );
  AND2_X1 U12509 ( .A1(n17289), .A2(n9984), .ZN(n9818) );
  NOR2_X1 U12510 ( .A1(n13003), .A2(n13916), .ZN(n9819) );
  AND2_X1 U12511 ( .A1(n13590), .A2(n13664), .ZN(n9820) );
  OR2_X1 U12512 ( .A1(n10027), .A2(n10028), .ZN(n9821) );
  NOR2_X1 U12513 ( .A1(n14874), .A2(n12738), .ZN(n12762) );
  NAND2_X1 U12514 ( .A1(n11465), .A2(n13243), .ZN(n9822) );
  INV_X1 U12515 ( .A(n16441), .ZN(n16448) );
  NAND2_X1 U12516 ( .A1(n15695), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16441) );
  OR3_X1 U12517 ( .A1(n16394), .A2(n18874), .A3(n15770), .ZN(n9823) );
  XNOR2_X1 U12518 ( .A(n10799), .B(n10800), .ZN(n10791) );
  NAND2_X1 U12519 ( .A1(n15016), .A2(n10708), .ZN(n15161) );
  AND2_X1 U12520 ( .A1(n15106), .A2(n10020), .ZN(n16273) );
  INV_X1 U12521 ( .A(n16462), .ZN(n16442) );
  NAND2_X1 U12522 ( .A1(n12531), .A2(n12530), .ZN(n13259) );
  NAND2_X1 U12523 ( .A1(n10039), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15088) );
  INV_X1 U12524 ( .A(n13815), .ZN(n10483) );
  AND4_X1 U12525 ( .A1(n10473), .A2(n10472), .A3(n10471), .A4(n10470), .ZN(
        n9824) );
  OR2_X1 U12526 ( .A1(n10676), .A2(n10671), .ZN(n9825) );
  AND2_X1 U12527 ( .A1(n10119), .A2(n10116), .ZN(n9826) );
  AND3_X1 U12528 ( .A1(n15070), .A2(n16230), .A3(n15078), .ZN(n9827) );
  AND2_X1 U12529 ( .A1(n9820), .A2(n9963), .ZN(n9828) );
  AND2_X1 U12530 ( .A1(n15624), .A2(n10100), .ZN(n9829) );
  AND2_X1 U12531 ( .A1(n9804), .A2(n17812), .ZN(n9830) );
  INV_X1 U12532 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15384) );
  OAI21_X1 U12533 ( .B1(n10332), .B2(n15384), .A(n10315), .ZN(n10345) );
  AND2_X1 U12534 ( .A1(n9938), .A2(n15187), .ZN(n9831) );
  OR2_X1 U12535 ( .A1(n10064), .A2(n15331), .ZN(n9832) );
  AND2_X1 U12536 ( .A1(n10111), .A2(n14993), .ZN(n9834) );
  NAND2_X1 U12537 ( .A1(n14263), .A2(n14252), .ZN(n14239) );
  NOR2_X1 U12538 ( .A1(n14211), .A2(n14212), .ZN(n12277) );
  NAND2_X1 U12539 ( .A1(n14504), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13965) );
  NAND2_X1 U12540 ( .A1(n9920), .A2(n10650), .ZN(n16240) );
  AND3_X1 U12541 ( .A1(n12966), .A2(n12965), .A3(n9972), .ZN(n9835) );
  AND2_X1 U12542 ( .A1(n10014), .A2(n12538), .ZN(n13603) );
  AND2_X1 U12543 ( .A1(n10564), .A2(n10559), .ZN(n9837) );
  AND2_X1 U12544 ( .A1(n11301), .A2(n9827), .ZN(n9838) );
  AND2_X1 U12545 ( .A1(n10097), .A2(n16442), .ZN(n9839) );
  NAND2_X1 U12546 ( .A1(n12784), .A2(n12783), .ZN(n14863) );
  NAND2_X1 U12547 ( .A1(n10513), .A2(n10515), .ZN(n10799) );
  NAND3_X1 U12548 ( .A1(n13016), .A2(n15418), .A3(n18227), .ZN(n9840) );
  INV_X1 U12549 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11310) );
  OR2_X1 U12550 ( .A1(n18086), .A2(n17754), .ZN(n17779) );
  OR2_X1 U12551 ( .A1(n13710), .A2(n9961), .ZN(n9841) );
  NAND2_X1 U12552 ( .A1(n13604), .A2(n12539), .ZN(n13609) );
  NOR2_X1 U12553 ( .A1(n14780), .A2(n14781), .ZN(n14766) );
  NAND2_X1 U12554 ( .A1(n13609), .A2(n13608), .ZN(n13380) );
  NAND2_X1 U12555 ( .A1(n13839), .A2(n10043), .ZN(n9842) );
  INV_X1 U12556 ( .A(n9891), .ZN(n14324) );
  OR2_X1 U12557 ( .A1(n13749), .A2(n10078), .ZN(n9843) );
  AND2_X1 U12558 ( .A1(n14685), .A2(n10066), .ZN(n9844) );
  AND2_X1 U12559 ( .A1(n14692), .A2(n10060), .ZN(n9845) );
  AND2_X1 U12560 ( .A1(n10571), .A2(n10564), .ZN(n9846) );
  AND2_X1 U12561 ( .A1(n10059), .A2(n14767), .ZN(n9847) );
  AND2_X1 U12562 ( .A1(n14886), .A2(n14878), .ZN(n13944) );
  NOR2_X1 U12563 ( .A1(n13888), .A2(n15234), .ZN(n14970) );
  NOR3_X1 U12564 ( .A1(n13709), .A2(n9841), .A3(n13807), .ZN(n13806) );
  NOR3_X1 U12565 ( .A1(n13888), .A2(n10052), .A3(n12498), .ZN(n12497) );
  INV_X1 U12566 ( .A(n14082), .ZN(n10083) );
  AND2_X1 U12567 ( .A1(n11294), .A2(n9966), .ZN(n9848) );
  NAND2_X1 U12568 ( .A1(n15941), .A2(n11701), .ZN(n15935) );
  NAND2_X1 U12569 ( .A1(n11733), .A2(n11732), .ZN(n13897) );
  AND2_X1 U12570 ( .A1(n10018), .A2(n9775), .ZN(n9849) );
  AND2_X1 U12571 ( .A1(n11473), .A2(n11456), .ZN(n13234) );
  OR2_X1 U12572 ( .A1(n11304), .A2(n15026), .ZN(n9850) );
  OR2_X1 U12573 ( .A1(n10714), .A2(n15167), .ZN(n9851) );
  NAND2_X1 U12574 ( .A1(n10277), .A2(n10992), .ZN(n11001) );
  AND2_X1 U12575 ( .A1(n12807), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n9852) );
  NAND2_X1 U12576 ( .A1(n10077), .A2(n11902), .ZN(n13787) );
  NAND2_X1 U12577 ( .A1(n11293), .A2(n11294), .ZN(n11292) );
  AND3_X1 U12578 ( .A1(n10475), .A2(n10474), .A3(n9824), .ZN(n10787) );
  OR2_X1 U12579 ( .A1(n11677), .A2(n11777), .ZN(n9853) );
  NOR2_X1 U12580 ( .A1(n14882), .A2(n12714), .ZN(n9854) );
  NOR2_X1 U12581 ( .A1(n9958), .A2(n14907), .ZN(n11293) );
  NAND2_X1 U12582 ( .A1(n10119), .A2(n10114), .ZN(n15092) );
  AND2_X1 U12583 ( .A1(n10650), .A2(n9923), .ZN(n9855) );
  NOR2_X1 U12584 ( .A1(n11195), .A2(n11055), .ZN(n9856) );
  OR2_X1 U12585 ( .A1(n10640), .A2(n9948), .ZN(n9857) );
  INV_X1 U12586 ( .A(n9913), .ZN(n9912) );
  NAND2_X1 U12587 ( .A1(n16229), .A2(n9916), .ZN(n9913) );
  OR2_X1 U12588 ( .A1(n9992), .A2(n14567), .ZN(n9858) );
  NOR2_X1 U12589 ( .A1(n13709), .A2(n13710), .ZN(n13711) );
  AND2_X1 U12590 ( .A1(n9810), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n9859)
         );
  INV_X1 U12591 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n19041) );
  OR2_X1 U12592 ( .A1(n14450), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9860) );
  NAND2_X1 U12593 ( .A1(n14886), .A2(n9969), .ZN(n14045) );
  AND2_X1 U12594 ( .A1(n14886), .A2(n9970), .ZN(n13943) );
  AND2_X1 U12595 ( .A1(n10425), .A2(n9924), .ZN(n9861) );
  INV_X1 U12596 ( .A(n13168), .ZN(n14901) );
  NOR2_X1 U12597 ( .A1(n16076), .A2(n16075), .ZN(n9862) );
  AND2_X1 U12598 ( .A1(n13609), .A2(n9810), .ZN(n13373) );
  NOR2_X1 U12599 ( .A1(n13374), .A2(n10842), .ZN(n13577) );
  NOR2_X1 U12600 ( .A1(n14780), .A2(n10057), .ZN(n14752) );
  NAND2_X1 U12601 ( .A1(n13760), .A2(n9968), .ZN(n13375) );
  NOR2_X1 U12602 ( .A1(n13780), .A2(n13879), .ZN(n13830) );
  NAND2_X1 U12603 ( .A1(n16076), .A2(n13791), .ZN(n13790) );
  AND2_X1 U12604 ( .A1(n13256), .A2(n13250), .ZN(n20076) );
  AND2_X1 U12605 ( .A1(n14681), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14041) );
  INV_X1 U12606 ( .A(n15069), .ZN(n9916) );
  AND2_X1 U12607 ( .A1(n19212), .A2(n14123), .ZN(n19203) );
  AND2_X1 U12608 ( .A1(n13577), .A2(n13590), .ZN(n13589) );
  INV_X1 U12609 ( .A(n17674), .ZN(n17781) );
  NOR2_X2 U12610 ( .A1(n17374), .A2(n16445), .ZN(n17674) );
  NOR2_X1 U12611 ( .A1(n13581), .A2(n12581), .ZN(n13803) );
  AND2_X1 U12612 ( .A1(n10044), .A2(n14906), .ZN(n9863) );
  AND2_X1 U12613 ( .A1(n13577), .A2(n9828), .ZN(n13700) );
  NAND2_X1 U12614 ( .A1(n10090), .A2(n9830), .ZN(n17811) );
  AND2_X1 U12615 ( .A1(n10808), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9864) );
  NOR2_X1 U12616 ( .A1(n14844), .A2(n10030), .ZN(n10029) );
  AND2_X1 U12617 ( .A1(n10072), .A2(n11245), .ZN(n9865) );
  OR2_X1 U12618 ( .A1(n14176), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9866) );
  NAND2_X1 U12619 ( .A1(n10642), .A2(n16248), .ZN(n9867) );
  INV_X1 U12620 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20105) );
  INV_X1 U12621 ( .A(n11055), .ZN(n10808) );
  AND3_X1 U12622 ( .A1(n10537), .A2(n10536), .A3(n10535), .ZN(n11055) );
  AND2_X1 U12623 ( .A1(n13863), .A2(n11052), .ZN(n9868) );
  AND2_X1 U12624 ( .A1(n17839), .A2(n10093), .ZN(n9869) );
  INV_X1 U12625 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n9896) );
  OR4_X1 U12626 ( .A1(n20931), .A2(n17421), .A3(n17428), .A4(n17467), .ZN(
        n9870) );
  INV_X1 U12627 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10100) );
  NAND2_X1 U12628 ( .A1(n11448), .A2(n13234), .ZN(n13241) );
  AND2_X1 U12629 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n9871) );
  XNOR2_X1 U12630 ( .A(n18227), .B(n18221), .ZN(n18884) );
  NAND2_X1 U12631 ( .A1(n17864), .A2(n17863), .ZN(n17862) );
  AND2_X1 U12632 ( .A1(n9795), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n9872) );
  AND2_X1 U12633 ( .A1(n12720), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n9873) );
  AND2_X1 U12634 ( .A1(n9795), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n9874)
         );
  AND2_X1 U12635 ( .A1(n12782), .A2(n12807), .ZN(n9875) );
  AND2_X1 U12636 ( .A1(n11933), .A2(n11932), .ZN(n9876) );
  OR2_X1 U12637 ( .A1(n13394), .A2(n9883), .ZN(n9877) );
  INV_X1 U12638 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n9943) );
  AND2_X1 U12639 ( .A1(n9811), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9878) );
  AND2_X1 U12640 ( .A1(n17627), .A2(n9894), .ZN(n9879) );
  NAND2_X1 U12641 ( .A1(n15144), .A2(n12471), .ZN(n9880) );
  INV_X1 U12642 ( .A(n14856), .ZN(n10034) );
  INV_X1 U12643 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n9982) );
  INV_X1 U12644 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10071) );
  NOR2_X1 U12645 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16112), .ZN(n20006) );
  OR2_X1 U12646 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n9881) );
  INV_X1 U12647 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n9985) );
  INV_X1 U12648 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10068) );
  INV_X1 U12649 ( .A(n9807), .ZN(n9882) );
  INV_X1 U12650 ( .A(n18939), .ZN(n19771) );
  OAI221_X1 U12651 ( .B1(n20317), .B2(n21100), .C1(n20317), .C2(n20300), .A(
        n20649), .ZN(n20319) );
  INV_X1 U12652 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18824) );
  NOR3_X2 U12653 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n9746), .A3(
        n18352), .ZN(n18280) );
  NOR3_X2 U12654 ( .A1(n9746), .A2(n18699), .A3(n18352), .ZN(n18325) );
  NOR3_X2 U12655 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n9746), .A3(
        n18445), .ZN(n18416) );
  NOR3_X2 U12656 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n9746), .A3(
        n18491), .ZN(n18462) );
  NOR3_X2 U12657 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n9746), .A3(
        n18399), .ZN(n18369) );
  AOI221_X2 U12658 ( .B1(n18565), .B2(n18566), .C1(n18564), .C2(n18566), .A(
        n18563), .ZN(n18600) );
  AND2_X1 U12659 ( .A1(n11319), .A2(n9883), .ZN(n11379) );
  AND2_X2 U12660 ( .A1(n14224), .A2(n14210), .ZN(n14208) );
  AND2_X2 U12661 ( .A1(n12440), .A2(n9884), .ZN(n14224) );
  NAND3_X1 U12662 ( .A1(n9886), .A2(n13569), .A3(n9885), .ZN(n16090) );
  NOR2_X2 U12663 ( .A1(n16092), .A2(n13730), .ZN(n16074) );
  NAND2_X1 U12664 ( .A1(n12382), .A2(n12381), .ZN(n16092) );
  INV_X1 U12665 ( .A(n9887), .ZN(n14575) );
  NOR2_X1 U12666 ( .A1(n14573), .A2(n14574), .ZN(n9888) );
  NAND2_X1 U12667 ( .A1(n14174), .A2(n14173), .ZN(n9889) );
  NAND3_X1 U12668 ( .A1(n12448), .A2(n10135), .A3(n12358), .ZN(n9892) );
  INV_X2 U12669 ( .A(n12460), .ZN(n12448) );
  NAND2_X1 U12670 ( .A1(n12361), .A2(n9892), .ZN(n12363) );
  CLKBUF_X1 U12671 ( .A(n16858), .Z(n9897) );
  AND2_X4 U12672 ( .A1(n10388), .A2(n9780), .ZN(n12838) );
  NAND2_X1 U12673 ( .A1(n10311), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10332) );
  OR2_X2 U12674 ( .A1(n9899), .A2(n10326), .ZN(n9906) );
  NAND2_X1 U12675 ( .A1(n9900), .A2(n10327), .ZN(n9899) );
  NAND2_X1 U12676 ( .A1(n10299), .A2(n9901), .ZN(n9900) );
  NAND2_X1 U12677 ( .A1(n9906), .A2(n9904), .ZN(n9902) );
  NAND3_X1 U12678 ( .A1(n10210), .A2(n10206), .A3(n10207), .ZN(n9917) );
  NAND2_X2 U12679 ( .A1(n10211), .A2(n9919), .ZN(n11014) );
  NAND3_X1 U12680 ( .A1(n9926), .A2(n9925), .A3(n9861), .ZN(n10514) );
  NAND4_X1 U12681 ( .A1(n10432), .A2(n10434), .A3(n10435), .A4(n10433), .ZN(
        n9925) );
  NAND4_X1 U12682 ( .A1(n10379), .A2(n10378), .A3(n10377), .A4(n10376), .ZN(
        n9926) );
  NAND2_X4 U12683 ( .A1(n10992), .A2(n9801), .ZN(n10905) );
  OAI22_X1 U12684 ( .A1(n12496), .A2(n19225), .B1(n16299), .B2(n18924), .ZN(
        n9927) );
  XNOR2_X1 U12685 ( .A(n15025), .B(n9850), .ZN(n12496) );
  NAND3_X1 U12686 ( .A1(n10563), .A2(n10571), .A3(n9837), .ZN(n9937) );
  NAND2_X1 U12687 ( .A1(n9846), .A2(n10563), .ZN(n10577) );
  NAND4_X1 U12688 ( .A1(n9940), .A2(n15024), .A3(n9838), .A4(n15023), .ZN(
        n9938) );
  OAI21_X2 U12689 ( .B1(n10738), .B2(n9947), .A(n9946), .ZN(n14985) );
  AND2_X1 U12690 ( .A1(n14842), .A2(n14841), .ZN(n10913) );
  INV_X1 U12691 ( .A(n14168), .ZN(n14717) );
  INV_X1 U12692 ( .A(n13836), .ZN(n9960) );
  NAND3_X1 U12693 ( .A1(n9967), .A2(n9968), .A3(n13760), .ZN(n13374) );
  NAND3_X1 U12694 ( .A1(n12964), .A2(n9973), .A3(n9835), .ZN(n9971) );
  INV_X1 U12695 ( .A(n18884), .ZN(n9977) );
  NAND2_X1 U12696 ( .A1(n9783), .A2(n9977), .ZN(n9975) );
  NAND3_X1 U12697 ( .A1(n9976), .A2(n9975), .A3(n9840), .ZN(n9974) );
  INV_X1 U12698 ( .A(n9978), .ZN(n16561) );
  AND2_X2 U12699 ( .A1(n11310), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11320) );
  NOR2_X1 U12700 ( .A1(n14092), .A2(n9992), .ZN(n14093) );
  AND2_X2 U12701 ( .A1(n14469), .A2(n13969), .ZN(n14092) );
  OR2_X1 U12702 ( .A1(n14092), .A2(n9858), .ZN(n9997) );
  INV_X1 U12703 ( .A(n14588), .ZN(n9998) );
  NAND2_X2 U12704 ( .A1(n9999), .A2(n11553), .ZN(n20188) );
  INV_X1 U12705 ( .A(n20258), .ZN(n9999) );
  OAI21_X1 U12706 ( .B1(n11565), .B2(n11549), .A(n11548), .ZN(n10000) );
  NAND2_X1 U12707 ( .A1(n13965), .A2(n10001), .ZN(n14477) );
  NAND3_X1 U12708 ( .A1(n10005), .A2(n11590), .A3(n11495), .ZN(n10004) );
  NAND3_X1 U12709 ( .A1(n10007), .A2(n11712), .A3(n10006), .ZN(n15929) );
  NAND2_X1 U12710 ( .A1(n11710), .A2(n10008), .ZN(n10006) );
  NAND3_X1 U12711 ( .A1(n15943), .A2(n11710), .A3(n15942), .ZN(n10007) );
  NAND2_X1 U12712 ( .A1(n11733), .A2(n10009), .ZN(n14553) );
  NAND2_X1 U12713 ( .A1(n13148), .A2(n13157), .ZN(n13133) );
  AND2_X2 U12714 ( .A1(n10010), .A2(n13241), .ZN(n11465) );
  NAND2_X1 U12715 ( .A1(n14526), .A2(n10012), .ZN(n11753) );
  AND2_X4 U12716 ( .A1(n10388), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12861) );
  NAND2_X1 U12717 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10364) );
  INV_X1 U12718 ( .A(n10312), .ZN(n13039) );
  INV_X1 U12719 ( .A(n10283), .ZN(n10013) );
  AND2_X2 U12720 ( .A1(n10958), .A2(n10269), .ZN(n10273) );
  NAND2_X1 U12721 ( .A1(n10789), .A2(n13866), .ZN(n10017) );
  NAND2_X1 U12722 ( .A1(n10794), .A2(n13855), .ZN(n10793) );
  NAND3_X1 U12723 ( .A1(n10018), .A2(n10017), .A3(n13854), .ZN(n10794) );
  NAND3_X1 U12724 ( .A1(n10020), .A2(n15106), .A3(n16274), .ZN(n10019) );
  NAND2_X2 U12725 ( .A1(n10455), .A2(n10454), .ZN(n10786) );
  NAND3_X1 U12726 ( .A1(n14848), .A2(n14857), .A3(n12852), .ZN(n10024) );
  NAND2_X1 U12727 ( .A1(n12714), .A2(n10038), .ZN(n10035) );
  CLKBUF_X1 U12728 ( .A(n9781), .Z(n10039) );
  AND2_X1 U12729 ( .A1(n9781), .A2(n10041), .ZN(n11284) );
  NAND2_X1 U12730 ( .A1(n9781), .A2(n10040), .ZN(n15006) );
  NAND2_X1 U12731 ( .A1(n13839), .A2(n10042), .ZN(n12712) );
  OAI21_X1 U12732 ( .B1(n10795), .B2(n9836), .A(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n10045) );
  NAND2_X1 U12733 ( .A1(n10046), .A2(n10797), .ZN(n15118) );
  NAND2_X1 U12734 ( .A1(n10798), .A2(n10795), .ZN(n10046) );
  INV_X1 U12735 ( .A(n10797), .ZN(n9836) );
  NOR3_X2 U12736 ( .A1(n13888), .A2(n10052), .A3(n10050), .ZN(n14742) );
  INV_X1 U12737 ( .A(n14780), .ZN(n10054) );
  NAND2_X1 U12738 ( .A1(n10054), .A2(n10055), .ZN(n15256) );
  OAI21_X2 U12739 ( .B1(n13601), .B2(n9832), .A(n10062), .ZN(n15324) );
  AOI22_X1 U12740 ( .A1(n9795), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12838), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12721) );
  AOI22_X1 U12741 ( .A1(n9795), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12838), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12745) );
  AOI22_X1 U12742 ( .A1(n9795), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12863), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12855) );
  NAND2_X1 U12743 ( .A1(n11874), .A2(n11873), .ZN(n13733) );
  INV_X1 U12744 ( .A(n13732), .ZN(n10073) );
  NOR2_X2 U12745 ( .A1(n14239), .A2(n14240), .ZN(n14221) );
  NOR2_X2 U12746 ( .A1(n14331), .A2(n14264), .ZN(n14263) );
  NAND2_X1 U12747 ( .A1(n11676), .A2(n11675), .ZN(n20107) );
  NAND4_X1 U12748 ( .A1(n11465), .A2(n11478), .A3(n11493), .A4(n13243), .ZN(
        n10076) );
  OAI21_X2 U12749 ( .B1(n11565), .B2(n11311), .A(n11479), .ZN(n11551) );
  NAND2_X2 U12750 ( .A1(n10076), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11565) );
  NOR2_X2 U12751 ( .A1(n13749), .A2(n9809), .ZN(n13909) );
  NAND2_X1 U12752 ( .A1(n17871), .A2(n15609), .ZN(n17863) );
  XNOR2_X1 U12753 ( .A(n15610), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n17864) );
  NOR2_X2 U12754 ( .A1(n17550), .A2(n15694), .ZN(n15695) );
  NAND2_X1 U12755 ( .A1(n17839), .A2(n10088), .ZN(n10090) );
  NAND2_X2 U12756 ( .A1(n17667), .A2(n17781), .ZN(n17635) );
  NAND2_X1 U12757 ( .A1(n16462), .A2(n10099), .ZN(n10095) );
  NOR2_X1 U12758 ( .A1(n17520), .A2(n10098), .ZN(n16443) );
  NAND3_X1 U12759 ( .A1(n9829), .A2(n17781), .A3(n17795), .ZN(n17765) );
  INV_X2 U12760 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13018) );
  AND2_X4 U12761 ( .A1(n10385), .A2(n9780), .ZN(n12853) );
  INV_X1 U12762 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10101) );
  NAND2_X1 U12763 ( .A1(n10102), .A2(n19043), .ZN(n10583) );
  NAND3_X1 U12764 ( .A1(n10517), .A2(n11055), .A3(n10799), .ZN(n10102) );
  NAND2_X1 U12765 ( .A1(n10283), .A2(n10270), .ZN(n10955) );
  INV_X1 U12766 ( .A(n10955), .ZN(n10103) );
  NAND2_X1 U12767 ( .A1(n10103), .A2(n19259), .ZN(n10965) );
  NAND3_X1 U12768 ( .A1(n10105), .A2(n15188), .A3(n10104), .ZN(n15015) );
  NAND3_X1 U12769 ( .A1(n11296), .A2(n10107), .A3(n15187), .ZN(n10105) );
  NAND2_X1 U12770 ( .A1(n10106), .A2(n10699), .ZN(n15186) );
  AND2_X1 U12771 ( .A1(n10113), .A2(n10111), .ZN(n12467) );
  OR2_X1 U12772 ( .A1(n13581), .A2(n13580), .ZN(n13583) );
  INV_X1 U12773 ( .A(n11451), .ZN(n13236) );
  NOR2_X1 U12774 ( .A1(n20145), .A2(n11451), .ZN(n11477) );
  CLKBUF_X1 U12775 ( .A(n14300), .Z(n20642) );
  NAND2_X1 U12776 ( .A1(n20160), .A2(n13244), .ZN(n11461) );
  AND3_X1 U12777 ( .A1(n11472), .A2(n12350), .A3(n13244), .ZN(n11393) );
  NAND2_X2 U12778 ( .A1(n10236), .A2(n10235), .ZN(n10266) );
  INV_X1 U12779 ( .A(n11837), .ZN(n11556) );
  AND2_X1 U12780 ( .A1(n11551), .A2(n11550), .ZN(n11552) );
  OAI21_X1 U12781 ( .B1(n11837), .B2(n13291), .A(n11662), .ZN(n11670) );
  AND4_X1 U12782 ( .A1(n10965), .A2(n10989), .A3(n10964), .A4(n10963), .ZN(
        n10985) );
  NAND2_X1 U12783 ( .A1(n10965), .A2(n10253), .ZN(n10988) );
  AND2_X1 U12784 ( .A1(n10539), .A2(n10267), .ZN(n10261) );
  NOR2_X1 U12785 ( .A1(n10266), .A2(n10265), .ZN(n10269) );
  INV_X1 U12786 ( .A(n10190), .ZN(n10191) );
  CLKBUF_X1 U12787 ( .A(n12853), .Z(n12863) );
  AND4_X1 U12788 ( .A1(n10367), .A2(n10366), .A3(n10365), .A4(n10364), .ZN(
        n10378) );
  OAI22_X1 U12789 ( .A1(n10905), .A2(n10325), .B1(n10329), .B2(n10324), .ZN(
        n10326) );
  NOR2_X1 U12790 ( .A1(n12924), .A2(n12923), .ZN(n15463) );
  INV_X2 U12791 ( .A(n15594), .ZN(n17209) );
  NOR2_X2 U12792 ( .A1(n13030), .A2(n12923), .ZN(n15593) );
  BUF_X4 U12793 ( .A(n15593), .Z(n17213) );
  AND2_X1 U12794 ( .A1(n20054), .A2(n13977), .ZN(n20081) );
  NAND2_X2 U12795 ( .A1(n20001), .A2(n13321), .ZN(n20004) );
  NAND2_X1 U12796 ( .A1(n12785), .A2(n9875), .ZN(n10121) );
  INV_X1 U12797 ( .A(n12763), .ZN(n12759) );
  AND2_X1 U12798 ( .A1(n14092), .A2(n13970), .ZN(n10122) );
  OR2_X1 U12799 ( .A1(n14460), .A2(n16059), .ZN(n10123) );
  INV_X1 U12800 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11766) );
  INV_X1 U12801 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20515) );
  AND2_X1 U12802 ( .A1(n15463), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10124) );
  AND4_X1 U12803 ( .A1(n11172), .A2(n11171), .A3(n11170), .A4(n11169), .ZN(
        n10125) );
  AND4_X1 U12804 ( .A1(n11066), .A2(n11065), .A3(n11064), .A4(n11063), .ZN(
        n10126) );
  AND2_X1 U12805 ( .A1(n11752), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10127) );
  AND2_X1 U12806 ( .A1(n17674), .A2(n15692), .ZN(n10128) );
  AND2_X1 U12807 ( .A1(n20000), .A2(n11456), .ZN(n19996) );
  INV_X2 U12808 ( .A(n19996), .ZN(n14389) );
  NAND2_X1 U12809 ( .A1(n13133), .A2(n13140), .ZN(n10129) );
  INV_X1 U12810 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15681) );
  AND2_X1 U12811 ( .A1(n15894), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10130) );
  AND2_X1 U12812 ( .A1(n10941), .A2(n10940), .ZN(n10131) );
  OR2_X1 U12813 ( .A1(n10140), .A2(n13582), .ZN(n10132) );
  AND3_X1 U12814 ( .A1(n18080), .A2(n18047), .A3(n15683), .ZN(n10133) );
  OR2_X1 U12815 ( .A1(n14176), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10134) );
  INV_X1 U12816 ( .A(n17394), .ZN(n17399) );
  INV_X1 U12817 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n10329) );
  INV_X1 U12818 ( .A(n11018), .ZN(n11196) );
  AND2_X1 U12819 ( .A1(n12355), .A2(n11464), .ZN(n10135) );
  AND4_X1 U12820 ( .A1(n11136), .A2(n11135), .A3(n11134), .A4(n11133), .ZN(
        n10136) );
  NAND2_X1 U12821 ( .A1(n20000), .A2(n14087), .ZN(n19986) );
  AND2_X1 U12822 ( .A1(n10943), .A2(n14983), .ZN(n10137) );
  INV_X1 U12823 ( .A(n14993), .ZN(n10732) );
  OR2_X1 U12824 ( .A1(n18834), .A2(n17881), .ZN(n18869) );
  INV_X1 U12825 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13219) );
  XOR2_X1 U12826 ( .A(n19235), .B(n10780), .Z(n10138) );
  AND2_X1 U12827 ( .A1(n9756), .A2(n17247), .ZN(n17254) );
  OR2_X1 U12828 ( .A1(n17634), .A2(n16458), .ZN(n10139) );
  OR2_X1 U12829 ( .A1(n12580), .A2(n13658), .ZN(n10140) );
  AND3_X1 U12830 ( .A1(n10488), .A2(n10487), .A3(n10486), .ZN(n10141) );
  NAND2_X1 U12831 ( .A1(n13167), .A2(n19768), .ZN(n13168) );
  OR2_X1 U12832 ( .A1(n18899), .A2(n9788), .ZN(n16263) );
  INV_X1 U12833 ( .A(n16263), .ZN(n11305) );
  INV_X1 U12834 ( .A(n11022), .ZN(n11198) );
  INV_X1 U12835 ( .A(n13644), .ZN(n19207) );
  NAND3_X2 U12836 ( .A1(n19856), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19683), 
        .ZN(n13644) );
  OR2_X1 U12837 ( .A1(n18893), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15334) );
  AND2_X1 U12838 ( .A1(n11353), .A2(n11352), .ZN(n10142) );
  AND3_X1 U12839 ( .A1(n11355), .A2(n11354), .A3(n10142), .ZN(n10143) );
  OR2_X2 U12840 ( .A1(n12357), .A2(n12356), .ZN(n20000) );
  INV_X1 U12841 ( .A(n20182), .ZN(n20299) );
  NAND2_X1 U12842 ( .A1(n11495), .A2(n20119), .ZN(n20182) );
  INV_X1 U12843 ( .A(n13427), .ZN(n13428) );
  INV_X1 U12844 ( .A(n13141), .ZN(n11449) );
  NAND2_X1 U12845 ( .A1(n20160), .A2(n11473), .ZN(n11452) );
  OAI22_X1 U12846 ( .A1(n13815), .A2(n12767), .B1(n21006), .B2(n10485), .ZN(
        n10430) );
  NAND2_X1 U12847 ( .A1(n11452), .A2(n13236), .ZN(n11453) );
  OR2_X1 U12848 ( .A1(n11633), .A2(n11632), .ZN(n11705) );
  INV_X1 U12849 ( .A(n11457), .ZN(n11458) );
  AND4_X1 U12850 ( .A1(n10589), .A2(n10588), .A3(n10587), .A4(n10586), .ZN(
        n10593) );
  INV_X1 U12851 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15683) );
  AND2_X1 U12852 ( .A1(n20611), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11785) );
  AND2_X1 U12853 ( .A1(n11635), .A2(n11634), .ZN(n11690) );
  AOI22_X1 U12854 ( .A1(n12266), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12096), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11368) );
  AND2_X2 U12855 ( .A1(n11320), .A2(n11319), .ZN(n11412) );
  AOI22_X1 U12856 ( .A1(n9751), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10243), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10147) );
  AND4_X1 U12857 ( .A1(n10530), .A2(n10529), .A3(n10528), .A4(n10527), .ZN(
        n10532) );
  AOI22_X1 U12858 ( .A1(n10243), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12862), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10224) );
  AOI22_X1 U12859 ( .A1(n9752), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10243), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10167) );
  OAI21_X1 U12860 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n13018), .A(
        n13019), .ZN(n13020) );
  INV_X1 U12861 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11566) );
  AND2_X1 U12862 ( .A1(n11813), .A2(n11811), .ZN(n13137) );
  OR2_X1 U12863 ( .A1(n11647), .A2(n11646), .ZN(n11718) );
  OR2_X1 U12864 ( .A1(n11539), .A2(n11538), .ZN(n11658) );
  AOI21_X1 U12865 ( .B1(n11772), .B2(n11771), .A(n11769), .ZN(n11813) );
  AOI21_X1 U12866 ( .B1(n11010), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10314), 
        .ZN(n10315) );
  OR2_X1 U12867 ( .A1(n12689), .A2(n10518), .ZN(n10522) );
  AND2_X1 U12868 ( .A1(n14109), .A2(n12345), .ZN(n12346) );
  NOR2_X1 U12869 ( .A1(n12291), .A2(n12290), .ZN(n12292) );
  NAND2_X1 U12870 ( .A1(n12157), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12158) );
  INV_X1 U12871 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14033) );
  INV_X1 U12872 ( .A(n13789), .ZN(n11902) );
  AND2_X1 U12873 ( .A1(n11649), .A2(n11648), .ZN(n11702) );
  INV_X1 U12874 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n13967) );
  INV_X1 U12875 ( .A(n14526), .ZN(n11755) );
  MUX2_X1 U12876 ( .A(n10768), .B(n10325), .S(n19265), .Z(n10564) );
  OR2_X1 U12877 ( .A1(n10132), .A2(n13580), .ZN(n12581) );
  NAND4_X1 U12878 ( .A1(n10258), .A2(n19259), .A3(n19279), .A4(n12509), .ZN(
        n10254) );
  INV_X1 U12879 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14057) );
  INV_X1 U12880 ( .A(n14070), .ZN(n14071) );
  OR2_X1 U12881 ( .A1(n16170), .A2(n11055), .ZN(n10714) );
  AND2_X1 U12882 ( .A1(n18931), .A2(n10808), .ZN(n10695) );
  INV_X1 U12883 ( .A(n9782), .ZN(n10874) );
  NAND2_X1 U12884 ( .A1(n10802), .A2(n10801), .ZN(n10810) );
  NAND2_X1 U12885 ( .A1(n10794), .A2(n10791), .ZN(n10795) );
  NOR2_X1 U12886 ( .A1(n12921), .A2(n12919), .ZN(n15560) );
  NAND2_X1 U12887 ( .A1(n17674), .A2(n18023), .ZN(n15686) );
  NOR2_X1 U12888 ( .A1(n17388), .A2(n15612), .ZN(n15591) );
  OAI22_X1 U12889 ( .A1(n13018), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18704), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13023) );
  INV_X1 U12890 ( .A(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n20954) );
  INV_X1 U12891 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11951) );
  AND2_X1 U12892 ( .A1(n13680), .A2(n15741), .ZN(n13687) );
  OR2_X1 U12893 ( .A1(n14188), .A2(n12448), .ZN(n14174) );
  AND2_X1 U12894 ( .A1(n12388), .A2(n12387), .ZN(n16073) );
  INV_X1 U12895 ( .A(n12343), .ZN(n14084) );
  OR2_X1 U12896 ( .A1(n13674), .A2(n13973), .ZN(n13675) );
  NAND2_X1 U12897 ( .A1(n12201), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12202) );
  AND2_X1 U12898 ( .A1(n12071), .A2(n14276), .ZN(n12072) );
  AND2_X1 U12899 ( .A1(n14275), .A2(n14274), .ZN(n14276) );
  NOR2_X1 U12900 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13671) );
  INV_X1 U12901 ( .A(n13247), .ZN(n14176) );
  INV_X1 U12902 ( .A(n14460), .ZN(n14014) );
  NAND2_X1 U12903 ( .A1(n9787), .A2(n13459), .ZN(n12437) );
  INV_X1 U12904 ( .A(n13455), .ZN(n12369) );
  OAI21_X1 U12905 ( .B1(n20843), .B2(n16110), .A(n20821), .ZN(n20119) );
  INV_X1 U12906 ( .A(n11253), .ZN(n13073) );
  AND2_X1 U12907 ( .A1(n12514), .A2(n10251), .ZN(n12807) );
  INV_X1 U12908 ( .A(n14059), .ZN(n11277) );
  OR2_X1 U12909 ( .A1(n10705), .A2(n15192), .ZN(n15188) );
  OR2_X1 U12910 ( .A1(n10696), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15227) );
  OR2_X1 U12911 ( .A1(n10698), .A2(n15279), .ZN(n15078) );
  INV_X1 U12912 ( .A(n10485), .ZN(n19417) );
  AND2_X1 U12913 ( .A1(n17600), .A2(n16731), .ZN(n16590) );
  BUF_X1 U12914 ( .A(n15560), .Z(n17216) );
  AND3_X1 U12915 ( .A1(n16462), .A2(n16458), .A3(n17781), .ZN(n15754) );
  INV_X1 U12916 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18058) );
  NAND2_X1 U12917 ( .A1(n15618), .A2(n15650), .ZN(n16445) );
  AOI21_X1 U12918 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n18708), .A(
        n13027), .ZN(n13926) );
  OAI211_X1 U12919 ( .C1(n13024), .C2(n13023), .A(n13923), .B(n13022), .ZN(
        n15633) );
  INV_X1 U12920 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14265) );
  AND2_X1 U12921 ( .A1(n12132), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12133) );
  NOR2_X1 U12922 ( .A1(n12004), .A2(n15839), .ZN(n11986) );
  INV_X1 U12923 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19921) );
  INV_X1 U12924 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n21005) );
  AND2_X1 U12925 ( .A1(n15776), .A2(n13679), .ZN(n13688) );
  NAND2_X1 U12926 ( .A1(n13688), .A2(n13682), .ZN(n19977) );
  INV_X1 U12927 ( .A(n12441), .ZN(n12456) );
  AND2_X1 U12928 ( .A1(n13413), .A2(n13182), .ZN(n13318) );
  INV_X1 U12929 ( .A(n12184), .ZN(n12201) );
  NAND2_X1 U12930 ( .A1(n11986), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11970) );
  OR2_X1 U12931 ( .A1(n12063), .A2(n11950), .ZN(n12035) );
  NAND2_X1 U12932 ( .A1(n19904), .A2(n12281), .ZN(n14518) );
  AND2_X1 U12933 ( .A1(n12432), .A2(n12431), .ZN(n14325) );
  OR2_X1 U12934 ( .A1(n14641), .A2(n14642), .ZN(n15957) );
  AND2_X1 U12935 ( .A1(n13256), .A2(n13391), .ZN(n16024) );
  NOR2_X2 U12936 ( .A1(n15867), .A2(n15868), .ZN(n15866) );
  INV_X1 U12937 ( .A(n15975), .ZN(n20093) );
  NAND2_X1 U12938 ( .A1(n20160), .A2(n12355), .ZN(n11770) );
  NOR2_X1 U12939 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n11484) );
  NOR2_X2 U12940 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20613) );
  INV_X1 U12941 ( .A(n20173), .ZN(n20174) );
  OR2_X1 U12942 ( .A1(n13410), .A2(n13409), .ZN(n15737) );
  AND2_X1 U12943 ( .A1(n10922), .A2(n10756), .ZN(n10757) );
  AND4_X1 U12944 ( .A1(n11070), .A2(n10126), .A3(n11069), .A4(n11068), .ZN(
        n13582) );
  INV_X1 U12945 ( .A(n12807), .ZN(n12541) );
  AND2_X1 U12946 ( .A1(n13773), .A2(n13706), .ZN(n13774) );
  OR2_X1 U12947 ( .A1(n11017), .A2(n10258), .ZN(n11195) );
  OAI21_X1 U12948 ( .B1(n14132), .B2(n16262), .A(n14060), .ZN(n14061) );
  INV_X1 U12949 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16155) );
  INV_X1 U12950 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18975) );
  INV_X1 U12951 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10815) );
  AND2_X1 U12952 ( .A1(n15231), .A2(n11273), .ZN(n15203) );
  OR2_X1 U12953 ( .A1(n10647), .A2(n15308), .ZN(n16252) );
  AND2_X1 U12954 ( .A1(n10977), .A2(n19768), .ZN(n11259) );
  NAND2_X1 U12955 ( .A1(n11259), .A2(n11012), .ZN(n16299) );
  INV_X1 U12956 ( .A(n19316), .ZN(n19419) );
  INV_X1 U12957 ( .A(n19509), .ZN(n19511) );
  INV_X1 U12958 ( .A(n19850), .ZN(n19578) );
  NAND2_X1 U12959 ( .A1(n15394), .A2(n19852), .ZN(n19451) );
  NOR2_X1 U12960 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16865), .ZN(n16843) );
  INV_X1 U12961 ( .A(n18733), .ZN(n16926) );
  NOR2_X1 U12962 ( .A1(n17524), .A2(n10139), .ZN(n17525) );
  OR2_X1 U12963 ( .A1(n18001), .A2(n16440), .ZN(n17597) );
  AOI21_X1 U12964 ( .B1(n16389), .B2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n18607), .ZN(n17716) );
  NAND2_X1 U12965 ( .A1(n15677), .A2(n17787), .ZN(n18084) );
  INV_X1 U12966 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17844) );
  NAND2_X1 U12967 ( .A1(n17713), .A2(n17882), .ZN(n17602) );
  INV_X1 U12968 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16458) );
  NOR2_X1 U12969 ( .A1(n18206), .A2(n18692), .ZN(n18173) );
  OAI21_X1 U12970 ( .B1(n13028), .B2(n15633), .A(n13926), .ZN(n18660) );
  INV_X1 U12971 ( .A(n15621), .ZN(n15622) );
  INV_X1 U12972 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15608) );
  INV_X1 U12973 ( .A(n18849), .ZN(n18836) );
  INV_X1 U12974 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18699) );
  INV_X1 U12975 ( .A(n18875), .ZN(n18870) );
  NAND2_X1 U12976 ( .A1(n12133), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12156) );
  NOR2_X1 U12977 ( .A1(n14027), .A2(n15855), .ZN(n15844) );
  NOR2_X1 U12978 ( .A1(n14026), .A2(n19954), .ZN(n19923) );
  AND2_X1 U12979 ( .A1(n13688), .A2(n13684), .ZN(n19974) );
  AND2_X1 U12980 ( .A1(n15776), .A2(n13690), .ZN(n15861) );
  AND2_X1 U12981 ( .A1(n12450), .A2(n12449), .ZN(n14210) );
  INV_X1 U12982 ( .A(n19986), .ZN(n19995) );
  AND2_X1 U12983 ( .A1(n14378), .A2(n14377), .ZN(n15850) );
  NAND2_X1 U12984 ( .A1(n11935), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12063) );
  NOR2_X1 U12985 ( .A1(n11823), .A2(n13564), .ZN(n11860) );
  INV_X1 U12986 ( .A(n19904), .ZN(n20046) );
  INV_X1 U12987 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14094) );
  AND2_X1 U12988 ( .A1(n14569), .A2(n13996), .ZN(n14595) );
  AND2_X1 U12989 ( .A1(n15955), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14630) );
  NOR2_X1 U12990 ( .A1(n15957), .A2(n11756), .ZN(n15955) );
  OR2_X1 U12991 ( .A1(n20054), .A2(n16024), .ZN(n15975) );
  NAND2_X1 U12992 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n13232), .ZN(n20821) );
  OAI22_X1 U12993 ( .A1(n20126), .A2(n20125), .B1(n20471), .B2(n20296), .ZN(
        n20183) );
  OAI22_X1 U12994 ( .A1(n20225), .A2(n20224), .B1(n20223), .B2(n20471), .ZN(
        n20249) );
  OAI21_X1 U12995 ( .B1(n20265), .B2(n20263), .A(n20262), .ZN(n20291) );
  NAND2_X1 U12996 ( .A1(n20107), .A2(n20106), .ZN(n20257) );
  INV_X1 U12997 ( .A(n20348), .ZN(n20340) );
  INV_X1 U12998 ( .A(n20383), .ZN(n20371) );
  INV_X1 U12999 ( .A(n20415), .ZN(n20407) );
  AND2_X1 U13000 ( .A1(n13420), .A2(n13474), .ZN(n20389) );
  INV_X1 U13001 ( .A(n20459), .ZN(n20466) );
  INV_X1 U13002 ( .A(n20507), .ZN(n20503) );
  INV_X1 U13003 ( .A(n20546), .ZN(n20537) );
  INV_X1 U13004 ( .A(n20549), .ZN(n20604) );
  OAI21_X1 U13005 ( .B1(n20617), .B2(n20616), .A(n20684), .ZN(n20636) );
  INV_X1 U13006 ( .A(n20661), .ZN(n20670) );
  INV_X1 U13007 ( .A(n20737), .ZN(n20717) );
  AND2_X1 U13008 ( .A1(n20739), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15747) );
  INV_X1 U13009 ( .A(n16106), .ZN(n20838) );
  AND2_X1 U13010 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20800), .ZN(n20806) );
  NOR2_X1 U13011 ( .A1(n19032), .A2(n19771), .ZN(n19055) );
  INV_X1 U13012 ( .A(n19042), .ZN(n19060) );
  NOR2_X1 U13013 ( .A1(n9882), .A2(n19680), .ZN(n19003) );
  INV_X1 U13014 ( .A(n19063), .ZN(n18980) );
  INV_X1 U13015 ( .A(n15196), .ZN(n16217) );
  OR2_X1 U13016 ( .A1(n13583), .A2(n13582), .ZN(n13659) );
  INV_X1 U13017 ( .A(n14911), .ZN(n14894) );
  NOR2_X1 U13018 ( .A1(n13207), .A2(n13645), .ZN(n19077) );
  INV_X1 U13019 ( .A(n19110), .ZN(n19126) );
  INV_X1 U13020 ( .A(n19136), .ZN(n13130) );
  INV_X1 U13021 ( .A(n13101), .ZN(n13099) );
  NOR2_X1 U13023 ( .A1(n15232), .A2(n15233), .ZN(n15220) );
  INV_X1 U13024 ( .A(n15289), .ZN(n16307) );
  INV_X1 U13025 ( .A(n16299), .ZN(n19220) );
  INV_X1 U13026 ( .A(n19424), .ZN(n19683) );
  OAI21_X1 U13027 ( .B1(n19240), .B2(n19280), .A(n19683), .ZN(n19283) );
  NOR2_X1 U13028 ( .A1(n19291), .A2(n19289), .ZN(n19310) );
  INV_X1 U13029 ( .A(n19319), .ZN(n19341) );
  AND2_X1 U13030 ( .A1(n19448), .A2(n19850), .ZN(n19390) );
  AND2_X1 U13031 ( .A1(n13819), .A2(n13818), .ZN(n19389) );
  AND2_X1 U13032 ( .A1(n19448), .A2(n19644), .ZN(n19443) );
  NOR2_X1 U13033 ( .A1(n19451), .A2(n19419), .ZN(n19473) );
  OAI22_X1 U13034 ( .A1(n19487), .A2(n19486), .B1(n19485), .B2(n19484), .ZN(
        n19505) );
  INV_X1 U13035 ( .A(n19532), .ZN(n19535) );
  OAI21_X1 U13036 ( .B1(n19575), .B2(n19543), .A(n19542), .ZN(n19564) );
  NOR2_X2 U13037 ( .A1(n19651), .A2(n19578), .ZN(n19636) );
  NOR2_X1 U13038 ( .A1(n19864), .A2(n19852), .ZN(n19644) );
  NOR2_X1 U13039 ( .A1(n19477), .A2(n19451), .ZN(n19756) );
  AND3_X1 U13040 ( .A1(n10329), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n19768) );
  INV_X1 U13041 ( .A(n19787), .ZN(n19773) );
  INV_X1 U13042 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19792) );
  NAND2_X1 U13043 ( .A1(n18227), .A2(n17930), .ZN(n18664) );
  NOR2_X1 U13044 ( .A1(n16909), .A2(n16591), .ZN(n16622) );
  NOR2_X1 U13045 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16702), .ZN(n16686) );
  NOR2_X1 U13046 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16725), .ZN(n16708) );
  NOR2_X1 U13047 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16769), .ZN(n16750) );
  NOR2_X1 U13048 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16795), .ZN(n16774) );
  NOR2_X1 U13049 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16834), .ZN(n16823) );
  NOR2_X1 U13050 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16889), .ZN(n16870) );
  INV_X1 U13051 ( .A(n16920), .ZN(n16930) );
  NOR2_X2 U13052 ( .A1(n18718), .A2(n13034), .ZN(n16935) );
  NAND2_X1 U13053 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17115), .ZN(n17078) );
  INV_X1 U13054 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17158) );
  OAI221_X1 U13055 ( .B1(n15419), .B2(n15642), .C1(n15419), .C2(n18666), .A(
        n18868), .ZN(n15770) );
  NOR2_X1 U13056 ( .A1(n20931), .A2(n17325), .ZN(n17320) );
  INV_X1 U13057 ( .A(n17311), .ZN(n17336) );
  INV_X1 U13058 ( .A(n17348), .ZN(n17392) );
  NAND3_X1 U13059 ( .A1(n12933), .A2(n12932), .A3(n12931), .ZN(n18874) );
  NOR2_X1 U13060 ( .A1(n15692), .A2(n17565), .ZN(n17895) );
  INV_X1 U13061 ( .A(n17685), .ZN(n17613) );
  NAND2_X1 U13062 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17706), .ZN(
        n17945) );
  NAND2_X1 U13063 ( .A1(n18037), .A2(n18084), .ZN(n18063) );
  NAND2_X1 U13064 ( .A1(n15682), .A2(n15681), .ZN(n17761) );
  INV_X1 U13065 ( .A(n18260), .ZN(n18607) );
  INV_X1 U13066 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17875) );
  INV_X1 U13067 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17925) );
  INV_X1 U13068 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18001) );
  INV_X1 U13069 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18047) );
  NOR2_X2 U13070 ( .A1(n18205), .A2(n16446), .ZN(n18083) );
  INV_X1 U13071 ( .A(n18205), .ZN(n18184) );
  INV_X1 U13072 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18888) );
  NOR2_X1 U13073 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18824), .ZN(
        n18849) );
  NAND2_X1 U13074 ( .A1(n18331), .A2(n18470), .ZN(n18260) );
  INV_X1 U13075 ( .A(n18658), .ZN(n18303) );
  INV_X1 U13076 ( .A(n18284), .ZN(n18348) );
  INV_X1 U13077 ( .A(n18307), .ZN(n18370) );
  INV_X1 U13078 ( .A(n18398), .ZN(n18463) );
  INV_X1 U13079 ( .A(n18494), .ZN(n18536) );
  AND2_X1 U13080 ( .A1(n18222), .A2(n18467), .ZN(n18597) );
  AND2_X1 U13081 ( .A1(n18607), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18608) );
  AND2_X1 U13082 ( .A1(n18607), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18626) );
  OAI22_X1 U13083 ( .A1(n16437), .A2(n18661), .B1(n16380), .B2(n18664), .ZN(
        n18714) );
  NOR2_X1 U13084 ( .A1(n18888), .A2(n18729), .ZN(n18868) );
  INV_X1 U13085 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20643) );
  INV_X1 U13086 ( .A(n19960), .ZN(n19931) );
  INV_X1 U13087 ( .A(n19974), .ZN(n19945) );
  INV_X1 U13088 ( .A(n14100), .ZN(n14118) );
  INV_X1 U13089 ( .A(n15794), .ZN(n14422) );
  INV_X1 U13090 ( .A(n15850), .ZN(n14448) );
  AND2_X1 U13091 ( .A1(n13336), .A2(n13335), .ZN(n20168) );
  INV_X1 U13092 ( .A(n15883), .ZN(n20003) );
  NAND2_X1 U13093 ( .A1(n13331), .A2(n15742), .ZN(n13517) );
  INV_X2 U13094 ( .A(n20008), .ZN(n13553) );
  NOR2_X1 U13095 ( .A1(n19893), .A2(n13290), .ZN(n13356) );
  AOI21_X1 U13096 ( .B1(n14178), .B2(n20045), .A(n14098), .ZN(n14099) );
  OAI21_X1 U13097 ( .B1(n14388), .B2(n14008), .A(n14376), .ZN(n14039) );
  INV_X1 U13098 ( .A(n15919), .ZN(n20050) );
  NAND2_X1 U13099 ( .A1(n16016), .A2(n13986), .ZN(n16001) );
  INV_X1 U13100 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16059) );
  INV_X1 U13101 ( .A(n20076), .ZN(n20102) );
  INV_X1 U13102 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20611) );
  AOI211_X2 U13103 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20296), .A(n20419), 
        .B(n20113), .ZN(n20180) );
  OR2_X1 U13104 ( .A1(n20257), .A2(n20108), .ZN(n20213) );
  OR2_X1 U13105 ( .A1(n20257), .A2(n20215), .ZN(n20294) );
  OR2_X1 U13106 ( .A1(n20257), .A2(n20253), .ZN(n20311) );
  NAND2_X1 U13107 ( .A1(n20389), .A2(n20610), .ZN(n20383) );
  AOI22_X1 U13108 ( .A1(n20356), .A2(n20352), .B1(n20554), .B2(n20351), .ZN(
        n20388) );
  NAND2_X1 U13109 ( .A1(n20389), .A2(n20639), .ZN(n20415) );
  NAND2_X1 U13110 ( .A1(n20514), .A2(n20548), .ZN(n20459) );
  NAND2_X1 U13111 ( .A1(n20514), .A2(n20610), .ZN(n20507) );
  AOI22_X1 U13112 ( .A1(n20481), .A2(n20476), .B1(n20474), .B2(n20473), .ZN(
        n20512) );
  NAND2_X1 U13113 ( .A1(n20514), .A2(n20513), .ZN(n20549) );
  AOI22_X1 U13114 ( .A1(n20561), .A2(n20558), .B1(n20554), .B2(n20553), .ZN(
        n20609) );
  NAND2_X1 U13115 ( .A1(n20679), .A2(n20548), .ZN(n20630) );
  NAND2_X1 U13116 ( .A1(n20679), .A2(n20610), .ZN(n20661) );
  INV_X2 U13117 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20742) );
  INV_X1 U13118 ( .A(n20818), .ZN(n20814) );
  INV_X1 U13119 ( .A(n20805), .ZN(n20798) );
  INV_X1 U13120 ( .A(n20806), .ZN(n20803) );
  OR2_X1 U13121 ( .A1(n13072), .A2(n13040), .ZN(n13046) );
  INV_X1 U13122 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19420) );
  NAND2_X1 U13123 ( .A1(n18895), .A2(n14139), .ZN(n19042) );
  INV_X1 U13124 ( .A(n19066), .ZN(n19036) );
  INV_X1 U13125 ( .A(n14901), .ZN(n14909) );
  INV_X1 U13126 ( .A(n19127), .ZN(n19084) );
  NAND2_X1 U13127 ( .A1(n19169), .A2(n19140), .ZN(n19167) );
  INV_X1 U13128 ( .A(n19169), .ZN(n19201) );
  INV_X1 U13129 ( .A(n13047), .ZN(n13101) );
  NAND2_X1 U13130 ( .A1(n11306), .A2(n11305), .ZN(n11307) );
  INV_X1 U13131 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16271) );
  INV_X1 U13132 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16282) );
  INV_X1 U13133 ( .A(n19203), .ZN(n16262) );
  INV_X1 U13134 ( .A(n12483), .ZN(n12484) );
  AOI21_X1 U13135 ( .B1(n12506), .B2(n19233), .A(n12505), .ZN(n12507) );
  INV_X1 U13136 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19235) );
  INV_X1 U13137 ( .A(n16294), .ZN(n15321) );
  INV_X1 U13138 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15769) );
  NAND2_X1 U13139 ( .A1(n19509), .A2(n19316), .ZN(n19311) );
  NAND2_X1 U13140 ( .A1(n19316), .A2(n19850), .ZN(n19368) );
  INV_X1 U13141 ( .A(n19390), .ZN(n19387) );
  INV_X1 U13142 ( .A(n19443), .ZN(n19440) );
  INV_X1 U13143 ( .A(n19473), .ZN(n19470) );
  INV_X1 U13144 ( .A(n19504), .ZN(n19502) );
  NAND2_X1 U13145 ( .A1(n19607), .A2(n19509), .ZN(n19532) );
  INV_X1 U13146 ( .A(n19727), .ZN(n19588) );
  INV_X1 U13147 ( .A(n19698), .ZN(n19623) );
  INV_X1 U13148 ( .A(n19677), .ZN(n19655) );
  NAND2_X1 U13149 ( .A1(n19607), .A2(n19644), .ZN(n19667) );
  INV_X1 U13150 ( .A(n19713), .ZN(n19709) );
  INV_X1 U13151 ( .A(n19757), .ZN(n19724) );
  INV_X1 U13152 ( .A(n19595), .ZN(n19750) );
  INV_X1 U13153 ( .A(n19849), .ZN(n19772) );
  INV_X1 U13154 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18873) );
  INV_X1 U13155 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17062) );
  INV_X1 U13156 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n16868) );
  NAND2_X1 U13157 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n16945), .ZN(n16920) );
  NOR2_X1 U13158 ( .A1(n17158), .A2(n17186), .ZN(n17172) );
  NOR2_X1 U13159 ( .A1(n16868), .A2(n17231), .ZN(n17234) );
  AND2_X1 U13160 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n17249), .ZN(n17246) );
  INV_X1 U13161 ( .A(n16436), .ZN(n17374) );
  NOR2_X1 U13162 ( .A1(n15526), .A2(n15525), .ZN(n17381) );
  INV_X1 U13163 ( .A(n17433), .ZN(n17460) );
  INV_X1 U13164 ( .A(n17512), .ZN(n17507) );
  AOI21_X1 U13165 ( .B1(n17529), .B2(n17528), .A(n17527), .ZN(n17534) );
  INV_X1 U13166 ( .A(n17711), .ZN(n17789) );
  INV_X1 U13167 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17726) );
  NAND2_X1 U13168 ( .A1(n17832), .A2(n16436), .ZN(n17794) );
  INV_X1 U13169 ( .A(n17832), .ZN(n17885) );
  AOI21_X1 U13170 ( .B1(n16461), .B2(n16460), .A(n16459), .ZN(n16464) );
  INV_X1 U13171 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17987) );
  OAI21_X2 U13172 ( .B1(n15640), .B2(n15639), .A(n18868), .ZN(n18205) );
  INV_X1 U13173 ( .A(n18083), .ZN(n18121) );
  INV_X1 U13174 ( .A(n18204), .ZN(n18165) );
  NAND2_X1 U13175 ( .A1(n18662), .A2(n18184), .ZN(n18199) );
  INV_X1 U13176 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18226) );
  INV_X1 U13177 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18245) );
  INV_X1 U13178 ( .A(n18394), .ZN(n18377) );
  INV_X1 U13179 ( .A(n18417), .ZN(n18376) );
  INV_X1 U13180 ( .A(n18567), .ZN(n18611) );
  INV_X1 U13181 ( .A(n18582), .ZN(n18635) );
  INV_X1 U13182 ( .A(n18868), .ZN(n18724) );
  INV_X1 U13183 ( .A(n18821), .ZN(n18737) );
  INV_X1 U13184 ( .A(n18818), .ZN(n18821) );
  INV_X1 U13185 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18764) );
  NOR2_X1 U13186 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12915), .ZN(n16546)
         );
  INV_X1 U13187 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19798) );
  NAND2_X1 U13188 ( .A1(n12466), .A2(n12465), .ZN(P1_U2842) );
  NAND2_X1 U13189 ( .A1(n12508), .A2(n12507), .ZN(P2_U3026) );
  AND2_X4 U13190 ( .A1(n15384), .A2(n10144), .ZN(n12862) );
  AOI22_X1 U13191 ( .A1(n9749), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12862), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10148) );
  AOI22_X1 U13192 ( .A1(n12720), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12853), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10146) );
  AOI22_X1 U13193 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12861), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10145) );
  NAND4_X1 U13194 ( .A1(n10148), .A2(n10147), .A3(n10146), .A4(n10145), .ZN(
        n10149) );
  NAND2_X1 U13195 ( .A1(n10149), .A2(n15408), .ZN(n10157) );
  AOI22_X1 U13196 ( .A1(n12720), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12853), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10154) );
  AOI22_X1 U13197 ( .A1(n9751), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10243), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10153) );
  AOI21_X1 U13198 ( .B1(n9748), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A(
        n10150), .ZN(n10152) );
  AOI22_X1 U13199 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12861), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10151) );
  NAND4_X1 U13200 ( .A1(n10154), .A2(n10153), .A3(n10152), .A4(n10151), .ZN(
        n10155) );
  NAND2_X1 U13201 ( .A1(n10155), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10156) );
  AOI22_X1 U13202 ( .A1(n9795), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12853), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10162) );
  AOI22_X1 U13203 ( .A1(n9751), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10243), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10161) );
  AOI22_X1 U13204 ( .A1(n9749), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12862), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10160) );
  AOI22_X1 U13205 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12861), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10159) );
  NAND4_X1 U13206 ( .A1(n10162), .A2(n10161), .A3(n10160), .A4(n10159), .ZN(
        n10163) );
  NAND2_X1 U13207 ( .A1(n10163), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10170) );
  AOI22_X1 U13208 ( .A1(n12720), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12853), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10166) );
  AOI22_X1 U13209 ( .A1(n9748), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12862), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10165) );
  AOI22_X1 U13210 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12861), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10164) );
  NAND4_X1 U13211 ( .A1(n10167), .A2(n10166), .A3(n10165), .A4(n10164), .ZN(
        n10168) );
  NAND2_X1 U13212 ( .A1(n10168), .A2(n15408), .ZN(n10169) );
  AOI22_X1 U13213 ( .A1(n9753), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10243), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10175) );
  AOI22_X1 U13214 ( .A1(n9750), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n12862), .ZN(n10174) );
  AOI22_X1 U13215 ( .A1(n12720), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12838), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10173) );
  AOI22_X1 U13216 ( .A1(n12853), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12861), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10172) );
  NAND4_X1 U13217 ( .A1(n10175), .A2(n10174), .A3(n10173), .A4(n10172), .ZN(
        n10176) );
  NAND2_X1 U13218 ( .A1(n10176), .A2(n15408), .ZN(n10184) );
  AOI22_X1 U13219 ( .A1(n9752), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9750), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10177) );
  INV_X1 U13220 ( .A(n10177), .ZN(n10182) );
  AOI22_X1 U13221 ( .A1(n12720), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12838), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10180) );
  AOI22_X1 U13222 ( .A1(n10243), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12862), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10179) );
  AOI22_X1 U13223 ( .A1(n12853), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12861), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10178) );
  NAND3_X1 U13224 ( .A1(n10179), .A2(n10180), .A3(n10178), .ZN(n10181) );
  AOI22_X1 U13225 ( .A1(n12720), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12853), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10189) );
  AOI22_X1 U13226 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12861), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10188) );
  AOI21_X1 U13227 ( .B1(n9749), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A(
        n10186), .ZN(n10187) );
  NAND3_X1 U13228 ( .A1(n10189), .A2(n10188), .A3(n10187), .ZN(n10192) );
  AOI22_X1 U13229 ( .A1(n9752), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10243), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10190) );
  AOI22_X1 U13230 ( .A1(n9753), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10243), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10196) );
  AOI22_X1 U13231 ( .A1(n9749), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12862), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10195) );
  AOI22_X1 U13232 ( .A1(n12720), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12853), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10194) );
  AOI22_X1 U13233 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12861), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10193) );
  NAND4_X1 U13234 ( .A1(n10196), .A2(n10195), .A3(n10194), .A4(n10193), .ZN(
        n10197) );
  NAND2_X1 U13235 ( .A1(n10197), .A2(n15408), .ZN(n10198) );
  AOI22_X1 U13236 ( .A1(n9750), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12862), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10203) );
  AOI22_X1 U13237 ( .A1(n9753), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10243), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10202) );
  AOI22_X1 U13238 ( .A1(n12720), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12838), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10201) );
  AOI22_X1 U13239 ( .A1(n12853), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12861), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10200) );
  NAND4_X1 U13240 ( .A1(n10203), .A2(n10202), .A3(n10201), .A4(n10200), .ZN(
        n10204) );
  AOI22_X1 U13241 ( .A1(n12720), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12853), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10209) );
  AOI22_X1 U13242 ( .A1(n9751), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10243), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10208) );
  AOI22_X1 U13243 ( .A1(n9752), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(n9748), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10215) );
  AOI22_X1 U13244 ( .A1(n10243), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12862), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10214) );
  AOI22_X1 U13245 ( .A1(n9795), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12838), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10213) );
  AOI22_X1 U13246 ( .A1(n12853), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12861), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10212) );
  NAND4_X1 U13247 ( .A1(n10215), .A2(n10214), .A3(n10213), .A4(n10212), .ZN(
        n10216) );
  NAND2_X1 U13248 ( .A1(n10216), .A2(n15408), .ZN(n10223) );
  AOI22_X1 U13249 ( .A1(n9750), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12862), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10220) );
  AOI22_X1 U13250 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12861), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10218) );
  AOI22_X1 U13251 ( .A1(n9795), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12853), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10217) );
  NAND4_X1 U13252 ( .A1(n10220), .A2(n10219), .A3(n10218), .A4(n10217), .ZN(
        n10221) );
  NAND2_X1 U13253 ( .A1(n10221), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10222) );
  AOI22_X1 U13254 ( .A1(n9795), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12838), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10225) );
  NAND2_X1 U13255 ( .A1(n10225), .A2(n10224), .ZN(n10229) );
  AOI22_X1 U13256 ( .A1(n9751), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(n9748), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10227) );
  AOI22_X1 U13257 ( .A1(n12853), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12861), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10226) );
  NAND2_X1 U13258 ( .A1(n10227), .A2(n10226), .ZN(n10228) );
  AOI22_X1 U13259 ( .A1(n9751), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10243), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10233) );
  AOI22_X1 U13260 ( .A1(n9748), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12862), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10232) );
  AOI22_X1 U13261 ( .A1(n9795), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12838), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10231) );
  AOI22_X1 U13262 ( .A1(n12853), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12861), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10230) );
  NAND4_X1 U13263 ( .A1(n10233), .A2(n10232), .A3(n10231), .A4(n10230), .ZN(
        n10234) );
  AOI22_X1 U13264 ( .A1(n12720), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12853), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10239) );
  AOI22_X1 U13265 ( .A1(n9748), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12862), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10238) );
  AOI22_X1 U13266 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12861), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10237) );
  NAND4_X1 U13267 ( .A1(n10240), .A2(n10239), .A3(n10238), .A4(n10237), .ZN(
        n10241) );
  NAND2_X1 U13268 ( .A1(n10241), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10250) );
  AOI22_X1 U13269 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12861), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10242) );
  INV_X1 U13270 ( .A(n10242), .ZN(n10248) );
  AOI22_X1 U13271 ( .A1(n12720), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12853), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10246) );
  AOI22_X1 U13272 ( .A1(n9750), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12862), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10244) );
  NAND3_X1 U13273 ( .A1(n10246), .A2(n10245), .A3(n10244), .ZN(n10247) );
  AND2_X1 U13274 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n10278) );
  NAND2_X2 U13275 ( .A1(n10251), .A2(n10539), .ZN(n10281) );
  NAND2_X1 U13276 ( .A1(n10281), .A2(n10265), .ZN(n10961) );
  NAND2_X1 U13277 ( .A1(n10988), .A2(n10268), .ZN(n10256) );
  NAND2_X1 U13278 ( .A1(n10256), .A2(n10255), .ZN(n10301) );
  NAND2_X1 U13279 ( .A1(n10301), .A2(n10257), .ZN(n10276) );
  NAND3_X1 U13280 ( .A1(n10254), .A2(n11013), .A3(n10281), .ZN(n10300) );
  MUX2_X1 U13281 ( .A(n12509), .B(n9755), .S(n10265), .Z(n10264) );
  OR2_X1 U13282 ( .A1(n10266), .A2(n10258), .ZN(n10259) );
  NAND2_X1 U13283 ( .A1(n10259), .A2(n10282), .ZN(n10260) );
  NAND2_X1 U13284 ( .A1(n10260), .A2(n10281), .ZN(n10263) );
  NAND3_X1 U13285 ( .A1(n10282), .A2(n19259), .A3(n10261), .ZN(n10293) );
  NAND2_X1 U13286 ( .A1(n10293), .A2(n10266), .ZN(n10262) );
  NAND4_X1 U13287 ( .A1(n10262), .A2(n14666), .A3(n10263), .A4(n10264), .ZN(
        n10991) );
  INV_X1 U13289 ( .A(n10270), .ZN(n10271) );
  NAND2_X1 U13290 ( .A1(n10273), .A2(n10271), .ZN(n10772) );
  NOR2_X1 U13291 ( .A1(n10279), .A2(n10266), .ZN(n10272) );
  NAND2_X1 U13292 ( .A1(n10772), .A2(n10272), .ZN(n10275) );
  NAND2_X1 U13293 ( .A1(n10276), .A2(n10302), .ZN(n10311) );
  NOR2_X1 U13294 ( .A1(n10283), .A2(n10274), .ZN(n10284) );
  NAND2_X1 U13295 ( .A1(n10284), .A2(n10282), .ZN(n10285) );
  NAND2_X1 U13296 ( .A1(n10286), .A2(n10285), .ZN(n10287) );
  INV_X1 U13297 ( .A(n10297), .ZN(n10290) );
  NAND2_X1 U13298 ( .A1(n18894), .A2(n10329), .ZN(n16363) );
  NOR2_X1 U13299 ( .A1(n16363), .A2(n19886), .ZN(n10289) );
  AOI21_X1 U13300 ( .B1(n10290), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10289), 
        .ZN(n10291) );
  NAND2_X1 U13301 ( .A1(n10292), .A2(n10291), .ZN(n10336) );
  NAND2_X1 U13302 ( .A1(n13039), .A2(n9788), .ZN(n16362) );
  NAND3_X1 U13303 ( .A1(n14666), .A2(n10266), .A3(n12509), .ZN(n10294) );
  INV_X1 U13304 ( .A(n10926), .ZN(n10295) );
  NOR2_X1 U13305 ( .A1(n12882), .A2(n10251), .ZN(n10296) );
  NAND2_X1 U13306 ( .A1(n10993), .A2(n10296), .ZN(n10313) );
  NAND2_X1 U13307 ( .A1(n10301), .A2(n10300), .ZN(n10987) );
  NAND2_X1 U13308 ( .A1(n10987), .A2(n10302), .ZN(n10303) );
  NAND2_X1 U13309 ( .A1(n10303), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10310) );
  INV_X1 U13310 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n10538) );
  NOR2_X1 U13311 ( .A1(n10279), .A2(n18894), .ZN(n10304) );
  NAND2_X1 U13312 ( .A1(n10826), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10307) );
  NAND2_X1 U13313 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10305) );
  AND2_X1 U13314 ( .A1(n16363), .A2(n10305), .ZN(n10306) );
  OAI211_X1 U13315 ( .C1(n10905), .C2(n10538), .A(n10307), .B(n10306), .ZN(
        n10308) );
  INV_X1 U13316 ( .A(n10308), .ZN(n10309) );
  AND2_X2 U13317 ( .A1(n10336), .A2(n10338), .ZN(n10337) );
  NOR2_X1 U13318 ( .A1(n16363), .A2(n19877), .ZN(n10314) );
  INV_X1 U13319 ( .A(n10345), .ZN(n10321) );
  INV_X1 U13320 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n10540) );
  NAND2_X1 U13321 ( .A1(n10826), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n10317) );
  NAND2_X1 U13322 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10316) );
  OAI211_X1 U13323 ( .C1(n10905), .C2(n10540), .A(n10317), .B(n10316), .ZN(
        n10318) );
  INV_X1 U13324 ( .A(n10318), .ZN(n10319) );
  INV_X1 U13325 ( .A(n10346), .ZN(n10320) );
  NAND2_X1 U13326 ( .A1(n10321), .A2(n10320), .ZN(n10323) );
  AOI21_X2 U13327 ( .B1(n10337), .B2(n10323), .A(n10322), .ZN(n10341) );
  INV_X1 U13328 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n10325) );
  INV_X1 U13329 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10324) );
  NAND2_X1 U13330 ( .A1(n10826), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10327) );
  AOI21_X1 U13331 ( .B1(n18894), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10330) );
  AOI22_X1 U13332 ( .A1(n9762), .A2(P2_EBX_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10335) );
  NAND2_X1 U13333 ( .A1(n9782), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n10334) );
  XNOR2_X2 U13334 ( .A(n10818), .B(n10817), .ZN(n10357) );
  NAND2_X1 U13335 ( .A1(n10357), .A2(n14126), .ZN(n10371) );
  INV_X1 U13336 ( .A(n10371), .ZN(n10344) );
  NAND2_X4 U13337 ( .A1(n10343), .A2(n10342), .ZN(n13265) );
  NAND2_X1 U13338 ( .A1(n10344), .A2(n10353), .ZN(n10375) );
  INV_X1 U13339 ( .A(n10346), .ZN(n10347) );
  XNOR2_X2 U13340 ( .A(n10345), .B(n10347), .ZN(n10352) );
  INV_X1 U13342 ( .A(n10357), .ZN(n10351) );
  NAND2_X1 U13343 ( .A1(n10351), .A2(n14126), .ZN(n10369) );
  NAND2_X1 U13344 ( .A1(n13265), .A2(n9791), .ZN(n10370) );
  INV_X1 U13345 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12543) );
  INV_X1 U13346 ( .A(n10352), .ZN(n10349) );
  INV_X1 U13347 ( .A(n10359), .ZN(n10350) );
  NOR2_X1 U13348 ( .A1(n13265), .A2(n10350), .ZN(n10358) );
  INV_X1 U13349 ( .A(n10357), .ZN(n13626) );
  NAND2_X1 U13350 ( .A1(n13216), .A2(n10352), .ZN(n10360) );
  INV_X1 U13351 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n19723) );
  NAND2_X1 U13352 ( .A1(n10476), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10354) );
  OAI211_X1 U13353 ( .C1(n10484), .C2(n12543), .A(n10355), .B(n10354), .ZN(
        n10356) );
  BUF_X2 U13354 ( .A(n10357), .Z(n13617) );
  AOI22_X1 U13355 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19287), .B1(
        n13718), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10367) );
  NOR2_X1 U13356 ( .A1(n13265), .A2(n10360), .ZN(n10362) );
  AOI22_X1 U13357 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19573), .B1(
        n19640), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10366) );
  AOI22_X1 U13358 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19348), .B1(
        n10478), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10365) );
  NAND2_X1 U13359 ( .A1(n13265), .A2(n13313), .ZN(n10368) );
  OR2_X2 U13360 ( .A1(n10369), .A2(n10368), .ZN(n19608) );
  INV_X1 U13361 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12726) );
  INV_X1 U13362 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10372) );
  OAI22_X1 U13363 ( .A1(n19608), .A2(n12726), .B1(n10372), .B2(n10485), .ZN(
        n10373) );
  AOI21_X1 U13364 ( .B1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n10491), .A(
        n10373), .ZN(n10377) );
  OR2_X1 U13365 ( .A1(n13265), .A2(n9791), .ZN(n10374) );
  NOR2_X2 U13366 ( .A1(n10375), .A2(n9792), .ZN(n19242) );
  AOI22_X1 U13367 ( .A1(n19483), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n19242), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10376) );
  NAND3_X1 U13368 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10761) );
  NOR2_X1 U13369 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n10761), .ZN(
        n11099) );
  AOI22_X1 U13370 ( .A1(n10467), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11099), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10384) );
  INV_X1 U13371 ( .A(n10761), .ZN(n10380) );
  INV_X1 U13372 ( .A(n12699), .ZN(n11141) );
  AOI22_X1 U13373 ( .A1(n10456), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11141), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10383) );
  INV_X1 U13374 ( .A(n12689), .ZN(n11067) );
  AOI22_X1 U13375 ( .A1(n11067), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12706), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10382) );
  AND2_X1 U13376 ( .A1(n12862), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10462) );
  AOI22_X1 U13377 ( .A1(n12695), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10462), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10381) );
  NAND4_X1 U13378 ( .A1(n10384), .A2(n10383), .A3(n10382), .A4(n10381), .ZN(
        n10394) );
  AND2_X1 U13379 ( .A1(n10385), .A2(n12672), .ZN(n10500) );
  NOR2_X1 U13380 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10386) );
  AND2_X1 U13381 ( .A1(n12672), .A2(n10386), .ZN(n10414) );
  AOI22_X1 U13382 ( .A1(n10500), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10392) );
  AND2_X1 U13383 ( .A1(n10387), .A2(n12672), .ZN(n10413) );
  AND2_X1 U13384 ( .A1(n12672), .A2(n10388), .ZN(n10400) );
  AOI22_X1 U13385 ( .A1(n10413), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10400), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10391) );
  AOI22_X1 U13386 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10395), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10390) );
  AOI22_X1 U13387 ( .A1(n10401), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12690), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10389) );
  NAND4_X1 U13388 ( .A1(n10392), .A2(n10391), .A3(n10390), .A4(n10389), .ZN(
        n10393) );
  AOI22_X1 U13389 ( .A1(n11067), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n11141), .ZN(n10399) );
  AOI22_X1 U13390 ( .A1(n12695), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12696), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10398) );
  AOI22_X1 U13391 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10395), .B1(
        n10467), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10397) );
  AOI22_X1 U13392 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12706), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10396) );
  NAND4_X1 U13393 ( .A1(n10399), .A2(n10398), .A3(n10397), .A4(n10396), .ZN(
        n10407) );
  AOI22_X1 U13394 ( .A1(n10500), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10400), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10405) );
  AOI22_X1 U13395 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10413), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10404) );
  AOI22_X1 U13396 ( .A1(n10456), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12690), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10403) );
  AOI22_X1 U13397 ( .A1(n10401), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n10462), .ZN(n10402) );
  NAND4_X1 U13398 ( .A1(n10405), .A2(n10404), .A3(n10403), .A4(n10402), .ZN(
        n10406) );
  NOR2_X1 U13399 ( .A1(n10407), .A2(n10406), .ZN(n11024) );
  NOR2_X1 U13400 ( .A1(n13221), .A2(n11024), .ZN(n10408) );
  NAND2_X1 U13401 ( .A1(n9788), .A2(n10408), .ZN(n10779) );
  NAND2_X1 U13402 ( .A1(n10456), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n10412) );
  AOI22_X1 U13403 ( .A1(n10462), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10400), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10411) );
  NAND2_X1 U13404 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n10410) );
  NAND2_X1 U13405 ( .A1(n12706), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n10409) );
  AND4_X1 U13406 ( .A1(n10412), .A2(n10411), .A3(n10410), .A4(n10409), .ZN(
        n10424) );
  AOI22_X1 U13407 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10500), .B1(
        n10413), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10420) );
  NAND2_X1 U13408 ( .A1(n10395), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n10419) );
  NAND2_X1 U13409 ( .A1(n10401), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n10418) );
  INV_X1 U13410 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12521) );
  NAND2_X1 U13411 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n11099), .ZN(
        n10415) );
  OAI21_X1 U13412 ( .B1(n12699), .B2(n12521), .A(n10415), .ZN(n10416) );
  AOI21_X1 U13413 ( .B1(n10414), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n10416), .ZN(n10417) );
  AND4_X1 U13414 ( .A1(n10420), .A2(n10419), .A3(n10418), .A4(n10417), .ZN(
        n10423) );
  AOI22_X1 U13415 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10467), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10422) );
  AOI22_X1 U13416 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n11067), .B1(
        n12695), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10421) );
  NAND4_X1 U13417 ( .A1(n10424), .A2(n10423), .A3(n10422), .A4(n10421), .ZN(
        n10542) );
  INV_X1 U13418 ( .A(n10542), .ZN(n11034) );
  NAND2_X1 U13419 ( .A1(n10779), .A2(n11034), .ZN(n10425) );
  AOI22_X1 U13420 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19573), .B1(
        n19640), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10429) );
  AOI22_X1 U13421 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19348), .B1(
        n10476), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10428) );
  AOI22_X1 U13422 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19287), .B1(
        n10477), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10427) );
  AOI22_X1 U13423 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n13718), .B1(
        n10478), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10426) );
  AOI22_X1 U13424 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19483), .B1(
        n10491), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10434) );
  AOI22_X1 U13425 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19242), .B1(
        n10490), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10433) );
  INV_X1 U13426 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12774) );
  INV_X1 U13427 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12600) );
  INV_X1 U13428 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12767) );
  NOR2_X1 U13429 ( .A1(n10431), .A2(n10430), .ZN(n10432) );
  INV_X1 U13430 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10436) );
  OAI22_X1 U13431 ( .A1(n12689), .A2(n10436), .B1(n12654), .B2(n12774), .ZN(
        n10440) );
  INV_X1 U13432 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11114) );
  NAND2_X1 U13433 ( .A1(n10462), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n10438) );
  NAND2_X1 U13434 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n10437) );
  OAI211_X1 U13435 ( .C1(n15402), .C2(n11114), .A(n10438), .B(n10437), .ZN(
        n10439) );
  NOR2_X1 U13436 ( .A1(n10440), .A2(n10439), .ZN(n10451) );
  AOI22_X1 U13437 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10500), .B1(
        n10413), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10447) );
  NAND2_X1 U13438 ( .A1(n10467), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10446) );
  NAND2_X1 U13439 ( .A1(n10401), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n10445) );
  INV_X1 U13440 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10442) );
  NAND2_X1 U13441 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n12696), .ZN(
        n10441) );
  OAI21_X1 U13442 ( .B1(n12699), .B2(n10442), .A(n10441), .ZN(n10443) );
  AOI21_X1 U13443 ( .B1(n10414), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n10443), .ZN(n10444) );
  AND4_X1 U13444 ( .A1(n10447), .A2(n10446), .A3(n10445), .A4(n10444), .ZN(
        n10450) );
  AOI22_X1 U13445 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12695), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10449) );
  AOI22_X1 U13446 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n10456), .B1(
        n10395), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10448) );
  NAND4_X1 U13447 ( .A1(n10451), .A2(n10450), .A3(n10449), .A4(n10448), .ZN(
        n11039) );
  INV_X1 U13448 ( .A(n11039), .ZN(n10452) );
  NAND2_X1 U13449 ( .A1(n10452), .A2(n9788), .ZN(n10453) );
  OR2_X1 U13450 ( .A1(n11202), .A2(n20888), .ZN(n10460) );
  NAND2_X1 U13451 ( .A1(n10395), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10459) );
  NAND2_X1 U13452 ( .A1(n10456), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10458) );
  NAND2_X1 U13453 ( .A1(n10401), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10457) );
  INV_X1 U13454 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10461) );
  INV_X1 U13455 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12794) );
  OAI22_X1 U13456 ( .A1(n12689), .A2(n10461), .B1(n12654), .B2(n12794), .ZN(
        n10466) );
  INV_X1 U13457 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11132) );
  NAND2_X1 U13458 ( .A1(n10462), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10464) );
  NAND2_X1 U13459 ( .A1(n10413), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10463) );
  OAI211_X1 U13460 ( .C1(n15402), .C2(n11132), .A(n10464), .B(n10463), .ZN(
        n10465) );
  NOR2_X1 U13461 ( .A1(n10466), .A2(n10465), .ZN(n10474) );
  NAND2_X1 U13462 ( .A1(n10467), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10473) );
  NAND2_X1 U13463 ( .A1(n12695), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10472) );
  AOI22_X1 U13464 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10414), .B1(
        n10400), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10471) );
  INV_X1 U13465 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12540) );
  NAND2_X1 U13466 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n12696), .ZN(
        n10468) );
  OAI21_X1 U13467 ( .B1(n12699), .B2(n12540), .A(n10468), .ZN(n10469) );
  AOI21_X1 U13468 ( .B1(n10500), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n10469), .ZN(n10470) );
  AOI22_X1 U13469 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19348), .B1(
        n13718), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10482) );
  AOI22_X1 U13470 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19640), .B1(
        n10476), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10481) );
  INV_X1 U13471 ( .A(n10477), .ZN(n19514) );
  AOI22_X1 U13472 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19287), .B1(
        n10477), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10480) );
  AOI22_X1 U13473 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n10478), .B1(
        n19573), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10479) );
  AND4_X1 U13474 ( .A1(n10482), .A2(n10481), .A3(n10480), .A4(n10479), .ZN(
        n10488) );
  AOI22_X1 U13475 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n10483), .B1(
        n19687), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10487) );
  INV_X1 U13476 ( .A(n19608), .ZN(n10590) );
  AOI22_X1 U13477 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19417), .B1(
        n10590), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10486) );
  INV_X1 U13478 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12542) );
  INV_X1 U13479 ( .A(n19242), .ZN(n10595) );
  INV_X1 U13480 ( .A(n19483), .ZN(n10594) );
  INV_X1 U13481 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11161) );
  OAI22_X1 U13482 ( .A1(n12542), .A2(n10595), .B1(n10594), .B2(n11161), .ZN(
        n10489) );
  INV_X1 U13483 ( .A(n10489), .ZN(n10494) );
  INV_X1 U13484 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12643) );
  INV_X1 U13485 ( .A(n10490), .ZN(n10597) );
  INV_X1 U13486 ( .A(n10491), .ZN(n10596) );
  INV_X1 U13487 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12639) );
  OAI22_X1 U13488 ( .A1(n12643), .A2(n10597), .B1(n10596), .B2(n12639), .ZN(
        n10492) );
  INV_X1 U13489 ( .A(n10492), .ZN(n10493) );
  NAND3_X1 U13490 ( .A1(n10141), .A2(n10494), .A3(n10493), .ZN(n10512) );
  INV_X1 U13491 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10495) );
  INV_X1 U13492 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12821) );
  OAI22_X1 U13493 ( .A1(n12689), .A2(n10495), .B1(n12654), .B2(n12821), .ZN(
        n10499) );
  NAND2_X1 U13494 ( .A1(n10462), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10497) );
  NAND2_X1 U13495 ( .A1(n10413), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n10496) );
  OAI211_X1 U13496 ( .C1(n11161), .C2(n15402), .A(n10497), .B(n10496), .ZN(
        n10498) );
  NOR2_X1 U13497 ( .A1(n10499), .A2(n10498), .ZN(n10510) );
  NAND2_X1 U13498 ( .A1(n10467), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10506) );
  NAND2_X1 U13499 ( .A1(n12695), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n10505) );
  AOI22_X1 U13500 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10504) );
  NAND2_X1 U13501 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n12696), .ZN(
        n10501) );
  OAI21_X1 U13502 ( .B1(n12699), .B2(n12542), .A(n10501), .ZN(n10502) );
  AOI21_X1 U13503 ( .B1(n10500), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n10502), .ZN(n10503) );
  AND4_X1 U13504 ( .A1(n10506), .A2(n10505), .A3(n10504), .A4(n10503), .ZN(
        n10509) );
  AOI22_X1 U13505 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10395), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10508) );
  AOI22_X1 U13506 ( .A1(n10456), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10401), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10507) );
  NAND4_X1 U13507 ( .A1(n10510), .A2(n10509), .A3(n10508), .A4(n10507), .ZN(
        n11048) );
  OR2_X1 U13508 ( .A1(n9790), .A2(n11048), .ZN(n10511) );
  INV_X1 U13509 ( .A(n10515), .ZN(n10516) );
  NAND2_X1 U13510 ( .A1(n10514), .A2(n10516), .ZN(n10517) );
  INV_X1 U13511 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10518) );
  AOI22_X1 U13512 ( .A1(n10462), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10413), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10521) );
  NAND2_X1 U13513 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10520) );
  NAND2_X1 U13514 ( .A1(n10456), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10519) );
  NAND2_X1 U13515 ( .A1(n12695), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10526) );
  NAND2_X1 U13516 ( .A1(n10401), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10525) );
  NAND2_X1 U13517 ( .A1(n10395), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10524) );
  NAND2_X1 U13518 ( .A1(n12706), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10523) );
  INV_X1 U13519 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10533) );
  NAND2_X1 U13520 ( .A1(n10500), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10530) );
  NAND2_X1 U13521 ( .A1(n10414), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10529) );
  NAND2_X1 U13522 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10528) );
  AOI22_X1 U13523 ( .A1(n11141), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n12696), .ZN(n10527) );
  NAND2_X1 U13524 ( .A1(n10467), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10531) );
  OAI211_X1 U13525 ( .C1(n11202), .C2(n10533), .A(n10532), .B(n10531), .ZN(
        n10534) );
  INV_X1 U13526 ( .A(n10534), .ZN(n10535) );
  OR2_X1 U13527 ( .A1(n11024), .A2(n19265), .ZN(n10541) );
  NAND2_X1 U13528 ( .A1(n19265), .A2(n10538), .ZN(n10566) );
  NOR2_X1 U13529 ( .A1(n10742), .A2(n10540), .ZN(n10569) );
  AOI21_X1 U13530 ( .B1(n10541), .B2(n10566), .A(n10569), .ZN(n10571) );
  NAND2_X1 U13531 ( .A1(n10257), .A2(n10542), .ZN(n10546) );
  INV_X1 U13532 ( .A(n10755), .ZN(n10543) );
  NAND2_X1 U13533 ( .A1(n10765), .A2(n10543), .ZN(n10545) );
  NAND2_X1 U13534 ( .A1(n19877), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10544) );
  NAND2_X1 U13535 ( .A1(n10545), .A2(n10544), .ZN(n10549) );
  XNOR2_X1 U13536 ( .A(n10549), .B(n10547), .ZN(n10919) );
  NAND2_X1 U13537 ( .A1(n10279), .A2(n10919), .ZN(n10918) );
  NAND2_X1 U13538 ( .A1(n10546), .A2(n10918), .ZN(n10768) );
  INV_X1 U13539 ( .A(n10547), .ZN(n10548) );
  NAND2_X1 U13540 ( .A1(n10549), .A2(n10548), .ZN(n10551) );
  NAND2_X1 U13541 ( .A1(n19868), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10550) );
  XNOR2_X1 U13542 ( .A(n10553), .B(n10554), .ZN(n10752) );
  MUX2_X1 U13543 ( .A(n11039), .B(n10752), .S(n10279), .Z(n10767) );
  INV_X1 U13544 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n10552) );
  MUX2_X1 U13545 ( .A(n10767), .B(n10552), .S(n19265), .Z(n10563) );
  NAND3_X1 U13546 ( .A1(n15505), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(
        n10754), .ZN(n10766) );
  INV_X1 U13547 ( .A(n10787), .ZN(n11044) );
  MUX2_X1 U13548 ( .A(n10766), .B(n11044), .S(n10257), .Z(n10557) );
  INV_X1 U13549 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n14127) );
  MUX2_X1 U13550 ( .A(n10557), .B(n14127), .S(n19265), .Z(n10558) );
  INV_X1 U13551 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n13386) );
  MUX2_X1 U13552 ( .A(n13386), .B(n11048), .S(n10742), .Z(n10559) );
  NOR2_X1 U13553 ( .A1(n10575), .A2(n10559), .ZN(n10560) );
  OR2_X1 U13554 ( .A1(n10631), .A2(n10560), .ZN(n19043) );
  INV_X1 U13555 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13867) );
  XNOR2_X1 U13556 ( .A(n10583), .B(n13867), .ZN(n13852) );
  OAI21_X1 U13557 ( .B1(n9846), .B2(n10563), .A(n10577), .ZN(n14163) );
  NOR2_X1 U13558 ( .A1(n10571), .A2(n10564), .ZN(n10565) );
  OR2_X1 U13559 ( .A1(n9846), .A2(n10565), .ZN(n14825) );
  OAI21_X1 U13560 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19886), .A(
        n10755), .ZN(n10921) );
  MUX2_X1 U13561 ( .A(n10921), .B(n13221), .S(n10257), .Z(n10568) );
  INV_X1 U13562 ( .A(n10566), .ZN(n10567) );
  AOI21_X1 U13563 ( .B1(n10568), .B2(n10742), .A(n10567), .ZN(n19059) );
  NAND2_X1 U13564 ( .A1(n19059), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13305) );
  AND2_X1 U13565 ( .A1(n10569), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10570) );
  OR2_X1 U13566 ( .A1(n10571), .A2(n10570), .ZN(n14836) );
  NOR2_X1 U13567 ( .A1(n13305), .A2(n14836), .ZN(n10572) );
  NAND2_X1 U13568 ( .A1(n13305), .A2(n14836), .ZN(n13304) );
  OAI21_X1 U13569 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n10572), .A(
        n13304), .ZN(n13280) );
  XNOR2_X1 U13570 ( .A(n14825), .B(n19235), .ZN(n13279) );
  OR2_X1 U13571 ( .A1(n13280), .A2(n13279), .ZN(n13282) );
  OAI21_X1 U13572 ( .B1(n14825), .B2(n19235), .A(n13282), .ZN(n13615) );
  OAI21_X1 U13573 ( .B1(n13614), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n13615), .ZN(n10574) );
  NAND2_X1 U13574 ( .A1(n13614), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10573) );
  NAND2_X1 U13575 ( .A1(n10574), .A2(n10573), .ZN(n13753) );
  INV_X1 U13576 ( .A(n10575), .ZN(n10579) );
  NAND2_X1 U13577 ( .A1(n10577), .A2(n10576), .ZN(n10578) );
  NAND2_X1 U13578 ( .A1(n10579), .A2(n10578), .ZN(n10580) );
  XNOR2_X1 U13579 ( .A(n10580), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13754) );
  NAND2_X1 U13580 ( .A1(n13753), .A2(n13754), .ZN(n10582) );
  INV_X1 U13581 ( .A(n10580), .ZN(n14150) );
  NAND2_X1 U13582 ( .A1(n14150), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10581) );
  NAND2_X1 U13583 ( .A1(n13852), .A2(n13853), .ZN(n10585) );
  NAND2_X1 U13584 ( .A1(n10583), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10584) );
  NAND2_X1 U13585 ( .A1(n10585), .A2(n10584), .ZN(n15119) );
  AOI22_X1 U13586 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19287), .B1(
        n10477), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10589) );
  AOI22_X1 U13587 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n13718), .B1(
        n10478), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10588) );
  AOI22_X1 U13588 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19573), .B1(
        n19640), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10587) );
  AOI22_X1 U13589 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19348), .B1(
        n10476), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10586) );
  AOI22_X1 U13590 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19417), .B1(
        n10590), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10592) );
  AOI22_X1 U13591 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10483), .B1(
        n19687), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10591) );
  NAND3_X1 U13592 ( .A1(n10593), .A2(n10592), .A3(n10591), .ZN(n10600) );
  INV_X1 U13593 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10607) );
  INV_X1 U13594 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11178) );
  OAI22_X1 U13595 ( .A1(n10607), .A2(n10595), .B1(n10594), .B2(n11178), .ZN(
        n10599) );
  INV_X1 U13596 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12662) );
  INV_X1 U13597 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12658) );
  OAI22_X1 U13598 ( .A1(n12662), .A2(n10597), .B1(n10596), .B2(n12658), .ZN(
        n10598) );
  INV_X1 U13599 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10601) );
  OR2_X1 U13600 ( .A1(n12689), .A2(n10601), .ZN(n10605) );
  AOI22_X1 U13601 ( .A1(n10462), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10400), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10604) );
  NAND2_X1 U13602 ( .A1(n10456), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n10603) );
  NAND2_X1 U13603 ( .A1(n12706), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10602) );
  AOI22_X1 U13604 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10500), .B1(
        n10413), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10612) );
  NAND2_X1 U13605 ( .A1(n10395), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n10611) );
  NAND2_X1 U13606 ( .A1(n10401), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n10610) );
  NAND2_X1 U13607 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n12696), .ZN(
        n10606) );
  OAI21_X1 U13608 ( .B1(n12699), .B2(n10607), .A(n10606), .ZN(n10608) );
  AOI21_X1 U13609 ( .B1(n10414), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n10608), .ZN(n10609) );
  AOI22_X1 U13610 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10467), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10614) );
  AOI22_X1 U13611 ( .A1(n12695), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12690), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10613) );
  NAND4_X1 U13612 ( .A1(n10616), .A2(n10615), .A3(n10614), .A4(n10613), .ZN(
        n11051) );
  INV_X1 U13613 ( .A(n11051), .ZN(n10617) );
  NAND2_X1 U13614 ( .A1(n10617), .A2(n9788), .ZN(n10618) );
  MUX2_X1 U13615 ( .A(n20987), .B(n11051), .S(n10742), .Z(n10627) );
  XNOR2_X1 U13616 ( .A(n10631), .B(n10627), .ZN(n19027) );
  INV_X1 U13617 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n20863) );
  XNOR2_X1 U13618 ( .A(n10622), .B(n20863), .ZN(n15120) );
  NAND2_X1 U13619 ( .A1(n15119), .A2(n15120), .ZN(n15110) );
  NAND2_X1 U13620 ( .A1(n10631), .A2(n10627), .ZN(n10621) );
  MUX2_X1 U13621 ( .A(P2_EBX_REG_7__SCAN_IN), .B(n11055), .S(n10742), .Z(
        n10628) );
  INV_X1 U13622 ( .A(n10628), .ZN(n10620) );
  XNOR2_X1 U13623 ( .A(n10621), .B(n10620), .ZN(n19019) );
  AND2_X1 U13624 ( .A1(n19019), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15108) );
  INV_X1 U13625 ( .A(n15108), .ZN(n10623) );
  NAND2_X1 U13626 ( .A1(n10622), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15111) );
  AND2_X1 U13627 ( .A1(n10623), .A2(n15111), .ZN(n10624) );
  NAND2_X1 U13628 ( .A1(n15110), .A2(n10624), .ZN(n10626) );
  INV_X1 U13629 ( .A(n19019), .ZN(n10625) );
  INV_X1 U13630 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16326) );
  NAND2_X1 U13631 ( .A1(n10625), .A2(n16326), .ZN(n10634) );
  NAND2_X1 U13632 ( .A1(n10626), .A2(n10634), .ZN(n16275) );
  INV_X1 U13633 ( .A(n10627), .ZN(n10629) );
  NOR2_X1 U13634 ( .A1(n10629), .A2(n10628), .ZN(n10630) );
  INV_X1 U13635 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n10836) );
  NOR2_X1 U13636 ( .A1(n10742), .A2(n10836), .ZN(n10632) );
  AND2_X1 U13637 ( .A1(n10640), .A2(n10632), .ZN(n10633) );
  OR2_X1 U13638 ( .A1(n10639), .A2(n10633), .ZN(n14814) );
  NOR2_X1 U13639 ( .A1(n14814), .A2(n11055), .ZN(n10635) );
  NAND2_X1 U13640 ( .A1(n10635), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16276) );
  INV_X1 U13641 ( .A(n10634), .ZN(n15109) );
  OR2_X1 U13642 ( .A1(n16276), .A2(n15109), .ZN(n10637) );
  INV_X1 U13643 ( .A(n10635), .ZN(n10636) );
  INV_X1 U13644 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16327) );
  INV_X1 U13645 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10845) );
  NOR2_X1 U13646 ( .A1(n10742), .A2(n10845), .ZN(n10638) );
  XNOR2_X1 U13647 ( .A(n10639), .B(n10638), .ZN(n19009) );
  NAND2_X1 U13648 ( .A1(n19009), .A2(n10808), .ZN(n10647) );
  INV_X1 U13649 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15308) );
  NAND2_X1 U13650 ( .A1(n10647), .A2(n15308), .ZN(n15304) );
  NAND3_X1 U13651 ( .A1(n9857), .A2(n19265), .A3(P2_EBX_REG_10__SCAN_IN), .ZN(
        n10641) );
  OAI211_X1 U13652 ( .C1(n9857), .C2(P2_EBX_REG_10__SCAN_IN), .A(n10729), .B(
        n10641), .ZN(n14799) );
  OR2_X1 U13653 ( .A1(n14799), .A2(n11055), .ZN(n10642) );
  INV_X1 U13654 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16248) );
  INV_X1 U13655 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13704) );
  NAND2_X1 U13656 ( .A1(n10729), .A2(n10652), .ZN(n10651) );
  INV_X1 U13657 ( .A(n10651), .ZN(n10646) );
  INV_X1 U13658 ( .A(n10643), .ZN(n10644) );
  NAND3_X1 U13659 ( .A1(n19265), .A2(P2_EBX_REG_11__SCAN_IN), .A3(n10644), 
        .ZN(n10645) );
  NAND2_X1 U13660 ( .A1(n10646), .A2(n10645), .ZN(n10649) );
  INV_X1 U13661 ( .A(n10649), .ZN(n18998) );
  AOI21_X1 U13662 ( .B1(n18998), .B2(n10808), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15095) );
  OR3_X1 U13663 ( .A1(n14799), .A2(n11055), .A3(n16248), .ZN(n16253) );
  NAND2_X1 U13664 ( .A1(n10808), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10648) );
  OR2_X1 U13665 ( .A1(n10649), .A2(n10648), .ZN(n15093) );
  AND3_X1 U13666 ( .A1(n16252), .A2(n16253), .A3(n15093), .ZN(n10650) );
  NAND2_X1 U13667 ( .A1(n19265), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10654) );
  INV_X1 U13668 ( .A(n10652), .ZN(n10653) );
  OR2_X1 U13669 ( .A1(n10654), .A2(n10653), .ZN(n10655) );
  NAND2_X1 U13670 ( .A1(n10680), .A2(n10655), .ZN(n14784) );
  NAND2_X1 U13671 ( .A1(n10808), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10656) );
  NOR2_X1 U13672 ( .A1(n14784), .A2(n10656), .ZN(n16238) );
  INV_X1 U13673 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n10657) );
  NOR2_X1 U13674 ( .A1(n10742), .A2(n10657), .ZN(n10678) );
  OAI21_X1 U13675 ( .B1(P2_EBX_REG_15__SCAN_IN), .B2(P2_EBX_REG_14__SCAN_IN), 
        .A(n19265), .ZN(n10658) );
  NAND3_X1 U13676 ( .A1(n10664), .A2(n19265), .A3(P2_EBX_REG_16__SCAN_IN), 
        .ZN(n10659) );
  NAND3_X1 U13677 ( .A1(n10666), .A2(n10729), .A3(n10659), .ZN(n18976) );
  NOR2_X1 U13678 ( .A1(n11055), .A2(n18976), .ZN(n10691) );
  XOR2_X1 U13679 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n10691), .Z(
        n15059) );
  NAND2_X1 U13680 ( .A1(n19265), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10660) );
  MUX2_X1 U13681 ( .A(n10660), .B(n19265), .S(n9816), .Z(n10662) );
  INV_X1 U13682 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n10661) );
  NAND2_X1 U13683 ( .A1(n9816), .A2(n10661), .ZN(n10663) );
  NAND2_X1 U13684 ( .A1(n10662), .A2(n10663), .ZN(n14761) );
  NOR2_X1 U13685 ( .A1(n11055), .A2(n14761), .ZN(n10693) );
  OR2_X1 U13686 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n10693), .ZN(
        n16229) );
  NAND3_X1 U13687 ( .A1(n10663), .A2(P2_EBX_REG_15__SCAN_IN), .A3(n19265), 
        .ZN(n10665) );
  NAND2_X1 U13688 ( .A1(n10665), .A2(n10664), .ZN(n18984) );
  NOR2_X1 U13689 ( .A1(n11055), .A2(n18984), .ZN(n10694) );
  NOR2_X1 U13690 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n10694), .ZN(
        n15069) );
  NAND2_X1 U13691 ( .A1(n19265), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10667) );
  NAND2_X1 U13692 ( .A1(n19265), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10673) );
  MUX2_X1 U13693 ( .A(n19265), .B(n10667), .S(n10676), .Z(n10668) );
  OR2_X1 U13694 ( .A1(n10676), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10669) );
  NAND3_X1 U13695 ( .A1(n10669), .A2(n19265), .A3(P2_EBX_REG_19__SCAN_IN), 
        .ZN(n10672) );
  NOR2_X1 U13696 ( .A1(P2_EBX_REG_19__SCAN_IN), .A2(P2_EBX_REG_18__SCAN_IN), 
        .ZN(n10670) );
  NOR2_X1 U13697 ( .A1(n10742), .A2(n10670), .ZN(n10671) );
  AND2_X1 U13698 ( .A1(n10672), .A2(n9825), .ZN(n18931) );
  AND2_X1 U13699 ( .A1(n15227), .A2(n15036), .ZN(n11302) );
  OR2_X1 U13700 ( .A1(n10674), .A2(n10673), .ZN(n10675) );
  NAND2_X1 U13701 ( .A1(n10676), .A2(n10675), .ZN(n18955) );
  NOR2_X1 U13702 ( .A1(n18955), .A2(n11055), .ZN(n10692) );
  OR2_X1 U13703 ( .A1(n10692), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15050) );
  OR2_X1 U13704 ( .A1(n14784), .A2(n11055), .ZN(n10677) );
  INV_X1 U13705 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16305) );
  INV_X1 U13706 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15279) );
  INV_X1 U13707 ( .A(n10678), .ZN(n10679) );
  XNOR2_X1 U13708 ( .A(n10680), .B(n10679), .ZN(n14768) );
  NAND2_X1 U13709 ( .A1(n14768), .A2(n10808), .ZN(n10698) );
  AND2_X1 U13710 ( .A1(n15279), .A2(n10698), .ZN(n15079) );
  NOR2_X1 U13711 ( .A1(n16239), .A2(n15079), .ZN(n11297) );
  AND2_X1 U13712 ( .A1(n15050), .A2(n11297), .ZN(n10687) );
  INV_X1 U13713 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n14903) );
  NAND2_X1 U13714 ( .A1(n10703), .A2(n10729), .ZN(n10701) );
  NAND2_X1 U13715 ( .A1(n19265), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10681) );
  NOR2_X1 U13716 ( .A1(n10682), .A2(n10681), .ZN(n10683) );
  OR2_X1 U13717 ( .A1(n14748), .A2(n11055), .ZN(n10684) );
  INV_X1 U13718 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10812) );
  NAND2_X1 U13719 ( .A1(n10684), .A2(n10812), .ZN(n15022) );
  NAND2_X1 U13720 ( .A1(n19265), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10685) );
  XNOR2_X1 U13721 ( .A(n9825), .B(n10685), .ZN(n18922) );
  NAND2_X1 U13722 ( .A1(n18922), .A2(n10808), .ZN(n10697) );
  INV_X1 U13723 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12500) );
  INV_X1 U13724 ( .A(n15026), .ZN(n10686) );
  NAND4_X1 U13725 ( .A1(n11302), .A2(n10687), .A3(n15022), .A4(n10686), .ZN(
        n10688) );
  NOR2_X1 U13726 ( .A1(n15069), .A2(n10688), .ZN(n10689) );
  AND3_X1 U13727 ( .A1(n15059), .A2(n16229), .A3(n10689), .ZN(n10690) );
  NAND2_X1 U13728 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n10691), .ZN(
        n15049) );
  NAND2_X1 U13729 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n10692), .ZN(
        n15051) );
  AND2_X1 U13730 ( .A1(n15049), .A2(n15051), .ZN(n11301) );
  NAND2_X1 U13731 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n10693), .ZN(
        n16230) );
  NAND2_X1 U13732 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n10694), .ZN(
        n15070) );
  NAND2_X1 U13733 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n10695), .ZN(
        n15037) );
  NAND2_X1 U13734 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n10696), .ZN(
        n15226) );
  INV_X1 U13735 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n14900) );
  NOR2_X1 U13736 ( .A1(n10742), .A2(n14900), .ZN(n10702) );
  INV_X1 U13737 ( .A(n10702), .ZN(n10700) );
  NAND2_X1 U13738 ( .A1(n10701), .A2(n10700), .ZN(n10710) );
  NAND2_X1 U13739 ( .A1(n10703), .A2(n10702), .ZN(n10704) );
  NAND2_X1 U13740 ( .A1(n10710), .A2(n10704), .ZN(n15708) );
  OR2_X1 U13741 ( .A1(n15708), .A2(n11055), .ZN(n10705) );
  INV_X1 U13742 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15192) );
  NAND2_X1 U13743 ( .A1(n10705), .A2(n15192), .ZN(n15187) );
  INV_X1 U13744 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n10888) );
  NOR2_X1 U13745 ( .A1(n10742), .A2(n10888), .ZN(n10709) );
  INV_X1 U13746 ( .A(n10709), .ZN(n10706) );
  XNOR2_X1 U13747 ( .A(n10710), .B(n10706), .ZN(n16178) );
  NAND2_X1 U13748 ( .A1(n16178), .A2(n10808), .ZN(n10707) );
  XNOR2_X1 U13749 ( .A(n10707), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15014) );
  NAND2_X1 U13750 ( .A1(n15015), .A2(n15014), .ZN(n15016) );
  INV_X1 U13751 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15180) );
  OR2_X1 U13752 ( .A1(n10707), .A2(n15180), .ZN(n10708) );
  NAND3_X1 U13753 ( .A1(n10711), .A2(P2_EBX_REG_24__SCAN_IN), .A3(n19265), 
        .ZN(n10712) );
  NAND2_X1 U13754 ( .A1(n10712), .A2(n10729), .ZN(n10713) );
  OR2_X1 U13755 ( .A1(n10726), .A2(n10713), .ZN(n16170) );
  INV_X1 U13756 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15167) );
  NAND2_X1 U13757 ( .A1(n10714), .A2(n15167), .ZN(n15162) );
  INV_X1 U13758 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n14872) );
  NAND2_X1 U13759 ( .A1(n10726), .A2(n14872), .ZN(n10731) );
  NAND3_X1 U13760 ( .A1(n19265), .A2(P2_EBX_REG_26__SCAN_IN), .A3(n10731), 
        .ZN(n10716) );
  INV_X1 U13761 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15153) );
  NOR2_X1 U13762 ( .A1(n11055), .A2(n15153), .ZN(n10717) );
  NAND2_X1 U13763 ( .A1(n16144), .A2(n10717), .ZN(n10740) );
  INV_X1 U13764 ( .A(n16144), .ZN(n10718) );
  OAI21_X1 U13765 ( .B1(n10718), .B2(n11055), .A(n15153), .ZN(n10719) );
  NAND2_X1 U13766 ( .A1(n10740), .A2(n10719), .ZN(n14996) );
  NAND2_X1 U13767 ( .A1(n19265), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10721) );
  INV_X1 U13768 ( .A(n10721), .ZN(n10724) );
  INV_X1 U13769 ( .A(n10722), .ZN(n10723) );
  NAND2_X1 U13770 ( .A1(n10724), .A2(n10723), .ZN(n10725) );
  NAND2_X1 U13771 ( .A1(n10736), .A2(n10725), .ZN(n16135) );
  NOR2_X1 U13772 ( .A1(n10726), .A2(n14872), .ZN(n10727) );
  NAND2_X1 U13773 ( .A1(n19265), .A2(n10727), .ZN(n10728) );
  AND2_X1 U13774 ( .A1(n10729), .A2(n10728), .ZN(n10730) );
  NAND2_X1 U13775 ( .A1(n10731), .A2(n10730), .ZN(n16156) );
  INV_X1 U13776 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n10896) );
  NAND2_X1 U13777 ( .A1(n10739), .A2(n10896), .ZN(n14993) );
  NAND2_X1 U13778 ( .A1(n12467), .A2(n10734), .ZN(n10738) );
  INV_X1 U13779 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15144) );
  INV_X1 U13780 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12471) );
  INV_X1 U13781 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n10904) );
  NOR2_X1 U13782 ( .A1(n10742), .A2(n10904), .ZN(n10735) );
  NAND2_X1 U13783 ( .A1(n10736), .A2(n10735), .ZN(n10737) );
  NAND2_X1 U13784 ( .A1(n10745), .A2(n10737), .ZN(n14731) );
  NOR2_X1 U13785 ( .A1(n14731), .A2(n11055), .ZN(n12472) );
  INV_X1 U13786 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n10741) );
  NOR2_X1 U13787 ( .A1(n10742), .A2(n10741), .ZN(n10744) );
  XNOR2_X1 U13788 ( .A(n10745), .B(n10744), .ZN(n10743) );
  INV_X1 U13789 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n10910) );
  OAI21_X1 U13790 ( .B1(n10743), .B2(n11055), .A(n10910), .ZN(n14984) );
  NAND2_X1 U13791 ( .A1(n14985), .A2(n14984), .ZN(n10945) );
  INV_X1 U13792 ( .A(n10743), .ZN(n16121) );
  NAND3_X1 U13793 ( .A1(n16121), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n10808), .ZN(n14983) );
  NAND2_X1 U13794 ( .A1(n10945), .A2(n14983), .ZN(n10751) );
  INV_X1 U13795 ( .A(n10947), .ZN(n10747) );
  NAND2_X1 U13796 ( .A1(n19265), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10746) );
  XNOR2_X1 U13797 ( .A(n10747), .B(n10746), .ZN(n14676) );
  AOI21_X1 U13798 ( .B1(n14676), .B2(n10808), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10944) );
  NOR2_X1 U13799 ( .A1(n11055), .A2(n10815), .ZN(n10748) );
  NAND2_X1 U13800 ( .A1(n14676), .A2(n10748), .ZN(n10943) );
  INV_X1 U13801 ( .A(n10943), .ZN(n10749) );
  NOR2_X1 U13802 ( .A1(n10944), .A2(n10749), .ZN(n10750) );
  XNOR2_X1 U13803 ( .A(n10751), .B(n10750), .ZN(n14080) );
  NAND2_X1 U13804 ( .A1(n10919), .A2(n10932), .ZN(n10759) );
  XNOR2_X1 U13805 ( .A(n10765), .B(n10755), .ZN(n10922) );
  INV_X1 U13806 ( .A(n10759), .ZN(n10756) );
  INV_X1 U13807 ( .A(n13072), .ZN(n10758) );
  OAI21_X1 U13808 ( .B1(n10921), .B2(n10759), .A(n10758), .ZN(n10760) );
  INV_X1 U13809 ( .A(n10760), .ZN(n10764) );
  AND2_X1 U13810 ( .A1(n15505), .A2(n10761), .ZN(n16346) );
  NAND2_X1 U13811 ( .A1(n11202), .A2(n16346), .ZN(n10763) );
  INV_X1 U13812 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n10762) );
  NAND2_X1 U13813 ( .A1(n10763), .A2(n10762), .ZN(n19878) );
  MUX2_X1 U13814 ( .A(n10764), .B(n19878), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n16361) );
  NOR2_X1 U13815 ( .A1(n10772), .A2(n15768), .ZN(n10775) );
  INV_X1 U13816 ( .A(n10765), .ZN(n10920) );
  NOR2_X1 U13817 ( .A1(n10920), .A2(n10921), .ZN(n10769) );
  OAI211_X1 U13818 ( .C1(n10769), .C2(n10768), .A(n10767), .B(n10766), .ZN(
        n10770) );
  INV_X1 U13819 ( .A(n10770), .ZN(n10771) );
  OR2_X1 U13820 ( .A1(n10936), .A2(n10771), .ZN(n13069) );
  INV_X1 U13821 ( .A(n10772), .ZN(n10773) );
  NAND2_X1 U13822 ( .A1(n10773), .A2(n10274), .ZN(n16351) );
  NOR2_X1 U13823 ( .A1(n13069), .A2(n16351), .ZN(n10774) );
  MUX2_X1 U13824 ( .A(n10775), .B(n10774), .S(n9788), .Z(n10971) );
  AND2_X1 U13825 ( .A1(n10274), .A2(n19768), .ZN(n10776) );
  INV_X1 U13826 ( .A(n13622), .ZN(n10783) );
  NAND2_X1 U13827 ( .A1(n13221), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13220) );
  NOR2_X1 U13828 ( .A1(n11024), .A2(n13220), .ZN(n10778) );
  AND2_X1 U13829 ( .A1(n13221), .A2(n13219), .ZN(n10777) );
  XNOR2_X1 U13830 ( .A(n10777), .B(n11024), .ZN(n13308) );
  NOR2_X1 U13831 ( .A1(n15370), .A2(n13308), .ZN(n13307) );
  NOR2_X1 U13832 ( .A1(n10778), .A2(n13307), .ZN(n10780) );
  XNOR2_X1 U13833 ( .A(n10779), .B(n11034), .ZN(n13285) );
  NAND2_X1 U13834 ( .A1(n10138), .A2(n13285), .ZN(n13284) );
  OR2_X1 U13835 ( .A1(n10780), .A2(n19235), .ZN(n10781) );
  NAND2_X1 U13836 ( .A1(n13284), .A2(n10781), .ZN(n10784) );
  XNOR2_X1 U13837 ( .A(n10784), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13623) );
  INV_X1 U13838 ( .A(n13623), .ZN(n10782) );
  NAND2_X1 U13839 ( .A1(n10784), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10785) );
  NAND2_X1 U13840 ( .A1(n10786), .A2(n10787), .ZN(n10788) );
  INV_X1 U13841 ( .A(n13757), .ZN(n10789) );
  INV_X1 U13842 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13866) );
  NAND2_X1 U13843 ( .A1(n10790), .A2(n13867), .ZN(n13854) );
  NAND2_X1 U13844 ( .A1(n10793), .A2(n10792), .ZN(n10798) );
  INV_X1 U13845 ( .A(n13855), .ZN(n10796) );
  NAND2_X1 U13846 ( .A1(n10796), .A2(n10800), .ZN(n10797) );
  INV_X1 U13847 ( .A(n10800), .ZN(n10801) );
  XNOR2_X1 U13848 ( .A(n10810), .B(n10808), .ZN(n10804) );
  NAND2_X1 U13849 ( .A1(n10803), .A2(n10804), .ZN(n15105) );
  INV_X1 U13850 ( .A(n10803), .ZN(n10806) );
  INV_X1 U13851 ( .A(n10804), .ZN(n10805) );
  NAND2_X1 U13852 ( .A1(n10808), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10809) );
  NAND3_X1 U13853 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16295) );
  NOR2_X1 U13854 ( .A1(n16295), .A2(n16305), .ZN(n11264) );
  INV_X1 U13855 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16233) );
  NAND2_X1 U13856 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15209) );
  NOR2_X1 U13857 ( .A1(n15209), .A2(n10812), .ZN(n11272) );
  AND2_X1 U13858 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11285) );
  AND2_X1 U13859 ( .A1(n11272), .A2(n11285), .ZN(n10813) );
  NAND2_X1 U13860 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11005) );
  INV_X1 U13861 ( .A(n11005), .ZN(n15241) );
  AND2_X1 U13862 ( .A1(n10813), .A2(n15241), .ZN(n15020) );
  AND2_X1 U13863 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n15020), .ZN(
        n10814) );
  NAND3_X1 U13864 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14067) );
  XNOR2_X1 U13865 ( .A(n10979), .B(n10815), .ZN(n14078) );
  NOR2_X2 U13866 ( .A1(n18899), .A2(n9790), .ZN(n19204) );
  NAND2_X1 U13867 ( .A1(n14078), .A2(n19204), .ZN(n10942) );
  NOR2_X1 U13868 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19764) );
  OR2_X1 U13869 ( .A1(n19856), .A2(n19764), .ZN(n19869) );
  NAND2_X1 U13870 ( .A1(n19869), .A2(n18894), .ZN(n10816) );
  NAND2_X1 U13871 ( .A1(n19856), .A2(n10329), .ZN(n18893) );
  INV_X2 U13872 ( .A(n15334), .ZN(n19030) );
  INV_X1 U13873 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n19836) );
  NOR2_X1 U13874 ( .A1(n18957), .A2(n19836), .ZN(n14070) );
  INV_X1 U13875 ( .A(n10817), .ZN(n10822) );
  NOR2_X1 U13876 ( .A1(n10820), .A2(n10819), .ZN(n10821) );
  AOI22_X1 U13877 ( .A1(n10823), .A2(P2_EBX_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10825) );
  NAND2_X1 U13878 ( .A1(n9782), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n10824) );
  OAI211_X1 U13879 ( .C1(n10333), .C2(n13866), .A(n10825), .B(n10824), .ZN(
        n13759) );
  NAND2_X1 U13880 ( .A1(n9782), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n10828) );
  NAND2_X1 U13881 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10827) );
  OAI211_X1 U13882 ( .C1(n10905), .C2(n13386), .A(n10828), .B(n10827), .ZN(
        n10829) );
  INV_X1 U13883 ( .A(n10829), .ZN(n10830) );
  OAI21_X1 U13884 ( .B1(n10333), .B2(n13867), .A(n10830), .ZN(n13383) );
  NAND2_X1 U13885 ( .A1(n9782), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n10832) );
  NAND2_X1 U13886 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10831) );
  OAI211_X1 U13887 ( .C1(n10905), .C2(n20987), .A(n10832), .B(n10831), .ZN(
        n10833) );
  AOI21_X1 U13888 ( .B1(n10907), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n10833), .ZN(n13376) );
  NAND2_X1 U13889 ( .A1(n9782), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n10835) );
  NAND2_X1 U13890 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10834) );
  OAI211_X1 U13891 ( .C1(n10905), .C2(n10836), .A(n10835), .B(n10834), .ZN(
        n10837) );
  AOI21_X1 U13892 ( .B1(n10907), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n10837), .ZN(n13579) );
  INV_X1 U13893 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n10840) );
  NAND2_X1 U13894 ( .A1(n9782), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n10839) );
  NAND2_X1 U13895 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10838) );
  OAI211_X1 U13896 ( .C1(n10905), .C2(n10840), .A(n10839), .B(n10838), .ZN(
        n10841) );
  AOI21_X1 U13897 ( .B1(n10907), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n10841), .ZN(n13519) );
  OR2_X1 U13898 ( .A1(n13579), .A2(n13519), .ZN(n10842) );
  NAND2_X1 U13899 ( .A1(n9782), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n10844) );
  NAND2_X1 U13900 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10843) );
  OAI211_X1 U13901 ( .C1(n10905), .C2(n10845), .A(n10844), .B(n10843), .ZN(
        n10846) );
  INV_X1 U13902 ( .A(n10846), .ZN(n10847) );
  OAI21_X1 U13903 ( .B1(n10333), .B2(n15308), .A(n10847), .ZN(n13590) );
  AOI22_X1 U13904 ( .A1(n10823), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n10849) );
  NAND2_X1 U13905 ( .A1(n9782), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n10848) );
  OAI211_X1 U13906 ( .C1(n10333), .C2(n16248), .A(n10849), .B(n10848), .ZN(
        n13664) );
  INV_X1 U13907 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n15101) );
  AOI22_X1 U13908 ( .A1(n10823), .A2(P2_EBX_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n10850) );
  OAI21_X1 U13909 ( .B1(n10874), .B2(n15101), .A(n10850), .ZN(n10851) );
  AOI21_X1 U13910 ( .B1(n10907), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n10851), .ZN(n13701) );
  AOI22_X1 U13911 ( .A1(n10823), .A2(P2_EBX_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n10853) );
  NAND2_X1 U13912 ( .A1(n9782), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n10852) );
  OAI211_X1 U13913 ( .C1(n10333), .C2(n16305), .A(n10853), .B(n10852), .ZN(
        n13781) );
  INV_X1 U13914 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n10855) );
  AOI22_X1 U13915 ( .A1(n10823), .A2(P2_EBX_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n10854) );
  OAI21_X1 U13916 ( .B1(n10874), .B2(n10855), .A(n10854), .ZN(n10856) );
  AOI21_X1 U13917 ( .B1(n10907), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n10856), .ZN(n13879) );
  AOI22_X1 U13918 ( .A1(n10823), .A2(P2_EBX_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n10858) );
  NAND2_X1 U13919 ( .A1(n9782), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n10857) );
  OAI211_X1 U13920 ( .C1(n10333), .C2(n16233), .A(n10858), .B(n10857), .ZN(
        n13831) );
  INV_X1 U13921 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n10861) );
  NAND2_X1 U13922 ( .A1(n9782), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n10860) );
  NAND2_X1 U13923 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10859) );
  OAI211_X1 U13924 ( .C1(n10905), .C2(n10861), .A(n10860), .B(n10859), .ZN(
        n10862) );
  AOI21_X1 U13925 ( .B1(n10907), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n10862), .ZN(n13710) );
  INV_X1 U13926 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10865) );
  AOI22_X1 U13927 ( .A1(n10823), .A2(P2_EBX_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n10864) );
  NAND2_X1 U13928 ( .A1(n9782), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n10863) );
  OAI211_X1 U13929 ( .C1(n10333), .C2(n10865), .A(n10864), .B(n10863), .ZN(
        n13771) );
  INV_X1 U13930 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n10867) );
  INV_X1 U13931 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10866) );
  OAI22_X1 U13932 ( .A1(n10905), .A2(n10867), .B1(n10329), .B2(n10866), .ZN(
        n10869) );
  INV_X1 U13933 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15251) );
  NOR2_X1 U13934 ( .A1(n10333), .A2(n15251), .ZN(n10868) );
  AOI211_X1 U13935 ( .C1(n9782), .C2(P2_REIP_REG_17__SCAN_IN), .A(n10869), .B(
        n10868), .ZN(n13807) );
  INV_X1 U13936 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15232) );
  AOI22_X1 U13937 ( .A1(n10823), .A2(P2_EBX_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n10871) );
  NAND2_X1 U13938 ( .A1(n9782), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n10870) );
  OAI211_X1 U13939 ( .C1(n10333), .C2(n15232), .A(n10871), .B(n10870), .ZN(
        n13836) );
  INV_X1 U13940 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n10873) );
  AOI22_X1 U13941 ( .A1(n10823), .A2(P2_EBX_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n10872) );
  OAI21_X1 U13942 ( .B1(n10874), .B2(n10873), .A(n10872), .ZN(n10875) );
  AOI21_X1 U13943 ( .B1(n10907), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n10875), .ZN(n14907) );
  NAND2_X1 U13944 ( .A1(n9782), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n10877) );
  NAND2_X1 U13945 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10876) );
  OAI211_X1 U13946 ( .C1(n10905), .C2(n9943), .A(n10877), .B(n10876), .ZN(
        n10878) );
  INV_X1 U13947 ( .A(n10878), .ZN(n10879) );
  OAI21_X1 U13948 ( .B1(n10333), .B2(n12500), .A(n10879), .ZN(n11294) );
  NAND2_X1 U13949 ( .A1(n10826), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n10881) );
  NAND2_X1 U13950 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10880) );
  OAI211_X1 U13951 ( .C1(n10905), .C2(n14903), .A(n10881), .B(n10880), .ZN(
        n10882) );
  AOI21_X1 U13952 ( .B1(n10907), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n10882), .ZN(n14739) );
  NAND2_X1 U13953 ( .A1(n10826), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n10884) );
  NAND2_X1 U13954 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10883) );
  OAI211_X1 U13955 ( .C1(n10905), .C2(n14900), .A(n10884), .B(n10883), .ZN(
        n10885) );
  AOI21_X1 U13956 ( .B1(n10907), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n10885), .ZN(n14895) );
  NAND2_X1 U13957 ( .A1(n10826), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n10887) );
  NAND2_X1 U13958 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10886) );
  OAI211_X1 U13959 ( .C1(n10905), .C2(n10888), .A(n10887), .B(n10886), .ZN(
        n10889) );
  AOI21_X1 U13960 ( .B1(n10907), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n10889), .ZN(n14887) );
  AOI22_X1 U13961 ( .A1(n10823), .A2(P2_EBX_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n10891) );
  NAND2_X1 U13962 ( .A1(n10826), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n10890) );
  OAI211_X1 U13963 ( .C1(n10333), .C2(n15167), .A(n10891), .B(n10890), .ZN(
        n14878) );
  NAND2_X1 U13964 ( .A1(n9782), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n10893) );
  NAND2_X1 U13965 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n10892) );
  OAI211_X1 U13966 ( .C1(n10905), .C2(n14872), .A(n10893), .B(n10892), .ZN(
        n10894) );
  INV_X1 U13967 ( .A(n10894), .ZN(n10895) );
  OAI21_X1 U13968 ( .B1(n10333), .B2(n10896), .A(n10895), .ZN(n13945) );
  AOI22_X1 U13969 ( .A1(n10823), .A2(P2_EBX_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n10898) );
  NAND2_X1 U13970 ( .A1(n9782), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n10897) );
  OAI211_X1 U13971 ( .C1(n10333), .C2(n15153), .A(n10898), .B(n10897), .ZN(
        n14861) );
  INV_X1 U13972 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n20953) );
  NAND2_X1 U13973 ( .A1(n10826), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n10900) );
  NAND2_X1 U13974 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n10899) );
  OAI211_X1 U13975 ( .C1(n10905), .C2(n20953), .A(n10900), .B(n10899), .ZN(
        n10901) );
  AOI21_X1 U13976 ( .B1(n10907), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n10901), .ZN(n14046) );
  NAND2_X1 U13977 ( .A1(n9782), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n10903) );
  NAND2_X1 U13978 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10902) );
  OAI211_X1 U13979 ( .C1(n10905), .C2(n10904), .A(n10903), .B(n10902), .ZN(
        n10906) );
  AOI21_X1 U13980 ( .B1(n10907), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n10906), .ZN(n12475) );
  AOI22_X1 U13981 ( .A1(n10823), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n10909) );
  NAND2_X1 U13982 ( .A1(n10826), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n10908) );
  OAI211_X1 U13983 ( .C1(n10333), .C2(n10910), .A(n10909), .B(n10908), .ZN(
        n14841) );
  AOI22_X1 U13984 ( .A1(n10823), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n10912) );
  NAND2_X1 U13985 ( .A1(n9782), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n10911) );
  OAI211_X1 U13986 ( .C1(n10333), .C2(n10815), .A(n10912), .B(n10911), .ZN(
        n10914) );
  INV_X1 U13987 ( .A(n10913), .ZN(n10916) );
  INV_X1 U13988 ( .A(n10914), .ZN(n10915) );
  NAND2_X1 U13989 ( .A1(n10916), .A2(n10915), .ZN(n10917) );
  NAND2_X1 U13990 ( .A1(n10329), .A2(n19544), .ZN(n14670) );
  NAND2_X1 U13991 ( .A1(n10274), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10935) );
  AOI21_X1 U13992 ( .B1(n10935), .B2(n9790), .A(n10919), .ZN(n10930) );
  INV_X1 U13993 ( .A(n10918), .ZN(n10929) );
  INV_X1 U13994 ( .A(n10919), .ZN(n10927) );
  OAI21_X1 U13995 ( .B1(n10920), .B2(n10921), .A(n10257), .ZN(n10925) );
  INV_X1 U13996 ( .A(n10921), .ZN(n10923) );
  OAI211_X1 U13997 ( .C1(n9790), .C2(n10923), .A(n14666), .B(n10922), .ZN(
        n10924) );
  OAI211_X1 U13998 ( .C1(n10927), .C2(n10926), .A(n10925), .B(n10924), .ZN(
        n10928) );
  OAI211_X1 U13999 ( .C1(n10930), .C2(n10929), .A(n10932), .B(n10928), .ZN(
        n10931) );
  OAI21_X1 U14000 ( .B1(n10932), .B2(n10279), .A(n10931), .ZN(n10933) );
  OR2_X1 U14001 ( .A1(n10936), .A2(n10933), .ZN(n10934) );
  MUX2_X1 U14002 ( .A(n10934), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n18894), .Z(n10972) );
  NAND2_X1 U14003 ( .A1(n10936), .A2(n19140), .ZN(n10937) );
  NAND2_X1 U14004 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n15363) );
  NOR2_X1 U14005 ( .A1(n14168), .A2(n13644), .ZN(n10938) );
  INV_X1 U14006 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15029) );
  NAND2_X1 U14007 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n13618), .ZN(
        n14131) );
  INV_X1 U14008 ( .A(n14687), .ZN(n14693) );
  NAND2_X1 U14009 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n14696), .ZN(
        n14686) );
  NAND2_X1 U14010 ( .A1(n14699), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14698) );
  NAND2_X1 U14011 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n14701), .ZN(
        n14700) );
  NAND2_X1 U14012 ( .A1(n14705), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14706) );
  NAND2_X1 U14013 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n14709), .ZN(
        n14708) );
  INV_X1 U14014 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14679) );
  XNOR2_X1 U14015 ( .A(n14677), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14710) );
  NAND2_X1 U14016 ( .A1(n18894), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12523) );
  NAND2_X1 U14017 ( .A1(n19420), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n10939) );
  NAND2_X1 U14018 ( .A1(n12523), .A2(n10939), .ZN(n14123) );
  OR2_X1 U14019 ( .A1(n14710), .A2(n16262), .ZN(n10940) );
  OAI211_X1 U14020 ( .C1(n14080), .C2(n16263), .A(n10942), .B(n10131), .ZN(
        P2_U2984) );
  INV_X1 U14021 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n10946) );
  NAND2_X1 U14022 ( .A1(n10947), .A2(n10946), .ZN(n10948) );
  MUX2_X1 U14023 ( .A(n10949), .B(n10948), .S(n19265), .Z(n16114) );
  XOR2_X1 U14024 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n10950), .Z(
        n10951) );
  XNOR2_X1 U14025 ( .A(n10952), .B(n10951), .ZN(n14066) );
  NAND2_X1 U14026 ( .A1(n13074), .A2(n9790), .ZN(n19138) );
  NAND2_X1 U14027 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19765) );
  INV_X1 U14028 ( .A(n19765), .ZN(n19785) );
  INV_X1 U14029 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n18896) );
  NOR2_X1 U14030 ( .A1(n18896), .A2(n19792), .ZN(n19784) );
  NAND2_X1 U14031 ( .A1(n18896), .A2(n19792), .ZN(n19787) );
  NOR3_X1 U14032 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19784), .A3(n19773), 
        .ZN(n19778) );
  INV_X1 U14033 ( .A(n19778), .ZN(n14667) );
  NAND2_X1 U14034 ( .A1(n10266), .A2(n15359), .ZN(n10976) );
  NAND2_X1 U14035 ( .A1(n10953), .A2(n15359), .ZN(n10954) );
  OR2_X1 U14036 ( .A1(n13072), .A2(n10954), .ZN(n10966) );
  NAND2_X1 U14037 ( .A1(n10955), .A2(n9755), .ZN(n10957) );
  AND2_X1 U14038 ( .A1(n9788), .A2(n10274), .ZN(n10956) );
  NAND2_X1 U14039 ( .A1(n10957), .A2(n10956), .ZN(n10989) );
  NAND2_X1 U14040 ( .A1(n9788), .A2(n10265), .ZN(n10983) );
  NAND2_X1 U14041 ( .A1(n10983), .A2(n14666), .ZN(n10959) );
  NAND2_X1 U14042 ( .A1(n10959), .A2(n10958), .ZN(n10960) );
  INV_X1 U14043 ( .A(n10266), .ZN(n11255) );
  NAND2_X1 U14044 ( .A1(n10960), .A2(n11255), .ZN(n10964) );
  NAND2_X1 U14045 ( .A1(n10961), .A2(n11255), .ZN(n10962) );
  NAND2_X1 U14046 ( .A1(n15502), .A2(n10962), .ZN(n10963) );
  AND2_X1 U14047 ( .A1(n10966), .A2(n10985), .ZN(n15356) );
  MUX2_X1 U14048 ( .A(n10953), .B(n10266), .S(n9788), .Z(n10967) );
  NAND2_X1 U14049 ( .A1(n10967), .A2(n19765), .ZN(n10968) );
  OR2_X1 U14050 ( .A1(n10968), .A2(n13072), .ZN(n10969) );
  NAND2_X1 U14051 ( .A1(n15356), .A2(n10969), .ZN(n10970) );
  NOR2_X1 U14052 ( .A1(n10971), .A2(n10970), .ZN(n10975) );
  AOI21_X1 U14053 ( .B1(n10972), .B2(n14666), .A(n19259), .ZN(n10973) );
  NAND2_X1 U14054 ( .A1(n19138), .A2(n10973), .ZN(n10974) );
  OAI211_X1 U14055 ( .C1(n19138), .C2(n10976), .A(n10975), .B(n10974), .ZN(
        n10977) );
  INV_X1 U14056 ( .A(n16351), .ZN(n10978) );
  NAND2_X1 U14057 ( .A1(n10982), .A2(n9790), .ZN(n19225) );
  INV_X1 U14058 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10980) );
  XNOR2_X1 U14059 ( .A(n10981), .B(n10980), .ZN(n14064) );
  NAND2_X1 U14060 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19217) );
  NOR2_X1 U14061 ( .A1(n19235), .A2(n19217), .ZN(n11003) );
  INV_X1 U14062 ( .A(n10983), .ZN(n10984) );
  INV_X1 U14063 ( .A(n19217), .ZN(n19221) );
  NOR2_X1 U14064 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19221), .ZN(
        n13627) );
  INV_X1 U14065 ( .A(n13627), .ZN(n11262) );
  NAND2_X1 U14066 ( .A1(n10987), .A2(n10986), .ZN(n11000) );
  NAND2_X1 U14067 ( .A1(n10988), .A2(n9790), .ZN(n15352) );
  NAND2_X1 U14068 ( .A1(n15352), .A2(n10989), .ZN(n10990) );
  NAND2_X1 U14069 ( .A1(n10990), .A2(n10268), .ZN(n10997) );
  OAI21_X1 U14070 ( .B1(n14666), .B2(n10266), .A(n10991), .ZN(n10994) );
  NAND2_X1 U14071 ( .A1(n10993), .A2(n10992), .ZN(n12876) );
  OAI211_X1 U14072 ( .C1(n19259), .C2(n10986), .A(n10994), .B(n12876), .ZN(
        n10995) );
  INV_X1 U14073 ( .A(n10995), .ZN(n10996) );
  NAND2_X1 U14074 ( .A1(n10997), .A2(n10996), .ZN(n10998) );
  AOI21_X1 U14075 ( .B1(n11000), .B2(n10999), .A(n10998), .ZN(n15400) );
  NAND2_X1 U14076 ( .A1(n15400), .A2(n11001), .ZN(n11002) );
  NAND2_X1 U14077 ( .A1(n11259), .A2(n11002), .ZN(n19213) );
  OAI211_X1 U14078 ( .C1(n11003), .C2(n15245), .A(n11262), .B(n16294), .ZN(
        n11004) );
  INV_X1 U14079 ( .A(n11004), .ZN(n13763) );
  NAND3_X1 U14080 ( .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15317) );
  NOR2_X1 U14081 ( .A1(n13758), .A2(n15317), .ZN(n15320) );
  AND3_X1 U14082 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n15320), .ZN(n11263) );
  NAND3_X1 U14083 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n11264), .A3(
        n16307), .ZN(n16292) );
  NOR2_X1 U14084 ( .A1(n15251), .A2(n11005), .ZN(n11268) );
  NAND2_X1 U14085 ( .A1(n15272), .A2(n11268), .ZN(n15233) );
  NAND2_X1 U14086 ( .A1(n11272), .A2(n15220), .ZN(n15193) );
  NAND2_X1 U14087 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11260) );
  NOR2_X1 U14088 ( .A1(n15193), .A2(n11260), .ZN(n15168) );
  NAND2_X1 U14089 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15150) );
  NOR2_X1 U14090 ( .A1(n15167), .A2(n15150), .ZN(n11258) );
  NAND2_X1 U14091 ( .A1(n15168), .A2(n11258), .ZN(n14068) );
  NOR4_X1 U14092 ( .A1(n14068), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n10815), .A4(n14067), .ZN(n11282) );
  AOI22_X1 U14093 ( .A1(n10823), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n11007) );
  NAND2_X1 U14094 ( .A1(n10826), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n11006) );
  OAI211_X1 U14095 ( .C1(n10333), .C2(n10980), .A(n11007), .B(n11006), .ZN(
        n11008) );
  NAND2_X1 U14096 ( .A1(n11010), .A2(n9788), .ZN(n11011) );
  NAND2_X1 U14097 ( .A1(n11011), .A2(n10297), .ZN(n11012) );
  NAND2_X1 U14098 ( .A1(n11013), .A2(n19680), .ZN(n11017) );
  INV_X1 U14099 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18912) );
  AND2_X2 U14100 ( .A1(n9790), .A2(n19680), .ZN(n11018) );
  INV_X1 U14101 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n13050) );
  OAI21_X1 U14102 ( .B1(n9755), .B2(n13050), .A(n19680), .ZN(n11015) );
  AOI21_X1 U14103 ( .B1(n11018), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n11015), .ZN(n11016) );
  NAND2_X1 U14104 ( .A1(n12878), .A2(n11018), .ZN(n11032) );
  OAI22_X1 U14105 ( .A1(n9755), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n19886), 
        .B2(n19680), .ZN(n11019) );
  INV_X1 U14106 ( .A(n11019), .ZN(n11020) );
  AND2_X1 U14107 ( .A1(n11032), .A2(n11020), .ZN(n11021) );
  INV_X1 U14108 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19793) );
  NOR2_X1 U14109 ( .A1(n9755), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11022) );
  AOI22_X1 U14110 ( .A1(n11022), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n11018), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11023) );
  OAI21_X1 U14111 ( .B1(n11249), .B2(n19793), .A(n11023), .ZN(n11029) );
  OR2_X1 U14112 ( .A1(n11024), .A2(n11195), .ZN(n11027) );
  AND2_X1 U14113 ( .A1(n9755), .A2(n19680), .ZN(n11025) );
  AOI22_X1 U14114 ( .A1(n10281), .A2(n11025), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11026) );
  NAND2_X1 U14115 ( .A1(n11027), .A2(n11026), .ZN(n13445) );
  NOR2_X1 U14116 ( .A1(n13446), .A2(n13445), .ZN(n11031) );
  NOR2_X1 U14117 ( .A1(n11028), .A2(n11029), .ZN(n11030) );
  NAND2_X1 U14118 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11033) );
  OAI211_X1 U14119 ( .C1(n11195), .C2(n11034), .A(n11033), .B(n11032), .ZN(
        n11036) );
  XNOR2_X1 U14120 ( .A(n11037), .B(n11036), .ZN(n13441) );
  INV_X1 U14121 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19795) );
  INV_X2 U14122 ( .A(n11198), .ZN(n11250) );
  AOI22_X1 U14123 ( .A1(n11250), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n11018), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11035) );
  OAI21_X1 U14124 ( .B1(n11249), .B2(n19795), .A(n11035), .ZN(n13440) );
  NOR2_X1 U14125 ( .A1(n13441), .A2(n13440), .ZN(n13442) );
  NOR2_X1 U14126 ( .A1(n11037), .A2(n11036), .ZN(n11038) );
  NOR2_X2 U14127 ( .A1(n13442), .A2(n11038), .ZN(n13600) );
  NAND2_X1 U14128 ( .A1(n11251), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11043) );
  NAND2_X1 U14129 ( .A1(n11223), .A2(n11039), .ZN(n11042) );
  AOI22_X1 U14130 ( .A1(n11018), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11041) );
  NAND2_X1 U14131 ( .A1(n11250), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11040) );
  NAND4_X1 U14132 ( .A1(n11043), .A2(n11042), .A3(n11041), .A4(n11040), .ZN(
        n13599) );
  NAND2_X1 U14133 ( .A1(n13600), .A2(n13599), .ZN(n13601) );
  NAND2_X1 U14134 ( .A1(n11251), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11047) );
  NAND2_X1 U14135 ( .A1(n11223), .A2(n11044), .ZN(n11046) );
  AOI22_X1 U14136 ( .A1(n11250), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n11018), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11045) );
  AOI22_X1 U14137 ( .A1(n11251), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n11250), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n11050) );
  AOI22_X1 U14138 ( .A1(n11223), .A2(n11048), .B1(n11018), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11049) );
  NAND2_X1 U14139 ( .A1(n11050), .A2(n11049), .ZN(n13864) );
  NAND2_X1 U14140 ( .A1(n11223), .A2(n11051), .ZN(n11052) );
  INV_X1 U14141 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19801) );
  AOI22_X1 U14142 ( .A1(n11250), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n11018), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11053) );
  OAI21_X1 U14143 ( .B1(n11249), .B2(n19801), .A(n11053), .ZN(n11054) );
  INV_X1 U14144 ( .A(n11054), .ZN(n15331) );
  INV_X1 U14145 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19185) );
  INV_X1 U14146 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19803) );
  OAI222_X1 U14147 ( .A1(n16326), .A2(n11196), .B1(n11198), .B2(n19185), .C1(
        n11249), .C2(n19803), .ZN(n15323) );
  NAND2_X1 U14148 ( .A1(n11251), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11073) );
  INV_X1 U14149 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13649) );
  NAND2_X1 U14150 ( .A1(n10500), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11059) );
  NAND2_X1 U14151 ( .A1(n10413), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11058) );
  AOI22_X1 U14152 ( .A1(n11141), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11099), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11057) );
  NAND2_X1 U14153 ( .A1(n10414), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11056) );
  AND4_X1 U14154 ( .A1(n11059), .A2(n11058), .A3(n11057), .A4(n11056), .ZN(
        n11061) );
  NAND2_X1 U14155 ( .A1(n10467), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11060) );
  OAI211_X1 U14156 ( .C1(n13649), .C2(n11202), .A(n11061), .B(n11060), .ZN(
        n11062) );
  INV_X1 U14157 ( .A(n11062), .ZN(n11070) );
  NAND2_X1 U14158 ( .A1(n10456), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11066) );
  AOI22_X1 U14159 ( .A1(n10462), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10400), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11065) );
  NAND2_X1 U14160 ( .A1(n12706), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11064) );
  NAND2_X1 U14161 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11063) );
  AOI22_X1 U14162 ( .A1(n12695), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10401), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11069) );
  AOI22_X1 U14163 ( .A1(n11067), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10395), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11068) );
  INV_X1 U14164 ( .A(n13582), .ZN(n13584) );
  NAND2_X1 U14165 ( .A1(n11223), .A2(n13584), .ZN(n11072) );
  AOI22_X1 U14166 ( .A1(n11250), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n11018), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11071) );
  INV_X1 U14167 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11075) );
  INV_X1 U14168 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11074) );
  OAI22_X1 U14169 ( .A1(n12689), .A2(n11075), .B1(n12654), .B2(n11074), .ZN(
        n11079) );
  INV_X1 U14170 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12544) );
  NAND2_X1 U14171 ( .A1(n10462), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11077) );
  NAND2_X1 U14172 ( .A1(n10413), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11076) );
  OAI211_X1 U14173 ( .C1(n15402), .C2(n12544), .A(n11077), .B(n11076), .ZN(
        n11078) );
  NOR2_X1 U14174 ( .A1(n11079), .A2(n11078), .ZN(n11090) );
  NAND2_X1 U14175 ( .A1(n10467), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11086) );
  NAND2_X1 U14176 ( .A1(n12695), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11085) );
  AOI22_X1 U14177 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10400), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11084) );
  INV_X1 U14178 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11081) );
  NAND2_X1 U14179 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n11099), .ZN(
        n11080) );
  OAI21_X1 U14180 ( .B1(n12699), .B2(n11081), .A(n11080), .ZN(n11082) );
  AOI21_X1 U14181 ( .B1(n10500), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A(
        n11082), .ZN(n11083) );
  AND4_X1 U14182 ( .A1(n11086), .A2(n11085), .A3(n11084), .A4(n11083), .ZN(
        n11089) );
  AOI22_X1 U14183 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10395), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11088) );
  AOI22_X1 U14184 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10456), .B1(
        n10401), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11087) );
  NAND4_X1 U14185 ( .A1(n11090), .A2(n11089), .A3(n11088), .A4(n11087), .ZN(
        n13588) );
  AOI22_X1 U14186 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n11251), .B1(n11223), 
        .B2(n13588), .ZN(n11092) );
  AOI22_X1 U14187 ( .A1(n11250), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n11018), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11091) );
  NAND2_X1 U14188 ( .A1(n11092), .A2(n11091), .ZN(n15310) );
  NAND2_X1 U14189 ( .A1(n14809), .A2(n15310), .ZN(n14790) );
  INV_X1 U14190 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11094) );
  INV_X1 U14191 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11093) );
  OAI22_X1 U14192 ( .A1(n12689), .A2(n11094), .B1(n12654), .B2(n11093), .ZN(
        n11098) );
  INV_X1 U14193 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12583) );
  NAND2_X1 U14194 ( .A1(n10462), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11096) );
  NAND2_X1 U14195 ( .A1(n10413), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11095) );
  OAI211_X1 U14196 ( .C1(n15402), .C2(n12583), .A(n11096), .B(n11095), .ZN(
        n11097) );
  NOR2_X1 U14197 ( .A1(n11098), .A2(n11097), .ZN(n11110) );
  NAND2_X1 U14198 ( .A1(n12695), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n11106) );
  NAND2_X1 U14199 ( .A1(n10401), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11105) );
  AOI22_X1 U14200 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10400), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11104) );
  INV_X1 U14201 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11101) );
  NAND2_X1 U14202 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n11099), .ZN(
        n11100) );
  OAI21_X1 U14203 ( .B1(n12699), .B2(n11101), .A(n11100), .ZN(n11102) );
  AOI21_X1 U14204 ( .B1(n10500), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A(
        n11102), .ZN(n11103) );
  AND4_X1 U14205 ( .A1(n11106), .A2(n11105), .A3(n11104), .A4(n11103), .ZN(
        n11109) );
  AOI22_X1 U14206 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10467), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11108) );
  AOI22_X1 U14207 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n10456), .B1(
        n10395), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11107) );
  NAND4_X1 U14208 ( .A1(n11110), .A2(n11109), .A3(n11108), .A4(n11107), .ZN(
        n13661) );
  AOI22_X1 U14209 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n11251), .B1(n11223), 
        .B2(n13661), .ZN(n11112) );
  AOI22_X1 U14210 ( .A1(n11250), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n11018), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11111) );
  INV_X1 U14211 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11113) );
  OAI22_X1 U14212 ( .A1(n12689), .A2(n11114), .B1(n12654), .B2(n11113), .ZN(
        n11118) );
  INV_X1 U14213 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12601) );
  NAND2_X1 U14214 ( .A1(n10462), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11116) );
  NAND2_X1 U14215 ( .A1(n10413), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11115) );
  OAI211_X1 U14216 ( .C1(n15402), .C2(n12601), .A(n11116), .B(n11115), .ZN(
        n11117) );
  NOR2_X1 U14217 ( .A1(n11118), .A2(n11117), .ZN(n11129) );
  NAND2_X1 U14218 ( .A1(n10467), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n11125) );
  NAND2_X1 U14219 ( .A1(n12695), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11124) );
  AOI22_X1 U14220 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10400), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11123) );
  INV_X1 U14221 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11120) );
  NAND2_X1 U14222 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n12696), .ZN(
        n11119) );
  OAI21_X1 U14223 ( .B1(n12699), .B2(n11120), .A(n11119), .ZN(n11121) );
  AOI21_X1 U14224 ( .B1(n10500), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A(
        n11121), .ZN(n11122) );
  AND4_X1 U14225 ( .A1(n11125), .A2(n11124), .A3(n11123), .A4(n11122), .ZN(
        n11128) );
  AOI22_X1 U14226 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10395), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11127) );
  AOI22_X1 U14227 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n10456), .B1(
        n10401), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11126) );
  NAND4_X1 U14228 ( .A1(n11129), .A2(n11128), .A3(n11127), .A4(n11126), .ZN(
        n13699) );
  NAND2_X1 U14229 ( .A1(n11223), .A2(n13699), .ZN(n11131) );
  AOI22_X1 U14230 ( .A1(n11250), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n11018), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11130) );
  OAI211_X1 U14231 ( .C1(n15101), .C2(n11249), .A(n11131), .B(n11130), .ZN(
        n15287) );
  NAND2_X1 U14232 ( .A1(n14791), .A2(n15287), .ZN(n14780) );
  NAND2_X1 U14233 ( .A1(n11251), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11154) );
  OR2_X1 U14234 ( .A1(n12689), .A2(n11132), .ZN(n11136) );
  AOI22_X1 U14235 ( .A1(n10462), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10413), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11135) );
  NAND2_X1 U14236 ( .A1(n10456), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11134) );
  NAND2_X1 U14237 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11133) );
  NAND2_X1 U14238 ( .A1(n10467), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11140) );
  NAND2_X1 U14239 ( .A1(n12695), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11139) );
  NAND2_X1 U14240 ( .A1(n10401), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11138) );
  NAND2_X1 U14241 ( .A1(n12706), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11137) );
  AND4_X1 U14242 ( .A1(n11140), .A2(n11139), .A3(n11138), .A4(n11137), .ZN(
        n11151) );
  INV_X1 U14243 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11148) );
  NAND2_X1 U14244 ( .A1(n10500), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11145) );
  NAND2_X1 U14245 ( .A1(n10414), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11144) );
  NAND2_X1 U14246 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11143) );
  AOI22_X1 U14247 ( .A1(n11141), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n12696), .ZN(n11142) );
  AND4_X1 U14248 ( .A1(n11145), .A2(n11144), .A3(n11143), .A4(n11142), .ZN(
        n11147) );
  NAND2_X1 U14249 ( .A1(n10395), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11146) );
  OAI211_X1 U14250 ( .C1(n11202), .C2(n11148), .A(n11147), .B(n11146), .ZN(
        n11149) );
  INV_X1 U14251 ( .A(n11149), .ZN(n11150) );
  INV_X1 U14252 ( .A(n13782), .ZN(n13784) );
  NAND2_X1 U14253 ( .A1(n11223), .A2(n13784), .ZN(n11153) );
  AOI22_X1 U14254 ( .A1(n11250), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n11018), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11152) );
  INV_X1 U14255 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11155) );
  OR2_X1 U14256 ( .A1(n11202), .A2(n11155), .ZN(n11159) );
  NAND2_X1 U14257 ( .A1(n10395), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11158) );
  NAND2_X1 U14258 ( .A1(n10456), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11157) );
  NAND2_X1 U14259 ( .A1(n10401), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11156) );
  AND4_X1 U14260 ( .A1(n11159), .A2(n11158), .A3(n11157), .A4(n11156), .ZN(
        n11174) );
  INV_X1 U14261 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11160) );
  OAI22_X1 U14262 ( .A1(n12689), .A2(n11161), .B1(n12654), .B2(n11160), .ZN(
        n11165) );
  INV_X1 U14263 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12636) );
  NAND2_X1 U14264 ( .A1(n10462), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11163) );
  NAND2_X1 U14265 ( .A1(n10413), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11162) );
  OAI211_X1 U14266 ( .C1(n12636), .C2(n15402), .A(n11163), .B(n11162), .ZN(
        n11164) );
  NOR2_X1 U14267 ( .A1(n11165), .A2(n11164), .ZN(n11173) );
  NAND2_X1 U14268 ( .A1(n10467), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11172) );
  NAND2_X1 U14269 ( .A1(n12695), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11171) );
  AOI22_X1 U14270 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11170) );
  INV_X1 U14271 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11167) );
  NAND2_X1 U14272 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n12696), .ZN(
        n11166) );
  OAI21_X1 U14273 ( .B1(n12699), .B2(n11167), .A(n11166), .ZN(n11168) );
  AOI21_X1 U14274 ( .B1(n10500), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A(
        n11168), .ZN(n11169) );
  AND3_X1 U14275 ( .A1(n11174), .A2(n11173), .A3(n10125), .ZN(n13882) );
  NAND2_X1 U14276 ( .A1(n11251), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11176) );
  AOI22_X1 U14277 ( .A1(n11250), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n11018), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11175) );
  OAI211_X1 U14278 ( .C1(n13882), .C2(n11195), .A(n11176), .B(n11175), .ZN(
        n14767) );
  INV_X1 U14279 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11177) );
  OAI22_X1 U14280 ( .A1(n12689), .A2(n11178), .B1(n12654), .B2(n11177), .ZN(
        n11182) );
  INV_X1 U14281 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12655) );
  NAND2_X1 U14282 ( .A1(n10462), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11180) );
  NAND2_X1 U14283 ( .A1(n10413), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11179) );
  OAI211_X1 U14284 ( .C1(n15402), .C2(n12655), .A(n11180), .B(n11179), .ZN(
        n11181) );
  NOR2_X1 U14285 ( .A1(n11182), .A2(n11181), .ZN(n11193) );
  NAND2_X1 U14286 ( .A1(n10467), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11189) );
  NAND2_X1 U14287 ( .A1(n12695), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11188) );
  AOI22_X1 U14288 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10400), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11187) );
  INV_X1 U14289 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11184) );
  NAND2_X1 U14290 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n12696), .ZN(
        n11183) );
  OAI21_X1 U14291 ( .B1(n12699), .B2(n11184), .A(n11183), .ZN(n11185) );
  AOI21_X1 U14292 ( .B1(n10500), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A(
        n11185), .ZN(n11186) );
  AND4_X1 U14293 ( .A1(n11189), .A2(n11188), .A3(n11187), .A4(n11186), .ZN(
        n11192) );
  INV_X1 U14294 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n20880) );
  AOI22_X1 U14295 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10395), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11191) );
  AOI22_X1 U14296 ( .A1(n10456), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10401), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11190) );
  NAND4_X1 U14297 ( .A1(n11193), .A2(n11192), .A3(n11191), .A4(n11190), .ZN(
        n13829) );
  INV_X1 U14298 ( .A(n13829), .ZN(n11194) );
  NOR2_X1 U14299 ( .A1(n11195), .A2(n11194), .ZN(n11200) );
  INV_X1 U14300 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n11197) );
  OAI22_X1 U14301 ( .A1(n11198), .A2(n11197), .B1(n11196), .B2(n16233), .ZN(
        n11199) );
  AOI211_X1 U14302 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n11251), .A(n11200), 
        .B(n11199), .ZN(n14754) );
  AOI22_X1 U14303 ( .A1(n11251), .A2(P2_REIP_REG_15__SCAN_IN), .B1(n11018), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11225) );
  INV_X1 U14304 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11201) );
  OR2_X1 U14305 ( .A1(n11202), .A2(n11201), .ZN(n11206) );
  NAND2_X1 U14306 ( .A1(n10395), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11205) );
  NAND2_X1 U14307 ( .A1(n10456), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11204) );
  NAND2_X1 U14308 ( .A1(n10401), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11203) );
  AND4_X1 U14309 ( .A1(n11206), .A2(n11205), .A3(n11204), .A4(n11203), .ZN(
        n11222) );
  INV_X1 U14310 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11208) );
  INV_X1 U14311 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11207) );
  OAI22_X1 U14312 ( .A1(n12689), .A2(n11208), .B1(n12654), .B2(n11207), .ZN(
        n11212) );
  INV_X1 U14313 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12688) );
  NAND2_X1 U14314 ( .A1(n10462), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11210) );
  NAND2_X1 U14315 ( .A1(n10413), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11209) );
  OAI211_X1 U14316 ( .C1(n15402), .C2(n12688), .A(n11210), .B(n11209), .ZN(
        n11211) );
  NOR2_X1 U14317 ( .A1(n11212), .A2(n11211), .ZN(n11221) );
  NAND2_X1 U14318 ( .A1(n10467), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11219) );
  NAND2_X1 U14319 ( .A1(n12695), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11218) );
  AOI22_X1 U14320 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10400), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11217) );
  INV_X1 U14321 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11214) );
  NAND2_X1 U14322 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n12696), .ZN(
        n11213) );
  OAI21_X1 U14323 ( .B1(n12699), .B2(n11214), .A(n11213), .ZN(n11215) );
  AOI21_X1 U14324 ( .B1(n10500), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A(
        n11215), .ZN(n11216) );
  AND4_X1 U14325 ( .A1(n11219), .A2(n11218), .A3(n11217), .A4(n11216), .ZN(
        n11220) );
  NAND3_X1 U14326 ( .A1(n11222), .A2(n11221), .A3(n11220), .ZN(n13707) );
  AOI22_X1 U14327 ( .A1(n11223), .A2(n13707), .B1(P2_EAX_REG_15__SCAN_IN), 
        .B2(n11250), .ZN(n11224) );
  NAND2_X1 U14328 ( .A1(n11225), .A2(n11224), .ZN(n15267) );
  NAND2_X1 U14329 ( .A1(n11251), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11227) );
  AOI22_X1 U14330 ( .A1(n11250), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n11018), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11226) );
  INV_X1 U14331 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19818) );
  AOI22_X1 U14332 ( .A1(n11250), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n11018), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11228) );
  OAI21_X1 U14333 ( .B1(n11249), .B2(n19818), .A(n11228), .ZN(n13887) );
  NAND2_X1 U14334 ( .A1(n13886), .A2(n13887), .ZN(n13888) );
  NAND2_X1 U14335 ( .A1(n11251), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11230) );
  AOI22_X1 U14336 ( .A1(n11250), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n11018), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11229) );
  AOI22_X1 U14337 ( .A1(n11250), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n11018), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11231) );
  OAI21_X1 U14338 ( .B1(n11249), .B2(n10873), .A(n11231), .ZN(n14971) );
  NAND2_X1 U14339 ( .A1(n11251), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11233) );
  AOI22_X1 U14340 ( .A1(n11250), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n11018), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11232) );
  INV_X1 U14341 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19823) );
  AOI22_X1 U14342 ( .A1(n11250), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n11018), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11234) );
  OAI21_X1 U14343 ( .B1(n11249), .B2(n19823), .A(n11234), .ZN(n14741) );
  INV_X1 U14344 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n11236) );
  AOI22_X1 U14345 ( .A1(n11250), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n11018), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11235) );
  OAI21_X1 U14346 ( .B1(n11249), .B2(n11236), .A(n11235), .ZN(n15195) );
  NAND2_X1 U14347 ( .A1(n14742), .A2(n15195), .ZN(n14956) );
  INV_X1 U14348 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19825) );
  AOI22_X1 U14349 ( .A1(n11250), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n11018), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11237) );
  OAI21_X1 U14350 ( .B1(n11249), .B2(n19825), .A(n11237), .ZN(n11238) );
  INV_X1 U14351 ( .A(n11238), .ZN(n14957) );
  OR2_X2 U14352 ( .A1(n14956), .A2(n14957), .ZN(n14949) );
  INV_X1 U14353 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n11240) );
  AOI22_X1 U14354 ( .A1(n11250), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n11018), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11239) );
  OAI21_X1 U14355 ( .B1(n11249), .B2(n11240), .A(n11239), .ZN(n11241) );
  INV_X1 U14356 ( .A(n11241), .ZN(n14948) );
  NOR2_X4 U14357 ( .A1(n14949), .A2(n14948), .ZN(n14950) );
  INV_X1 U14358 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n21016) );
  AOI22_X1 U14359 ( .A1(n11250), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n11018), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11242) );
  OAI21_X1 U14360 ( .B1(n11249), .B2(n21016), .A(n11242), .ZN(n13947) );
  INV_X1 U14361 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n15000) );
  AOI22_X1 U14362 ( .A1(n11250), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n11018), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11243) );
  OAI21_X1 U14363 ( .B1(n11249), .B2(n15000), .A(n11243), .ZN(n14934) );
  INV_X1 U14364 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19831) );
  AOI22_X1 U14365 ( .A1(n11250), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n11018), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11244) );
  OAI21_X1 U14366 ( .B1(n11249), .B2(n19831), .A(n11244), .ZN(n11245) );
  INV_X1 U14367 ( .A(n11245), .ZN(n14926) );
  INV_X1 U14368 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n12478) );
  AOI22_X1 U14369 ( .A1(n11250), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n11018), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11246) );
  OAI21_X1 U14370 ( .B1(n11249), .B2(n12478), .A(n11246), .ZN(n11247) );
  INV_X1 U14371 ( .A(n11247), .ZN(n12477) );
  INV_X1 U14372 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19833) );
  AOI22_X1 U14373 ( .A1(n11250), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n11018), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11248) );
  OAI21_X1 U14374 ( .B1(n11249), .B2(n19833), .A(n11248), .ZN(n14913) );
  NAND2_X1 U14375 ( .A1(n14914), .A2(n14913), .ZN(n12879) );
  AOI222_X1 U14376 ( .A1(n11251), .A2(P2_REIP_REG_30__SCAN_IN), .B1(n11250), 
        .B2(P2_EAX_REG_30__SCAN_IN), .C1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), 
        .C2(n11018), .ZN(n12881) );
  NOR2_X2 U14377 ( .A1(n12879), .A2(n12881), .ZN(n12880) );
  AOI222_X1 U14378 ( .A1(n11251), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n11250), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n11018), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11252) );
  XNOR2_X1 U14379 ( .A(n12880), .B(n11252), .ZN(n16116) );
  AND2_X1 U14380 ( .A1(n9790), .A2(n11255), .ZN(n11256) );
  NAND2_X1 U14381 ( .A1(n11254), .A2(n11256), .ZN(n13071) );
  OAI21_X1 U14382 ( .B1(n11253), .B2(n9788), .A(n13071), .ZN(n11257) );
  INV_X1 U14383 ( .A(n14067), .ZN(n11275) );
  INV_X1 U14384 ( .A(n11258), .ZN(n11274) );
  NOR2_X1 U14385 ( .A1(n11259), .A2(n19030), .ZN(n19216) );
  INV_X1 U14386 ( .A(n19216), .ZN(n13214) );
  NAND2_X1 U14387 ( .A1(n15321), .A2(n13214), .ZN(n15292) );
  INV_X1 U14388 ( .A(n11260), .ZN(n15175) );
  AOI21_X1 U14389 ( .B1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n19221), .A(
        n19213), .ZN(n11261) );
  NOR2_X1 U14390 ( .A1(n19216), .A2(n11261), .ZN(n13628) );
  OAI221_X1 U14391 ( .B1(n15321), .B2(n11263), .C1(n15321), .C2(n11262), .A(
        n13628), .ZN(n16293) );
  NAND2_X1 U14392 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n11264), .ZN(
        n11265) );
  OAI21_X1 U14393 ( .B1(n11265), .B2(n16233), .A(n16294), .ZN(n11266) );
  INV_X1 U14394 ( .A(n11266), .ZN(n11267) );
  OR2_X1 U14395 ( .A1(n16293), .A2(n11267), .ZN(n15270) );
  NAND2_X1 U14396 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n11268), .ZN(
        n11269) );
  AND2_X1 U14397 ( .A1(n16294), .A2(n11269), .ZN(n11270) );
  NOR2_X1 U14398 ( .A1(n15270), .A2(n11270), .ZN(n15231) );
  INV_X1 U14399 ( .A(n15292), .ZN(n11271) );
  OR2_X1 U14400 ( .A1(n11272), .A2(n11271), .ZN(n11273) );
  OAI21_X1 U14401 ( .B1(n15321), .B2(n15175), .A(n15203), .ZN(n15166) );
  AOI21_X1 U14402 ( .B1(n11274), .B2(n15292), .A(n15166), .ZN(n15145) );
  OAI21_X1 U14403 ( .B1(n11275), .B2(n15321), .A(n15145), .ZN(n14069) );
  NOR2_X1 U14404 ( .A1(n15321), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11276) );
  OAI21_X1 U14405 ( .B1(n14069), .B2(n11276), .A(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11278) );
  INV_X1 U14406 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19838) );
  NOR2_X1 U14407 ( .A1(n18957), .A2(n19838), .ZN(n14059) );
  AND2_X1 U14408 ( .A1(n11278), .A2(n11277), .ZN(n11279) );
  AOI211_X1 U14409 ( .C1(n14064), .C2(n19233), .A(n11282), .B(n11281), .ZN(
        n11283) );
  OAI21_X1 U14410 ( .B1(n14066), .B2(n19225), .A(n11283), .ZN(P2_U3015) );
  NAND2_X1 U14411 ( .A1(n15225), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15035) );
  NAND2_X1 U14412 ( .A1(n15035), .A2(n12500), .ZN(n11287) );
  OAI21_X1 U14413 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n9844), .A(
        n14684), .ZN(n11288) );
  INV_X1 U14414 ( .A(n11288), .ZN(n18923) );
  NAND2_X1 U14415 ( .A1(n18923), .A2(n19203), .ZN(n11290) );
  INV_X1 U14416 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n11289) );
  OR2_X1 U14417 ( .A1(n18957), .A2(n11289), .ZN(n12502) );
  OAI211_X1 U14418 ( .C1(n19212), .C2(n10068), .A(n11290), .B(n12502), .ZN(
        n11291) );
  AOI21_X1 U14419 ( .B1(n12506), .B2(n19204), .A(n11291), .ZN(n11309) );
  OR2_X1 U14420 ( .A1(n11294), .A2(n11293), .ZN(n11295) );
  NAND2_X1 U14421 ( .A1(n11292), .A2(n11295), .ZN(n18924) );
  OR2_X1 U14422 ( .A1(n18924), .A2(n13644), .ZN(n11308) );
  INV_X1 U14423 ( .A(n11297), .ZN(n11298) );
  OAI21_X2 U14424 ( .B1(n15077), .B2(n11298), .A(n15078), .ZN(n16232) );
  INV_X1 U14425 ( .A(n16230), .ZN(n11299) );
  INV_X1 U14426 ( .A(n15050), .ZN(n11300) );
  OAI21_X1 U14427 ( .B1(n15038), .B2(n11303), .A(n11302), .ZN(n15025) );
  INV_X1 U14428 ( .A(n15024), .ZN(n11304) );
  INV_X1 U14429 ( .A(n12496), .ZN(n11306) );
  NAND3_X1 U14430 ( .A1(n11309), .A2(n11308), .A3(n11307), .ZN(P2_U2994) );
  NOR2_X2 U14431 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11310), .ZN(
        n11318) );
  NOR2_X4 U14432 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13411) );
  AOI22_X1 U14433 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11371), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11317) );
  AND2_X2 U14434 ( .A1(n11320), .A2(n13411), .ZN(n11496) );
  AOI22_X1 U14435 ( .A1(n11496), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9785), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11316) );
  AOI22_X1 U14436 ( .A1(n11438), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11501), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11315) );
  AOI22_X1 U14437 ( .A1(n11379), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9747), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11314) );
  AND2_X4 U14438 ( .A1(n11320), .A2(n13393), .ZN(n12318) );
  AND2_X2 U14439 ( .A1(n11318), .A2(n13393), .ZN(n11372) );
  AOI22_X1 U14440 ( .A1(n12318), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11372), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11325) );
  AOI22_X1 U14441 ( .A1(n12266), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12096), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11324) );
  AND2_X2 U14442 ( .A1(n11318), .A2(n11319), .ZN(n11533) );
  AOI22_X1 U14443 ( .A1(n11533), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11380), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11323) );
  AND2_X2 U14444 ( .A1(n11321), .A2(n13392), .ZN(n11528) );
  AOI22_X1 U14445 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11528), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11322) );
  INV_X2 U14446 ( .A(n20160), .ZN(n11472) );
  NAND2_X1 U14447 ( .A1(n11496), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11331) );
  NAND2_X1 U14448 ( .A1(n11438), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11330) );
  NAND2_X1 U14449 ( .A1(n9785), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11329) );
  NAND2_X1 U14450 ( .A1(n11501), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11328) );
  NAND2_X1 U14451 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11335) );
  NAND2_X1 U14452 ( .A1(n12318), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11334) );
  NAND2_X1 U14453 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11333) );
  NAND2_X1 U14454 ( .A1(n11528), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11332) );
  NAND2_X1 U14455 ( .A1(n11533), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n11339) );
  NAND2_X1 U14456 ( .A1(n11371), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n11338) );
  NAND2_X1 U14457 ( .A1(n12266), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11337) );
  NAND2_X1 U14458 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11336) );
  NAND2_X1 U14459 ( .A1(n11372), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n11343) );
  NAND2_X1 U14460 ( .A1(n11379), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n11342) );
  NAND2_X1 U14461 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11341) );
  NAND2_X1 U14462 ( .A1(n11380), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11340) );
  NAND2_X1 U14463 ( .A1(n11533), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11351) );
  NAND2_X1 U14464 ( .A1(n11372), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11350) );
  NAND2_X1 U14465 ( .A1(n11379), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11349) );
  NAND2_X1 U14466 ( .A1(n11380), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11348) );
  NAND2_X1 U14467 ( .A1(n11501), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11355) );
  NAND2_X1 U14468 ( .A1(n11496), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11354) );
  NAND2_X1 U14469 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11353) );
  NAND2_X1 U14470 ( .A1(n11438), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11352) );
  NAND2_X1 U14471 ( .A1(n12318), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11359) );
  NAND2_X1 U14472 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11358) );
  NAND2_X1 U14473 ( .A1(n11371), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11357) );
  NAND2_X1 U14474 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11356) );
  NAND2_X1 U14475 ( .A1(n12266), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11363) );
  NAND2_X1 U14476 ( .A1(n11528), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11362) );
  NAND2_X1 U14477 ( .A1(n9785), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11361) );
  NAND2_X1 U14478 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11360) );
  NAND4_X2 U14479 ( .A1(n11366), .A2(n10143), .A3(n11365), .A4(n11364), .ZN(
        n11455) );
  AOI22_X1 U14480 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11496), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11370) );
  AOI22_X1 U14481 ( .A1(n11528), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9785), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11369) );
  AOI22_X1 U14482 ( .A1(n11438), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9772), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11367) );
  NAND4_X1 U14483 ( .A1(n11370), .A2(n11369), .A3(n11368), .A4(n11367), .ZN(
        n11378) );
  AOI22_X1 U14484 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11371), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11376) );
  AOI22_X1 U14485 ( .A1(n11533), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11379), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11375) );
  AOI22_X1 U14486 ( .A1(n11372), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11380), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11374) );
  AOI22_X1 U14487 ( .A1(n12318), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9747), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11373) );
  NAND4_X1 U14488 ( .A1(n11376), .A2(n11375), .A3(n11374), .A4(n11373), .ZN(
        n11377) );
  INV_X1 U14489 ( .A(n11451), .ZN(n11391) );
  AOI22_X1 U14490 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11371), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11384) );
  AOI22_X1 U14491 ( .A1(n11533), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11379), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11383) );
  AOI22_X1 U14492 ( .A1(n11372), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11380), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11382) );
  AOI22_X1 U14493 ( .A1(n12318), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9747), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11381) );
  NAND4_X1 U14494 ( .A1(n11384), .A2(n11383), .A3(n11382), .A4(n11381), .ZN(
        n11390) );
  AOI22_X1 U14495 ( .A1(n12266), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12096), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11388) );
  AOI22_X1 U14496 ( .A1(n11528), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11417), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11387) );
  AOI22_X1 U14497 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11496), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11386) );
  AOI22_X1 U14498 ( .A1(n11438), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9757), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11385) );
  NAND4_X1 U14499 ( .A1(n11388), .A2(n11387), .A3(n11386), .A4(n11385), .ZN(
        n11389) );
  NAND2_X1 U14500 ( .A1(n11391), .A2(n20145), .ZN(n11659) );
  INV_X1 U14501 ( .A(n11659), .ZN(n11392) );
  NAND2_X1 U14502 ( .A1(n11393), .A2(n11392), .ZN(n13144) );
  AOI22_X1 U14503 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11371), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11397) );
  AOI22_X1 U14504 ( .A1(n11533), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11379), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11396) );
  AOI22_X1 U14505 ( .A1(n11372), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11380), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11395) );
  AOI22_X1 U14506 ( .A1(n12318), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9747), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11394) );
  NAND4_X1 U14507 ( .A1(n11397), .A2(n11396), .A3(n11395), .A4(n11394), .ZN(
        n11403) );
  AOI22_X1 U14508 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11496), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11401) );
  AOI22_X1 U14509 ( .A1(n11438), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11501), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11400) );
  AOI22_X1 U14510 ( .A1(n11528), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11417), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11399) );
  AOI22_X1 U14511 ( .A1(n12266), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12096), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11398) );
  NAND4_X1 U14512 ( .A1(n11401), .A2(n11400), .A3(n11399), .A4(n11398), .ZN(
        n11402) );
  NAND2_X1 U14513 ( .A1(n11533), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11407) );
  NAND2_X1 U14514 ( .A1(n11372), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11406) );
  NAND2_X1 U14515 ( .A1(n11379), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11405) );
  NAND2_X1 U14516 ( .A1(n11380), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11404) );
  NAND2_X1 U14517 ( .A1(n12318), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11411) );
  NAND2_X1 U14518 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11410) );
  NAND2_X1 U14519 ( .A1(n11371), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11409) );
  NAND2_X1 U14520 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11408) );
  NAND2_X1 U14521 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11416) );
  NAND2_X1 U14522 ( .A1(n11496), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11415) );
  NAND2_X1 U14523 ( .A1(n11501), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11414) );
  NAND2_X1 U14524 ( .A1(n11438), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11413) );
  NAND2_X1 U14525 ( .A1(n12266), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11421) );
  NAND2_X1 U14526 ( .A1(n11528), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11420) );
  NAND2_X1 U14527 ( .A1(n9785), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11419) );
  NAND2_X1 U14528 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11418) );
  NAND4_X4 U14529 ( .A1(n11425), .A2(n11424), .A3(n11423), .A4(n11422), .ZN(
        n11464) );
  NAND2_X1 U14530 ( .A1(n13175), .A2(n11464), .ZN(n13157) );
  NAND2_X1 U14531 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20750) );
  OAI21_X1 U14532 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(P1_STATE_REG_2__SCAN_IN), 
        .A(n20750), .ZN(n13141) );
  NAND2_X1 U14533 ( .A1(n11472), .A2(n9786), .ZN(n12354) );
  INV_X1 U14534 ( .A(n12354), .ZN(n11447) );
  NAND2_X1 U14535 ( .A1(n11533), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11429) );
  NAND2_X1 U14536 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11428) );
  NAND2_X1 U14537 ( .A1(n11379), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11427) );
  NAND2_X1 U14538 ( .A1(n11380), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11426) );
  NAND2_X1 U14539 ( .A1(n11371), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11433) );
  NAND2_X1 U14540 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11432) );
  NAND2_X1 U14541 ( .A1(n12266), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11431) );
  NAND2_X1 U14542 ( .A1(n9785), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11430) );
  NAND2_X1 U14543 ( .A1(n12318), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11437) );
  NAND2_X1 U14544 ( .A1(n11372), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11436) );
  NAND2_X1 U14545 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11435) );
  NAND2_X1 U14546 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11434) );
  NAND2_X1 U14547 ( .A1(n11496), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11442) );
  NAND2_X1 U14548 ( .A1(n11528), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11441) );
  NAND2_X1 U14549 ( .A1(n11438), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11440) );
  NAND2_X1 U14550 ( .A1(n11501), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11439) );
  NAND4_X4 U14551 ( .A1(n11446), .A2(n11445), .A3(n11444), .A4(n11443), .ZN(
        n12355) );
  NAND2_X1 U14552 ( .A1(n11447), .A2(n13677), .ZN(n13193) );
  INV_X1 U14553 ( .A(n13193), .ZN(n11448) );
  INV_X1 U14554 ( .A(n11461), .ZN(n11450) );
  NAND2_X1 U14555 ( .A1(n11450), .A2(n20136), .ZN(n11454) );
  NAND2_X1 U14556 ( .A1(n11454), .A2(n11453), .ZN(n11460) );
  NAND2_X1 U14557 ( .A1(n11481), .A2(n12352), .ZN(n11476) );
  NAND2_X1 U14558 ( .A1(n11476), .A2(n20145), .ZN(n11459) );
  OAI21_X1 U14559 ( .B1(n20152), .B2(n11473), .A(n11456), .ZN(n11457) );
  NAND3_X1 U14560 ( .A1(n11460), .A2(n11459), .A3(n11458), .ZN(n11468) );
  INV_X1 U14561 ( .A(n11468), .ZN(n11463) );
  NOR2_X1 U14562 ( .A1(n11466), .A2(n11464), .ZN(n11462) );
  NAND2_X1 U14563 ( .A1(n11463), .A2(n11462), .ZN(n13148) );
  INV_X1 U14564 ( .A(n11464), .ZN(n13183) );
  NAND2_X1 U14565 ( .A1(n11822), .A2(n12448), .ZN(n11467) );
  OAI211_X1 U14566 ( .C1(n13244), .C2(n20842), .A(n11467), .B(n13685), .ZN(
        n11471) );
  NAND2_X1 U14567 ( .A1(n11468), .A2(n13183), .ZN(n11470) );
  NAND2_X1 U14568 ( .A1(n11464), .A2(n20136), .ZN(n11469) );
  NAND2_X1 U14569 ( .A1(n11470), .A2(n11469), .ZN(n13198) );
  NAND2_X1 U14570 ( .A1(n11472), .A2(n11473), .ZN(n11474) );
  NAND2_X1 U14571 ( .A1(n11820), .A2(n13244), .ZN(n11480) );
  AOI21_X1 U14572 ( .B1(n11480), .B2(n14652), .A(n9786), .ZN(n11478) );
  MUX2_X1 U14573 ( .A(n20835), .B(n15747), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n11479) );
  AND2_X1 U14574 ( .A1(n14652), .A2(n12355), .ZN(n11491) );
  INV_X1 U14575 ( .A(n13677), .ZN(n11776) );
  AND2_X1 U14576 ( .A1(n11776), .A2(n9787), .ZN(n13162) );
  INV_X1 U14577 ( .A(n11481), .ZN(n11482) );
  NAND2_X1 U14578 ( .A1(n11482), .A2(n20145), .ZN(n11483) );
  NAND2_X1 U14579 ( .A1(n13162), .A2(n11483), .ZN(n11489) );
  INV_X1 U14580 ( .A(n11484), .ZN(n20822) );
  NOR2_X1 U14581 ( .A1(n20822), .A2(n11495), .ZN(n11488) );
  NAND2_X1 U14582 ( .A1(n9786), .A2(n12350), .ZN(n13251) );
  INV_X1 U14583 ( .A(n11485), .ZN(n11486) );
  NAND2_X1 U14584 ( .A1(n11486), .A2(n15742), .ZN(n11487) );
  NAND4_X1 U14585 ( .A1(n11489), .A2(n11488), .A3(n13251), .A4(n11487), .ZN(
        n11490) );
  AOI21_X1 U14586 ( .B1(n11480), .B2(n11491), .A(n11490), .ZN(n11492) );
  NAND2_X1 U14587 ( .A1(n11493), .A2(n11492), .ZN(n11550) );
  INV_X1 U14588 ( .A(n11550), .ZN(n11494) );
  XNOR2_X1 U14589 ( .A(n11551), .B(n11494), .ZN(n11848) );
  NAND2_X1 U14590 ( .A1(n11848), .A2(n11495), .ZN(n11520) );
  AOI22_X1 U14591 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12299), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11500) );
  AOI22_X1 U14592 ( .A1(n12318), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12329), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11499) );
  AOI22_X1 U14593 ( .A1(n12325), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12328), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11498) );
  AOI22_X1 U14594 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12317), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11497) );
  NAND4_X1 U14595 ( .A1(n11500), .A2(n11499), .A3(n11498), .A4(n11497), .ZN(
        n11507) );
  AOI22_X1 U14596 ( .A1(n12323), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11505) );
  AOI22_X1 U14597 ( .A1(n12266), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12327), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11504) );
  AOI22_X1 U14598 ( .A1(n12144), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11503) );
  AOI22_X1 U14599 ( .A1(n12326), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11501), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11502) );
  NAND4_X1 U14600 ( .A1(n11505), .A2(n11504), .A3(n11503), .A4(n11502), .ZN(
        n11506) );
  NOR2_X1 U14601 ( .A1(n11777), .A2(n11720), .ZN(n11527) );
  AOI22_X1 U14602 ( .A1(n12323), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11371), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11511) );
  AOI22_X1 U14603 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12329), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11510) );
  AOI22_X1 U14604 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12144), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11509) );
  AOI22_X1 U14605 ( .A1(n12316), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12328), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11508) );
  NAND4_X1 U14606 ( .A1(n11511), .A2(n11510), .A3(n11509), .A4(n11508), .ZN(
        n11517) );
  AOI22_X1 U14607 ( .A1(n12325), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12327), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11515) );
  AOI22_X1 U14608 ( .A1(n12266), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11514) );
  AOI22_X1 U14609 ( .A1(n12326), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9772), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11513) );
  AOI22_X1 U14610 ( .A1(n12248), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12317), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11512) );
  NAND4_X1 U14611 ( .A1(n11515), .A2(n11514), .A3(n11513), .A4(n11512), .ZN(
        n11516) );
  MUX2_X1 U14612 ( .A(n11650), .B(n11527), .S(n11666), .Z(n11518) );
  INV_X1 U14613 ( .A(n11518), .ZN(n11519) );
  INV_X1 U14614 ( .A(n11666), .ZN(n11522) );
  NAND2_X1 U14615 ( .A1(n20152), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11521) );
  MUX2_X1 U14616 ( .A(n11522), .B(n11521), .S(n11464), .Z(n11524) );
  AOI21_X1 U14617 ( .B1(n13244), .B2(n11720), .A(n11495), .ZN(n11523) );
  NAND2_X1 U14618 ( .A1(n11524), .A2(n11523), .ZN(n11663) );
  NAND2_X1 U14619 ( .A1(n11664), .A2(n11663), .ZN(n11526) );
  INV_X1 U14620 ( .A(n11650), .ZN(n11525) );
  NAND2_X1 U14621 ( .A1(n11526), .A2(n11525), .ZN(n11545) );
  INV_X1 U14622 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11543) );
  INV_X1 U14623 ( .A(n11527), .ZN(n11542) );
  INV_X1 U14624 ( .A(n11597), .ZN(n11540) );
  AOI22_X1 U14625 ( .A1(n12323), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11532) );
  AOI22_X1 U14626 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12327), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11531) );
  AOI22_X1 U14627 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12144), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11530) );
  AOI22_X1 U14628 ( .A1(n12329), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12317), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11529) );
  NAND4_X1 U14629 ( .A1(n11532), .A2(n11531), .A3(n11530), .A4(n11529), .ZN(
        n11539) );
  AOI22_X1 U14630 ( .A1(n12248), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11537) );
  AOI22_X1 U14631 ( .A1(n12325), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12328), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11536) );
  AOI22_X1 U14632 ( .A1(n12324), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11535) );
  AOI22_X1 U14633 ( .A1(n12326), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9772), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11534) );
  NAND4_X1 U14634 ( .A1(n11537), .A2(n11536), .A3(n11535), .A4(n11534), .ZN(
        n11538) );
  NAND2_X1 U14635 ( .A1(n11540), .A2(n11658), .ZN(n11541) );
  OAI211_X1 U14636 ( .C1(n11809), .C2(n11543), .A(n11542), .B(n11541), .ZN(
        n11544) );
  NAND2_X1 U14637 ( .A1(n11545), .A2(n11544), .ZN(n11546) );
  INV_X1 U14638 ( .A(n11838), .ZN(n11557) );
  NAND2_X1 U14639 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11568) );
  OAI21_X1 U14640 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n11568), .ZN(n20472) );
  OR2_X1 U14641 ( .A1(n15747), .A2(n20555), .ZN(n11559) );
  OAI21_X1 U14642 ( .B1(n20835), .B2(n20472), .A(n11559), .ZN(n11547) );
  INV_X1 U14643 ( .A(n11547), .ZN(n11548) );
  INV_X1 U14644 ( .A(n11552), .ZN(n11553) );
  INV_X1 U14645 ( .A(n11777), .ZN(n11554) );
  NAND2_X1 U14646 ( .A1(n11554), .A2(n11658), .ZN(n11555) );
  NAND2_X1 U14647 ( .A1(n11840), .A2(n9769), .ZN(n11653) );
  INV_X1 U14648 ( .A(n11653), .ZN(n11589) );
  INV_X1 U14649 ( .A(n11559), .ZN(n11562) );
  INV_X1 U14650 ( .A(n11560), .ZN(n11561) );
  OAI21_X1 U14651 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n11562), .A(
        n11561), .ZN(n11563) );
  INV_X1 U14652 ( .A(n20835), .ZN(n11570) );
  INV_X1 U14653 ( .A(n11568), .ZN(n11567) );
  NAND2_X1 U14654 ( .A1(n11567), .A2(n11766), .ZN(n20516) );
  NAND2_X1 U14655 ( .A1(n11568), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11569) );
  NAND2_X1 U14656 ( .A1(n20516), .A2(n11569), .ZN(n20123) );
  NAND2_X1 U14657 ( .A1(n11570), .A2(n20123), .ZN(n11573) );
  INV_X1 U14658 ( .A(n15747), .ZN(n11571) );
  NAND2_X1 U14659 ( .A1(n11571), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11572) );
  AOI22_X1 U14660 ( .A1(n12323), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11371), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11579) );
  AOI22_X1 U14661 ( .A1(n12316), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12329), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11578) );
  AOI22_X1 U14662 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11577) );
  AOI22_X1 U14663 ( .A1(n12318), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12317), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11576) );
  NAND4_X1 U14664 ( .A1(n11579), .A2(n11578), .A3(n11577), .A4(n11576), .ZN(
        n11585) );
  INV_X1 U14665 ( .A(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n21003) );
  AOI22_X1 U14666 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11583) );
  AOI22_X1 U14667 ( .A1(n12327), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12144), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11582) );
  AOI22_X1 U14668 ( .A1(n12266), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12328), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11581) );
  AOI22_X1 U14669 ( .A1(n12326), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9757), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11580) );
  NAND4_X1 U14670 ( .A1(n11583), .A2(n11582), .A3(n11581), .A4(n11580), .ZN(
        n11584) );
  INV_X1 U14671 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n20143) );
  OAI22_X1 U14672 ( .A1(n11809), .A2(n20143), .B1(n11677), .B2(n11597), .ZN(
        n11586) );
  INV_X1 U14673 ( .A(n11586), .ZN(n11587) );
  XNOR2_X2 U14674 ( .A(n11588), .B(n11587), .ZN(n11652) );
  INV_X1 U14675 ( .A(n11565), .ZN(n11591) );
  NAND2_X1 U14676 ( .A1(n11591), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11596) );
  NOR3_X1 U14677 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n11766), .A3(
        n20555), .ZN(n20394) );
  NAND2_X1 U14678 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20394), .ZN(
        n20392) );
  NAND2_X1 U14679 ( .A1(n20515), .A2(n20392), .ZN(n11593) );
  NAND3_X1 U14680 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20681) );
  INV_X1 U14681 ( .A(n20681), .ZN(n11592) );
  NAND2_X1 U14682 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n11592), .ZN(
        n20674) );
  NAND2_X1 U14683 ( .A1(n11593), .A2(n20674), .ZN(n20417) );
  OAI22_X1 U14684 ( .A1(n20835), .A2(n20417), .B1(n15747), .B2(n20515), .ZN(
        n11594) );
  INV_X1 U14685 ( .A(n11594), .ZN(n11595) );
  XNOR2_X2 U14686 ( .A(n11590), .B(n20295), .ZN(n20416) );
  INV_X1 U14687 ( .A(n11809), .ZN(n11791) );
  AOI22_X1 U14688 ( .A1(n12323), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11371), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11601) );
  AOI22_X1 U14689 ( .A1(n12316), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12329), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11600) );
  AOI22_X1 U14690 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11599) );
  AOI22_X1 U14691 ( .A1(n12248), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12317), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11598) );
  NAND4_X1 U14692 ( .A1(n11601), .A2(n11600), .A3(n11599), .A4(n11598), .ZN(
        n11607) );
  AOI22_X1 U14693 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11605) );
  AOI22_X1 U14694 ( .A1(n12327), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12144), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11604) );
  AOI22_X1 U14695 ( .A1(n12324), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12328), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11603) );
  AOI22_X1 U14696 ( .A1(n12326), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11501), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11602) );
  NAND4_X1 U14697 ( .A1(n11605), .A2(n11604), .A3(n11603), .A4(n11602), .ZN(
        n11606) );
  AOI22_X1 U14698 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11814), .B2(n11694), .ZN(n11608) );
  NAND2_X1 U14699 ( .A1(n9767), .A2(n11589), .ZN(n11675) );
  INV_X1 U14700 ( .A(n11675), .ZN(n11622) );
  AOI22_X1 U14701 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11613) );
  AOI22_X1 U14702 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12248), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11612) );
  AOI22_X1 U14703 ( .A1(n12326), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9772), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11611) );
  AOI22_X1 U14704 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n12299), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11610) );
  NAND4_X1 U14705 ( .A1(n11613), .A2(n11612), .A3(n11611), .A4(n11610), .ZN(
        n11619) );
  AOI22_X1 U14706 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12316), .B1(
        n12329), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11617) );
  AOI22_X1 U14707 ( .A1(n12327), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12144), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11616) );
  AOI22_X1 U14708 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n12324), .B1(
        n12328), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11615) );
  AOI22_X1 U14709 ( .A1(n12323), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12317), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11614) );
  NAND4_X1 U14710 ( .A1(n11617), .A2(n11616), .A3(n11615), .A4(n11614), .ZN(
        n11618) );
  NAND2_X1 U14711 ( .A1(n11814), .A2(n11693), .ZN(n11621) );
  INV_X1 U14712 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n20159) );
  OR2_X1 U14713 ( .A1(n11809), .A2(n20159), .ZN(n11620) );
  NAND2_X1 U14714 ( .A1(n11621), .A2(n11620), .ZN(n11682) );
  INV_X1 U14715 ( .A(n11691), .ZN(n11637) );
  INV_X1 U14716 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11623) );
  OR2_X1 U14717 ( .A1(n11809), .A2(n11623), .ZN(n11635) );
  AOI22_X1 U14718 ( .A1(n12323), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11371), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11627) );
  AOI22_X1 U14719 ( .A1(n12316), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12329), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11626) );
  AOI22_X1 U14720 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11625) );
  AOI22_X1 U14721 ( .A1(n12248), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12317), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11624) );
  NAND4_X1 U14722 ( .A1(n11627), .A2(n11626), .A3(n11625), .A4(n11624), .ZN(
        n11633) );
  AOI22_X1 U14723 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11631) );
  AOI22_X1 U14724 ( .A1(n12327), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12144), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11630) );
  AOI22_X1 U14725 ( .A1(n12324), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12328), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11629) );
  AOI22_X1 U14726 ( .A1(n12326), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9757), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11628) );
  NAND4_X1 U14727 ( .A1(n11631), .A2(n11630), .A3(n11629), .A4(n11628), .ZN(
        n11632) );
  NAND2_X1 U14728 ( .A1(n11814), .A2(n11705), .ZN(n11634) );
  INV_X1 U14729 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n20171) );
  OR2_X1 U14730 ( .A1(n11809), .A2(n20171), .ZN(n11649) );
  AOI22_X1 U14731 ( .A1(n12248), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12323), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11641) );
  AOI22_X1 U14732 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12299), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11640) );
  AOI22_X1 U14733 ( .A1(n12326), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9772), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11639) );
  AOI22_X1 U14734 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12317), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11638) );
  NAND4_X1 U14735 ( .A1(n11641), .A2(n11640), .A3(n11639), .A4(n11638), .ZN(
        n11647) );
  AOI22_X1 U14736 ( .A1(n12316), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12324), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11645) );
  AOI22_X1 U14737 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12327), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11644) );
  AOI22_X1 U14738 ( .A1(n12325), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12144), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11643) );
  AOI22_X1 U14739 ( .A1(n12329), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11642) );
  NAND4_X1 U14740 ( .A1(n11645), .A2(n11644), .A3(n11643), .A4(n11642), .ZN(
        n11646) );
  NAND2_X1 U14741 ( .A1(n11814), .A2(n11718), .ZN(n11648) );
  NAND2_X4 U14742 ( .A1(n11716), .A2(n11651), .ZN(n14460) );
  NAND3_X1 U14743 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14603) );
  XNOR2_X2 U14744 ( .A(n11653), .B(n11652), .ZN(n13420) );
  NAND2_X1 U14745 ( .A1(n13420), .A2(n12351), .ZN(n11657) );
  NAND2_X1 U14746 ( .A1(n11666), .A2(n11658), .ZN(n11678) );
  XNOR2_X1 U14747 ( .A(n11678), .B(n11677), .ZN(n11655) );
  NAND2_X1 U14748 ( .A1(n13183), .A2(n20145), .ZN(n11665) );
  INV_X1 U14749 ( .A(n11665), .ZN(n11654) );
  AOI21_X1 U14750 ( .B1(n11655), .B2(n15742), .A(n11654), .ZN(n11656) );
  NAND2_X1 U14751 ( .A1(n11657), .A2(n11656), .ZN(n13426) );
  XNOR2_X1 U14752 ( .A(n11666), .B(n11658), .ZN(n11660) );
  OAI211_X1 U14753 ( .C1(n11660), .C2(n20842), .A(n11392), .B(n20160), .ZN(
        n11661) );
  INV_X1 U14754 ( .A(n11661), .ZN(n11662) );
  XNOR2_X1 U14755 ( .A(n11664), .B(n11663), .ZN(n11845) );
  OAI21_X1 U14756 ( .B1(n20842), .B2(n11666), .A(n11665), .ZN(n11667) );
  INV_X1 U14757 ( .A(n11667), .ZN(n11668) );
  OAI21_X2 U14758 ( .B1(n11845), .B2(n11770), .A(n11668), .ZN(n13246) );
  XNOR2_X1 U14759 ( .A(n11670), .B(n11669), .ZN(n13299) );
  NAND2_X1 U14760 ( .A1(n13299), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13300) );
  INV_X1 U14761 ( .A(n11670), .ZN(n11671) );
  NAND2_X1 U14762 ( .A1(n13300), .A2(n11672), .ZN(n11673) );
  INV_X1 U14763 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20082) );
  XNOR2_X1 U14764 ( .A(n11673), .B(n20082), .ZN(n13424) );
  NAND2_X1 U14765 ( .A1(n13426), .A2(n13424), .ZN(n13425) );
  NAND2_X1 U14766 ( .A1(n11673), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11674) );
  INV_X1 U14767 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20069) );
  INV_X1 U14768 ( .A(n13471), .ZN(n13474) );
  NAND2_X1 U14769 ( .A1(n9768), .A2(n13474), .ZN(n11676) );
  NAND2_X1 U14770 ( .A1(n11678), .A2(n11677), .ZN(n11696) );
  XNOR2_X1 U14771 ( .A(n11696), .B(n11694), .ZN(n11679) );
  OAI22_X1 U14772 ( .A1(n20107), .A2(n11770), .B1(n20842), .B2(n11679), .ZN(
        n13559) );
  NAND2_X1 U14773 ( .A1(n13560), .A2(n13559), .ZN(n13558) );
  NAND2_X1 U14774 ( .A1(n11680), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11681) );
  NAND2_X1 U14775 ( .A1(n13558), .A2(n11681), .ZN(n20042) );
  INV_X1 U14776 ( .A(n11682), .ZN(n11683) );
  NAND2_X1 U14777 ( .A1(n11684), .A2(n11691), .ZN(n11858) );
  NAND2_X1 U14778 ( .A1(n11696), .A2(n11694), .ZN(n11685) );
  XNOR2_X1 U14779 ( .A(n11685), .B(n11693), .ZN(n11686) );
  NAND2_X1 U14780 ( .A1(n11686), .A2(n15742), .ZN(n11687) );
  INV_X1 U14781 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20062) );
  XNOR2_X1 U14782 ( .A(n11688), .B(n20062), .ZN(n20041) );
  NAND2_X1 U14783 ( .A1(n20042), .A2(n20041), .ZN(n20040) );
  NAND2_X1 U14784 ( .A1(n11688), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11689) );
  NAND2_X1 U14785 ( .A1(n11691), .A2(n11690), .ZN(n11692) );
  NAND2_X1 U14786 ( .A1(n11872), .A2(n12351), .ZN(n11699) );
  AND2_X1 U14787 ( .A1(n11694), .A2(n11693), .ZN(n11695) );
  NAND2_X1 U14788 ( .A1(n11696), .A2(n11695), .ZN(n11704) );
  XNOR2_X1 U14789 ( .A(n11704), .B(n11705), .ZN(n11697) );
  NAND2_X1 U14790 ( .A1(n11697), .A2(n15742), .ZN(n11698) );
  NAND2_X1 U14791 ( .A1(n11699), .A2(n11698), .ZN(n11700) );
  INV_X1 U14792 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16060) );
  XNOR2_X1 U14793 ( .A(n11700), .B(n16060), .ZN(n15942) );
  NAND2_X1 U14794 ( .A1(n11700), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11701) );
  NAND2_X1 U14795 ( .A1(n11703), .A2(n11702), .ZN(n11879) );
  NAND3_X1 U14796 ( .A1(n11716), .A2(n12351), .A3(n11879), .ZN(n11709) );
  INV_X1 U14797 ( .A(n11704), .ZN(n11706) );
  NAND2_X1 U14798 ( .A1(n11706), .A2(n11705), .ZN(n11717) );
  XNOR2_X1 U14799 ( .A(n11717), .B(n11718), .ZN(n11707) );
  NAND2_X1 U14800 ( .A1(n11707), .A2(n15742), .ZN(n11708) );
  INV_X1 U14801 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15936) );
  NAND2_X1 U14802 ( .A1(n15937), .A2(n15936), .ZN(n11710) );
  INV_X1 U14803 ( .A(n15937), .ZN(n11711) );
  NAND2_X1 U14804 ( .A1(n11711), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11712) );
  INV_X1 U14805 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11714) );
  NAND2_X1 U14806 ( .A1(n11814), .A2(n11720), .ZN(n11713) );
  OAI21_X1 U14807 ( .B1(n11714), .B2(n11809), .A(n11713), .ZN(n11715) );
  INV_X1 U14808 ( .A(n11717), .ZN(n11719) );
  NAND2_X1 U14809 ( .A1(n11719), .A2(n11718), .ZN(n11727) );
  XNOR2_X1 U14810 ( .A(n11727), .B(n11720), .ZN(n11721) );
  AND2_X1 U14811 ( .A1(n11721), .A2(n15742), .ZN(n11722) );
  AOI21_X1 U14812 ( .B1(n11880), .B2(n12351), .A(n11722), .ZN(n11723) );
  INV_X1 U14813 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16082) );
  NAND2_X1 U14814 ( .A1(n11723), .A2(n16082), .ZN(n15931) );
  NAND2_X1 U14815 ( .A1(n15929), .A2(n15931), .ZN(n11725) );
  INV_X1 U14816 ( .A(n11723), .ZN(n11724) );
  NAND2_X1 U14817 ( .A1(n11724), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15930) );
  NAND2_X1 U14818 ( .A1(n11725), .A2(n15930), .ZN(n13844) );
  OR3_X1 U14819 ( .A1(n11727), .A2(n11726), .A3(n20842), .ZN(n11728) );
  INV_X1 U14820 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11729) );
  NAND2_X1 U14821 ( .A1(n13845), .A2(n11729), .ZN(n11730) );
  NAND2_X1 U14822 ( .A1(n13844), .A2(n11730), .ZN(n11733) );
  INV_X1 U14823 ( .A(n13845), .ZN(n11731) );
  NAND2_X1 U14824 ( .A1(n11731), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11732) );
  NAND2_X1 U14825 ( .A1(n14460), .A2(n16059), .ZN(n11734) );
  INV_X1 U14826 ( .A(n14009), .ZN(n11747) );
  NAND2_X1 U14827 ( .A1(n14014), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14545) );
  INV_X1 U14828 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16017) );
  NAND2_X1 U14829 ( .A1(n14460), .A2(n16017), .ZN(n11735) );
  NAND2_X1 U14830 ( .A1(n14545), .A2(n11735), .ZN(n14016) );
  NAND2_X1 U14831 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11736) );
  AND2_X1 U14832 ( .A1(n14460), .A2(n11736), .ZN(n14011) );
  NOR2_X1 U14833 ( .A1(n14016), .A2(n14011), .ZN(n14544) );
  INV_X1 U14834 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11742) );
  NAND2_X1 U14835 ( .A1(n14460), .A2(n11742), .ZN(n14543) );
  INV_X1 U14836 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16008) );
  NAND2_X1 U14837 ( .A1(n14460), .A2(n16008), .ZN(n11737) );
  AND2_X1 U14838 ( .A1(n14543), .A2(n11737), .ZN(n11738) );
  NAND2_X1 U14839 ( .A1(n15893), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11739) );
  NAND2_X1 U14840 ( .A1(n14545), .A2(n11739), .ZN(n11744) );
  INV_X1 U14841 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11740) );
  NOR2_X1 U14842 ( .A1(n14460), .A2(n11740), .ZN(n11745) );
  NOR2_X1 U14843 ( .A1(n11744), .A2(n11745), .ZN(n15896) );
  XNOR2_X1 U14844 ( .A(n14460), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14536) );
  NAND2_X1 U14845 ( .A1(n14460), .A2(n11740), .ZN(n14534) );
  NAND2_X1 U14846 ( .A1(n14536), .A2(n14534), .ZN(n11741) );
  AOI21_X1 U14847 ( .B1(n14532), .B2(n15896), .A(n11741), .ZN(n15894) );
  NOR2_X1 U14848 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14010) );
  AND2_X1 U14849 ( .A1(n14010), .A2(n11742), .ZN(n11743) );
  NOR2_X1 U14850 ( .A1(n14460), .A2(n11743), .ZN(n14542) );
  NOR2_X1 U14851 ( .A1(n11744), .A2(n14542), .ZN(n14531) );
  INV_X1 U14852 ( .A(n11745), .ZN(n14533) );
  NAND2_X1 U14853 ( .A1(n14531), .A2(n14533), .ZN(n11746) );
  AOI21_X1 U14854 ( .B1(n11747), .B2(n10130), .A(n11746), .ZN(n11751) );
  NOR2_X1 U14855 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11748) );
  NAND2_X1 U14856 ( .A1(n14009), .A2(n11748), .ZN(n11749) );
  NAND2_X1 U14857 ( .A1(n11749), .A2(n15893), .ZN(n11750) );
  XNOR2_X1 U14858 ( .A(n14460), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14525) );
  NAND2_X1 U14859 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14642) );
  INV_X1 U14860 ( .A(n14642), .ZN(n11752) );
  NAND2_X1 U14861 ( .A1(n11753), .A2(n14460), .ZN(n14504) );
  NOR2_X1 U14862 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11754) );
  INV_X1 U14863 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11756) );
  INV_X1 U14864 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14521) );
  INV_X1 U14865 ( .A(n13966), .ZN(n14487) );
  INV_X1 U14866 ( .A(n11759), .ZN(n11762) );
  INV_X1 U14867 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14606) );
  MUX2_X1 U14868 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n14606), .S(
        n14460), .Z(n11757) );
  INV_X1 U14869 ( .A(n11757), .ZN(n11761) );
  INV_X1 U14870 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n21048) );
  INV_X1 U14871 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n13995) );
  NAND2_X1 U14872 ( .A1(n21048), .A2(n13995), .ZN(n13968) );
  NOR3_X1 U14873 ( .A1(n13968), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11758) );
  OAI211_X1 U14874 ( .C1(n11762), .C2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n11761), .B(n11760), .ZN(n11763) );
  INV_X1 U14875 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12451) );
  XNOR2_X1 U14876 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11786) );
  NAND2_X1 U14877 ( .A1(n11785), .A2(n11786), .ZN(n11765) );
  NAND2_X1 U14878 ( .A1(n20555), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11764) );
  NAND2_X1 U14879 ( .A1(n11765), .A2(n11764), .ZN(n11790) );
  MUX2_X1 U14880 ( .A(n11766), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n11789) );
  NAND2_X1 U14881 ( .A1(n11790), .A2(n11789), .ZN(n11768) );
  NAND2_X1 U14882 ( .A1(n11766), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11767) );
  MUX2_X1 U14883 ( .A(n20515), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n11771) );
  NOR2_X1 U14884 ( .A1(n13387), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11769) );
  XNOR2_X1 U14885 ( .A(n11772), .B(n11771), .ZN(n13134) );
  INV_X1 U14886 ( .A(n11814), .ZN(n11794) );
  NAND2_X1 U14887 ( .A1(n11472), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11773) );
  NAND2_X1 U14888 ( .A1(n11794), .A2(n11773), .ZN(n11788) );
  INV_X1 U14889 ( .A(n11788), .ZN(n11774) );
  NAND2_X1 U14890 ( .A1(n11774), .A2(n12355), .ZN(n11795) );
  INV_X1 U14891 ( .A(n13137), .ZN(n11775) );
  NOR2_X1 U14892 ( .A1(n11795), .A2(n11775), .ZN(n11807) );
  NAND2_X1 U14893 ( .A1(n13291), .A2(n20160), .ZN(n11787) );
  NAND2_X1 U14894 ( .A1(n11776), .A2(n11787), .ZN(n11803) );
  NOR3_X1 U14895 ( .A1(n11472), .A2(n11777), .A3(n13183), .ZN(n11780) );
  INV_X1 U14896 ( .A(n11785), .ZN(n11779) );
  NAND2_X1 U14897 ( .A1(n11311), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11778) );
  NAND2_X1 U14898 ( .A1(n11779), .A2(n11778), .ZN(n11781) );
  NOR3_X1 U14899 ( .A1(n11803), .A2(n11780), .A3(n11781), .ZN(n11784) );
  INV_X1 U14900 ( .A(n11781), .ZN(n11782) );
  AOI21_X1 U14901 ( .B1(n11782), .B2(n11814), .A(n11817), .ZN(n11783) );
  NOR2_X1 U14902 ( .A1(n11784), .A2(n11783), .ZN(n11801) );
  XNOR2_X1 U14903 ( .A(n11786), .B(n11785), .ZN(n13136) );
  AOI22_X1 U14904 ( .A1(n11788), .A2(n11787), .B1(n11791), .B2(n13136), .ZN(
        n11796) );
  INV_X1 U14905 ( .A(n11796), .ZN(n11800) );
  XNOR2_X1 U14906 ( .A(n11790), .B(n11789), .ZN(n13135) );
  INV_X1 U14907 ( .A(n11803), .ZN(n11793) );
  NAND2_X1 U14908 ( .A1(n11791), .A2(n13135), .ZN(n11792) );
  OAI211_X1 U14909 ( .C1(n11794), .C2(n13135), .A(n11793), .B(n11792), .ZN(
        n11799) );
  INV_X1 U14910 ( .A(n11801), .ZN(n11797) );
  OAI211_X1 U14911 ( .C1(n11797), .C2(n11796), .A(n13136), .B(n11795), .ZN(
        n11798) );
  OAI211_X1 U14912 ( .C1(n11801), .C2(n11800), .A(n11799), .B(n11798), .ZN(
        n11805) );
  INV_X1 U14913 ( .A(n13135), .ZN(n11802) );
  NAND3_X1 U14914 ( .A1(n11803), .A2(n11802), .A3(n11814), .ZN(n11804) );
  AOI22_X1 U14915 ( .A1(n11805), .A2(n11804), .B1(n11809), .B2(n13134), .ZN(
        n11806) );
  AOI211_X1 U14916 ( .C1(n11817), .C2(n13134), .A(n11807), .B(n11806), .ZN(
        n11808) );
  AOI21_X1 U14917 ( .B1(n13137), .B2(n11809), .A(n11808), .ZN(n11810) );
  AOI21_X1 U14918 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n11495), .A(
        n11810), .ZN(n11816) );
  NAND2_X1 U14919 ( .A1(n20105), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11812) );
  NAND2_X1 U14920 ( .A1(n13139), .A2(n11814), .ZN(n11815) );
  NAND2_X1 U14921 ( .A1(n11816), .A2(n11815), .ZN(n11819) );
  NAND2_X1 U14922 ( .A1(n11817), .A2(n13139), .ZN(n11818) );
  AOI21_X1 U14923 ( .B1(n14652), .B2(n13183), .A(n11659), .ZN(n11821) );
  NAND2_X1 U14924 ( .A1(n13185), .A2(n11822), .ZN(n15735) );
  NAND2_X1 U14925 ( .A1(n14586), .A2(n20046), .ZN(n12289) );
  INV_X1 U14926 ( .A(n12044), .ZN(n12062) );
  AND2_X1 U14927 ( .A1(n13234), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11850) );
  INV_X1 U14928 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n11827) );
  NAND2_X1 U14929 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11823) );
  INV_X1 U14930 ( .A(n11823), .ZN(n11825) );
  INV_X1 U14931 ( .A(n11860), .ZN(n11824) );
  OAI21_X1 U14932 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11825), .A(
        n11824), .ZN(n13562) );
  AOI22_X1 U14933 ( .A1(n12345), .A2(n13562), .B1(n14083), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11826) );
  OAI21_X1 U14934 ( .B1(n12343), .B2(n11827), .A(n11826), .ZN(n11828) );
  AOI21_X1 U14935 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n11850), .A(
        n11828), .ZN(n11829) );
  NAND2_X1 U14936 ( .A1(n14083), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11857) );
  INV_X1 U14937 ( .A(n11857), .ZN(n11834) );
  INV_X1 U14938 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n11831) );
  XNOR2_X1 U14939 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13736) );
  AOI21_X1 U14940 ( .B1(n12345), .B2(n13736), .A(n14083), .ZN(n11830) );
  OAI21_X1 U14941 ( .B1(n12343), .B2(n11831), .A(n11830), .ZN(n11832) );
  AOI21_X1 U14942 ( .B1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n11850), .A(
        n11832), .ZN(n11833) );
  NOR2_X1 U14943 ( .A1(n11834), .A2(n11833), .ZN(n11835) );
  NAND2_X1 U14944 ( .A1(n11838), .A2(n11837), .ZN(n11839) );
  NAND2_X1 U14945 ( .A1(n20214), .A2(n12044), .ZN(n11844) );
  INV_X1 U14946 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n11841) );
  INV_X1 U14947 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13298) );
  OAI22_X1 U14948 ( .A1(n12343), .A2(n11841), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13298), .ZN(n11842) );
  AOI21_X1 U14949 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n11850), .A(
        n11842), .ZN(n11843) );
  NAND2_X1 U14950 ( .A1(n11846), .A2(n12350), .ZN(n11847) );
  NAND2_X1 U14951 ( .A1(n11847), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13269) );
  INV_X1 U14952 ( .A(n11850), .ZN(n11863) );
  NAND2_X1 U14953 ( .A1(n14084), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11852) );
  NAND2_X1 U14954 ( .A1(n20742), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11851) );
  OAI211_X1 U14955 ( .C1(n11863), .C2(n11311), .A(n11852), .B(n11851), .ZN(
        n11853) );
  AOI21_X1 U14956 ( .B1(n11849), .B2(n12044), .A(n11853), .ZN(n13268) );
  OR2_X1 U14957 ( .A1(n13269), .A2(n13268), .ZN(n13271) );
  INV_X1 U14958 ( .A(n13268), .ZN(n11854) );
  OR2_X1 U14959 ( .A1(n11854), .A2(n12340), .ZN(n11855) );
  NAND2_X1 U14960 ( .A1(n13271), .A2(n11855), .ZN(n13295) );
  NAND2_X1 U14961 ( .A1(n13296), .A2(n13295), .ZN(n13431) );
  INV_X1 U14962 ( .A(n11858), .ZN(n11859) );
  NAND2_X1 U14963 ( .A1(n11859), .A2(n12044), .ZN(n11866) );
  NAND2_X1 U14964 ( .A1(n11860), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11867) );
  OAI21_X1 U14965 ( .B1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n11860), .A(
        n11867), .ZN(n20049) );
  INV_X1 U14966 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16101) );
  OAI21_X1 U14967 ( .B1(n20643), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20742), .ZN(n11862) );
  NAND2_X1 U14968 ( .A1(n14084), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n11861) );
  OAI211_X1 U14969 ( .C1(n11863), .C2(n16101), .A(n11862), .B(n11861), .ZN(
        n11864) );
  OAI21_X1 U14970 ( .B1(n12340), .B2(n20049), .A(n11864), .ZN(n11865) );
  NAND2_X1 U14971 ( .A1(n11866), .A2(n11865), .ZN(n13572) );
  NAND2_X1 U14972 ( .A1(n13574), .A2(n13572), .ZN(n13595) );
  INV_X1 U14973 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n11870) );
  INV_X1 U14974 ( .A(n11867), .ZN(n11868) );
  OAI21_X1 U14975 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n11868), .A(
        n11875), .ZN(n19959) );
  AOI22_X1 U14976 ( .A1(n12345), .A2(n19959), .B1(n14083), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11869) );
  OAI21_X1 U14977 ( .B1(n12343), .B2(n11870), .A(n11869), .ZN(n11871) );
  AOI21_X1 U14978 ( .B1(n11872), .B2(n12044), .A(n11871), .ZN(n13594) );
  INV_X1 U14979 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n13748) );
  OAI21_X1 U14980 ( .B1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n11876), .A(
        n11881), .ZN(n19953) );
  AOI22_X1 U14981 ( .A1(n12345), .A2(n19953), .B1(n14083), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11877) );
  OAI21_X1 U14982 ( .B1(n12343), .B2(n13748), .A(n11877), .ZN(n11878) );
  NAND2_X1 U14983 ( .A1(n11880), .A2(n12044), .ZN(n11888) );
  INV_X1 U14984 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n11885) );
  INV_X1 U14985 ( .A(n11881), .ZN(n11883) );
  INV_X1 U14986 ( .A(n11903), .ZN(n11882) );
  OAI21_X1 U14987 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n11883), .A(
        n11882), .ZN(n19940) );
  AOI22_X1 U14988 ( .A1(n12345), .A2(n19940), .B1(n14083), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11884) );
  OAI21_X1 U14989 ( .B1(n12343), .B2(n11885), .A(n11884), .ZN(n11886) );
  INV_X1 U14990 ( .A(n11886), .ZN(n11887) );
  NAND2_X1 U14991 ( .A1(n11888), .A2(n11887), .ZN(n13750) );
  NAND2_X1 U14992 ( .A1(n9803), .A2(n13750), .ZN(n13749) );
  AOI22_X1 U14993 ( .A1(n12323), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12316), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11892) );
  AOI22_X1 U14994 ( .A1(n12325), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12328), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11891) );
  AOI22_X1 U14995 ( .A1(n12144), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11890) );
  AOI22_X1 U14996 ( .A1(n12326), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9772), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11889) );
  NAND4_X1 U14997 ( .A1(n11892), .A2(n11891), .A3(n11890), .A4(n11889), .ZN(
        n11898) );
  AOI22_X1 U14998 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12324), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11896) );
  AOI22_X1 U14999 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12329), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11895) );
  AOI22_X1 U15000 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12327), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11894) );
  AOI22_X1 U15001 ( .A1(n12248), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12317), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11893) );
  NAND4_X1 U15002 ( .A1(n11896), .A2(n11895), .A3(n11894), .A4(n11893), .ZN(
        n11897) );
  OAI21_X1 U15003 ( .B1(n11898), .B2(n11897), .A(n12044), .ZN(n11901) );
  NAND2_X1 U15004 ( .A1(n14084), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11900) );
  XNOR2_X1 U15005 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n11903), .ZN(
        n13848) );
  AOI22_X1 U15006 ( .A1(n12345), .A2(n13848), .B1(n14083), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11899) );
  XNOR2_X1 U15007 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n11918), .ZN(
        n13901) );
  INV_X1 U15008 ( .A(n13901), .ZN(n19925) );
  AOI22_X1 U15009 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11907) );
  AOI22_X1 U15010 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12324), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11906) );
  AOI22_X1 U15011 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12329), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11905) );
  AOI22_X1 U15012 ( .A1(n12326), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11501), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11904) );
  NAND4_X1 U15013 ( .A1(n11907), .A2(n11906), .A3(n11905), .A4(n11904), .ZN(
        n11913) );
  AOI22_X1 U15014 ( .A1(n12248), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12323), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11911) );
  AOI22_X1 U15015 ( .A1(n12144), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12328), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11910) );
  AOI22_X1 U15016 ( .A1(n12316), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11909) );
  AOI22_X1 U15017 ( .A1(n12327), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12317), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11908) );
  NAND4_X1 U15018 ( .A1(n11911), .A2(n11910), .A3(n11909), .A4(n11908), .ZN(
        n11912) );
  OAI21_X1 U15019 ( .B1(n11913), .B2(n11912), .A(n12044), .ZN(n11916) );
  NAND2_X1 U15020 ( .A1(n14084), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11915) );
  NAND2_X1 U15021 ( .A1(n14083), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11914) );
  NAND3_X1 U15022 ( .A1(n11916), .A2(n11915), .A3(n11914), .ZN(n11917) );
  AOI21_X1 U15023 ( .B1(n19925), .B2(n12345), .A(n11917), .ZN(n13876) );
  XNOR2_X1 U15024 ( .A(n11934), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14561) );
  NAND2_X1 U15025 ( .A1(n14561), .A2(n13671), .ZN(n11933) );
  AOI22_X1 U15026 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12327), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11922) );
  AOI22_X1 U15027 ( .A1(n12144), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11921) );
  AOI22_X1 U15028 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12328), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11920) );
  AOI22_X1 U15029 ( .A1(n12326), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9757), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11919) );
  NAND4_X1 U15030 ( .A1(n11922), .A2(n11921), .A3(n11920), .A4(n11919), .ZN(
        n11928) );
  AOI22_X1 U15031 ( .A1(n12325), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12299), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11926) );
  AOI22_X1 U15032 ( .A1(n12316), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12324), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11925) );
  AOI22_X1 U15033 ( .A1(n12248), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12329), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11924) );
  AOI22_X1 U15034 ( .A1(n12323), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12317), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11923) );
  NAND4_X1 U15035 ( .A1(n11926), .A2(n11925), .A3(n11924), .A4(n11923), .ZN(
        n11927) );
  OAI21_X1 U15036 ( .B1(n11928), .B2(n11927), .A(n12044), .ZN(n11931) );
  NAND2_X1 U15037 ( .A1(n14084), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n11930) );
  NAND2_X1 U15038 ( .A1(n14083), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11929) );
  INV_X1 U15039 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n11937) );
  OAI21_X1 U15040 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11935), .A(
        n12063), .ZN(n15928) );
  AOI22_X1 U15041 ( .A1(n12345), .A2(n15928), .B1(n14083), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11936) );
  OAI21_X1 U15042 ( .B1(n12343), .B2(n11937), .A(n11936), .ZN(n14003) );
  NAND2_X1 U15043 ( .A1(n13909), .A2(n14003), .ZN(n14002) );
  AOI22_X1 U15044 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11941) );
  AOI22_X1 U15045 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12324), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11940) );
  AOI22_X1 U15046 ( .A1(n12327), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12144), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11939) );
  AOI22_X1 U15047 ( .A1(n12326), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9757), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11938) );
  NAND4_X1 U15048 ( .A1(n11941), .A2(n11940), .A3(n11939), .A4(n11938), .ZN(
        n11947) );
  AOI22_X1 U15049 ( .A1(n12323), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11371), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11945) );
  AOI22_X1 U15050 ( .A1(n12316), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12328), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11944) );
  AOI22_X1 U15051 ( .A1(n12329), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11943) );
  AOI22_X1 U15052 ( .A1(n12248), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12317), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11942) );
  NAND4_X1 U15053 ( .A1(n11945), .A2(n11944), .A3(n11943), .A4(n11942), .ZN(
        n11946) );
  OR2_X1 U15054 ( .A1(n11947), .A2(n11946), .ZN(n11948) );
  NAND2_X1 U15055 ( .A1(n13909), .A2(n15874), .ZN(n11949) );
  INV_X1 U15056 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11952) );
  XNOR2_X1 U15057 ( .A(n12088), .B(n11952), .ZN(n15824) );
  NAND2_X1 U15058 ( .A1(n15824), .A2(n13671), .ZN(n11969) );
  AOI22_X1 U15059 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12324), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11956) );
  AOI22_X1 U15060 ( .A1(n12316), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12144), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11955) );
  AOI22_X1 U15061 ( .A1(n12327), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12326), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11954) );
  AOI22_X1 U15062 ( .A1(n12328), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12317), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11953) );
  NAND4_X1 U15063 ( .A1(n11956), .A2(n11955), .A3(n11954), .A4(n11953), .ZN(
        n11964) );
  AOI22_X1 U15064 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11371), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11962) );
  AOI22_X1 U15065 ( .A1(n12325), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12329), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11961) );
  AOI22_X1 U15066 ( .A1(n12248), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11380), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11960) );
  NAND2_X1 U15067 ( .A1(n12323), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n11958) );
  AOI21_X1 U15068 ( .B1(n9772), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A(n13671), .ZN(n11957) );
  AND2_X1 U15069 ( .A1(n11958), .A2(n11957), .ZN(n11959) );
  NAND4_X1 U15070 ( .A1(n11962), .A2(n11961), .A3(n11960), .A4(n11959), .ZN(
        n11963) );
  NAND2_X1 U15071 ( .A1(n12310), .A2(n12340), .ZN(n12110) );
  OAI21_X1 U15072 ( .B1(n11964), .B2(n11963), .A(n12110), .ZN(n11967) );
  NAND2_X1 U15073 ( .A1(n14084), .A2(P1_EAX_REG_18__SCAN_IN), .ZN(n11966) );
  NAND2_X1 U15074 ( .A1(n20742), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11965) );
  NAND3_X1 U15075 ( .A1(n11967), .A2(n11966), .A3(n11965), .ZN(n11968) );
  NAND2_X1 U15076 ( .A1(n11969), .A2(n11968), .ZN(n14351) );
  INV_X1 U15077 ( .A(n14351), .ZN(n12071) );
  XNOR2_X1 U15078 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n11970), .ZN(
        n15901) );
  INV_X1 U15079 ( .A(n12310), .ZN(n12338) );
  AOI22_X1 U15080 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12329), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11974) );
  AOI22_X1 U15081 ( .A1(n12325), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12327), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11973) );
  AOI22_X1 U15082 ( .A1(n12324), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12096), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11972) );
  AOI22_X1 U15083 ( .A1(n12326), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9772), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11971) );
  NAND4_X1 U15084 ( .A1(n11974), .A2(n11973), .A3(n11972), .A4(n11971), .ZN(
        n11980) );
  AOI22_X1 U15085 ( .A1(n12323), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11978) );
  AOI22_X1 U15086 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12144), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11977) );
  AOI22_X1 U15087 ( .A1(n12316), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11380), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11976) );
  AOI22_X1 U15088 ( .A1(n12318), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12317), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11975) );
  NAND4_X1 U15089 ( .A1(n11978), .A2(n11977), .A3(n11976), .A4(n11975), .ZN(
        n11979) );
  OR2_X1 U15090 ( .A1(n11980), .A2(n11979), .ZN(n11984) );
  INV_X1 U15091 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n11982) );
  INV_X1 U15092 ( .A(n14083), .ZN(n11981) );
  OAI22_X1 U15093 ( .A1(n12343), .A2(n11982), .B1(n11981), .B2(n11951), .ZN(
        n11983) );
  AOI21_X1 U15094 ( .B1(n12338), .B2(n11984), .A(n11983), .ZN(n11985) );
  OAI21_X1 U15095 ( .B1(n15901), .B2(n12340), .A(n11985), .ZN(n14275) );
  INV_X1 U15096 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15829) );
  XNOR2_X1 U15097 ( .A(n11986), .B(n15829), .ZN(n15835) );
  NAND2_X1 U15098 ( .A1(n15835), .A2(n13671), .ZN(n12003) );
  AOI22_X1 U15099 ( .A1(n12323), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11371), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11990) );
  AOI22_X1 U15100 ( .A1(n12144), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12328), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11989) );
  AOI22_X1 U15101 ( .A1(n12248), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11988) );
  AOI22_X1 U15102 ( .A1(n12327), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12326), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11987) );
  NAND4_X1 U15103 ( .A1(n11990), .A2(n11989), .A3(n11988), .A4(n11987), .ZN(
        n11998) );
  AOI22_X1 U15104 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11996) );
  AOI22_X1 U15105 ( .A1(n12316), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12299), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11995) );
  AOI22_X1 U15106 ( .A1(n12324), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12329), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11994) );
  NAND2_X1 U15107 ( .A1(n12317), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11992) );
  NAND2_X1 U15108 ( .A1(n11501), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11991) );
  AND3_X1 U15109 ( .A1(n11992), .A2(n11991), .A3(n12340), .ZN(n11993) );
  NAND4_X1 U15110 ( .A1(n11996), .A2(n11995), .A3(n11994), .A4(n11993), .ZN(
        n11997) );
  OAI21_X1 U15111 ( .B1(n11998), .B2(n11997), .A(n12110), .ZN(n12001) );
  NAND2_X1 U15112 ( .A1(n14084), .A2(P1_EAX_REG_16__SCAN_IN), .ZN(n12000) );
  NAND2_X1 U15113 ( .A1(n20742), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11999) );
  NAND3_X1 U15114 ( .A1(n12001), .A2(n12000), .A3(n11999), .ZN(n12002) );
  NAND2_X1 U15115 ( .A1(n12003), .A2(n12002), .ZN(n14360) );
  INV_X1 U15116 ( .A(n14360), .ZN(n12070) );
  XNOR2_X1 U15117 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n12004), .ZN(
        n15909) );
  INV_X1 U15118 ( .A(n15909), .ZN(n12019) );
  AOI22_X1 U15119 ( .A1(n12248), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12008) );
  AOI22_X1 U15120 ( .A1(n12316), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12327), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12007) );
  AOI22_X1 U15121 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11380), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12006) );
  AOI22_X1 U15122 ( .A1(n12326), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9757), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12005) );
  NAND4_X1 U15123 ( .A1(n12008), .A2(n12007), .A3(n12006), .A4(n12005), .ZN(
        n12014) );
  AOI22_X1 U15124 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12012) );
  AOI22_X1 U15125 ( .A1(n12324), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12144), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12011) );
  AOI22_X1 U15126 ( .A1(n12329), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12328), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12010) );
  AOI22_X1 U15127 ( .A1(n12323), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12317), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12009) );
  NAND4_X1 U15128 ( .A1(n12012), .A2(n12011), .A3(n12010), .A4(n12009), .ZN(
        n12013) );
  OAI21_X1 U15129 ( .B1(n12014), .B2(n12013), .A(n12044), .ZN(n12017) );
  NAND2_X1 U15130 ( .A1(n14084), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12016) );
  NAND2_X1 U15131 ( .A1(n14083), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12015) );
  NAND3_X1 U15132 ( .A1(n12017), .A2(n12016), .A3(n12015), .ZN(n12018) );
  AOI21_X1 U15133 ( .B1(n12019), .B2(n12345), .A(n12018), .ZN(n14369) );
  INV_X1 U15134 ( .A(n14369), .ZN(n12069) );
  XNOR2_X1 U15135 ( .A(n12020), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15848) );
  AOI22_X1 U15136 ( .A1(n12324), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12327), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12024) );
  AOI22_X1 U15137 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12144), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12023) );
  AOI22_X1 U15138 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12328), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12022) );
  AOI22_X1 U15139 ( .A1(n12326), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9772), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12021) );
  NAND4_X1 U15140 ( .A1(n12024), .A2(n12023), .A3(n12022), .A4(n12021), .ZN(
        n12030) );
  AOI22_X1 U15141 ( .A1(n12248), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12323), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12028) );
  AOI22_X1 U15142 ( .A1(n12325), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12316), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12027) );
  AOI22_X1 U15143 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12317), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12026) );
  AOI22_X1 U15144 ( .A1(n12329), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11380), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12025) );
  NAND4_X1 U15145 ( .A1(n12028), .A2(n12027), .A3(n12026), .A4(n12025), .ZN(
        n12029) );
  OAI21_X1 U15146 ( .B1(n12030), .B2(n12029), .A(n12044), .ZN(n12033) );
  NAND2_X1 U15147 ( .A1(n14084), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12032) );
  NAND2_X1 U15148 ( .A1(n14083), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12031) );
  NAND3_X1 U15149 ( .A1(n12033), .A2(n12032), .A3(n12031), .ZN(n12034) );
  AOI21_X1 U15150 ( .B1(n15848), .B2(n12345), .A(n12034), .ZN(n14375) );
  INV_X1 U15151 ( .A(n14375), .ZN(n12068) );
  XNOR2_X1 U15152 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n12035), .ZN(
        n14030) );
  AOI22_X1 U15153 ( .A1(n12316), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12299), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12039) );
  AOI22_X1 U15154 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12329), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12038) );
  AOI22_X1 U15155 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12327), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12037) );
  AOI22_X1 U15156 ( .A1(n12326), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11501), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12036) );
  NAND4_X1 U15157 ( .A1(n12039), .A2(n12038), .A3(n12037), .A4(n12036), .ZN(
        n12046) );
  AOI22_X1 U15158 ( .A1(n12325), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12318), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12043) );
  AOI22_X1 U15159 ( .A1(n12324), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12144), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12042) );
  AOI22_X1 U15160 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12041) );
  AOI22_X1 U15161 ( .A1(n12323), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12317), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12040) );
  NAND4_X1 U15162 ( .A1(n12043), .A2(n12042), .A3(n12041), .A4(n12040), .ZN(
        n12045) );
  OAI21_X1 U15163 ( .B1(n12046), .B2(n12045), .A(n12044), .ZN(n12049) );
  NAND2_X1 U15164 ( .A1(n14084), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n12048) );
  NAND2_X1 U15165 ( .A1(n14083), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12047) );
  AND3_X1 U15166 ( .A1(n12049), .A2(n12048), .A3(n12047), .ZN(n12050) );
  OAI21_X1 U15167 ( .B1(n14030), .B2(n12340), .A(n12050), .ZN(n14008) );
  INV_X1 U15168 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n12067) );
  AOI22_X1 U15169 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12248), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12054) );
  AOI22_X1 U15170 ( .A1(n12316), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12328), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12053) );
  AOI22_X1 U15171 ( .A1(n12329), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12052) );
  AOI22_X1 U15172 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12317), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12051) );
  NAND4_X1 U15173 ( .A1(n12054), .A2(n12053), .A3(n12052), .A4(n12051), .ZN(
        n12060) );
  AOI22_X1 U15174 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12323), .B1(
        n12324), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12058) );
  AOI22_X1 U15175 ( .A1(n12325), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12327), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12057) );
  AOI22_X1 U15176 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12299), .B1(
        n12144), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12056) );
  AOI22_X1 U15177 ( .A1(n12326), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9757), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12055) );
  NAND4_X1 U15178 ( .A1(n12058), .A2(n12057), .A3(n12056), .A4(n12055), .ZN(
        n12059) );
  NOR2_X1 U15179 ( .A1(n12060), .A2(n12059), .ZN(n12061) );
  OR2_X1 U15180 ( .A1(n12062), .A2(n12061), .ZN(n12066) );
  XNOR2_X1 U15181 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n12063), .ZN(
        n15918) );
  INV_X1 U15182 ( .A(n15918), .ZN(n12064) );
  AOI22_X1 U15183 ( .A1(n14083), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n12345), .B2(n12064), .ZN(n12065) );
  OAI211_X1 U15184 ( .C1(n12067), .C2(n12343), .A(n12066), .B(n12065), .ZN(
        n14385) );
  AND2_X1 U15185 ( .A1(n14008), .A2(n14385), .ZN(n14007) );
  AND2_X1 U15186 ( .A1(n12068), .A2(n14007), .ZN(n14366) );
  AOI22_X1 U15187 ( .A1(n12316), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12324), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12076) );
  AOI22_X1 U15188 ( .A1(n12323), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12075) );
  AOI22_X1 U15189 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12329), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12074) );
  AOI22_X1 U15190 ( .A1(n12325), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12144), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12073) );
  NAND4_X1 U15191 ( .A1(n12076), .A2(n12075), .A3(n12074), .A4(n12073), .ZN(
        n12082) );
  AOI22_X1 U15192 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12327), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12080) );
  AOI22_X1 U15193 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11380), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12079) );
  AOI22_X1 U15194 ( .A1(n12326), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9757), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12078) );
  AOI22_X1 U15195 ( .A1(n12248), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12317), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12077) );
  NAND4_X1 U15196 ( .A1(n12080), .A2(n12079), .A3(n12078), .A4(n12077), .ZN(
        n12081) );
  NOR2_X1 U15197 ( .A1(n12082), .A2(n12081), .ZN(n12087) );
  INV_X1 U15198 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n12084) );
  NAND2_X1 U15199 ( .A1(n20742), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12083) );
  OAI211_X1 U15200 ( .C1(n12343), .C2(n12084), .A(n12340), .B(n12083), .ZN(
        n12085) );
  INV_X1 U15201 ( .A(n12085), .ZN(n12086) );
  OAI21_X1 U15202 ( .B1(n12310), .B2(n12087), .A(n12086), .ZN(n12095) );
  INV_X1 U15203 ( .A(n12132), .ZN(n12093) );
  INV_X1 U15204 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n12091) );
  INV_X1 U15205 ( .A(n12089), .ZN(n12090) );
  NAND2_X1 U15206 ( .A1(n12091), .A2(n12090), .ZN(n12092) );
  NAND2_X1 U15207 ( .A1(n12093), .A2(n12092), .ZN(n15892) );
  NAND2_X1 U15208 ( .A1(n12095), .A2(n12094), .ZN(n14346) );
  AOI22_X1 U15209 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12102) );
  AOI22_X1 U15210 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12327), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12101) );
  AOI22_X1 U15211 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12317), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12100) );
  NAND2_X1 U15212 ( .A1(n12323), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n12098) );
  AOI21_X1 U15213 ( .B1(n9757), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A(n13671), .ZN(n12097) );
  AND2_X1 U15214 ( .A1(n12098), .A2(n12097), .ZN(n12099) );
  NAND4_X1 U15215 ( .A1(n12102), .A2(n12101), .A3(n12100), .A4(n12099), .ZN(
        n12108) );
  AOI22_X1 U15216 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n12316), .B1(
        n12329), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12106) );
  AOI22_X1 U15217 ( .A1(n12324), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12144), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12105) );
  AOI22_X1 U15218 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n12248), .B1(
        n11380), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12104) );
  AOI22_X1 U15219 ( .A1(n12325), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12326), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12103) );
  NAND4_X1 U15220 ( .A1(n12106), .A2(n12105), .A3(n12104), .A4(n12103), .ZN(
        n12107) );
  OR2_X1 U15221 ( .A1(n12108), .A2(n12107), .ZN(n12109) );
  NAND2_X1 U15222 ( .A1(n12110), .A2(n12109), .ZN(n12115) );
  INV_X1 U15223 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n12111) );
  INV_X1 U15224 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15807) );
  OAI22_X1 U15225 ( .A1(n12343), .A2(n12111), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15807), .ZN(n12112) );
  INV_X1 U15226 ( .A(n12112), .ZN(n12114) );
  XNOR2_X1 U15227 ( .A(n12132), .B(n15807), .ZN(n15798) );
  AND2_X1 U15228 ( .A1(n15798), .A2(n12345), .ZN(n12113) );
  AOI21_X1 U15229 ( .B1(n12115), .B2(n12114), .A(n12113), .ZN(n14343) );
  AOI22_X1 U15230 ( .A1(n12323), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12120) );
  AOI22_X1 U15231 ( .A1(n12325), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12329), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12119) );
  AOI22_X1 U15232 ( .A1(n12316), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11380), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12118) );
  AOI22_X1 U15233 ( .A1(n12248), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12317), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12117) );
  NAND4_X1 U15234 ( .A1(n12120), .A2(n12119), .A3(n12118), .A4(n12117), .ZN(
        n12126) );
  AOI22_X1 U15235 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12324), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12124) );
  AOI22_X1 U15236 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12327), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12123) );
  AOI22_X1 U15237 ( .A1(n12144), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12328), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12122) );
  AOI22_X1 U15238 ( .A1(n12326), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9757), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12121) );
  NAND4_X1 U15239 ( .A1(n12124), .A2(n12123), .A3(n12122), .A4(n12121), .ZN(
        n12125) );
  NOR2_X1 U15240 ( .A1(n12126), .A2(n12125), .ZN(n12131) );
  INV_X1 U15241 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n12128) );
  NAND2_X1 U15242 ( .A1(n20742), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12127) );
  OAI211_X1 U15243 ( .C1(n12343), .C2(n12128), .A(n12340), .B(n12127), .ZN(
        n12129) );
  INV_X1 U15244 ( .A(n12129), .ZN(n12130) );
  OAI21_X1 U15245 ( .B1(n12310), .B2(n12131), .A(n12130), .ZN(n12138) );
  INV_X1 U15246 ( .A(n12133), .ZN(n12135) );
  INV_X1 U15247 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12134) );
  NAND2_X1 U15248 ( .A1(n12135), .A2(n12134), .ZN(n12136) );
  NAND2_X1 U15249 ( .A1(n12156), .A2(n12136), .ZN(n15797) );
  NAND2_X1 U15250 ( .A1(n14334), .A2(n14335), .ZN(n14328) );
  AOI22_X1 U15251 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12329), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12143) );
  AOI22_X1 U15252 ( .A1(n11372), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12324), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12142) );
  AOI22_X1 U15253 ( .A1(n12326), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9772), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12141) );
  AOI22_X1 U15254 ( .A1(n12323), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12140) );
  NAND4_X1 U15255 ( .A1(n12143), .A2(n12142), .A3(n12141), .A4(n12140), .ZN(
        n12150) );
  AOI22_X1 U15256 ( .A1(n12248), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12327), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12148) );
  AOI22_X1 U15257 ( .A1(n12325), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12144), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12147) );
  AOI22_X1 U15258 ( .A1(n12316), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12328), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12146) );
  AOI22_X1 U15259 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12317), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12145) );
  NAND4_X1 U15260 ( .A1(n12148), .A2(n12147), .A3(n12146), .A4(n12145), .ZN(
        n12149) );
  NOR2_X1 U15261 ( .A1(n12150), .A2(n12149), .ZN(n12153) );
  INV_X1 U15262 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15779) );
  AOI21_X1 U15263 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15779), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12151) );
  AOI21_X1 U15264 ( .B1(n14084), .B2(P1_EAX_REG_22__SCAN_IN), .A(n12151), .ZN(
        n12152) );
  OAI21_X1 U15265 ( .B1(n12310), .B2(n12153), .A(n12152), .ZN(n12155) );
  XNOR2_X1 U15266 ( .A(n12156), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15783) );
  NAND2_X1 U15267 ( .A1(n15783), .A2(n13671), .ZN(n12154) );
  NAND2_X1 U15268 ( .A1(n12155), .A2(n12154), .ZN(n14329) );
  INV_X1 U15269 ( .A(n12156), .ZN(n12157) );
  NAND2_X1 U15270 ( .A1(n12158), .A2(n14265), .ZN(n12159) );
  NAND2_X1 U15271 ( .A1(n12184), .A2(n12159), .ZN(n14499) );
  AOI22_X1 U15272 ( .A1(n12323), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12299), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12163) );
  AOI22_X1 U15273 ( .A1(n12316), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12329), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12162) );
  AOI22_X1 U15274 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12144), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12161) );
  AOI22_X1 U15275 ( .A1(n12326), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9757), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12160) );
  NAND4_X1 U15276 ( .A1(n12163), .A2(n12162), .A3(n12161), .A4(n12160), .ZN(
        n12169) );
  AOI22_X1 U15277 ( .A1(n12325), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12327), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12167) );
  AOI22_X1 U15278 ( .A1(n12324), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12328), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12166) );
  AOI22_X1 U15279 ( .A1(n12318), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12165) );
  AOI22_X1 U15280 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12317), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12164) );
  NAND4_X1 U15281 ( .A1(n12167), .A2(n12166), .A3(n12165), .A4(n12164), .ZN(
        n12168) );
  NOR2_X1 U15282 ( .A1(n12169), .A2(n12168), .ZN(n12186) );
  AOI22_X1 U15283 ( .A1(n12325), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12324), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12173) );
  AOI22_X1 U15284 ( .A1(n12316), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12329), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12172) );
  AOI22_X1 U15285 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9772), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12171) );
  AOI22_X1 U15286 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12170) );
  NAND4_X1 U15287 ( .A1(n12173), .A2(n12172), .A3(n12171), .A4(n12170), .ZN(
        n12179) );
  AOI22_X1 U15288 ( .A1(n12318), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12299), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12177) );
  AOI22_X1 U15289 ( .A1(n12144), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12328), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12176) );
  AOI22_X1 U15290 ( .A1(n12327), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12326), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12175) );
  AOI22_X1 U15291 ( .A1(n12323), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12317), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12174) );
  NAND4_X1 U15292 ( .A1(n12177), .A2(n12176), .A3(n12175), .A4(n12174), .ZN(
        n12178) );
  NOR2_X1 U15293 ( .A1(n12179), .A2(n12178), .ZN(n12185) );
  XNOR2_X1 U15294 ( .A(n12186), .B(n12185), .ZN(n12182) );
  OAI21_X1 U15295 ( .B1(n20643), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n20742), .ZN(n12181) );
  NAND2_X1 U15296 ( .A1(n14084), .A2(P1_EAX_REG_23__SCAN_IN), .ZN(n12180) );
  OAI211_X1 U15297 ( .C1(n12182), .C2(n12310), .A(n12181), .B(n12180), .ZN(
        n12183) );
  OAI21_X1 U15298 ( .B1(n12340), .B2(n14499), .A(n12183), .ZN(n14264) );
  XOR2_X1 U15299 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B(n12201), .Z(
        n14495) );
  INV_X1 U15300 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14491) );
  OAI21_X1 U15301 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n14491), .A(n12340), 
        .ZN(n12199) );
  NOR2_X1 U15302 ( .A1(n12186), .A2(n12185), .ZN(n12216) );
  AOI22_X1 U15303 ( .A1(n12323), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11371), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12190) );
  AOI22_X1 U15304 ( .A1(n12316), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12329), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12189) );
  AOI22_X1 U15305 ( .A1(n11372), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12188) );
  AOI22_X1 U15306 ( .A1(n12318), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12317), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12187) );
  NAND4_X1 U15307 ( .A1(n12190), .A2(n12189), .A3(n12188), .A4(n12187), .ZN(
        n12196) );
  AOI22_X1 U15308 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12194) );
  AOI22_X1 U15309 ( .A1(n12327), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12144), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12193) );
  AOI22_X1 U15310 ( .A1(n12266), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12328), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12192) );
  AOI22_X1 U15311 ( .A1(n12326), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9772), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12191) );
  NAND4_X1 U15312 ( .A1(n12194), .A2(n12193), .A3(n12192), .A4(n12191), .ZN(
        n12195) );
  OR2_X1 U15313 ( .A1(n12196), .A2(n12195), .ZN(n12215) );
  XNOR2_X1 U15314 ( .A(n12216), .B(n12215), .ZN(n12197) );
  NOR2_X1 U15315 ( .A1(n12197), .A2(n12310), .ZN(n12198) );
  AOI211_X1 U15316 ( .C1(n14084), .C2(P1_EAX_REG_24__SCAN_IN), .A(n12199), .B(
        n12198), .ZN(n12200) );
  AOI21_X1 U15317 ( .B1(n12345), .B2(n14495), .A(n12200), .ZN(n14252) );
  NAND2_X1 U15318 ( .A1(n12202), .A2(n21030), .ZN(n12203) );
  NAND2_X1 U15319 ( .A1(n12237), .A2(n12203), .ZN(n14483) );
  AOI22_X1 U15320 ( .A1(n12325), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12324), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12207) );
  AOI22_X1 U15321 ( .A1(n11372), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12328), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12206) );
  AOI22_X1 U15322 ( .A1(n12327), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12326), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12205) );
  AOI22_X1 U15323 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12317), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12204) );
  NAND4_X1 U15324 ( .A1(n12207), .A2(n12206), .A3(n12205), .A4(n12204), .ZN(
        n12214) );
  AOI22_X1 U15325 ( .A1(n12318), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12323), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12212) );
  AOI22_X1 U15326 ( .A1(n12316), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12144), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12211) );
  AOI22_X1 U15327 ( .A1(n12329), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12210) );
  AOI22_X1 U15328 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9772), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12209) );
  NAND4_X1 U15329 ( .A1(n12212), .A2(n12211), .A3(n12210), .A4(n12209), .ZN(
        n12213) );
  NOR2_X1 U15330 ( .A1(n12214), .A2(n12213), .ZN(n12222) );
  NAND2_X1 U15331 ( .A1(n12216), .A2(n12215), .ZN(n12221) );
  XNOR2_X1 U15332 ( .A(n12222), .B(n12221), .ZN(n12219) );
  NOR2_X1 U15333 ( .A1(n21030), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12217) );
  AOI211_X1 U15334 ( .C1(n14084), .C2(P1_EAX_REG_25__SCAN_IN), .A(n13671), .B(
        n12217), .ZN(n12218) );
  OAI21_X1 U15335 ( .B1(n12219), .B2(n12310), .A(n12218), .ZN(n12220) );
  OAI21_X1 U15336 ( .B1(n12340), .B2(n14483), .A(n12220), .ZN(n14240) );
  XNOR2_X1 U15337 ( .A(n12237), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14475) );
  INV_X1 U15338 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14471) );
  OAI21_X1 U15339 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n14471), .A(n12340), 
        .ZN(n12235) );
  NOR2_X1 U15340 ( .A1(n12222), .A2(n12221), .ZN(n12242) );
  INV_X1 U15341 ( .A(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n20958) );
  AOI22_X1 U15342 ( .A1(n12323), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12226) );
  AOI22_X1 U15343 ( .A1(n12316), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12329), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12225) );
  AOI22_X1 U15344 ( .A1(n11372), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12224) );
  AOI22_X1 U15345 ( .A1(n12318), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12317), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12223) );
  NAND4_X1 U15346 ( .A1(n12226), .A2(n12225), .A3(n12224), .A4(n12223), .ZN(
        n12232) );
  AOI22_X1 U15347 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12230) );
  AOI22_X1 U15348 ( .A1(n12327), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12144), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12229) );
  AOI22_X1 U15349 ( .A1(n12266), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12328), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12228) );
  AOI22_X1 U15350 ( .A1(n12326), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9757), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12227) );
  NAND4_X1 U15351 ( .A1(n12230), .A2(n12229), .A3(n12228), .A4(n12227), .ZN(
        n12231) );
  OR2_X1 U15352 ( .A1(n12232), .A2(n12231), .ZN(n12241) );
  XNOR2_X1 U15353 ( .A(n12242), .B(n12241), .ZN(n12233) );
  NOR2_X1 U15354 ( .A1(n12233), .A2(n12310), .ZN(n12234) );
  AOI211_X1 U15355 ( .C1(n14084), .C2(P1_EAX_REG_26__SCAN_IN), .A(n12235), .B(
        n12234), .ZN(n12236) );
  AOI21_X1 U15356 ( .B1(n12345), .B2(n14475), .A(n12236), .ZN(n14222) );
  INV_X1 U15357 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14214) );
  NAND2_X1 U15358 ( .A1(n12239), .A2(n14214), .ZN(n12240) );
  NAND2_X1 U15359 ( .A1(n12291), .A2(n12240), .ZN(n14464) );
  NAND2_X1 U15360 ( .A1(n12242), .A2(n12241), .ZN(n12260) );
  AOI22_X1 U15361 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n12323), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12247) );
  AOI22_X1 U15362 ( .A1(n12266), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12328), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12246) );
  AOI22_X1 U15363 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12326), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12245) );
  AOI22_X1 U15364 ( .A1(n12329), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12317), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12244) );
  NAND4_X1 U15365 ( .A1(n12247), .A2(n12246), .A3(n12245), .A4(n12244), .ZN(
        n12254) );
  AOI22_X1 U15366 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n12248), .B1(
        n12299), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12252) );
  AOI22_X1 U15367 ( .A1(n12325), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12144), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12251) );
  AOI22_X1 U15368 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12316), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12250) );
  AOI22_X1 U15369 ( .A1(n12327), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11501), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12249) );
  NAND4_X1 U15370 ( .A1(n12252), .A2(n12251), .A3(n12250), .A4(n12249), .ZN(
        n12253) );
  NOR2_X1 U15371 ( .A1(n12254), .A2(n12253), .ZN(n12261) );
  XNOR2_X1 U15372 ( .A(n12260), .B(n12261), .ZN(n12257) );
  OAI21_X1 U15373 ( .B1(n20643), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n20742), .ZN(n12256) );
  NAND2_X1 U15374 ( .A1(n14084), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n12255) );
  OAI211_X1 U15375 ( .C1(n12257), .C2(n12310), .A(n12256), .B(n12255), .ZN(
        n12258) );
  OAI21_X1 U15376 ( .B1(n12340), .B2(n14464), .A(n12258), .ZN(n14212) );
  INV_X1 U15377 ( .A(n12291), .ZN(n12259) );
  XOR2_X1 U15378 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B(n12259), .Z(
        n14203) );
  INV_X1 U15379 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12290) );
  AOI21_X1 U15380 ( .B1(n12290), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12275) );
  NOR2_X1 U15381 ( .A1(n12261), .A2(n12260), .ZN(n12307) );
  AOI22_X1 U15382 ( .A1(n12323), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12265) );
  AOI22_X1 U15383 ( .A1(n12316), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12329), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12264) );
  AOI22_X1 U15384 ( .A1(n11372), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12263) );
  AOI22_X1 U15385 ( .A1(n12318), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12317), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12262) );
  NAND4_X1 U15386 ( .A1(n12265), .A2(n12264), .A3(n12263), .A4(n12262), .ZN(
        n12272) );
  AOI22_X1 U15387 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12270) );
  AOI22_X1 U15388 ( .A1(n12327), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12144), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12269) );
  AOI22_X1 U15389 ( .A1(n12266), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12328), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12268) );
  AOI22_X1 U15390 ( .A1(n12326), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9772), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12267) );
  NAND4_X1 U15391 ( .A1(n12270), .A2(n12269), .A3(n12268), .A4(n12267), .ZN(
        n12271) );
  OR2_X1 U15392 ( .A1(n12272), .A2(n12271), .ZN(n12306) );
  XNOR2_X1 U15393 ( .A(n12307), .B(n12306), .ZN(n12273) );
  NOR2_X1 U15394 ( .A1(n12273), .A2(n12310), .ZN(n12274) );
  AOI211_X1 U15395 ( .C1(n14084), .C2(P1_EAX_REG_28__SCAN_IN), .A(n12275), .B(
        n12274), .ZN(n12276) );
  AOI21_X1 U15396 ( .B1(n12345), .B2(n14203), .A(n12276), .ZN(n12278) );
  OAI21_X1 U15397 ( .B1(n12277), .B2(n12278), .A(n12313), .ZN(n14396) );
  NAND3_X1 U15398 ( .A1(n11495), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16103) );
  INV_X1 U15399 ( .A(n16103), .ZN(n12279) );
  NAND2_X1 U15400 ( .A1(n20836), .A2(n20835), .ZN(n12280) );
  NAND2_X1 U15401 ( .A1(n12280), .A2(n11495), .ZN(n12281) );
  NOR2_X1 U15402 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20742), .ZN(n15740) );
  INV_X1 U15403 ( .A(n15740), .ZN(n12283) );
  NAND2_X1 U15404 ( .A1(n20643), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12282) );
  AND2_X1 U15405 ( .A1(n12283), .A2(n12282), .ZN(n13272) );
  INV_X1 U15406 ( .A(n13272), .ZN(n12284) );
  INV_X1 U15407 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n20802) );
  NOR2_X1 U15408 ( .A1(n16045), .A2(n20802), .ZN(n14587) );
  NOR2_X1 U15409 ( .A1(n14518), .A2(n12290), .ZN(n12285) );
  AOI211_X1 U15410 ( .C1(n15919), .C2(n14203), .A(n14587), .B(n12285), .ZN(
        n12286) );
  INV_X1 U15411 ( .A(n12287), .ZN(n12288) );
  NAND2_X1 U15412 ( .A1(n12289), .A2(n12288), .ZN(P1_U2971) );
  INV_X1 U15413 ( .A(n12292), .ZN(n12293) );
  INV_X1 U15414 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14190) );
  NAND2_X1 U15415 ( .A1(n12293), .A2(n14190), .ZN(n12294) );
  NAND2_X1 U15416 ( .A1(n13674), .A2(n12294), .ZN(n14454) );
  AOI22_X1 U15417 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12327), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12298) );
  AOI22_X1 U15418 ( .A1(n12329), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12144), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12297) );
  AOI22_X1 U15419 ( .A1(n12318), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12296) );
  AOI22_X1 U15420 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12317), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12295) );
  NAND4_X1 U15421 ( .A1(n12298), .A2(n12297), .A3(n12296), .A4(n12295), .ZN(
        n12305) );
  AOI22_X1 U15422 ( .A1(n12323), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12299), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12303) );
  AOI22_X1 U15423 ( .A1(n12325), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12324), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12302) );
  AOI22_X1 U15424 ( .A1(n12326), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9757), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12301) );
  AOI22_X1 U15425 ( .A1(n12316), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12328), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12300) );
  NAND4_X1 U15426 ( .A1(n12303), .A2(n12302), .A3(n12301), .A4(n12300), .ZN(
        n12304) );
  NOR2_X1 U15427 ( .A1(n12305), .A2(n12304), .ZN(n12315) );
  NAND2_X1 U15428 ( .A1(n12307), .A2(n12306), .ZN(n12314) );
  XNOR2_X1 U15429 ( .A(n12315), .B(n12314), .ZN(n12311) );
  AOI21_X1 U15430 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20742), .A(
        n13671), .ZN(n12309) );
  NAND2_X1 U15431 ( .A1(n14084), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n12308) );
  OAI211_X1 U15432 ( .C1(n12311), .C2(n12310), .A(n12309), .B(n12308), .ZN(
        n12312) );
  OAI21_X1 U15433 ( .B1(n12340), .B2(n14454), .A(n12312), .ZN(n14187) );
  NOR2_X1 U15434 ( .A1(n12315), .A2(n12314), .ZN(n12337) );
  AOI22_X1 U15435 ( .A1(n12316), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12144), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12322) );
  AOI22_X1 U15436 ( .A1(n11372), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12321) );
  AOI22_X1 U15437 ( .A1(n12139), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11501), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12320) );
  AOI22_X1 U15438 ( .A1(n12318), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12317), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12319) );
  NAND4_X1 U15439 ( .A1(n12322), .A2(n12321), .A3(n12320), .A4(n12319), .ZN(
        n12335) );
  AOI22_X1 U15440 ( .A1(n12323), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12333) );
  AOI22_X1 U15441 ( .A1(n12325), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12324), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12332) );
  AOI22_X1 U15442 ( .A1(n12327), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12326), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12331) );
  AOI22_X1 U15443 ( .A1(n12329), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12328), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12330) );
  NAND4_X1 U15444 ( .A1(n12333), .A2(n12332), .A3(n12331), .A4(n12330), .ZN(
        n12334) );
  NOR2_X1 U15445 ( .A1(n12335), .A2(n12334), .ZN(n12336) );
  XNOR2_X1 U15446 ( .A(n12337), .B(n12336), .ZN(n12339) );
  NAND2_X1 U15447 ( .A1(n12339), .A2(n12338), .ZN(n12348) );
  INV_X1 U15448 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n12342) );
  NAND2_X1 U15449 ( .A1(n20742), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12341) );
  OAI211_X1 U15450 ( .C1(n12343), .C2(n12342), .A(n12341), .B(n12340), .ZN(
        n12344) );
  INV_X1 U15451 ( .A(n12344), .ZN(n12347) );
  XNOR2_X1 U15452 ( .A(n13674), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14109) );
  AOI21_X1 U15453 ( .B1(n12348), .B2(n12347), .A(n12346), .ZN(n14082) );
  XNOR2_X1 U15454 ( .A(n14186), .B(n10083), .ZN(n14100) );
  INV_X1 U15455 ( .A(n20145), .ZN(n12349) );
  NAND2_X1 U15456 ( .A1(n12349), .A2(n11464), .ZN(n12374) );
  OAI22_X1 U15457 ( .A1(n13247), .A2(n11392), .B1(n11822), .B2(n13685), .ZN(
        n13195) );
  NAND2_X1 U15458 ( .A1(n13225), .A2(n12352), .ZN(n12353) );
  INV_X1 U15459 ( .A(n13317), .ZN(n19899) );
  NAND4_X1 U15460 ( .A1(n14087), .A2(n13244), .A3(n13317), .A4(n11473), .ZN(
        n13315) );
  INV_X2 U15461 ( .A(n10135), .ZN(n14175) );
  NOR3_X1 U15462 ( .A1(n12354), .A2(n13315), .A3(n14175), .ZN(n12356) );
  NAND2_X1 U15463 ( .A1(n14100), .A2(n19996), .ZN(n12466) );
  INV_X1 U15464 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n12358) );
  INV_X1 U15465 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20090) );
  NAND2_X1 U15466 ( .A1(n12374), .A2(n20090), .ZN(n12360) );
  NAND2_X1 U15467 ( .A1(n10135), .A2(n12358), .ZN(n12359) );
  NAND3_X1 U15468 ( .A1(n12360), .A2(n9787), .A3(n12359), .ZN(n12361) );
  NAND2_X1 U15469 ( .A1(n12374), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12362) );
  OAI21_X1 U15470 ( .B1(n12448), .B2(P1_EBX_REG_0__SCAN_IN), .A(n12362), .ZN(
        n13248) );
  XNOR2_X1 U15471 ( .A(n12363), .B(n13248), .ZN(n13460) );
  NAND2_X1 U15472 ( .A1(n13460), .A2(n13459), .ZN(n13461) );
  NAND2_X1 U15473 ( .A1(n13461), .A2(n12363), .ZN(n13456) );
  INV_X1 U15474 ( .A(n13456), .ZN(n12370) );
  INV_X1 U15475 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n12364) );
  NAND2_X1 U15476 ( .A1(n12441), .A2(n12364), .ZN(n12368) );
  NAND2_X1 U15477 ( .A1(n12452), .A2(n20082), .ZN(n12366) );
  NAND2_X1 U15478 ( .A1(n13459), .A2(n12364), .ZN(n12365) );
  NAND3_X1 U15479 ( .A1(n12366), .A2(n9787), .A3(n12365), .ZN(n12367) );
  AND2_X1 U15480 ( .A1(n12368), .A2(n12367), .ZN(n13455) );
  INV_X1 U15481 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n12371) );
  NAND2_X1 U15482 ( .A1(n13459), .A2(n12371), .ZN(n12372) );
  OAI211_X1 U15483 ( .C1(n12448), .C2(n20069), .A(n12372), .B(n12452), .ZN(
        n12373) );
  OAI21_X1 U15484 ( .B1(n12437), .B2(P1_EBX_REG_3__SCAN_IN), .A(n12373), .ZN(
        n13467) );
  MUX2_X1 U15485 ( .A(n12456), .B(n12452), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n12378) );
  INV_X1 U15486 ( .A(n12374), .ZN(n12375) );
  NAND2_X1 U15487 ( .A1(n12375), .A2(n14175), .ZN(n12430) );
  NAND2_X1 U15488 ( .A1(n14175), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12376) );
  AND2_X1 U15489 ( .A1(n12430), .A2(n12376), .ZN(n12377) );
  NAND2_X1 U15490 ( .A1(n12378), .A2(n12377), .ZN(n13569) );
  INV_X1 U15491 ( .A(n16090), .ZN(n12382) );
  INV_X1 U15492 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n19999) );
  NAND2_X1 U15493 ( .A1(n13459), .A2(n19999), .ZN(n12379) );
  OAI211_X1 U15494 ( .C1(n12448), .C2(n16060), .A(n12379), .B(n12452), .ZN(
        n12380) );
  OAI21_X1 U15495 ( .B1(n12437), .B2(P1_EBX_REG_5__SCAN_IN), .A(n12380), .ZN(
        n16089) );
  MUX2_X1 U15496 ( .A(n12456), .B(n12452), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n12385) );
  NAND2_X1 U15497 ( .A1(n14175), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12383) );
  AND2_X1 U15498 ( .A1(n12430), .A2(n12383), .ZN(n12384) );
  AND2_X1 U15499 ( .A1(n12385), .A2(n12384), .ZN(n13730) );
  INV_X1 U15500 ( .A(n12437), .ZN(n12446) );
  INV_X1 U15501 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n19993) );
  NAND2_X1 U15502 ( .A1(n12446), .A2(n19993), .ZN(n12388) );
  NAND2_X1 U15503 ( .A1(n13459), .A2(n19993), .ZN(n12386) );
  OAI211_X1 U15504 ( .C1(n12448), .C2(n16082), .A(n12386), .B(n12452), .ZN(
        n12387) );
  MUX2_X1 U15505 ( .A(n12456), .B(n12452), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n12391) );
  NAND2_X1 U15506 ( .A1(n14175), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12389) );
  AND2_X1 U15507 ( .A1(n12430), .A2(n12389), .ZN(n12390) );
  NAND2_X1 U15508 ( .A1(n12391), .A2(n12390), .ZN(n13791) );
  INV_X1 U15509 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n19990) );
  NAND2_X1 U15510 ( .A1(n13459), .A2(n19990), .ZN(n12392) );
  OAI211_X1 U15511 ( .C1(n12448), .C2(n16059), .A(n12392), .B(n12452), .ZN(
        n12393) );
  OAI21_X1 U15512 ( .B1(n12437), .B2(P1_EBX_REG_9__SCAN_IN), .A(n12393), .ZN(
        n16051) );
  INV_X1 U15513 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n13912) );
  NAND2_X1 U15514 ( .A1(n12441), .A2(n13912), .ZN(n12399) );
  INV_X1 U15515 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14557) );
  NAND2_X1 U15516 ( .A1(n12452), .A2(n14557), .ZN(n12397) );
  NAND2_X1 U15517 ( .A1(n13459), .A2(n13912), .ZN(n12396) );
  NAND3_X1 U15518 ( .A1(n12397), .A2(n9787), .A3(n12396), .ZN(n12398) );
  INV_X1 U15519 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16021) );
  INV_X1 U15520 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15879) );
  NAND2_X1 U15521 ( .A1(n13459), .A2(n15879), .ZN(n12400) );
  OAI211_X1 U15522 ( .C1(n12448), .C2(n16021), .A(n12400), .B(n12452), .ZN(
        n12401) );
  OAI21_X1 U15523 ( .B1(n12437), .B2(P1_EBX_REG_11__SCAN_IN), .A(n12401), .ZN(
        n15868) );
  MUX2_X1 U15524 ( .A(n12456), .B(n12452), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n12404) );
  NAND2_X1 U15525 ( .A1(n14175), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12402) );
  AND2_X1 U15526 ( .A1(n12430), .A2(n12402), .ZN(n12403) );
  NAND2_X1 U15527 ( .A1(n12404), .A2(n12403), .ZN(n14383) );
  NAND2_X1 U15528 ( .A1(n15866), .A2(n14383), .ZN(n14022) );
  INV_X1 U15529 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n14031) );
  NAND2_X1 U15530 ( .A1(n13459), .A2(n14031), .ZN(n12405) );
  OAI211_X1 U15531 ( .C1(n12448), .C2(n16017), .A(n12405), .B(n12452), .ZN(
        n12406) );
  OAI21_X1 U15532 ( .B1(n12437), .B2(P1_EBX_REG_13__SCAN_IN), .A(n12406), .ZN(
        n14023) );
  OR2_X2 U15533 ( .A1(n14022), .A2(n14023), .ZN(n14380) );
  NAND2_X1 U15534 ( .A1(n13247), .A2(n11740), .ZN(n12408) );
  MUX2_X1 U15535 ( .A(n12437), .B(n9787), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n12407) );
  AND2_X1 U15536 ( .A1(n12408), .A2(n12407), .ZN(n14370) );
  INV_X1 U15537 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n15845) );
  NAND2_X1 U15538 ( .A1(n12441), .A2(n15845), .ZN(n12412) );
  NAND2_X1 U15539 ( .A1(n12452), .A2(n16008), .ZN(n12410) );
  NAND2_X1 U15540 ( .A1(n13459), .A2(n15845), .ZN(n12409) );
  NAND3_X1 U15541 ( .A1(n12410), .A2(n9787), .A3(n12409), .ZN(n12411) );
  NAND2_X1 U15542 ( .A1(n12412), .A2(n12411), .ZN(n14379) );
  NAND2_X1 U15543 ( .A1(n14370), .A2(n14379), .ZN(n12413) );
  INV_X1 U15544 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15998) );
  NAND2_X1 U15545 ( .A1(n12452), .A2(n15998), .ZN(n12415) );
  INV_X1 U15546 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14363) );
  NAND2_X1 U15547 ( .A1(n13459), .A2(n14363), .ZN(n12414) );
  NAND3_X1 U15548 ( .A1(n12415), .A2(n9787), .A3(n12414), .ZN(n12416) );
  OAI21_X1 U15549 ( .B1(n12456), .B2(P1_EBX_REG_16__SCAN_IN), .A(n12416), .ZN(
        n14361) );
  INV_X1 U15550 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15984) );
  NAND2_X1 U15551 ( .A1(n13247), .A2(n15984), .ZN(n12418) );
  MUX2_X1 U15552 ( .A(n12437), .B(n9787), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n12417) );
  AND2_X1 U15553 ( .A1(n12418), .A2(n12417), .ZN(n14285) );
  INV_X1 U15554 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n15821) );
  NAND2_X1 U15555 ( .A1(n12441), .A2(n15821), .ZN(n12422) );
  INV_X1 U15556 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15971) );
  NAND2_X1 U15557 ( .A1(n12452), .A2(n15971), .ZN(n12420) );
  NAND2_X1 U15558 ( .A1(n13459), .A2(n15821), .ZN(n12419) );
  NAND3_X1 U15559 ( .A1(n12420), .A2(n9787), .A3(n12419), .ZN(n12421) );
  MUX2_X1 U15560 ( .A(n12437), .B(n9787), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n12423) );
  NAND2_X1 U15561 ( .A1(n10134), .A2(n12423), .ZN(n14348) );
  MUX2_X1 U15562 ( .A(n12456), .B(n12452), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n12426) );
  NAND2_X1 U15563 ( .A1(n14175), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12424) );
  AND2_X1 U15564 ( .A1(n12430), .A2(n12424), .ZN(n12425) );
  NAND2_X1 U15565 ( .A1(n12426), .A2(n12425), .ZN(n14338) );
  NAND2_X1 U15566 ( .A1(n14347), .A2(n14338), .ZN(n14340) );
  MUX2_X1 U15567 ( .A(n12437), .B(n9787), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n12428) );
  NAND2_X1 U15568 ( .A1(n13247), .A2(n11756), .ZN(n12427) );
  NAND2_X1 U15569 ( .A1(n12428), .A2(n12427), .ZN(n14332) );
  MUX2_X1 U15570 ( .A(n12456), .B(n12452), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n12432) );
  NAND2_X1 U15571 ( .A1(n14175), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12429) );
  AND2_X1 U15572 ( .A1(n12430), .A2(n12429), .ZN(n12431) );
  MUX2_X1 U15573 ( .A(n12437), .B(n9787), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n12433) );
  NAND2_X1 U15574 ( .A1(n9866), .A2(n12433), .ZN(n14260) );
  NAND2_X1 U15575 ( .A1(n12452), .A2(n21048), .ZN(n12435) );
  INV_X1 U15576 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14322) );
  NAND2_X1 U15577 ( .A1(n13459), .A2(n14322), .ZN(n12434) );
  NAND3_X1 U15578 ( .A1(n12435), .A2(n9787), .A3(n12434), .ZN(n12436) );
  OAI21_X1 U15579 ( .B1(n12456), .B2(P1_EBX_REG_24__SCAN_IN), .A(n12436), .ZN(
        n14256) );
  NAND2_X1 U15580 ( .A1(n14261), .A2(n14256), .ZN(n14235) );
  MUX2_X1 U15581 ( .A(n12437), .B(n9787), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n12439) );
  NAND2_X1 U15582 ( .A1(n13247), .A2(n13995), .ZN(n12438) );
  NAND2_X1 U15583 ( .A1(n12439), .A2(n12438), .ZN(n14236) );
  NOR2_X2 U15584 ( .A1(n14235), .A2(n14236), .ZN(n12440) );
  INV_X1 U15585 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14320) );
  NAND2_X1 U15586 ( .A1(n12441), .A2(n14320), .ZN(n12445) );
  NAND2_X1 U15587 ( .A1(n12452), .A2(n14606), .ZN(n12443) );
  NAND2_X1 U15588 ( .A1(n13459), .A2(n14320), .ZN(n12442) );
  NAND3_X1 U15589 ( .A1(n12443), .A2(n9787), .A3(n12442), .ZN(n12444) );
  INV_X1 U15590 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14319) );
  NAND2_X1 U15591 ( .A1(n12446), .A2(n14319), .ZN(n12450) );
  INV_X1 U15592 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14599) );
  NAND2_X1 U15593 ( .A1(n13459), .A2(n14319), .ZN(n12447) );
  OAI211_X1 U15594 ( .C1(n12448), .C2(n14599), .A(n12447), .B(n12452), .ZN(
        n12449) );
  NAND2_X1 U15595 ( .A1(n12452), .A2(n12451), .ZN(n12454) );
  INV_X1 U15596 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14318) );
  NAND2_X1 U15597 ( .A1(n13459), .A2(n14318), .ZN(n12453) );
  NAND3_X1 U15598 ( .A1(n12454), .A2(n9787), .A3(n12453), .ZN(n12455) );
  OAI21_X1 U15599 ( .B1(n12456), .B2(P1_EBX_REG_28__SCAN_IN), .A(n12455), .ZN(
        n14197) );
  INV_X1 U15600 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n12457) );
  NAND2_X1 U15601 ( .A1(n13459), .A2(n12457), .ZN(n12458) );
  OAI21_X1 U15602 ( .B1(n14176), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n12458), .ZN(n12459) );
  MUX2_X1 U15603 ( .A(n12458), .B(n12459), .S(n9787), .Z(n14189) );
  NOR2_X2 U15604 ( .A1(n14199), .A2(n14189), .ZN(n14188) );
  OAI22_X1 U15605 ( .A1(n14188), .A2(n9787), .B1(n12459), .B2(n14199), .ZN(
        n12462) );
  INV_X1 U15606 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14567) );
  NOR2_X1 U15607 ( .A1(n13459), .A2(n14567), .ZN(n12461) );
  AOI21_X1 U15608 ( .B1(n14176), .B2(P1_EBX_REG_30__SCAN_IN), .A(n12461), .ZN(
        n14172) );
  XNOR2_X1 U15609 ( .A(n12462), .B(n14172), .ZN(n14114) );
  INV_X1 U15610 ( .A(n14114), .ZN(n12463) );
  INV_X1 U15611 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14112) );
  INV_X1 U15612 ( .A(n12464), .ZN(n12465) );
  XNOR2_X1 U15613 ( .A(n12468), .B(n12470), .ZN(n14040) );
  INV_X1 U15614 ( .A(n12468), .ZN(n12469) );
  AOI22_X1 U15615 ( .A1(n14040), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n12470), .B2(n12469), .ZN(n12474) );
  XNOR2_X1 U15616 ( .A(n12472), .B(n12471), .ZN(n12473) );
  XNOR2_X1 U15617 ( .A(n12474), .B(n12473), .ZN(n12486) );
  NAND2_X1 U15618 ( .A1(n12486), .A2(n16323), .ZN(n12485) );
  NOR2_X2 U15619 ( .A1(n14050), .A2(n15144), .ZN(n15137) );
  XNOR2_X1 U15620 ( .A(n15137), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12492) );
  INV_X1 U15621 ( .A(n14068), .ZN(n15128) );
  NAND2_X1 U15622 ( .A1(n15128), .A2(n15144), .ZN(n15143) );
  NAND2_X1 U15623 ( .A1(n15143), .A2(n15145), .ZN(n15133) );
  AND2_X1 U15624 ( .A1(n9815), .A2(n12475), .ZN(n12476) );
  OR2_X1 U15625 ( .A1(n12476), .A2(n14842), .ZN(n14852) );
  AOI21_X1 U15626 ( .B1(n12477), .B2(n14928), .A(n14914), .ZN(n14922) );
  NOR2_X1 U15627 ( .A1(n18957), .A2(n12478), .ZN(n12487) );
  AOI21_X1 U15628 ( .B1(n19228), .B2(n14922), .A(n12487), .ZN(n12479) );
  OAI21_X1 U15629 ( .B1(n14852), .B2(n16299), .A(n12479), .ZN(n12481) );
  NOR3_X1 U15630 ( .A1(n14068), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n15144), .ZN(n12480) );
  AOI211_X1 U15631 ( .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n15133), .A(
        n12481), .B(n12480), .ZN(n12482) );
  OAI21_X1 U15632 ( .B1(n12492), .B2(n16318), .A(n12482), .ZN(n12483) );
  NAND2_X1 U15633 ( .A1(n12485), .A2(n12484), .ZN(P2_U3018) );
  NAND2_X1 U15634 ( .A1(n12486), .A2(n11305), .ZN(n12495) );
  OAI21_X1 U15635 ( .B1(n14042), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n14678), .ZN(n14722) );
  INV_X1 U15636 ( .A(n14722), .ZN(n12490) );
  AOI21_X1 U15637 ( .B1(n16247), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n12487), .ZN(n12488) );
  OAI21_X1 U15638 ( .B1(n14852), .B2(n13644), .A(n12488), .ZN(n12489) );
  AOI21_X1 U15639 ( .B1(n12490), .B2(n19203), .A(n12489), .ZN(n12491) );
  OAI21_X1 U15640 ( .B1(n12492), .B2(n16265), .A(n12491), .ZN(n12493) );
  INV_X1 U15641 ( .A(n12493), .ZN(n12494) );
  NAND2_X1 U15642 ( .A1(n12495), .A2(n12494), .ZN(P2_U2986) );
  AOI21_X1 U15643 ( .B1(n12498), .B2(n9798), .A(n12497), .ZN(n18926) );
  INV_X1 U15644 ( .A(n18926), .ZN(n12499) );
  OAI22_X1 U15645 ( .A1(n15231), .A2(n12500), .B1(n15346), .B2(n12499), .ZN(
        n12501) );
  INV_X1 U15646 ( .A(n12501), .ZN(n12504) );
  OAI211_X1 U15647 ( .C1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(n15220), .B(n15209), .ZN(
        n12503) );
  NAND3_X1 U15648 ( .A1(n12504), .A2(n12503), .A3(n12502), .ZN(n12505) );
  NAND2_X1 U15649 ( .A1(n12509), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12535) );
  NAND2_X1 U15650 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19415) );
  INV_X1 U15651 ( .A(n19415), .ZN(n12510) );
  NAND2_X1 U15652 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12510), .ZN(
        n12516) );
  INV_X1 U15653 ( .A(n12516), .ZN(n12511) );
  NAND2_X1 U15654 ( .A1(n12511), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19239) );
  OAI211_X1 U15655 ( .C1(n12511), .C2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n19239), .B(n19856), .ZN(n12512) );
  INV_X1 U15656 ( .A(n12512), .ZN(n12513) );
  AOI21_X1 U15657 ( .B1(n12524), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n12513), .ZN(n12515) );
  AND2_X1 U15658 ( .A1(n9790), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12514) );
  NAND2_X1 U15659 ( .A1(n10016), .A2(n9852), .ZN(n12538) );
  INV_X1 U15660 ( .A(n12523), .ZN(n12527) );
  NAND2_X1 U15661 ( .A1(n13265), .A2(n12527), .ZN(n12520) );
  INV_X1 U15662 ( .A(n19856), .ZN(n19513) );
  NAND2_X1 U15663 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19570) );
  NAND2_X1 U15664 ( .A1(n19570), .A2(n19868), .ZN(n12517) );
  NAND2_X1 U15665 ( .A1(n12517), .A2(n12516), .ZN(n13811) );
  NOR2_X1 U15666 ( .A1(n19513), .A2(n13811), .ZN(n12518) );
  AOI21_X1 U15667 ( .B1(n12524), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12518), .ZN(n12519) );
  NAND2_X1 U15668 ( .A1(n12520), .A2(n12519), .ZN(n12532) );
  XNOR2_X1 U15669 ( .A(n12532), .B(n12533), .ZN(n13260) );
  INV_X1 U15670 ( .A(n13260), .ZN(n12531) );
  AOI22_X1 U15671 ( .A1(n12524), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19856), .B2(n19886), .ZN(n12522) );
  NAND2_X1 U15672 ( .A1(n12807), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12529) );
  NAND2_X1 U15673 ( .A1(n12524), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12525) );
  XNOR2_X1 U15674 ( .A(n19877), .B(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n13810) );
  NAND2_X1 U15675 ( .A1(n13810), .A2(n19856), .ZN(n19543) );
  NAND2_X1 U15676 ( .A1(n12525), .A2(n19543), .ZN(n12526) );
  INV_X1 U15677 ( .A(n15355), .ZN(n13165) );
  NAND2_X1 U15678 ( .A1(n13165), .A2(n12529), .ZN(n13261) );
  NAND2_X1 U15679 ( .A1(n12532), .A2(n12533), .ZN(n12534) );
  NAND2_X1 U15680 ( .A1(n13603), .A2(n13605), .ZN(n13604) );
  INV_X1 U15681 ( .A(n12535), .ZN(n12536) );
  NAND2_X1 U15682 ( .A1(n12536), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12537) );
  AND2_X1 U15683 ( .A1(n12538), .A2(n12537), .ZN(n12539) );
  NOR2_X1 U15684 ( .A1(n12541), .A2(n12540), .ZN(n13608) );
  OAI22_X1 U15685 ( .A1(n12689), .A2(n12544), .B1(n12654), .B2(n12543), .ZN(
        n12549) );
  INV_X1 U15686 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12547) );
  NAND2_X1 U15687 ( .A1(n10462), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12546) );
  NAND2_X1 U15688 ( .A1(n10413), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12545) );
  OAI211_X1 U15689 ( .C1(n15402), .C2(n12547), .A(n12546), .B(n12545), .ZN(
        n12548) );
  NOR2_X1 U15690 ( .A1(n12549), .A2(n12548), .ZN(n12560) );
  NAND2_X1 U15691 ( .A1(n10467), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12556) );
  NAND2_X1 U15692 ( .A1(n12695), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12555) );
  AOI22_X1 U15693 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10414), .B1(
        n10400), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12554) );
  INV_X1 U15694 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12551) );
  NAND2_X1 U15695 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n12696), .ZN(
        n12550) );
  OAI21_X1 U15696 ( .B1(n12699), .B2(n12551), .A(n12550), .ZN(n12552) );
  AOI21_X1 U15697 ( .B1(n10500), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A(
        n12552), .ZN(n12553) );
  AND4_X1 U15698 ( .A1(n12556), .A2(n12555), .A3(n12554), .A4(n12553), .ZN(
        n12559) );
  AOI22_X1 U15699 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10395), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12558) );
  AOI22_X1 U15700 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n10456), .B1(
        n10401), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12557) );
  NAND4_X1 U15701 ( .A1(n12560), .A2(n12559), .A3(n12558), .A4(n12557), .ZN(
        n13804) );
  INV_X1 U15702 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12562) );
  INV_X1 U15703 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12561) );
  OAI22_X1 U15704 ( .A1(n12689), .A2(n12562), .B1(n12654), .B2(n12561), .ZN(
        n12567) );
  INV_X1 U15705 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12565) );
  NAND2_X1 U15706 ( .A1(n10462), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12564) );
  NAND2_X1 U15707 ( .A1(n10413), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12563) );
  OAI211_X1 U15708 ( .C1(n12565), .C2(n15402), .A(n12564), .B(n12563), .ZN(
        n12566) );
  NOR2_X1 U15709 ( .A1(n12567), .A2(n12566), .ZN(n12578) );
  NAND2_X1 U15710 ( .A1(n10467), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12574) );
  NAND2_X1 U15711 ( .A1(n12695), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12573) );
  AOI22_X1 U15712 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12572) );
  INV_X1 U15713 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12569) );
  NAND2_X1 U15714 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n12696), .ZN(
        n12568) );
  OAI21_X1 U15715 ( .B1(n12699), .B2(n12569), .A(n12568), .ZN(n12570) );
  AOI21_X1 U15716 ( .B1(n10500), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A(
        n12570), .ZN(n12571) );
  AND4_X1 U15717 ( .A1(n12574), .A2(n12573), .A3(n12572), .A4(n12571), .ZN(
        n12577) );
  AOI22_X1 U15718 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10395), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12576) );
  AOI22_X1 U15719 ( .A1(n10456), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10401), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12575) );
  NAND4_X1 U15720 ( .A1(n12578), .A2(n12577), .A3(n12576), .A4(n12575), .ZN(
        n13773) );
  NOR2_X1 U15721 ( .A1(n13882), .A2(n13782), .ZN(n13827) );
  AND2_X1 U15722 ( .A1(n13829), .A2(n13827), .ZN(n12579) );
  AND2_X1 U15723 ( .A1(n12579), .A2(n13699), .ZN(n13705) );
  NAND2_X1 U15724 ( .A1(n13804), .A2(n13774), .ZN(n12580) );
  NAND2_X1 U15725 ( .A1(n13588), .A2(n13661), .ZN(n13658) );
  INV_X1 U15726 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13580) );
  INV_X1 U15727 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12582) );
  OAI22_X1 U15728 ( .A1(n12689), .A2(n12583), .B1(n12654), .B2(n12582), .ZN(
        n12588) );
  INV_X1 U15729 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12586) );
  NAND2_X1 U15730 ( .A1(n10462), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n12585) );
  NAND2_X1 U15731 ( .A1(n10413), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n12584) );
  OAI211_X1 U15732 ( .C1(n15402), .C2(n12586), .A(n12585), .B(n12584), .ZN(
        n12587) );
  NOR2_X1 U15733 ( .A1(n12588), .A2(n12587), .ZN(n12599) );
  NAND2_X1 U15734 ( .A1(n10467), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n12595) );
  NAND2_X1 U15735 ( .A1(n12695), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n12594) );
  AOI22_X1 U15736 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10414), .B1(
        n10400), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12593) );
  INV_X1 U15737 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12590) );
  NAND2_X1 U15738 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n12696), .ZN(
        n12589) );
  OAI21_X1 U15739 ( .B1(n12699), .B2(n12590), .A(n12589), .ZN(n12591) );
  AOI21_X1 U15740 ( .B1(n10500), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A(
        n12591), .ZN(n12592) );
  AND4_X1 U15741 ( .A1(n12595), .A2(n12594), .A3(n12593), .A4(n12592), .ZN(
        n12598) );
  AOI22_X1 U15742 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10395), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12597) );
  AOI22_X1 U15743 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n10456), .B1(
        n10401), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12596) );
  NAND4_X1 U15744 ( .A1(n12599), .A2(n12598), .A3(n12597), .A4(n12596), .ZN(
        n13838) );
  OAI22_X1 U15745 ( .A1(n12689), .A2(n12601), .B1(n12654), .B2(n12600), .ZN(
        n12606) );
  INV_X1 U15746 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12604) );
  NAND2_X1 U15747 ( .A1(n10462), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n12603) );
  NAND2_X1 U15748 ( .A1(n10413), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n12602) );
  OAI211_X1 U15749 ( .C1(n15402), .C2(n12604), .A(n12603), .B(n12602), .ZN(
        n12605) );
  NOR2_X1 U15750 ( .A1(n12606), .A2(n12605), .ZN(n12617) );
  NAND2_X1 U15751 ( .A1(n10467), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n12613) );
  NAND2_X1 U15752 ( .A1(n12695), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n12612) );
  AOI22_X1 U15753 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10414), .B1(
        n10400), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12611) );
  INV_X1 U15754 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12608) );
  NAND2_X1 U15755 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n12696), .ZN(
        n12607) );
  OAI21_X1 U15756 ( .B1(n12699), .B2(n12608), .A(n12607), .ZN(n12609) );
  AOI21_X1 U15757 ( .B1(n10500), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n12609), .ZN(n12610) );
  AND4_X1 U15758 ( .A1(n12613), .A2(n12612), .A3(n12611), .A4(n12610), .ZN(
        n12616) );
  AOI22_X1 U15759 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10395), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12615) );
  AOI22_X1 U15760 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n10456), .B1(
        n10401), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12614) );
  NAND4_X1 U15761 ( .A1(n12617), .A2(n12616), .A3(n12615), .A4(n12614), .ZN(
        n14906) );
  INV_X1 U15762 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12618) );
  OAI22_X1 U15763 ( .A1(n12689), .A2(n12618), .B1(n12654), .B2(n20888), .ZN(
        n12623) );
  INV_X1 U15764 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12621) );
  NAND2_X1 U15765 ( .A1(n10462), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n12620) );
  NAND2_X1 U15766 ( .A1(n10413), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n12619) );
  OAI211_X1 U15767 ( .C1(n15402), .C2(n12621), .A(n12620), .B(n12619), .ZN(
        n12622) );
  NOR2_X1 U15768 ( .A1(n12623), .A2(n12622), .ZN(n12634) );
  NAND2_X1 U15769 ( .A1(n10467), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n12630) );
  NAND2_X1 U15770 ( .A1(n12695), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12629) );
  AOI22_X1 U15771 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10414), .B1(
        n10400), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12628) );
  INV_X1 U15772 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12625) );
  NAND2_X1 U15773 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n12696), .ZN(
        n12624) );
  OAI21_X1 U15774 ( .B1(n12699), .B2(n12625), .A(n12624), .ZN(n12626) );
  AOI21_X1 U15775 ( .B1(n10500), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A(
        n12626), .ZN(n12627) );
  AND4_X1 U15776 ( .A1(n12630), .A2(n12629), .A3(n12628), .A4(n12627), .ZN(
        n12633) );
  AOI22_X1 U15777 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10395), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12632) );
  AOI22_X1 U15778 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n10456), .B1(
        n10401), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12631) );
  INV_X1 U15779 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12635) );
  OAI22_X1 U15780 ( .A1(n12689), .A2(n12636), .B1(n12654), .B2(n12635), .ZN(
        n12641) );
  NAND2_X1 U15781 ( .A1(n10462), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n12638) );
  NAND2_X1 U15782 ( .A1(n10413), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n12637) );
  OAI211_X1 U15783 ( .C1(n12639), .C2(n15402), .A(n12638), .B(n12637), .ZN(
        n12640) );
  NOR2_X1 U15784 ( .A1(n12641), .A2(n12640), .ZN(n12652) );
  NAND2_X1 U15785 ( .A1(n10467), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n12648) );
  NAND2_X1 U15786 ( .A1(n12695), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n12647) );
  AOI22_X1 U15787 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12646) );
  NAND2_X1 U15788 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n12696), .ZN(
        n12642) );
  OAI21_X1 U15789 ( .B1(n12699), .B2(n12643), .A(n12642), .ZN(n12644) );
  AOI21_X1 U15790 ( .B1(n10500), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A(
        n12644), .ZN(n12645) );
  AND4_X1 U15791 ( .A1(n12648), .A2(n12647), .A3(n12646), .A4(n12645), .ZN(
        n12651) );
  AOI22_X1 U15792 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10395), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12650) );
  AOI22_X1 U15793 ( .A1(n10456), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10401), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12649) );
  NAND4_X1 U15794 ( .A1(n12652), .A2(n12651), .A3(n12650), .A4(n12649), .ZN(
        n14902) );
  INV_X1 U15795 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12653) );
  OAI22_X1 U15796 ( .A1(n12689), .A2(n12655), .B1(n12654), .B2(n12653), .ZN(
        n12660) );
  NAND2_X1 U15797 ( .A1(n10462), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n12657) );
  NAND2_X1 U15798 ( .A1(n10413), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n12656) );
  OAI211_X1 U15799 ( .C1(n15402), .C2(n12658), .A(n12657), .B(n12656), .ZN(
        n12659) );
  NOR2_X1 U15800 ( .A1(n12660), .A2(n12659), .ZN(n12671) );
  NAND2_X1 U15801 ( .A1(n10467), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n12667) );
  NAND2_X1 U15802 ( .A1(n12695), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n12666) );
  AOI22_X1 U15803 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10400), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12665) );
  NAND2_X1 U15804 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n12696), .ZN(
        n12661) );
  OAI21_X1 U15805 ( .B1(n12699), .B2(n12662), .A(n12661), .ZN(n12663) );
  AOI21_X1 U15806 ( .B1(n10500), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n12663), .ZN(n12664) );
  AND4_X1 U15807 ( .A1(n12667), .A2(n12666), .A3(n12665), .A4(n12664), .ZN(
        n12670) );
  AOI22_X1 U15808 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10395), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12669) );
  AOI22_X1 U15809 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n10456), .B1(
        n10401), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12668) );
  NAND4_X1 U15810 ( .A1(n12671), .A2(n12670), .A3(n12669), .A4(n12668), .ZN(
        n14891) );
  INV_X1 U15811 ( .A(n12862), .ZN(n12842) );
  INV_X1 U15812 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13825) );
  NAND2_X1 U15813 ( .A1(n9795), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12674) );
  AND2_X1 U15814 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12673) );
  OR2_X1 U15815 ( .A1(n12673), .A2(n12672), .ZN(n12864) );
  OAI211_X1 U15816 ( .C1(n12842), .C2(n13825), .A(n12674), .B(n12864), .ZN(
        n12675) );
  INV_X1 U15817 ( .A(n12675), .ZN(n12679) );
  AOI22_X1 U15818 ( .A1(n9759), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(n9749), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12678) );
  AOI22_X1 U15819 ( .A1(n9752), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12861), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12677) );
  AOI22_X1 U15820 ( .A1(n12863), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12838), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12676) );
  NAND4_X1 U15821 ( .A1(n12679), .A2(n12678), .A3(n12677), .A4(n12676), .ZN(
        n12687) );
  AOI22_X1 U15822 ( .A1(n9795), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12863), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12685) );
  AOI22_X1 U15823 ( .A1(n9751), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(n9748), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12684) );
  AOI22_X1 U15824 ( .A1(n9759), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12861), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12683) );
  INV_X1 U15825 ( .A(n12864), .ZN(n12840) );
  NAND2_X1 U15826 ( .A1(n12862), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12680) );
  AND3_X1 U15827 ( .A1(n12840), .A2(n12681), .A3(n12680), .ZN(n12682) );
  NAND4_X1 U15828 ( .A1(n12685), .A2(n12684), .A3(n12683), .A4(n12682), .ZN(
        n12686) );
  NAND2_X1 U15829 ( .A1(n12687), .A2(n12686), .ZN(n12736) );
  NOR2_X1 U15830 ( .A1(n9788), .A2(n12736), .ZN(n12711) );
  OR2_X1 U15831 ( .A1(n12689), .A2(n12688), .ZN(n12694) );
  AOI22_X1 U15832 ( .A1(n10462), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10400), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12693) );
  NAND2_X1 U15833 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12692) );
  NAND2_X1 U15834 ( .A1(n10456), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n12691) );
  AND4_X1 U15835 ( .A1(n12694), .A2(n12693), .A3(n12692), .A4(n12691), .ZN(
        n12710) );
  AOI22_X1 U15836 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10500), .B1(
        n10413), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12704) );
  NAND2_X1 U15837 ( .A1(n10467), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n12703) );
  NAND2_X1 U15838 ( .A1(n12695), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n12702) );
  INV_X1 U15839 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12698) );
  NAND2_X1 U15840 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n12696), .ZN(
        n12697) );
  OAI21_X1 U15841 ( .B1(n12699), .B2(n12698), .A(n12697), .ZN(n12700) );
  AOI21_X1 U15842 ( .B1(n10414), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n12700), .ZN(n12701) );
  AND4_X1 U15843 ( .A1(n12704), .A2(n12703), .A3(n12702), .A4(n12701), .ZN(
        n12709) );
  AOI22_X1 U15844 ( .A1(n12705), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10401), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12708) );
  AOI22_X1 U15845 ( .A1(n10395), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12706), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12707) );
  NAND4_X1 U15846 ( .A1(n12710), .A2(n12709), .A3(n12708), .A4(n12707), .ZN(
        n12716) );
  XNOR2_X1 U15847 ( .A(n12711), .B(n12716), .ZN(n12737) );
  INV_X1 U15848 ( .A(n12736), .ZN(n12715) );
  NAND2_X1 U15849 ( .A1(n9788), .A2(n12715), .ZN(n14883) );
  INV_X1 U15850 ( .A(n12712), .ZN(n14892) );
  INV_X1 U15851 ( .A(n12737), .ZN(n12713) );
  NAND2_X1 U15852 ( .A1(n12716), .A2(n12715), .ZN(n12739) );
  INV_X1 U15853 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12718) );
  NAND2_X1 U15854 ( .A1(n12863), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12717) );
  OAI211_X1 U15855 ( .C1(n12842), .C2(n12718), .A(n12717), .B(n12864), .ZN(
        n12719) );
  INV_X1 U15856 ( .A(n12719), .ZN(n12724) );
  AOI22_X1 U15857 ( .A1(n9753), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(n9748), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12723) );
  AOI22_X1 U15858 ( .A1(n9759), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12861), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12722) );
  NAND4_X1 U15859 ( .A1(n12724), .A2(n12723), .A3(n12722), .A4(n12721), .ZN(
        n12733) );
  NAND2_X1 U15860 ( .A1(n12863), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12725) );
  OAI211_X1 U15861 ( .C1(n12842), .C2(n12726), .A(n12725), .B(n12840), .ZN(
        n12727) );
  INV_X1 U15862 ( .A(n12727), .ZN(n12731) );
  AOI22_X1 U15863 ( .A1(n9751), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(n9750), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12730) );
  AOI22_X1 U15864 ( .A1(n9759), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12861), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12729) );
  AOI22_X1 U15865 ( .A1(n12720), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12838), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12728) );
  NAND4_X1 U15866 ( .A1(n12731), .A2(n12730), .A3(n12729), .A4(n12728), .ZN(
        n12732) );
  NAND2_X1 U15867 ( .A1(n12733), .A2(n12732), .ZN(n12735) );
  XOR2_X1 U15868 ( .A(n12739), .B(n12735), .Z(n12734) );
  NAND2_X1 U15869 ( .A1(n12734), .A2(n12807), .ZN(n14875) );
  INV_X1 U15870 ( .A(n12735), .ZN(n12740) );
  NAND2_X1 U15871 ( .A1(n9788), .A2(n12740), .ZN(n14877) );
  NOR3_X1 U15872 ( .A1(n12737), .A2(n12736), .A3(n14877), .ZN(n12738) );
  INV_X1 U15873 ( .A(n12739), .ZN(n12741) );
  AND2_X1 U15874 ( .A1(n12741), .A2(n12740), .ZN(n12758) );
  INV_X1 U15875 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12743) );
  NAND2_X1 U15876 ( .A1(n12863), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n12742) );
  OAI211_X1 U15877 ( .C1(n12842), .C2(n12743), .A(n12742), .B(n12864), .ZN(
        n12744) );
  INV_X1 U15878 ( .A(n12744), .ZN(n12748) );
  AOI22_X1 U15879 ( .A1(n9753), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(n9750), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12747) );
  AOI22_X1 U15880 ( .A1(n9759), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12861), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12746) );
  NAND4_X1 U15881 ( .A1(n12748), .A2(n12747), .A3(n12746), .A4(n12745), .ZN(
        n12757) );
  INV_X1 U15882 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12750) );
  NAND2_X1 U15883 ( .A1(n12863), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n12749) );
  OAI211_X1 U15884 ( .C1(n12842), .C2(n12750), .A(n12749), .B(n12840), .ZN(
        n12751) );
  INV_X1 U15885 ( .A(n12751), .ZN(n12755) );
  AOI22_X1 U15886 ( .A1(n9752), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(n9749), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12754) );
  AOI22_X1 U15887 ( .A1(n9759), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12861), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12753) );
  NAND4_X1 U15888 ( .A1(n12755), .A2(n12754), .A3(n12753), .A4(n12752), .ZN(
        n12756) );
  AND2_X1 U15889 ( .A1(n12757), .A2(n12756), .ZN(n12760) );
  NAND2_X1 U15890 ( .A1(n12758), .A2(n12760), .ZN(n12802) );
  OAI211_X1 U15891 ( .C1(n12758), .C2(n12760), .A(n12807), .B(n12802), .ZN(
        n12763) );
  XNOR2_X1 U15892 ( .A(n12762), .B(n12759), .ZN(n14871) );
  INV_X1 U15893 ( .A(n12760), .ZN(n12761) );
  NOR2_X1 U15894 ( .A1(n9790), .A2(n12761), .ZN(n14870) );
  NAND2_X1 U15895 ( .A1(n14871), .A2(n14870), .ZN(n14869) );
  INV_X1 U15896 ( .A(n12762), .ZN(n12764) );
  NAND2_X1 U15897 ( .A1(n12863), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n12766) );
  OAI211_X1 U15898 ( .C1(n12842), .C2(n12767), .A(n12766), .B(n12864), .ZN(
        n12768) );
  INV_X1 U15899 ( .A(n12768), .ZN(n12772) );
  AOI22_X1 U15900 ( .A1(n9752), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(n9749), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12771) );
  AOI22_X1 U15901 ( .A1(n9759), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12861), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12770) );
  NAND4_X1 U15902 ( .A1(n12772), .A2(n12771), .A3(n12770), .A4(n12769), .ZN(
        n12781) );
  NAND2_X1 U15903 ( .A1(n12863), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n12773) );
  OAI211_X1 U15904 ( .C1(n12842), .C2(n12774), .A(n12773), .B(n12840), .ZN(
        n12775) );
  INV_X1 U15905 ( .A(n12775), .ZN(n12779) );
  AOI22_X1 U15906 ( .A1(n9751), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(n9748), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12778) );
  AOI22_X1 U15907 ( .A1(n9759), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12861), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12777) );
  NAND4_X1 U15908 ( .A1(n12779), .A2(n12778), .A3(n12777), .A4(n12776), .ZN(
        n12780) );
  AND2_X1 U15909 ( .A1(n12781), .A2(n12780), .ZN(n12803) );
  XNOR2_X1 U15910 ( .A(n12802), .B(n12803), .ZN(n12782) );
  INV_X1 U15911 ( .A(n14866), .ZN(n12784) );
  NAND2_X1 U15912 ( .A1(n9788), .A2(n12803), .ZN(n14865) );
  INV_X1 U15913 ( .A(n14865), .ZN(n12783) );
  INV_X1 U15914 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12787) );
  NAND2_X1 U15915 ( .A1(n12863), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n12786) );
  OAI211_X1 U15916 ( .C1(n12842), .C2(n12787), .A(n12786), .B(n12864), .ZN(
        n12788) );
  INV_X1 U15917 ( .A(n12788), .ZN(n12792) );
  AOI22_X1 U15918 ( .A1(n9753), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(n9750), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12791) );
  AOI22_X1 U15919 ( .A1(n9759), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12861), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12790) );
  NAND4_X1 U15920 ( .A1(n12792), .A2(n12791), .A3(n12790), .A4(n12789), .ZN(
        n12801) );
  NAND2_X1 U15921 ( .A1(n12863), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12793) );
  OAI211_X1 U15922 ( .C1(n12842), .C2(n12794), .A(n12793), .B(n12840), .ZN(
        n12795) );
  INV_X1 U15923 ( .A(n12795), .ZN(n12799) );
  AOI22_X1 U15924 ( .A1(n9751), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(n9748), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12798) );
  AOI22_X1 U15925 ( .A1(n9759), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12861), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12797) );
  NAND4_X1 U15926 ( .A1(n12799), .A2(n12798), .A3(n12797), .A4(n12796), .ZN(
        n12800) );
  NAND2_X1 U15927 ( .A1(n12801), .A2(n12800), .ZN(n12805) );
  INV_X1 U15928 ( .A(n12805), .ZN(n12812) );
  INV_X1 U15929 ( .A(n12802), .ZN(n12804) );
  NAND2_X1 U15930 ( .A1(n12804), .A2(n12803), .ZN(n12806) );
  INV_X1 U15931 ( .A(n12806), .ZN(n12808) );
  OR2_X1 U15932 ( .A1(n12806), .A2(n12805), .ZN(n14849) );
  OAI211_X1 U15933 ( .C1(n12812), .C2(n12808), .A(n14849), .B(n12807), .ZN(
        n12809) );
  INV_X1 U15934 ( .A(n12809), .ZN(n12810) );
  NAND2_X1 U15935 ( .A1(n9788), .A2(n12812), .ZN(n14856) );
  INV_X1 U15936 ( .A(n14848), .ZN(n12829) );
  INV_X1 U15937 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12814) );
  NAND2_X1 U15938 ( .A1(n12863), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n12813) );
  OAI211_X1 U15939 ( .C1(n12842), .C2(n12814), .A(n12813), .B(n12864), .ZN(
        n12815) );
  INV_X1 U15940 ( .A(n12815), .ZN(n12819) );
  AOI22_X1 U15941 ( .A1(n9753), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(n9750), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12818) );
  AOI22_X1 U15942 ( .A1(n9759), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12861), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12817) );
  NAND4_X1 U15943 ( .A1(n12819), .A2(n12818), .A3(n12817), .A4(n12816), .ZN(
        n12828) );
  NAND2_X1 U15944 ( .A1(n12863), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n12820) );
  OAI211_X1 U15945 ( .C1(n12842), .C2(n12821), .A(n12820), .B(n12840), .ZN(
        n12822) );
  INV_X1 U15946 ( .A(n12822), .ZN(n12826) );
  AOI22_X1 U15947 ( .A1(n9752), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(n9749), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12825) );
  AOI22_X1 U15948 ( .A1(n9759), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12861), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12824) );
  NAND4_X1 U15949 ( .A1(n12826), .A2(n12825), .A3(n12824), .A4(n12823), .ZN(
        n12827) );
  AND2_X1 U15950 ( .A1(n12828), .A2(n12827), .ZN(n14850) );
  NAND2_X1 U15951 ( .A1(n11014), .A2(n14850), .ZN(n12830) );
  NOR2_X1 U15952 ( .A1(n14849), .A2(n12830), .ZN(n12851) );
  AOI22_X1 U15953 ( .A1(n9759), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(n9749), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12837) );
  INV_X1 U15954 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12832) );
  NAND2_X1 U15955 ( .A1(n9795), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n12831) );
  OAI211_X1 U15956 ( .C1(n12842), .C2(n12832), .A(n12831), .B(n12864), .ZN(
        n12833) );
  INV_X1 U15957 ( .A(n12833), .ZN(n12836) );
  AOI22_X1 U15958 ( .A1(n12863), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9751), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12835) );
  AOI22_X1 U15959 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12861), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12834) );
  NAND4_X1 U15960 ( .A1(n12837), .A2(n12836), .A3(n12835), .A4(n12834), .ZN(
        n12849) );
  AOI22_X1 U15961 ( .A1(n9752), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(n9748), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12847) );
  AOI22_X1 U15962 ( .A1(n12720), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12863), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12846) );
  INV_X1 U15963 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12841) );
  NAND2_X1 U15964 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n12839) );
  OAI211_X1 U15965 ( .C1(n12842), .C2(n12841), .A(n12840), .B(n12839), .ZN(
        n12843) );
  INV_X1 U15966 ( .A(n12843), .ZN(n12845) );
  AOI22_X1 U15967 ( .A1(n9759), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12861), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12844) );
  NAND4_X1 U15968 ( .A1(n12847), .A2(n12846), .A3(n12845), .A4(n12844), .ZN(
        n12848) );
  AND2_X1 U15969 ( .A1(n12849), .A2(n12848), .ZN(n12850) );
  NAND2_X1 U15970 ( .A1(n12851), .A2(n12850), .ZN(n12852) );
  OAI21_X1 U15971 ( .B1(n12851), .B2(n12850), .A(n12852), .ZN(n14844) );
  INV_X1 U15972 ( .A(n12861), .ZN(n15381) );
  INV_X1 U15973 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12856) );
  AOI21_X1 U15974 ( .B1(n12862), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n12864), .ZN(n12854) );
  OAI211_X1 U15975 ( .C1(n15381), .C2(n12856), .A(n12855), .B(n12854), .ZN(
        n12871) );
  AOI22_X1 U15976 ( .A1(n9751), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(n9750), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12858) );
  NAND2_X1 U15977 ( .A1(n12858), .A2(n12857), .ZN(n12870) );
  AOI22_X1 U15978 ( .A1(n9753), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(n9759), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12860) );
  NAND2_X1 U15979 ( .A1(n12860), .A2(n12859), .ZN(n12869) );
  AOI22_X1 U15980 ( .A1(n9795), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12861), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12867) );
  NAND2_X1 U15981 ( .A1(n12862), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n12866) );
  NAND2_X1 U15982 ( .A1(n12863), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n12865) );
  NAND4_X1 U15983 ( .A1(n12867), .A2(n12866), .A3(n12865), .A4(n12864), .ZN(
        n12868) );
  OAI22_X1 U15984 ( .A1(n12871), .A2(n12870), .B1(n12869), .B2(n12868), .ZN(
        n12872) );
  XNOR2_X1 U15985 ( .A(n12873), .B(n12872), .ZN(n14171) );
  AND2_X1 U15986 ( .A1(n10986), .A2(n19765), .ZN(n13066) );
  NAND2_X1 U15987 ( .A1(n13073), .A2(n13066), .ZN(n12874) );
  NOR2_X1 U15988 ( .A1(n13072), .A2(n12874), .ZN(n12875) );
  AOI21_X1 U15989 ( .B1(n13074), .B2(n15379), .A(n12875), .ZN(n15358) );
  NAND2_X1 U15990 ( .A1(n15358), .A2(n12876), .ZN(n12877) );
  AOI21_X1 U15991 ( .B1(n12881), .B2(n12879), .A(n12880), .ZN(n14712) );
  INV_X1 U15992 ( .A(n12882), .ZN(n12883) );
  NOR4_X1 U15993 ( .A1(P2_ADDRESS_REG_16__SCAN_IN), .A2(
        P2_ADDRESS_REG_15__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_13__SCAN_IN), .ZN(n12887) );
  NOR4_X1 U15994 ( .A1(P2_ADDRESS_REG_20__SCAN_IN), .A2(
        P2_ADDRESS_REG_19__SCAN_IN), .A3(P2_ADDRESS_REG_18__SCAN_IN), .A4(
        P2_ADDRESS_REG_17__SCAN_IN), .ZN(n12886) );
  NOR4_X1 U15995 ( .A1(P2_ADDRESS_REG_7__SCAN_IN), .A2(
        P2_ADDRESS_REG_6__SCAN_IN), .A3(P2_ADDRESS_REG_5__SCAN_IN), .A4(
        P2_ADDRESS_REG_4__SCAN_IN), .ZN(n12885) );
  NOR4_X1 U15996 ( .A1(P2_ADDRESS_REG_12__SCAN_IN), .A2(
        P2_ADDRESS_REG_11__SCAN_IN), .A3(P2_ADDRESS_REG_10__SCAN_IN), .A4(
        P2_ADDRESS_REG_9__SCAN_IN), .ZN(n12884) );
  NAND4_X1 U15997 ( .A1(n12887), .A2(n12886), .A3(n12885), .A4(n12884), .ZN(
        n12892) );
  NOR4_X1 U15998 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_21__SCAN_IN), .ZN(n12890) );
  NOR4_X1 U15999 ( .A1(P2_ADDRESS_REG_25__SCAN_IN), .A2(
        P2_ADDRESS_REG_24__SCAN_IN), .A3(P2_ADDRESS_REG_23__SCAN_IN), .A4(
        P2_ADDRESS_REG_22__SCAN_IN), .ZN(n12889) );
  NOR4_X1 U16000 ( .A1(P2_ADDRESS_REG_3__SCAN_IN), .A2(
        P2_ADDRESS_REG_28__SCAN_IN), .A3(P2_ADDRESS_REG_27__SCAN_IN), .A4(
        P2_ADDRESS_REG_26__SCAN_IN), .ZN(n12888) );
  NAND4_X1 U16001 ( .A1(n12890), .A2(n12889), .A3(n12888), .A4(n19798), .ZN(
        n12891) );
  MUX2_X1 U16002 ( .A(BUF1_REG_14__SCAN_IN), .B(BUF2_REG_14__SCAN_IN), .S(
        n13643), .Z(n19088) );
  INV_X1 U16003 ( .A(n19088), .ZN(n12895) );
  INV_X1 U16004 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n12894) );
  OAI22_X1 U16005 ( .A1(n14973), .A2(n12895), .B1(n19110), .B2(n12894), .ZN(
        n12896) );
  AOI21_X1 U16006 ( .B1(n14712), .B2(n19127), .A(n12896), .ZN(n12899) );
  AND2_X1 U16007 ( .A1(n12509), .A2(n9755), .ZN(n12897) );
  AOI22_X1 U16008 ( .A1(n19078), .A2(BUF1_REG_30__SCAN_IN), .B1(n19077), .B2(
        BUF2_REG_30__SCAN_IN), .ZN(n12898) );
  AND2_X1 U16009 ( .A1(n12899), .A2(n12898), .ZN(n12900) );
  OAI21_X1 U16010 ( .B1(n14171), .B2(n19112), .A(n12900), .ZN(P2_U2889) );
  NOR2_X1 U16011 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12902) );
  NOR4_X1 U16012 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12901) );
  NAND4_X1 U16013 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n12902), .A4(n12901), .ZN(n12915) );
  NOR4_X1 U16014 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(
        P1_ADDRESS_REG_16__SCAN_IN), .A3(P1_ADDRESS_REG_15__SCAN_IN), .A4(
        P1_ADDRESS_REG_14__SCAN_IN), .ZN(n12906) );
  NOR4_X1 U16015 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(
        P1_ADDRESS_REG_20__SCAN_IN), .A3(P1_ADDRESS_REG_19__SCAN_IN), .A4(
        P1_ADDRESS_REG_18__SCAN_IN), .ZN(n12905) );
  NOR4_X1 U16016 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(
        P1_ADDRESS_REG_6__SCAN_IN), .A3(P1_ADDRESS_REG_5__SCAN_IN), .A4(
        P1_ADDRESS_REG_4__SCAN_IN), .ZN(n12904) );
  NOR4_X1 U16017 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(
        P1_ADDRESS_REG_11__SCAN_IN), .A3(P1_ADDRESS_REG_10__SCAN_IN), .A4(
        P1_ADDRESS_REG_9__SCAN_IN), .ZN(n12903) );
  AND4_X1 U16018 ( .A1(n12906), .A2(n12905), .A3(n12904), .A4(n12903), .ZN(
        n12911) );
  NOR4_X1 U16019 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_13__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12909) );
  NOR4_X1 U16020 ( .A1(P1_ADDRESS_REG_25__SCAN_IN), .A2(
        P1_ADDRESS_REG_24__SCAN_IN), .A3(P1_ADDRESS_REG_23__SCAN_IN), .A4(
        P1_ADDRESS_REG_22__SCAN_IN), .ZN(n12908) );
  NOR4_X1 U16021 ( .A1(P1_ADDRESS_REG_8__SCAN_IN), .A2(
        P1_ADDRESS_REG_28__SCAN_IN), .A3(P1_ADDRESS_REG_27__SCAN_IN), .A4(
        P1_ADDRESS_REG_26__SCAN_IN), .ZN(n12907) );
  INV_X1 U16022 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20760) );
  AND4_X1 U16023 ( .A1(n12909), .A2(n12908), .A3(n12907), .A4(n20760), .ZN(
        n12910) );
  NAND2_X1 U16024 ( .A1(n12911), .A2(n12910), .ZN(n12912) );
  INV_X1 U16025 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20834) );
  NOR3_X1 U16026 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20834), .ZN(n12914) );
  NOR4_X1 U16027 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n12913) );
  NAND4_X1 U16028 ( .A1(n20116), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n12914), .A4(
        n12913), .ZN(U214) );
  NOR2_X1 U16029 ( .A1(n13643), .A2(n12915), .ZN(n16468) );
  NAND2_X1 U16030 ( .A1(n16468), .A2(U214), .ZN(U212) );
  INV_X1 U16031 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18855) );
  NAND2_X1 U16032 ( .A1(n18834), .A2(n18824), .ZN(n18837) );
  NOR2_X2 U16033 ( .A1(n13030), .A2(n12920), .ZN(n15552) );
  INV_X2 U16034 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12916) );
  AOI22_X1 U16035 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12933) );
  AOI22_X1 U16036 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n15550), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12932) );
  NOR2_X2 U16037 ( .A1(n12923), .A2(n12919), .ZN(n15553) );
  AOI22_X1 U16038 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12918) );
  OAI21_X1 U16039 ( .B1(n12993), .B2(n18226), .A(n12918), .ZN(n12930) );
  BUF_X4 U16040 ( .A(n15554), .Z(n17205) );
  AOI22_X1 U16041 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n15559), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12928) );
  NOR2_X2 U16042 ( .A1(n16921), .A2(n12921), .ZN(n17176) );
  AOI22_X1 U16043 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12927) );
  NOR2_X2 U16044 ( .A1(n12922), .A2(n13030), .ZN(n15435) );
  INV_X2 U16045 ( .A(n15562), .ZN(n17214) );
  AOI22_X1 U16046 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12926) );
  NOR2_X2 U16047 ( .A1(n18848), .A2(n13018), .ZN(n18685) );
  BUF_X4 U16048 ( .A(n15595), .Z(n17189) );
  AOI22_X1 U16049 ( .A1(n17207), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12925) );
  NAND4_X1 U16050 ( .A1(n12928), .A2(n12927), .A3(n12926), .A4(n12925), .ZN(
        n12929) );
  AOI22_X1 U16051 ( .A1(n9763), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12937) );
  AOI22_X1 U16052 ( .A1(n17209), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17205), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12936) );
  INV_X2 U16053 ( .A(n12993), .ZN(n17122) );
  AOI22_X1 U16054 ( .A1(n17122), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n15550), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12935) );
  AOI22_X1 U16055 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12934) );
  NAND4_X1 U16056 ( .A1(n12937), .A2(n12936), .A3(n12935), .A4(n12934), .ZN(
        n12943) );
  AOI22_X1 U16057 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9758), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12941) );
  AOI22_X1 U16058 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12940) );
  AOI22_X1 U16059 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12939) );
  AOI22_X1 U16060 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n17215), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12938) );
  NAND4_X1 U16061 ( .A1(n12941), .A2(n12940), .A3(n12939), .A4(n12938), .ZN(
        n12942) );
  INV_X1 U16062 ( .A(n18253), .ZN(n17259) );
  AOI22_X1 U16063 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12953) );
  AOI22_X1 U16064 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12952) );
  AOI22_X1 U16065 ( .A1(n17209), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12944) );
  OAI21_X1 U16066 ( .B1(n12917), .B2(n20954), .A(n12944), .ZN(n12950) );
  AOI22_X1 U16067 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n15550), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12948) );
  AOI22_X1 U16068 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12947) );
  AOI22_X1 U16069 ( .A1(n9758), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12946) );
  AOI22_X1 U16070 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12945) );
  NAND4_X1 U16071 ( .A1(n12948), .A2(n12947), .A3(n12946), .A4(n12945), .ZN(
        n12949) );
  NAND2_X1 U16072 ( .A1(n17259), .A2(n18247), .ZN(n13015) );
  AOI22_X1 U16073 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12957) );
  AOI22_X1 U16074 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12956) );
  AOI22_X1 U16075 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12955) );
  AOI22_X1 U16076 ( .A1(n17207), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12954) );
  NAND4_X1 U16077 ( .A1(n12957), .A2(n12956), .A3(n12955), .A4(n12954), .ZN(
        n12963) );
  AOI22_X1 U16078 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12961) );
  AOI22_X1 U16079 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12960) );
  AOI22_X1 U16080 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n15550), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12959) );
  AOI22_X1 U16081 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12958) );
  NAND4_X1 U16082 ( .A1(n12961), .A2(n12960), .A3(n12959), .A4(n12958), .ZN(
        n12962) );
  AOI22_X1 U16083 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12966) );
  AOI22_X1 U16084 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12965) );
  AOI22_X1 U16085 ( .A1(n17207), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12964) );
  AOI22_X1 U16086 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12970) );
  AOI22_X1 U16087 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12969) );
  AOI22_X1 U16088 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12968) );
  AOI22_X1 U16089 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17224), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12967) );
  NAND4_X1 U16090 ( .A1(n12970), .A2(n12969), .A3(n12968), .A4(n12967), .ZN(
        n12971) );
  AOI22_X1 U16091 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12975) );
  AOI22_X1 U16092 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12974) );
  AOI22_X1 U16093 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12973) );
  AOI22_X1 U16094 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12972) );
  NAND4_X1 U16095 ( .A1(n12975), .A2(n12974), .A3(n12973), .A4(n12972), .ZN(
        n12981) );
  AOI22_X1 U16096 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(n9763), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12979) );
  AOI22_X1 U16097 ( .A1(n9758), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n15550), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12978) );
  AOI22_X1 U16098 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12977) );
  AOI22_X1 U16099 ( .A1(n17207), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12976) );
  NAND4_X1 U16100 ( .A1(n12979), .A2(n12978), .A3(n12977), .A4(n12976), .ZN(
        n12980) );
  NOR2_X1 U16101 ( .A1(n9796), .A2(n18238), .ZN(n15643) );
  NAND2_X1 U16102 ( .A1(n13004), .A2(n15643), .ZN(n13917) );
  AOI22_X1 U16103 ( .A1(n17207), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12991) );
  AOI22_X1 U16104 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n15559), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12990) );
  AOI22_X1 U16105 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12982) );
  OAI21_X1 U16106 ( .B1(n12993), .B2(n18245), .A(n12982), .ZN(n12988) );
  AOI22_X1 U16107 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n15550), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12986) );
  AOI22_X1 U16108 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12985) );
  AOI22_X1 U16109 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12984) );
  AOI22_X1 U16110 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12983) );
  NAND4_X1 U16111 ( .A1(n12986), .A2(n12985), .A3(n12984), .A4(n12983), .ZN(
        n12987) );
  NOR2_X1 U16112 ( .A1(n18253), .A2(n18247), .ZN(n15634) );
  NAND4_X1 U16113 ( .A1(n18238), .A2(n18242), .A3(n13016), .A4(n15634), .ZN(
        n13014) );
  AOI22_X1 U16114 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n15559), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12992) );
  OAI21_X1 U16115 ( .B1(n12993), .B2(n18230), .A(n12992), .ZN(n12999) );
  AOI22_X1 U16116 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(n9763), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12997) );
  AOI22_X1 U16117 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n15552), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12996) );
  AOI22_X1 U16118 ( .A1(n17207), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n15550), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12995) );
  AOI22_X1 U16119 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12994) );
  NAND4_X1 U16120 ( .A1(n12997), .A2(n12996), .A3(n12995), .A4(n12994), .ZN(
        n12998) );
  NAND2_X1 U16121 ( .A1(n16394), .A2(n9783), .ZN(n13931) );
  INV_X1 U16122 ( .A(n13931), .ZN(n13003) );
  NAND2_X1 U16123 ( .A1(n18232), .A2(n17267), .ZN(n13929) );
  INV_X1 U16124 ( .A(n13929), .ZN(n15629) );
  NAND2_X1 U16125 ( .A1(n18253), .A2(n15635), .ZN(n18673) );
  AND2_X1 U16126 ( .A1(n13004), .A2(n18673), .ZN(n13012) );
  NAND2_X1 U16127 ( .A1(n18253), .A2(n17267), .ZN(n15773) );
  INV_X1 U16128 ( .A(n15773), .ZN(n18693) );
  OAI211_X1 U16129 ( .C1(n9796), .C2(n18693), .A(n18874), .B(n18227), .ZN(
        n13919) );
  OAI21_X1 U16130 ( .B1(n15629), .B2(n13012), .A(n13919), .ZN(n13005) );
  INV_X1 U16131 ( .A(n13005), .ZN(n13013) );
  INV_X1 U16132 ( .A(n18238), .ZN(n13006) );
  OAI22_X1 U16133 ( .A1(n13016), .A2(n13006), .B1(n15635), .B2(n15773), .ZN(
        n13011) );
  NOR2_X1 U16134 ( .A1(n9796), .A2(n15634), .ZN(n13009) );
  NOR2_X1 U16135 ( .A1(n18227), .A2(n18874), .ZN(n13918) );
  INV_X1 U16136 ( .A(n18232), .ZN(n13007) );
  NOR2_X1 U16137 ( .A1(n13918), .A2(n13007), .ZN(n13008) );
  OAI22_X1 U16138 ( .A1(n18242), .A2(n13009), .B1(n15634), .B2(n13008), .ZN(
        n13010) );
  AOI211_X1 U16139 ( .C1(n18221), .C2(n13012), .A(n13011), .B(n13010), .ZN(
        n13920) );
  OAI21_X1 U16140 ( .B1(n18238), .B2(n13013), .A(n13920), .ZN(n15644) );
  NAND2_X1 U16141 ( .A1(n18232), .A2(n18238), .ZN(n18672) );
  NOR2_X1 U16142 ( .A1(n13015), .A2(n18672), .ZN(n15418) );
  AOI22_X1 U16143 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n18699), .B2(n18848), .ZN(
        n13925) );
  NAND2_X1 U16144 ( .A1(n18217), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13924) );
  XNOR2_X1 U16145 ( .A(n13925), .B(n13924), .ZN(n13028) );
  NOR2_X1 U16146 ( .A1(n13925), .A2(n13924), .ZN(n13017) );
  OAI22_X1 U16147 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18708), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13020), .ZN(n13025) );
  NOR2_X1 U16148 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18708), .ZN(
        n13021) );
  NAND2_X1 U16149 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13020), .ZN(
        n13026) );
  AOI22_X1 U16150 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13025), .B1(
        n13021), .B2(n13026), .ZN(n13923) );
  NAND2_X1 U16151 ( .A1(n13024), .A2(n13023), .ZN(n13022) );
  AOI21_X1 U16152 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n13026), .A(
        n13025), .ZN(n13027) );
  INV_X1 U16153 ( .A(n18887), .ZN(n18885) );
  NOR4_X4 U16154 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .A4(n18834), .ZN(n18733) );
  INV_X1 U16155 ( .A(n18729), .ZN(n13029) );
  NAND2_X1 U16156 ( .A1(n13029), .A2(n9746), .ZN(n18722) );
  NAND2_X1 U16157 ( .A1(n13030), .A2(n16921), .ZN(n18841) );
  NOR2_X1 U16158 ( .A1(n18874), .A2(n18885), .ZN(n18891) );
  INV_X1 U16159 ( .A(n18891), .ZN(n16910) );
  OAI22_X1 U16160 ( .A1(n18855), .A2(n16945), .B1(n18841), .B2(n16910), .ZN(
        n13038) );
  INV_X1 U16161 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17252) );
  INV_X1 U16162 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n20849) );
  NAND2_X1 U16163 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n20849), .ZN(n18882) );
  INV_X1 U16164 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n20848) );
  NOR2_X1 U16165 ( .A1(n18882), .A2(n20848), .ZN(n18749) );
  OAI21_X1 U16166 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(P3_STATE_REG_2__SCAN_IN), 
        .A(n20849), .ZN(n18739) );
  NOR2_X1 U16167 ( .A1(n18749), .A2(n18739), .ZN(n15627) );
  INV_X1 U16168 ( .A(n15627), .ZN(n18872) );
  AOI211_X1 U16169 ( .C1(n18227), .C2(n18872), .A(n18870), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n13033) );
  NAND2_X1 U16170 ( .A1(n18887), .A2(n18874), .ZN(n13034) );
  AOI211_X4 U16171 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n16394), .A(n13033), .B(
        n13034), .ZN(n16947) );
  NAND2_X1 U16172 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17842) );
  NOR2_X1 U16173 ( .A1(n17842), .A2(n17844), .ZN(n17826) );
  NAND2_X1 U16174 ( .A1(n17826), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17814) );
  NAND2_X1 U16175 ( .A1(n17782), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16812) );
  NAND2_X1 U16176 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17717) );
  NAND2_X1 U16177 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17678) );
  NAND3_X1 U16178 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17630) );
  NOR2_X1 U16179 ( .A1(n17630), .A2(n17629), .ZN(n16583) );
  NAND2_X1 U16180 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17604) );
  NAND2_X1 U16181 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17562) );
  NAND2_X1 U16182 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17548), .ZN(
        n17530) );
  NAND2_X1 U16183 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17531) );
  NAND2_X1 U16184 ( .A1(n16412), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13031) );
  XOR2_X2 U16185 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(n13031), .Z(
        n16858) );
  INV_X1 U16186 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16731) );
  OAI21_X1 U16187 ( .B1(n16858), .B2(n16731), .A(n18733), .ZN(n16872) );
  OAI22_X1 U16188 ( .A1(n17252), .A2(n16911), .B1(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16872), .ZN(n13037) );
  NAND2_X1 U16189 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n16394), .ZN(n13032) );
  AOI211_X4 U16190 ( .C1(n18875), .C2(n18873), .A(n13034), .B(n13032), .ZN(
        n16946) );
  INV_X1 U16191 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17257) );
  NAND2_X1 U16192 ( .A1(n17257), .A2(n17252), .ZN(n16938) );
  OAI21_X1 U16193 ( .B1(n17252), .B2(n17257), .A(n16938), .ZN(n17253) );
  INV_X1 U16194 ( .A(n13033), .ZN(n18718) );
  OAI22_X1 U16195 ( .A1(n16937), .A2(n17253), .B1(n16909), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n13036) );
  NAND2_X1 U16196 ( .A1(n16907), .A2(n18733), .ZN(n16873) );
  AOI221_X1 U16197 ( .B1(n16920), .B2(n16873), .C1(n16920), .C2(n16731), .A(
        n17875), .ZN(n13035) );
  OR4_X1 U16198 ( .A1(n13038), .A2(n13037), .A3(n13036), .A4(n13035), .ZN(
        P3_U2670) );
  INV_X1 U16199 ( .A(n15502), .ZN(n16348) );
  NAND2_X1 U16200 ( .A1(n16348), .A2(n19768), .ZN(n19137) );
  OR2_X1 U16201 ( .A1(n13072), .A2(n19137), .ZN(n19068) );
  INV_X1 U16202 ( .A(n19068), .ZN(n13041) );
  INV_X1 U16203 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n19890) );
  NAND2_X1 U16204 ( .A1(n13039), .A2(n19768), .ZN(n13040) );
  OAI211_X1 U16205 ( .C1(n13041), .C2(n19890), .A(n18893), .B(n13046), .ZN(
        P2_U2814) );
  NAND2_X1 U16206 ( .A1(n13073), .A2(n19768), .ZN(n13042) );
  NOR2_X1 U16207 ( .A1(n18895), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n13044)
         );
  INV_X1 U16208 ( .A(n10986), .ZN(n13043) );
  AOI22_X1 U16209 ( .A1(n13044), .A2(n18893), .B1(n13043), .B2(n18895), .ZN(
        P2_U3612) );
  NOR3_X1 U16210 ( .A1(n13046), .A2(n9788), .A3(n19785), .ZN(n13045) );
  INV_X1 U16211 ( .A(n13118), .ZN(n13051) );
  INV_X1 U16212 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16513) );
  INV_X1 U16213 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18218) );
  AOI22_X1 U16214 ( .A1(n13645), .A2(n16513), .B1(n18218), .B2(n13643), .ZN(
        n19075) );
  INV_X1 U16215 ( .A(n19075), .ZN(n13642) );
  INV_X1 U16216 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n13048) );
  OAI21_X1 U16217 ( .B1(n9788), .B2(n19765), .A(n14143), .ZN(n13047) );
  INV_X1 U16218 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n19168) );
  OAI222_X1 U16219 ( .A1(n13051), .A2(n13642), .B1(n13048), .B2(n13101), .C1(
        n19136), .C2(n19168), .ZN(P2_U2952) );
  INV_X1 U16220 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n13049) );
  OAI222_X1 U16221 ( .A1(n13050), .A2(n19136), .B1(n13049), .B2(n13101), .C1(
        n13051), .C2(n13642), .ZN(P2_U2967) );
  INV_X1 U16222 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13053) );
  INV_X1 U16223 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13052) );
  AOI22_X1 U16224 ( .A1(n13645), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n13643), .ZN(n19085) );
  OAI222_X1 U16225 ( .A1(n13053), .A2(n19136), .B1(n13052), .B2(n13101), .C1(
        n13051), .C2(n19085), .ZN(P2_U2982) );
  NAND2_X1 U16226 ( .A1(n13118), .A2(n19088), .ZN(n13056) );
  NAND2_X1 U16227 ( .A1(n13099), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13054) );
  OAI211_X1 U16228 ( .C1(n12894), .C2(n19136), .A(n13056), .B(n13054), .ZN(
        P2_U2966) );
  NAND2_X1 U16229 ( .A1(n13099), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13055) );
  OAI211_X1 U16230 ( .C1(n11197), .C2(n19136), .A(n13056), .B(n13055), .ZN(
        P2_U2981) );
  INV_X1 U16231 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19180) );
  MUX2_X1 U16232 ( .A(BUF1_REG_10__SCAN_IN), .B(BUF2_REG_10__SCAN_IN), .S(
        n13643), .Z(n19099) );
  NAND2_X1 U16233 ( .A1(n13118), .A2(n19099), .ZN(n13065) );
  NAND2_X1 U16234 ( .A1(n13099), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13057) );
  OAI211_X1 U16235 ( .C1(n19180), .C2(n19136), .A(n13065), .B(n13057), .ZN(
        P2_U2977) );
  INV_X1 U16236 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19175) );
  MUX2_X1 U16237 ( .A(BUF1_REG_12__SCAN_IN), .B(BUF2_REG_12__SCAN_IN), .S(
        n13643), .Z(n19094) );
  NAND2_X1 U16238 ( .A1(n13118), .A2(n19094), .ZN(n13063) );
  NAND2_X1 U16239 ( .A1(n13099), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13058) );
  OAI211_X1 U16240 ( .C1(n19175), .C2(n19136), .A(n13063), .B(n13058), .ZN(
        P2_U2979) );
  INV_X1 U16241 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n21066) );
  NAND2_X1 U16242 ( .A1(n13643), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13060) );
  INV_X1 U16243 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16495) );
  OR2_X1 U16244 ( .A1(n13643), .A2(n16495), .ZN(n13059) );
  NAND2_X1 U16245 ( .A1(n13060), .A2(n13059), .ZN(n19103) );
  NAND2_X1 U16246 ( .A1(n13118), .A2(n19103), .ZN(n13115) );
  NAND2_X1 U16247 ( .A1(n13099), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n13061) );
  OAI211_X1 U16248 ( .C1(n21066), .C2(n19136), .A(n13115), .B(n13061), .ZN(
        P2_U2976) );
  INV_X1 U16249 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n20973) );
  NAND2_X1 U16250 ( .A1(n13099), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13062) );
  OAI211_X1 U16251 ( .C1(n20973), .C2(n19136), .A(n13063), .B(n13062), .ZN(
        P2_U2964) );
  INV_X1 U16252 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n20984) );
  NAND2_X1 U16253 ( .A1(n13099), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13064) );
  OAI211_X1 U16254 ( .C1(n20984), .C2(n19136), .A(n13065), .B(n13064), .ZN(
        P2_U2962) );
  NOR2_X1 U16255 ( .A1(n13066), .A2(n15359), .ZN(n13067) );
  NAND2_X1 U16256 ( .A1(n13073), .A2(n13067), .ZN(n13068) );
  NOR2_X1 U16257 ( .A1(n13072), .A2(n13068), .ZN(n16345) );
  INV_X1 U16258 ( .A(n19768), .ZN(n16375) );
  NOR2_X1 U16259 ( .A1(n16345), .A2(n16375), .ZN(n18900) );
  INV_X1 U16260 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n13080) );
  INV_X1 U16261 ( .A(n13069), .ZN(n13070) );
  MUX2_X1 U16262 ( .A(n13070), .B(n16361), .S(n9790), .Z(n13077) );
  INV_X1 U16263 ( .A(n13071), .ZN(n15378) );
  AOI22_X1 U16264 ( .A1(n13074), .A2(n15378), .B1(n13073), .B2(n13072), .ZN(
        n13076) );
  INV_X1 U16265 ( .A(n13074), .ZN(n13166) );
  NAND2_X1 U16266 ( .A1(n13166), .A2(n15379), .ZN(n13075) );
  AND2_X1 U16267 ( .A1(n13076), .A2(n13075), .ZN(n16352) );
  OAI21_X1 U16268 ( .B1(n13077), .B2(n16351), .A(n16352), .ZN(n13078) );
  NAND2_X1 U16269 ( .A1(n13078), .A2(n18900), .ZN(n13079) );
  OAI21_X1 U16270 ( .B1(n18900), .B2(n13080), .A(n13079), .ZN(P2_U3609) );
  AOI22_X1 U16271 ( .A1(n13130), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n13099), .B2(
        P2_LWORD_REG_6__SCAN_IN), .ZN(n13081) );
  OAI22_X1 U16272 ( .A1(n13643), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n13645), .ZN(n19271) );
  INV_X1 U16273 ( .A(n19271), .ZN(n16189) );
  NAND2_X1 U16274 ( .A1(n13118), .A2(n16189), .ZN(n13124) );
  NAND2_X1 U16275 ( .A1(n13081), .A2(n13124), .ZN(P2_U2973) );
  AOI22_X1 U16276 ( .A1(n13130), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n13099), .B2(
        P2_LWORD_REG_7__SCAN_IN), .ZN(n13083) );
  AOI22_X1 U16277 ( .A1(n13645), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n13643), .ZN(n19281) );
  INV_X1 U16278 ( .A(n19281), .ZN(n13082) );
  NAND2_X1 U16279 ( .A1(n13118), .A2(n13082), .ZN(n13126) );
  NAND2_X1 U16280 ( .A1(n13083), .A2(n13126), .ZN(P2_U2974) );
  AOI22_X1 U16281 ( .A1(n13130), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n13099), 
        .B2(P2_UWORD_REG_4__SCAN_IN), .ZN(n13084) );
  INV_X1 U16282 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16502) );
  INV_X1 U16283 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18241) );
  AOI22_X1 U16284 ( .A1(n13645), .A2(n16502), .B1(n18241), .B2(n13643), .ZN(
        n19260) );
  NAND2_X1 U16285 ( .A1(n13118), .A2(n19260), .ZN(n13106) );
  NAND2_X1 U16286 ( .A1(n13084), .A2(n13106), .ZN(P2_U2956) );
  AOI22_X1 U16287 ( .A1(n13130), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n13099), 
        .B2(P2_LWORD_REG_11__SCAN_IN), .ZN(n13089) );
  INV_X1 U16288 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n13085) );
  OR2_X1 U16289 ( .A1(n13643), .A2(n13085), .ZN(n13087) );
  NAND2_X1 U16290 ( .A1(n13643), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13086) );
  AND2_X1 U16291 ( .A1(n13087), .A2(n13086), .ZN(n19097) );
  INV_X1 U16292 ( .A(n19097), .ZN(n13088) );
  NAND2_X1 U16293 ( .A1(n13118), .A2(n13088), .ZN(n13131) );
  NAND2_X1 U16294 ( .A1(n13089), .A2(n13131), .ZN(P2_U2978) );
  AOI22_X1 U16295 ( .A1(n13130), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n13099), 
        .B2(P2_UWORD_REG_3__SCAN_IN), .ZN(n13091) );
  AOI22_X1 U16296 ( .A1(n13645), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n13643), .ZN(n19254) );
  INV_X1 U16297 ( .A(n19254), .ZN(n13090) );
  NAND2_X1 U16298 ( .A1(n13118), .A2(n13090), .ZN(n13104) );
  NAND2_X1 U16299 ( .A1(n13091), .A2(n13104), .ZN(P2_U2955) );
  AOI22_X1 U16300 ( .A1(n13130), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n13099), 
        .B2(P2_UWORD_REG_1__SCAN_IN), .ZN(n13093) );
  AOI22_X1 U16301 ( .A1(n13645), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n13643), .ZN(n19248) );
  INV_X1 U16302 ( .A(n19248), .ZN(n13092) );
  NAND2_X1 U16303 ( .A1(n13118), .A2(n13092), .ZN(n13120) );
  NAND2_X1 U16304 ( .A1(n13093), .A2(n13120), .ZN(P2_U2953) );
  AOI22_X1 U16305 ( .A1(n13130), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n13099), 
        .B2(P2_LWORD_REG_13__SCAN_IN), .ZN(n13098) );
  INV_X1 U16306 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n13094) );
  OR2_X1 U16307 ( .A1(n13643), .A2(n13094), .ZN(n13096) );
  NAND2_X1 U16308 ( .A1(n13643), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13095) );
  AND2_X1 U16309 ( .A1(n13096), .A2(n13095), .ZN(n19091) );
  INV_X1 U16310 ( .A(n19091), .ZN(n13097) );
  NAND2_X1 U16311 ( .A1(n13118), .A2(n13097), .ZN(n13113) );
  NAND2_X1 U16312 ( .A1(n13098), .A2(n13113), .ZN(P2_U2980) );
  AOI22_X1 U16313 ( .A1(n13130), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n13099), 
        .B2(P2_UWORD_REG_2__SCAN_IN), .ZN(n13100) );
  INV_X1 U16314 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16506) );
  INV_X1 U16315 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18231) );
  AOI22_X1 U16316 ( .A1(n13645), .A2(n16506), .B1(n18231), .B2(n13643), .ZN(
        n16199) );
  NAND2_X1 U16317 ( .A1(n13118), .A2(n16199), .ZN(n13102) );
  NAND2_X1 U16318 ( .A1(n13100), .A2(n13102), .ZN(P2_U2954) );
  AOI22_X1 U16319 ( .A1(n13130), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n13099), .B2(
        P2_LWORD_REG_2__SCAN_IN), .ZN(n13103) );
  NAND2_X1 U16320 ( .A1(n13103), .A2(n13102), .ZN(P2_U2969) );
  AOI22_X1 U16321 ( .A1(n13130), .A2(P2_EAX_REG_3__SCAN_IN), .B1(n13047), .B2(
        P2_LWORD_REG_3__SCAN_IN), .ZN(n13105) );
  NAND2_X1 U16322 ( .A1(n13105), .A2(n13104), .ZN(P2_U2970) );
  AOI22_X1 U16323 ( .A1(n13130), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n13047), .B2(
        P2_LWORD_REG_4__SCAN_IN), .ZN(n13107) );
  NAND2_X1 U16324 ( .A1(n13107), .A2(n13106), .ZN(P2_U2971) );
  AOI22_X1 U16325 ( .A1(n13130), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n13047), .B2(
        P2_LWORD_REG_8__SCAN_IN), .ZN(n13112) );
  INV_X1 U16326 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n13108) );
  OR2_X1 U16327 ( .A1(n13643), .A2(n13108), .ZN(n13110) );
  NAND2_X1 U16328 ( .A1(n13643), .A2(BUF2_REG_8__SCAN_IN), .ZN(n13109) );
  AND2_X1 U16329 ( .A1(n13110), .A2(n13109), .ZN(n19106) );
  INV_X1 U16330 ( .A(n19106), .ZN(n13111) );
  NAND2_X1 U16331 ( .A1(n13118), .A2(n13111), .ZN(n13128) );
  NAND2_X1 U16332 ( .A1(n13112), .A2(n13128), .ZN(P2_U2975) );
  AOI22_X1 U16333 ( .A1(n13130), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n13047), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13114) );
  NAND2_X1 U16334 ( .A1(n13114), .A2(n13113), .ZN(P2_U2965) );
  AOI22_X1 U16335 ( .A1(n13130), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n13047), 
        .B2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13116) );
  NAND2_X1 U16336 ( .A1(n13116), .A2(n13115), .ZN(P2_U2961) );
  AOI22_X1 U16337 ( .A1(n13130), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n13047), .B2(
        P2_LWORD_REG_5__SCAN_IN), .ZN(n13119) );
  AOI22_X1 U16338 ( .A1(n13645), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n13643), .ZN(n19266) );
  INV_X1 U16339 ( .A(n19266), .ZN(n13117) );
  NAND2_X1 U16340 ( .A1(n13118), .A2(n13117), .ZN(n13122) );
  NAND2_X1 U16341 ( .A1(n13119), .A2(n13122), .ZN(P2_U2972) );
  AOI22_X1 U16342 ( .A1(n13130), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n13047), .B2(
        P2_LWORD_REG_1__SCAN_IN), .ZN(n13121) );
  NAND2_X1 U16343 ( .A1(n13121), .A2(n13120), .ZN(P2_U2968) );
  AOI22_X1 U16344 ( .A1(n13130), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n13047), 
        .B2(P2_UWORD_REG_5__SCAN_IN), .ZN(n13123) );
  NAND2_X1 U16345 ( .A1(n13123), .A2(n13122), .ZN(P2_U2957) );
  AOI22_X1 U16346 ( .A1(n13130), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n13047), 
        .B2(P2_UWORD_REG_6__SCAN_IN), .ZN(n13125) );
  NAND2_X1 U16347 ( .A1(n13125), .A2(n13124), .ZN(P2_U2958) );
  AOI22_X1 U16348 ( .A1(n13130), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n13047), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n13127) );
  NAND2_X1 U16349 ( .A1(n13127), .A2(n13126), .ZN(P2_U2959) );
  AOI22_X1 U16350 ( .A1(n13130), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n13099), 
        .B2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13129) );
  NAND2_X1 U16351 ( .A1(n13129), .A2(n13128), .ZN(P2_U2960) );
  AOI22_X1 U16352 ( .A1(n13130), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n13099), 
        .B2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13132) );
  NAND2_X1 U16353 ( .A1(n13132), .A2(n13131), .ZN(P2_U2963) );
  NOR4_X1 U16354 ( .A1(n13137), .A2(n13136), .A3(n13135), .A4(n13134), .ZN(
        n13138) );
  OR2_X1 U16355 ( .A1(n13139), .A2(n13138), .ZN(n13228) );
  INV_X1 U16356 ( .A(n13228), .ZN(n13140) );
  INV_X1 U16357 ( .A(n13327), .ZN(n15763) );
  OR2_X1 U16358 ( .A1(n13142), .A2(n15763), .ZN(n13143) );
  NAND2_X1 U16359 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n16106) );
  AND2_X1 U16360 ( .A1(n13143), .A2(n16106), .ZN(n20841) );
  NOR2_X1 U16361 ( .A1(n10129), .A2(n20841), .ZN(n15732) );
  OR2_X1 U16362 ( .A1(n15732), .A2(n19899), .ZN(n13154) );
  INV_X1 U16363 ( .A(n13154), .ZN(n19906) );
  INV_X1 U16364 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13156) );
  NAND2_X1 U16365 ( .A1(n13185), .A2(n13677), .ZN(n13389) );
  AND2_X1 U16366 ( .A1(n13389), .A2(n15735), .ZN(n13242) );
  INV_X1 U16367 ( .A(n13144), .ZN(n13145) );
  NAND2_X1 U16368 ( .A1(n13145), .A2(n11464), .ZN(n13146) );
  AND2_X1 U16369 ( .A1(n13242), .A2(n13146), .ZN(n13152) );
  INV_X1 U16370 ( .A(n13147), .ZN(n13391) );
  NAND2_X1 U16371 ( .A1(n13232), .A2(n13391), .ZN(n13151) );
  INV_X1 U16372 ( .A(n13149), .ZN(n13159) );
  NAND2_X1 U16373 ( .A1(n13159), .A2(n13228), .ZN(n13150) );
  OAI211_X1 U16374 ( .C1(n13232), .C2(n13152), .A(n13151), .B(n13150), .ZN(
        n13153) );
  NAND2_X1 U16375 ( .A1(n13153), .A2(n11456), .ZN(n15733) );
  OR2_X1 U16376 ( .A1(n13154), .A2(n15733), .ZN(n13155) );
  OAI21_X1 U16377 ( .B1(n19906), .B2(n13156), .A(n13155), .ZN(P1_U3484) );
  NOR2_X1 U16378 ( .A1(n13228), .A2(n19899), .ZN(n13158) );
  NAND2_X1 U16379 ( .A1(n13159), .A2(n13158), .ZN(n19895) );
  INV_X1 U16380 ( .A(n20840), .ZN(n13161) );
  AND2_X1 U16381 ( .A1(n20613), .A2(n20739), .ZN(n19892) );
  OAI21_X1 U16382 ( .B1(n19892), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n13161), 
        .ZN(n13160) );
  OAI21_X1 U16383 ( .B1(n13162), .B2(n13161), .A(n13160), .ZN(P1_U3487) );
  NAND2_X1 U16384 ( .A1(n9790), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13163) );
  NAND4_X1 U16385 ( .A1(n10251), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n13163), 
        .A4(n19680), .ZN(n13164) );
  NAND2_X1 U16386 ( .A1(n13166), .A2(n15378), .ZN(n15357) );
  NAND2_X1 U16387 ( .A1(n15357), .A2(n11001), .ZN(n13167) );
  MUX2_X1 U16388 ( .A(n14126), .B(n10538), .S(n14909), .Z(n13169) );
  OAI21_X1 U16389 ( .B1(n19881), .B2(n14911), .A(n13169), .ZN(P2_U2887) );
  NOR2_X1 U16390 ( .A1(n13313), .A2(n13168), .ZN(n13173) );
  AOI21_X1 U16391 ( .B1(P2_EBX_REG_1__SCAN_IN), .B2(n14909), .A(n13173), .ZN(
        n13174) );
  OAI21_X1 U16392 ( .B1(n19871), .B2(n14911), .A(n13174), .ZN(P2_U2886) );
  NOR2_X1 U16393 ( .A1(n13149), .A2(n13291), .ZN(n13403) );
  INV_X1 U16394 ( .A(n13176), .ZN(n13177) );
  NAND2_X1 U16395 ( .A1(n13389), .A2(n13177), .ZN(n13180) );
  NAND3_X1 U16396 ( .A1(n13176), .A2(n13459), .A3(n16106), .ZN(n13178) );
  OAI21_X1 U16397 ( .B1(n20838), .B2(n13327), .A(n13314), .ZN(n13179) );
  OAI21_X1 U16398 ( .B1(n13403), .B2(n13180), .A(n13179), .ZN(n13181) );
  INV_X1 U16399 ( .A(n13181), .ZN(n13189) );
  NOR2_X1 U16400 ( .A1(n13149), .A2(n12355), .ZN(n13413) );
  NOR2_X1 U16401 ( .A1(n13228), .A2(n20838), .ZN(n13182) );
  NOR2_X1 U16402 ( .A1(n13225), .A2(n13183), .ZN(n13184) );
  NAND2_X1 U16403 ( .A1(n11480), .A2(n13184), .ZN(n13196) );
  NAND2_X1 U16404 ( .A1(n13196), .A2(n13185), .ZN(n13186) );
  NAND2_X1 U16405 ( .A1(n13186), .A2(n13149), .ZN(n13230) );
  OAI21_X1 U16406 ( .B1(n13685), .B2(n20136), .A(n13230), .ZN(n13187) );
  OR2_X1 U16407 ( .A1(n13318), .A2(n13187), .ZN(n13188) );
  AOI21_X1 U16408 ( .B1(n13232), .B2(n13189), .A(n13188), .ZN(n13191) );
  NAND2_X1 U16409 ( .A1(n13191), .A2(n13190), .ZN(n15719) );
  INV_X1 U16410 ( .A(n16110), .ZN(n16112) );
  NOR2_X1 U16411 ( .A1(n11495), .A2(n16112), .ZN(n13418) );
  AOI22_X1 U16412 ( .A1(n15719), .A2(n13317), .B1(P1_FLUSH_REG_SCAN_IN), .B2(
        n13418), .ZN(n13192) );
  OAI21_X1 U16413 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n21100), .A(n13192), 
        .ZN(n20824) );
  NOR2_X1 U16414 ( .A1(n13192), .A2(n20822), .ZN(n16098) );
  OR2_X1 U16415 ( .A1(n13176), .A2(n11448), .ZN(n13194) );
  NOR2_X1 U16416 ( .A1(n13413), .A2(n13194), .ZN(n13200) );
  INV_X1 U16417 ( .A(n13195), .ZN(n13197) );
  OAI211_X1 U16418 ( .C1(n11820), .C2(n9787), .A(n13197), .B(n13196), .ZN(
        n13199) );
  NOR2_X1 U16419 ( .A1(n13199), .A2(n13198), .ZN(n13252) );
  NAND2_X1 U16420 ( .A1(n13200), .A2(n13252), .ZN(n14655) );
  NAND2_X1 U16421 ( .A1(n11849), .A2(n14655), .ZN(n13204) );
  INV_X1 U16422 ( .A(n14652), .ZN(n13201) );
  MUX2_X1 U16423 ( .A(n13403), .B(n13201), .S(n11311), .Z(n13202) );
  INV_X1 U16424 ( .A(n13202), .ZN(n13203) );
  NAND2_X1 U16425 ( .A1(n13204), .A2(n13203), .ZN(n15717) );
  OAI22_X1 U16426 ( .A1(n20739), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20821), .ZN(n13205) );
  AOI22_X1 U16427 ( .A1(n16098), .A2(n15717), .B1(n20824), .B2(n13205), .ZN(
        n13206) );
  OAI21_X1 U16428 ( .B1(n11311), .B2(n20824), .A(n13206), .ZN(P1_U3474) );
  INV_X1 U16429 ( .A(n19102), .ZN(n19135) );
  NOR2_X1 U16430 ( .A1(n13209), .A2(n13208), .ZN(n13210) );
  NOR2_X1 U16431 ( .A1(n11028), .A2(n13210), .ZN(n13213) );
  NAND2_X1 U16432 ( .A1(n13724), .A2(n13213), .ZN(n19129) );
  OAI211_X1 U16433 ( .C1(n13724), .C2(n13213), .A(n19129), .B(n19131), .ZN(
        n13212) );
  AOI22_X1 U16434 ( .A1(n19127), .A2(n13213), .B1(n19126), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n13211) );
  OAI211_X1 U16435 ( .C1(n19135), .C2(n13642), .A(n13212), .B(n13211), .ZN(
        P2_U2919) );
  NOR2_X1 U16436 ( .A1(n15334), .A2(n18912), .ZN(n14121) );
  INV_X1 U16437 ( .A(n13213), .ZN(n19064) );
  OAI22_X1 U16438 ( .A1(n13214), .A2(n13219), .B1(n15346), .B2(n19064), .ZN(
        n13215) );
  AOI211_X1 U16439 ( .C1(n19220), .C2(n13216), .A(n14121), .B(n13215), .ZN(
        n13224) );
  INV_X1 U16440 ( .A(n19059), .ZN(n13218) );
  INV_X1 U16441 ( .A(n13305), .ZN(n13217) );
  AOI21_X1 U16442 ( .B1(n13219), .B2(n13218), .A(n13217), .ZN(n14122) );
  OAI21_X1 U16443 ( .B1(n13221), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13220), .ZN(n14119) );
  INV_X1 U16444 ( .A(n14119), .ZN(n13222) );
  AOI22_X1 U16445 ( .A1(n16323), .A2(n14122), .B1(n19233), .B2(n13222), .ZN(
        n13223) );
  OAI211_X1 U16446 ( .C1(n15321), .C2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13224), .B(n13223), .ZN(P2_U3046) );
  INV_X1 U16447 ( .A(n13225), .ZN(n13231) );
  NAND2_X1 U16448 ( .A1(n12355), .A2(n13327), .ZN(n13226) );
  NAND3_X1 U16449 ( .A1(n13226), .A2(n20136), .A3(n16106), .ZN(n13227) );
  OR2_X1 U16450 ( .A1(n13228), .A2(n13227), .ZN(n13229) );
  OAI211_X1 U16451 ( .C1(n13232), .C2(n13231), .A(n13230), .B(n13229), .ZN(
        n13233) );
  NAND2_X1 U16452 ( .A1(n13233), .A2(n13317), .ZN(n13240) );
  NAND2_X1 U16453 ( .A1(n13291), .A2(n13327), .ZN(n13680) );
  NAND3_X1 U16454 ( .A1(n13176), .A2(n13680), .A3(n16106), .ZN(n13235) );
  NAND3_X1 U16455 ( .A1(n13235), .A2(n11464), .A3(n14088), .ZN(n13237) );
  NAND2_X1 U16456 ( .A1(n13237), .A2(n13236), .ZN(n13238) );
  OAI211_X1 U16457 ( .C1(n13244), .C2(n13241), .A(n13243), .B(n13242), .ZN(
        n13245) );
  OAI21_X1 U16458 ( .B1(n13246), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n11669), .ZN(n13274) );
  INV_X1 U16459 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20095) );
  NAND2_X1 U16460 ( .A1(n13247), .A2(n20095), .ZN(n13249) );
  NAND2_X1 U16461 ( .A1(n13249), .A2(n13248), .ZN(n14307) );
  OAI22_X1 U16462 ( .A1(n9766), .A2(n12355), .B1(n13241), .B2(n20152), .ZN(
        n13250) );
  NAND2_X1 U16463 ( .A1(n13252), .A2(n13251), .ZN(n13253) );
  NAND2_X1 U16464 ( .A1(n13256), .A2(n13253), .ZN(n13994) );
  INV_X1 U16465 ( .A(n13994), .ZN(n13254) );
  OAI21_X1 U16466 ( .B1(n16024), .B2(n13254), .A(n20095), .ZN(n20092) );
  NAND2_X1 U16467 ( .A1(n20099), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13273) );
  OAI211_X1 U16468 ( .C1(n14307), .C2(n20102), .A(n20092), .B(n13273), .ZN(
        n13255) );
  INV_X1 U16469 ( .A(n13255), .ZN(n13258) );
  NAND2_X1 U16470 ( .A1(n13256), .A2(n13403), .ZN(n20094) );
  INV_X1 U16471 ( .A(n20094), .ZN(n13991) );
  NOR2_X1 U16472 ( .A1(n20099), .A2(n13256), .ZN(n20089) );
  OAI21_X1 U16473 ( .B1(n13991), .B2(n20089), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13257) );
  OAI211_X1 U16474 ( .C1(n20088), .C2(n13274), .A(n13258), .B(n13257), .ZN(
        P1_U3031) );
  NAND2_X1 U16475 ( .A1(n13262), .A2(n13261), .ZN(n13263) );
  NOR2_X1 U16476 ( .A1(n14901), .A2(n10325), .ZN(n13266) );
  AOI21_X1 U16477 ( .B1(n14901), .B2(n13265), .A(n13266), .ZN(n13267) );
  OAI21_X1 U16478 ( .B1(n19864), .B2(n14911), .A(n13267), .ZN(P2_U2885) );
  NAND2_X1 U16479 ( .A1(n13269), .A2(n13268), .ZN(n13270) );
  NAND2_X1 U16480 ( .A1(n13271), .A2(n13270), .ZN(n20005) );
  NAND2_X1 U16481 ( .A1(n13272), .A2(n14518), .ZN(n13277) );
  INV_X1 U16482 ( .A(n13273), .ZN(n13276) );
  NOR2_X1 U16483 ( .A1(n19904), .A2(n13274), .ZN(n13275) );
  AOI211_X1 U16484 ( .C1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n13277), .A(
        n13276), .B(n13275), .ZN(n13278) );
  OAI21_X1 U16485 ( .B1(n20115), .B2(n20005), .A(n13278), .ZN(P1_U2999) );
  AOI21_X1 U16486 ( .B1(n14833), .B2(n10324), .A(n13618), .ZN(n14820) );
  INV_X1 U16487 ( .A(n14820), .ZN(n13289) );
  NAND2_X1 U16488 ( .A1(n13280), .A2(n13279), .ZN(n13281) );
  NAND2_X1 U16489 ( .A1(n13282), .A2(n13281), .ZN(n19226) );
  OAI22_X1 U16490 ( .A1(n19226), .A2(n16263), .B1(n10324), .B2(n19212), .ZN(
        n13283) );
  AOI21_X1 U16491 ( .B1(n19207), .B2(n13265), .A(n13283), .ZN(n13288) );
  OAI21_X1 U16492 ( .B1(n10138), .B2(n13285), .A(n13284), .ZN(n13286) );
  INV_X1 U16493 ( .A(n13286), .ZN(n19232) );
  AOI22_X1 U16494 ( .A1(n19232), .A2(n19204), .B1(P2_REIP_REG_2__SCAN_IN), 
        .B2(n19030), .ZN(n13287) );
  OAI211_X1 U16495 ( .C1(n16262), .C2(n13289), .A(n13288), .B(n13287), .ZN(
        P2_U3012) );
  OR2_X1 U16496 ( .A1(n9761), .A2(n12355), .ZN(n13334) );
  INV_X1 U16497 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14444) );
  INV_X1 U16498 ( .A(n20022), .ZN(n13294) );
  INV_X1 U16499 ( .A(n20116), .ZN(n20114) );
  INV_X1 U16500 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13292) );
  NOR2_X1 U16501 ( .A1(n20114), .A2(n13292), .ZN(n13293) );
  AOI21_X1 U16502 ( .B1(DATAI_15_), .B2(n20114), .A(n13293), .ZN(n14445) );
  INV_X1 U16503 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20010) );
  OAI222_X1 U16504 ( .A1(n13334), .A2(n14444), .B1(n13294), .B2(n14445), .C1(
        n13356), .C2(n20010), .ZN(P1_U2967) );
  OAI21_X1 U16505 ( .B1(n13296), .B2(n13295), .A(n13431), .ZN(n14298) );
  INV_X1 U16506 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n13735) );
  OAI22_X1 U16507 ( .A1(n14518), .A2(n13298), .B1(n16045), .B2(n13735), .ZN(
        n13297) );
  AOI21_X1 U16508 ( .B1(n15919), .B2(n13298), .A(n13297), .ZN(n13303) );
  NOR2_X1 U16509 ( .A1(n13299), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20087) );
  INV_X1 U16510 ( .A(n20087), .ZN(n13301) );
  NAND3_X1 U16511 ( .A1(n13301), .A2(n20046), .A3(n13300), .ZN(n13302) );
  OAI211_X1 U16512 ( .C1(n20115), .C2(n14298), .A(n13303), .B(n13302), .ZN(
        P1_U2998) );
  OAI21_X1 U16513 ( .B1(n14836), .B2(n13305), .A(n13304), .ZN(n13306) );
  XNOR2_X1 U16514 ( .A(n13306), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15343) );
  INV_X1 U16515 ( .A(n15343), .ZN(n13310) );
  AOI21_X1 U16516 ( .B1(n15370), .B2(n13308), .A(n13307), .ZN(n15342) );
  AOI22_X1 U16517 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16247), .B1(
        n19204), .B2(n15342), .ZN(n13309) );
  NAND2_X1 U16518 ( .A1(n19030), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n15344) );
  OAI211_X1 U16519 ( .C1(n16263), .C2(n13310), .A(n13309), .B(n15344), .ZN(
        n13311) );
  AOI21_X1 U16520 ( .B1(n19203), .B2(n14833), .A(n13311), .ZN(n13312) );
  OAI21_X1 U16521 ( .B1(n13313), .B2(n13644), .A(n13312), .ZN(P2_U3013) );
  NOR2_X1 U16522 ( .A1(n13193), .A2(n13315), .ZN(n13316) );
  NAND2_X1 U16523 ( .A1(n11472), .A2(n11456), .ZN(n13324) );
  AND2_X1 U16524 ( .A1(n13324), .A2(n14088), .ZN(n13321) );
  NAND2_X1 U16525 ( .A1(n20114), .A2(DATAI_1_), .ZN(n13323) );
  NAND2_X1 U16526 ( .A1(n20116), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13322) );
  AND2_X1 U16527 ( .A1(n13323), .A2(n13322), .ZN(n20133) );
  INV_X1 U16528 ( .A(n13324), .ZN(n13325) );
  AND2_X1 U16529 ( .A1(n20001), .A2(n13234), .ZN(n13326) );
  OAI222_X1 U16530 ( .A1(n14298), .A2(n20004), .B1(n20133), .B2(n20003), .C1(
        n20001), .C2(n11841), .ZN(P1_U2903) );
  INV_X1 U16531 ( .A(n13133), .ZN(n13328) );
  INV_X1 U16532 ( .A(n13685), .ZN(n13330) );
  NAND2_X1 U16533 ( .A1(n13331), .A2(n13330), .ZN(n13332) );
  AOI222_X1 U16534 ( .A1(n20007), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n20008), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .C1(n20006), .C2(P1_LWORD_REG_4__SCAN_IN), .ZN(n13333) );
  INV_X1 U16535 ( .A(n13333), .ZN(P1_U2932) );
  AOI22_X1 U16536 ( .A1(n20036), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n9761), .ZN(n13337) );
  NAND2_X1 U16537 ( .A1(n20114), .A2(DATAI_6_), .ZN(n13336) );
  NAND2_X1 U16538 ( .A1(n20116), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13335) );
  INV_X1 U16539 ( .A(n20168), .ZN(n14416) );
  NAND2_X1 U16540 ( .A1(n20022), .A2(n14416), .ZN(n13369) );
  NAND2_X1 U16541 ( .A1(n13337), .A2(n13369), .ZN(P1_U2958) );
  AOI22_X1 U16542 ( .A1(n20036), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n9761), .ZN(n13339) );
  NAND2_X1 U16543 ( .A1(n20116), .A2(n16513), .ZN(n13338) );
  OAI21_X1 U16544 ( .B1(n20116), .B2(DATAI_0_), .A(n13338), .ZN(n20122) );
  INV_X1 U16545 ( .A(n20122), .ZN(n14439) );
  NAND2_X1 U16546 ( .A1(n20022), .A2(n14439), .ZN(n13359) );
  NAND2_X1 U16547 ( .A1(n13339), .A2(n13359), .ZN(P1_U2952) );
  AOI22_X1 U16548 ( .A1(n20036), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n9761), .ZN(n13340) );
  INV_X1 U16549 ( .A(n20133), .ZN(n14434) );
  NAND2_X1 U16550 ( .A1(n20022), .A2(n14434), .ZN(n13357) );
  NAND2_X1 U16551 ( .A1(n13340), .A2(n13357), .ZN(P1_U2953) );
  AOI22_X1 U16552 ( .A1(n20036), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n9761), .ZN(n13342) );
  INV_X1 U16553 ( .A(DATAI_7_), .ZN(n21076) );
  NAND2_X1 U16554 ( .A1(n20116), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13341) );
  OAI21_X1 U16555 ( .B1(n20116), .B2(n21076), .A(n13341), .ZN(n14412) );
  NAND2_X1 U16556 ( .A1(n20022), .A2(n14412), .ZN(n13365) );
  NAND2_X1 U16557 ( .A1(n13342), .A2(n13365), .ZN(P1_U2944) );
  AOI22_X1 U16558 ( .A1(n20036), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n9761), .ZN(n13345) );
  NAND2_X1 U16559 ( .A1(n20114), .A2(DATAI_3_), .ZN(n13344) );
  NAND2_X1 U16560 ( .A1(n20116), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13343) );
  AND2_X1 U16561 ( .A1(n13344), .A2(n13343), .ZN(n20147) );
  INV_X1 U16562 ( .A(n20147), .ZN(n14426) );
  NAND2_X1 U16563 ( .A1(n20022), .A2(n14426), .ZN(n13363) );
  NAND2_X1 U16564 ( .A1(n13345), .A2(n13363), .ZN(P1_U2955) );
  AOI22_X1 U16565 ( .A1(n20036), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n9761), .ZN(n13348) );
  NAND2_X1 U16566 ( .A1(n20114), .A2(DATAI_4_), .ZN(n13347) );
  NAND2_X1 U16567 ( .A1(n20116), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13346) );
  AND2_X1 U16568 ( .A1(n13347), .A2(n13346), .ZN(n20154) );
  INV_X1 U16569 ( .A(n20154), .ZN(n14423) );
  NAND2_X1 U16570 ( .A1(n20022), .A2(n14423), .ZN(n13371) );
  NAND2_X1 U16571 ( .A1(n13348), .A2(n13371), .ZN(P1_U2956) );
  AOI22_X1 U16572 ( .A1(n20036), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n9761), .ZN(n13351) );
  NAND2_X1 U16573 ( .A1(n20114), .A2(DATAI_5_), .ZN(n13350) );
  NAND2_X1 U16574 ( .A1(n20116), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13349) );
  AND2_X1 U16575 ( .A1(n13350), .A2(n13349), .ZN(n20162) );
  INV_X1 U16576 ( .A(n20162), .ZN(n14419) );
  NAND2_X1 U16577 ( .A1(n20022), .A2(n14419), .ZN(n13367) );
  NAND2_X1 U16578 ( .A1(n13351), .A2(n13367), .ZN(P1_U2957) );
  AOI22_X1 U16579 ( .A1(n20036), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n9761), .ZN(n13352) );
  MUX2_X1 U16580 ( .A(DATAI_11_), .B(BUF1_REG_11__SCAN_IN), .S(n20116), .Z(
        n15882) );
  NAND2_X1 U16581 ( .A1(n20022), .A2(n15882), .ZN(n20030) );
  NAND2_X1 U16582 ( .A1(n13352), .A2(n20030), .ZN(P1_U2948) );
  AOI22_X1 U16583 ( .A1(n20036), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n9761), .ZN(n13355) );
  NAND2_X1 U16584 ( .A1(n20114), .A2(DATAI_2_), .ZN(n13354) );
  NAND2_X1 U16585 ( .A1(n20116), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13353) );
  AND2_X1 U16586 ( .A1(n13354), .A2(n13353), .ZN(n20138) );
  INV_X1 U16587 ( .A(n20138), .ZN(n14430) );
  NAND2_X1 U16588 ( .A1(n20022), .A2(n14430), .ZN(n13361) );
  NAND2_X1 U16589 ( .A1(n13355), .A2(n13361), .ZN(P1_U2954) );
  AOI22_X1 U16590 ( .A1(n20036), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n9761), .ZN(n13358) );
  NAND2_X1 U16591 ( .A1(n13358), .A2(n13357), .ZN(P1_U2938) );
  AOI22_X1 U16592 ( .A1(n20036), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n9761), .ZN(n13360) );
  NAND2_X1 U16593 ( .A1(n13360), .A2(n13359), .ZN(P1_U2937) );
  AOI22_X1 U16594 ( .A1(n20036), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n9761), .ZN(n13362) );
  NAND2_X1 U16595 ( .A1(n13362), .A2(n13361), .ZN(P1_U2939) );
  AOI22_X1 U16596 ( .A1(n20036), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n9761), .ZN(n13364) );
  NAND2_X1 U16597 ( .A1(n13364), .A2(n13363), .ZN(P1_U2940) );
  AOI22_X1 U16598 ( .A1(n20036), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n9761), .ZN(n13366) );
  NAND2_X1 U16599 ( .A1(n13366), .A2(n13365), .ZN(P1_U2959) );
  AOI22_X1 U16600 ( .A1(n20036), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n9761), .ZN(n13368) );
  NAND2_X1 U16601 ( .A1(n13368), .A2(n13367), .ZN(P1_U2942) );
  AOI22_X1 U16602 ( .A1(n20036), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n9761), .ZN(n13370) );
  NAND2_X1 U16603 ( .A1(n13370), .A2(n13369), .ZN(P1_U2943) );
  AOI22_X1 U16604 ( .A1(n20036), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n9761), .ZN(n13372) );
  NAND2_X1 U16605 ( .A1(n13372), .A2(n13371), .ZN(P1_U2941) );
  XNOR2_X1 U16606 ( .A(n13373), .B(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13379) );
  NAND2_X1 U16607 ( .A1(n13375), .A2(n13376), .ZN(n13377) );
  NAND2_X1 U16608 ( .A1(n13374), .A2(n13377), .ZN(n19035) );
  MUX2_X1 U16609 ( .A(n20987), .B(n19035), .S(n14901), .Z(n13378) );
  OAI21_X1 U16610 ( .B1(n13379), .B2(n14911), .A(n13378), .ZN(P2_U2881) );
  INV_X1 U16611 ( .A(n13380), .ZN(n13382) );
  INV_X1 U16612 ( .A(n13373), .ZN(n13381) );
  OAI211_X1 U16613 ( .C1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .C2(n13382), .A(
        n13381), .B(n14894), .ZN(n13385) );
  OAI21_X1 U16614 ( .B1(n13762), .B2(n13383), .A(n13375), .ZN(n13858) );
  INV_X1 U16615 ( .A(n13858), .ZN(n19049) );
  NAND2_X1 U16616 ( .A1(n19049), .A2(n14901), .ZN(n13384) );
  OAI211_X1 U16617 ( .C1(n14901), .C2(n13386), .A(n13385), .B(n13384), .ZN(
        P2_U2882) );
  INV_X1 U16618 ( .A(n20416), .ZN(n13477) );
  INV_X1 U16619 ( .A(n14655), .ZN(n13400) );
  XNOR2_X1 U16620 ( .A(n13388), .B(n13387), .ZN(n13398) );
  INV_X1 U16621 ( .A(n13389), .ZN(n13390) );
  NOR2_X1 U16622 ( .A1(n13391), .A2(n13390), .ZN(n13405) );
  MUX2_X1 U16623 ( .A(n13392), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n13393), .Z(n13394) );
  INV_X1 U16624 ( .A(n9786), .ZN(n13401) );
  INV_X1 U16625 ( .A(n13392), .ZN(n13395) );
  OAI211_X1 U16626 ( .C1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C2(n13393), .A(
        n9784), .B(n13395), .ZN(n20820) );
  NOR3_X1 U16627 ( .A1(n14655), .A2(n13401), .A3(n20820), .ZN(n13396) );
  AOI211_X1 U16628 ( .C1(n13403), .C2(n13398), .A(n13397), .B(n13396), .ZN(
        n13399) );
  OAI21_X1 U16629 ( .B1(n13477), .B2(n13400), .A(n13399), .ZN(n20819) );
  MUX2_X1 U16630 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n20819), .S(
        n15719), .Z(n15730) );
  NOR2_X1 U16631 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n20739), .ZN(n13415) );
  AOI22_X1 U16632 ( .A1(n15730), .A2(n20739), .B1(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13415), .ZN(n13410) );
  INV_X1 U16633 ( .A(n20552), .ZN(n20111) );
  XNOR2_X1 U16634 ( .A(n13393), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13402) );
  NOR3_X1 U16635 ( .A1(n14655), .A2(n13401), .A3(n13402), .ZN(n13407) );
  INV_X1 U16636 ( .A(n13402), .ZN(n14660) );
  INV_X1 U16637 ( .A(n13403), .ZN(n14651) );
  XNOR2_X1 U16638 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13404) );
  OAI22_X1 U16639 ( .A1(n13405), .A2(n14660), .B1(n14651), .B2(n13404), .ZN(
        n13406) );
  AOI211_X1 U16640 ( .C1(n20111), .C2(n14655), .A(n13407), .B(n13406), .ZN(
        n14664) );
  NOR2_X1 U16641 ( .A1(n15719), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13408) );
  AOI21_X1 U16642 ( .B1(n14664), .B2(n15719), .A(n13408), .ZN(n15723) );
  AOI22_X1 U16643 ( .A1(n13415), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15723), .B2(n20739), .ZN(n13409) );
  INV_X1 U16644 ( .A(n20295), .ZN(n20551) );
  OR2_X1 U16645 ( .A1(n11590), .A2(n20551), .ZN(n13412) );
  XNOR2_X1 U16646 ( .A(n13412), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n19961) );
  NAND2_X1 U16647 ( .A1(n19961), .A2(n13413), .ZN(n16100) );
  NAND2_X1 U16648 ( .A1(n15719), .A2(n16100), .ZN(n13414) );
  OAI211_X1 U16649 ( .C1(n15719), .C2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n13414), .B(n20739), .ZN(n13417) );
  NAND2_X1 U16650 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n13415), .ZN(
        n13416) );
  AND2_X1 U16651 ( .A1(n13417), .A2(n13416), .ZN(n15736) );
  OAI21_X1 U16652 ( .B1(n15737), .B2(n13411), .A(n15736), .ZN(n13435) );
  OAI21_X1 U16653 ( .B1(n13435), .B2(P1_FLUSH_REG_SCAN_IN), .A(n13418), .ZN(
        n13419) );
  NAND2_X1 U16654 ( .A1(n20214), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20521) );
  XOR2_X1 U16655 ( .A(n20521), .B(n13420), .Z(n13421) );
  AND2_X1 U16656 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21100), .ZN(n14648) );
  OAI22_X1 U16657 ( .A1(n13421), .A2(n20836), .B1(n20552), .B2(n14648), .ZN(
        n13422) );
  NAND2_X1 U16658 ( .A1(n20104), .A2(n13422), .ZN(n13423) );
  OAI21_X1 U16659 ( .B1(n20104), .B2(n11766), .A(n13423), .ZN(P1_U3476) );
  OAI21_X1 U16660 ( .B1(n13424), .B2(n13426), .A(n13425), .ZN(n20077) );
  INV_X1 U16661 ( .A(n13429), .ZN(n13430) );
  AOI21_X1 U16662 ( .B1(n13428), .B2(n13431), .A(n13430), .ZN(n13439) );
  AOI22_X1 U16663 ( .A1(n20039), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20099), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13432) );
  OAI21_X1 U16664 ( .B1(n20050), .B2(n13736), .A(n13432), .ZN(n13433) );
  AOI21_X1 U16665 ( .B1(n13439), .B2(n20045), .A(n13433), .ZN(n13434) );
  OAI21_X1 U16666 ( .B1(n19904), .B2(n20077), .A(n13434), .ZN(P1_U2997) );
  NOR2_X1 U16667 ( .A1(n13435), .A2(n16112), .ZN(n15745) );
  INV_X1 U16668 ( .A(n11849), .ZN(n13436) );
  OAI22_X1 U16669 ( .A1(n11846), .A2(n20836), .B1(n13436), .B2(n14648), .ZN(
        n13437) );
  OAI21_X1 U16670 ( .B1(n15745), .B2(n13437), .A(n20104), .ZN(n13438) );
  OAI21_X1 U16671 ( .B1(n20104), .B2(n20611), .A(n13438), .ZN(P1_U3478) );
  INV_X1 U16672 ( .A(n13439), .ZN(n13745) );
  OAI222_X1 U16673 ( .A1(n13745), .A2(n20004), .B1(n20138), .B2(n20003), .C1(
        n20001), .C2(n11831), .ZN(P1_U2902) );
  NAND2_X1 U16674 ( .A1(n13441), .A2(n13440), .ZN(n13444) );
  INV_X1 U16675 ( .A(n13442), .ZN(n13443) );
  NAND2_X1 U16676 ( .A1(n13444), .A2(n13443), .ZN(n19866) );
  INV_X1 U16677 ( .A(n19866), .ZN(n13454) );
  XNOR2_X1 U16678 ( .A(n19864), .B(n19866), .ZN(n13450) );
  XNOR2_X1 U16679 ( .A(n13446), .B(n13445), .ZN(n19875) );
  NOR2_X1 U16680 ( .A1(n19852), .A2(n19875), .ZN(n13447) );
  AOI21_X1 U16681 ( .B1(n19875), .B2(n19852), .A(n13447), .ZN(n19130) );
  NAND2_X1 U16682 ( .A1(n19130), .A2(n19129), .ZN(n19128) );
  INV_X1 U16683 ( .A(n13447), .ZN(n13448) );
  NAND2_X1 U16684 ( .A1(n19128), .A2(n13448), .ZN(n13449) );
  NAND2_X1 U16685 ( .A1(n13449), .A2(n13450), .ZN(n13598) );
  OAI21_X1 U16686 ( .B1(n13450), .B2(n13449), .A(n13598), .ZN(n13451) );
  NAND2_X1 U16687 ( .A1(n13451), .A2(n19131), .ZN(n13453) );
  AOI22_X1 U16688 ( .A1(n19102), .A2(n16199), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19126), .ZN(n13452) );
  OAI211_X1 U16689 ( .C1(n13454), .C2(n19084), .A(n13453), .B(n13452), .ZN(
        P2_U2917) );
  NAND2_X1 U16690 ( .A1(n13456), .A2(n13455), .ZN(n13457) );
  AND2_X1 U16691 ( .A1(n13468), .A2(n13457), .ZN(n20075) );
  INV_X1 U16692 ( .A(n20000), .ZN(n14381) );
  AOI22_X1 U16693 ( .A1(n19995), .A2(n20075), .B1(n14381), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n13458) );
  OAI21_X1 U16694 ( .B1(n13745), .B2(n14389), .A(n13458), .ZN(P1_U2870) );
  OR2_X1 U16695 ( .A1(n13460), .A2(n13459), .ZN(n13462) );
  AND2_X1 U16696 ( .A1(n13462), .A2(n13461), .ZN(n20103) );
  INV_X1 U16697 ( .A(n20103), .ZN(n14301) );
  AOI22_X1 U16698 ( .A1(n19995), .A2(n14301), .B1(n14381), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13463) );
  OAI21_X1 U16699 ( .B1(n14389), .B2(n14298), .A(n13463), .ZN(P1_U2871) );
  INV_X1 U16700 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n14306) );
  OAI222_X1 U16701 ( .A1(n14307), .A2(n19986), .B1(n20000), .B2(n14306), .C1(
        n20005), .C2(n14389), .ZN(P1_U2872) );
  NOR2_X1 U16702 ( .A1(n13465), .A2(n13464), .ZN(n13466) );
  AND2_X1 U16703 ( .A1(n13468), .A2(n13467), .ZN(n13469) );
  NOR2_X1 U16704 ( .A1(n13570), .A2(n13469), .ZN(n20063) );
  AOI22_X1 U16705 ( .A1(n19995), .A2(n20063), .B1(n14381), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n13470) );
  OAI21_X1 U16706 ( .B1(n13566), .B2(n14389), .A(n13470), .ZN(P1_U2869) );
  OAI21_X1 U16707 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n20107), .A(n20522), 
        .ZN(n13473) );
  NAND2_X1 U16708 ( .A1(n20613), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13472) );
  NOR2_X1 U16709 ( .A1(n20214), .A2(n13472), .ZN(n20323) );
  AND2_X1 U16710 ( .A1(n20679), .A2(n20323), .ZN(n20616) );
  AOI21_X1 U16711 ( .B1(n20613), .B2(n13473), .A(n20616), .ZN(n13476) );
  NOR2_X1 U16712 ( .A1(n20521), .A2(n20836), .ZN(n20680) );
  AND2_X1 U16713 ( .A1(n20389), .A2(n20680), .ZN(n20393) );
  INV_X1 U16714 ( .A(n20393), .ZN(n13475) );
  OAI211_X1 U16715 ( .C1(n13477), .C2(n14648), .A(n13476), .B(n13475), .ZN(
        n13478) );
  NAND2_X1 U16716 ( .A1(n20104), .A2(n13478), .ZN(n13479) );
  OAI21_X1 U16717 ( .B1(n20104), .B2(n20515), .A(n13479), .ZN(P1_U3475) );
  INV_X1 U16718 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n13481) );
  INV_X1 U16719 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14409) );
  INV_X2 U16720 ( .A(n20006), .ZN(n20837) );
  INV_X1 U16721 ( .A(P1_UWORD_REG_7__SCAN_IN), .ZN(n13480) );
  OAI222_X1 U16722 ( .A1(n13481), .A2(n13553), .B1(n13517), .B2(n14409), .C1(
        n20837), .C2(n13480), .ZN(P1_U2913) );
  INV_X1 U16723 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13483) );
  INV_X1 U16724 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n14397) );
  INV_X1 U16725 ( .A(P1_UWORD_REG_11__SCAN_IN), .ZN(n13482) );
  OAI222_X1 U16726 ( .A1(n13483), .A2(n13553), .B1(n13517), .B2(n14397), .C1(
        n20837), .C2(n13482), .ZN(P1_U2909) );
  OAI222_X1 U16727 ( .A1(n13566), .A2(n20004), .B1(n20147), .B2(n20003), .C1(
        n20001), .C2(n11827), .ZN(P1_U2901) );
  INV_X1 U16728 ( .A(P1_UWORD_REG_12__SCAN_IN), .ZN(n13486) );
  INV_X1 U16729 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13485) );
  INV_X1 U16730 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13484) );
  OAI222_X1 U16731 ( .A1(n13486), .A2(n20837), .B1(n13517), .B2(n13485), .C1(
        n13553), .C2(n13484), .ZN(P1_U2908) );
  INV_X1 U16732 ( .A(P1_UWORD_REG_3__SCAN_IN), .ZN(n13488) );
  INV_X1 U16733 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n13487) );
  OAI222_X1 U16734 ( .A1(n13488), .A2(n20837), .B1(n13517), .B2(n12084), .C1(
        n13553), .C2(n13487), .ZN(P1_U2917) );
  INV_X1 U16735 ( .A(P1_UWORD_REG_9__SCAN_IN), .ZN(n13491) );
  INV_X1 U16736 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13490) );
  INV_X1 U16737 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13489) );
  OAI222_X1 U16738 ( .A1(n13491), .A2(n20837), .B1(n13517), .B2(n13490), .C1(
        n13553), .C2(n13489), .ZN(P1_U2911) );
  INV_X1 U16739 ( .A(P1_UWORD_REG_0__SCAN_IN), .ZN(n13494) );
  INV_X1 U16740 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13493) );
  INV_X1 U16741 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n13492) );
  OAI222_X1 U16742 ( .A1(n13494), .A2(n20837), .B1(n13517), .B2(n13493), .C1(
        n13553), .C2(n13492), .ZN(P1_U2920) );
  INV_X1 U16743 ( .A(P1_UWORD_REG_14__SCAN_IN), .ZN(n13496) );
  INV_X1 U16744 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13495) );
  OAI222_X1 U16745 ( .A1(n13496), .A2(n20837), .B1(n13517), .B2(n12342), .C1(
        n13553), .C2(n13495), .ZN(P1_U2906) );
  INV_X1 U16746 ( .A(P1_UWORD_REG_1__SCAN_IN), .ZN(n13498) );
  INV_X1 U16747 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n13497) );
  OAI222_X1 U16748 ( .A1(n13498), .A2(n20837), .B1(n13517), .B2(n11982), .C1(
        n13553), .C2(n13497), .ZN(P1_U2919) );
  INV_X1 U16749 ( .A(P1_UWORD_REG_13__SCAN_IN), .ZN(n13501) );
  INV_X1 U16750 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13500) );
  INV_X1 U16751 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13499) );
  OAI222_X1 U16752 ( .A1(n13501), .A2(n20837), .B1(n13517), .B2(n13500), .C1(
        n13553), .C2(n13499), .ZN(P1_U2907) );
  INV_X1 U16753 ( .A(P1_UWORD_REG_6__SCAN_IN), .ZN(n13504) );
  INV_X1 U16754 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13503) );
  INV_X1 U16755 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n13502) );
  OAI222_X1 U16756 ( .A1(n13504), .A2(n20837), .B1(n13517), .B2(n13503), .C1(
        n13553), .C2(n13502), .ZN(P1_U2914) );
  INV_X1 U16757 ( .A(P1_UWORD_REG_5__SCAN_IN), .ZN(n13506) );
  INV_X1 U16758 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n13505) );
  OAI222_X1 U16759 ( .A1(n13506), .A2(n20837), .B1(n13517), .B2(n12128), .C1(
        n13553), .C2(n13505), .ZN(P1_U2915) );
  INV_X1 U16760 ( .A(P1_UWORD_REG_2__SCAN_IN), .ZN(n13509) );
  INV_X1 U16761 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13508) );
  INV_X1 U16762 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n13507) );
  OAI222_X1 U16763 ( .A1(n13509), .A2(n20837), .B1(n13517), .B2(n13508), .C1(
        n13553), .C2(n13507), .ZN(P1_U2918) );
  INV_X1 U16764 ( .A(P1_UWORD_REG_10__SCAN_IN), .ZN(n13512) );
  INV_X1 U16765 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13511) );
  INV_X1 U16766 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13510) );
  OAI222_X1 U16767 ( .A1(n13512), .A2(n20837), .B1(n13517), .B2(n13511), .C1(
        n13553), .C2(n13510), .ZN(P1_U2910) );
  INV_X1 U16768 ( .A(P1_UWORD_REG_8__SCAN_IN), .ZN(n13515) );
  INV_X1 U16769 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13514) );
  INV_X1 U16770 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n13513) );
  OAI222_X1 U16771 ( .A1(n13515), .A2(n20837), .B1(n13517), .B2(n13514), .C1(
        n13553), .C2(n13513), .ZN(P1_U2912) );
  INV_X1 U16772 ( .A(P1_UWORD_REG_4__SCAN_IN), .ZN(n13518) );
  INV_X1 U16773 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n13516) );
  OAI222_X1 U16774 ( .A1(n13518), .A2(n20837), .B1(n13517), .B2(n12111), .C1(
        n13553), .C2(n13516), .ZN(P1_U2916) );
  XOR2_X1 U16775 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(n13581), .Z(n13522)
         );
  OR2_X1 U16776 ( .A1(n13374), .A2(n13519), .ZN(n13578) );
  NAND2_X1 U16777 ( .A1(n13374), .A2(n13519), .ZN(n13520) );
  NAND2_X1 U16778 ( .A1(n13578), .A2(n13520), .ZN(n19021) );
  MUX2_X1 U16779 ( .A(n19021), .B(n10840), .S(n13168), .Z(n13521) );
  OAI21_X1 U16780 ( .B1(n13522), .B2(n14911), .A(n13521), .ZN(P2_U2880) );
  INV_X1 U16781 ( .A(P1_LWORD_REG_9__SCAN_IN), .ZN(n13525) );
  INV_X1 U16782 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n13524) );
  INV_X1 U16783 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n13523) );
  OAI222_X1 U16784 ( .A1(n13525), .A2(n20837), .B1(n13556), .B2(n13524), .C1(
        n13523), .C2(n13553), .ZN(P1_U2927) );
  INV_X1 U16785 ( .A(P1_LWORD_REG_2__SCAN_IN), .ZN(n13527) );
  INV_X1 U16786 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n13526) );
  OAI222_X1 U16787 ( .A1(n13527), .A2(n20837), .B1(n11831), .B2(n13556), .C1(
        n13526), .C2(n13553), .ZN(P1_U2934) );
  INV_X1 U16788 ( .A(P1_LWORD_REG_14__SCAN_IN), .ZN(n13530) );
  INV_X1 U16789 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n13529) );
  INV_X1 U16790 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n13528) );
  OAI222_X1 U16791 ( .A1(n13530), .A2(n20837), .B1(n13556), .B2(n13529), .C1(
        n13528), .C2(n13553), .ZN(P1_U2922) );
  INV_X1 U16792 ( .A(P1_LWORD_REG_6__SCAN_IN), .ZN(n13532) );
  INV_X1 U16793 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n13531) );
  OAI222_X1 U16794 ( .A1(n13532), .A2(n20837), .B1(n13556), .B2(n13748), .C1(
        n13531), .C2(n13553), .ZN(P1_U2930) );
  INV_X1 U16795 ( .A(P1_LWORD_REG_5__SCAN_IN), .ZN(n13534) );
  INV_X1 U16796 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n13533) );
  OAI222_X1 U16797 ( .A1(n13534), .A2(n20837), .B1(n11870), .B2(n13556), .C1(
        n13533), .C2(n13553), .ZN(P1_U2931) );
  INV_X1 U16798 ( .A(P1_LWORD_REG_12__SCAN_IN), .ZN(n13536) );
  INV_X1 U16799 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n13535) );
  OAI222_X1 U16800 ( .A1(n13536), .A2(n20837), .B1(n13556), .B2(n12067), .C1(
        n13535), .C2(n13553), .ZN(P1_U2924) );
  INV_X1 U16801 ( .A(P1_LWORD_REG_13__SCAN_IN), .ZN(n13539) );
  INV_X1 U16802 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n13538) );
  INV_X1 U16803 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n13537) );
  OAI222_X1 U16804 ( .A1(n13539), .A2(n20837), .B1(n13556), .B2(n13538), .C1(
        n13537), .C2(n13553), .ZN(P1_U2923) );
  INV_X1 U16805 ( .A(P1_LWORD_REG_11__SCAN_IN), .ZN(n13541) );
  INV_X1 U16806 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n13540) );
  OAI222_X1 U16807 ( .A1(n13541), .A2(n20837), .B1(n13556), .B2(n11937), .C1(
        n13540), .C2(n13553), .ZN(P1_U2925) );
  INV_X1 U16808 ( .A(P1_LWORD_REG_7__SCAN_IN), .ZN(n13543) );
  INV_X1 U16809 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n13542) );
  OAI222_X1 U16810 ( .A1(n13543), .A2(n20837), .B1(n11885), .B2(n13556), .C1(
        n13542), .C2(n13553), .ZN(P1_U2929) );
  INV_X1 U16811 ( .A(P1_LWORD_REG_0__SCAN_IN), .ZN(n13545) );
  INV_X1 U16812 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20002) );
  INV_X1 U16813 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n13544) );
  OAI222_X1 U16814 ( .A1(n13545), .A2(n20837), .B1(n13556), .B2(n20002), .C1(
        n13544), .C2(n13553), .ZN(P1_U2936) );
  INV_X1 U16815 ( .A(P1_LWORD_REG_3__SCAN_IN), .ZN(n13547) );
  INV_X1 U16816 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n13546) );
  OAI222_X1 U16817 ( .A1(n13547), .A2(n20837), .B1(n11827), .B2(n13556), .C1(
        n13546), .C2(n13553), .ZN(P1_U2933) );
  INV_X1 U16818 ( .A(P1_LWORD_REG_8__SCAN_IN), .ZN(n13550) );
  INV_X1 U16819 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n13549) );
  INV_X1 U16820 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n13548) );
  OAI222_X1 U16821 ( .A1(n13550), .A2(n20837), .B1(n13556), .B2(n13549), .C1(
        n13548), .C2(n13553), .ZN(P1_U2928) );
  INV_X1 U16822 ( .A(P1_LWORD_REG_1__SCAN_IN), .ZN(n13552) );
  INV_X1 U16823 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n13551) );
  OAI222_X1 U16824 ( .A1(n13552), .A2(n20837), .B1(n11841), .B2(n13556), .C1(
        n13551), .C2(n13553), .ZN(P1_U2935) );
  INV_X1 U16825 ( .A(P1_LWORD_REG_10__SCAN_IN), .ZN(n13557) );
  INV_X1 U16826 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n13555) );
  INV_X1 U16827 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n13554) );
  OAI222_X1 U16828 ( .A1(n13557), .A2(n20837), .B1(n13556), .B2(n13555), .C1(
        n13554), .C2(n13553), .ZN(P1_U2926) );
  OR2_X1 U16829 ( .A1(n13560), .A2(n13559), .ZN(n13561) );
  NAND2_X1 U16830 ( .A1(n9765), .A2(n13561), .ZN(n20064) );
  INV_X1 U16831 ( .A(n13562), .ZN(n13691) );
  INV_X1 U16832 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n13563) );
  OAI22_X1 U16833 ( .A1(n14518), .A2(n13564), .B1(n16045), .B2(n13563), .ZN(
        n13565) );
  AOI21_X1 U16834 ( .B1(n13691), .B2(n15919), .A(n13565), .ZN(n13568) );
  INV_X1 U16835 ( .A(n13566), .ZN(n13697) );
  NAND2_X1 U16836 ( .A1(n13697), .A2(n20045), .ZN(n13567) );
  OAI211_X1 U16837 ( .C1(n20064), .C2(n19904), .A(n13568), .B(n13567), .ZN(
        P1_U2996) );
  OR2_X1 U16838 ( .A1(n13570), .A2(n13569), .ZN(n13571) );
  NAND2_X1 U16839 ( .A1(n16090), .A2(n13571), .ZN(n20058) );
  INV_X1 U16840 ( .A(n13572), .ZN(n13573) );
  XNOR2_X1 U16841 ( .A(n13574), .B(n13573), .ZN(n20044) );
  INV_X1 U16842 ( .A(n20044), .ZN(n13575) );
  INV_X1 U16843 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n19978) );
  OAI222_X1 U16844 ( .A1(n20058), .A2(n19986), .B1(n14389), .B2(n13575), .C1(
        n20000), .C2(n19978), .ZN(P1_U2868) );
  INV_X1 U16845 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n13576) );
  OAI222_X1 U16846 ( .A1(n20001), .A2(n13576), .B1(n20154), .B2(n20003), .C1(
        n20004), .C2(n13575), .ZN(P1_U2900) );
  AOI21_X1 U16847 ( .B1(n13579), .B2(n13578), .A(n13577), .ZN(n16321) );
  INV_X1 U16848 ( .A(n16321), .ZN(n14818) );
  INV_X1 U16849 ( .A(n13583), .ZN(n13585) );
  OAI211_X1 U16850 ( .C1(n13585), .C2(n13584), .A(n14894), .B(n13659), .ZN(
        n13587) );
  NAND2_X1 U16851 ( .A1(n13168), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13586) );
  OAI211_X1 U16852 ( .C1(n14818), .C2(n14909), .A(n13587), .B(n13586), .ZN(
        P2_U2879) );
  INV_X1 U16853 ( .A(n13588), .ZN(n13657) );
  XNOR2_X1 U16854 ( .A(n13659), .B(n13657), .ZN(n13593) );
  NOR2_X1 U16855 ( .A1(n13577), .A2(n13590), .ZN(n13591) );
  OR2_X1 U16856 ( .A1(n13589), .A2(n13591), .ZN(n19011) );
  MUX2_X1 U16857 ( .A(n19011), .B(n10845), .S(n13168), .Z(n13592) );
  OAI21_X1 U16858 ( .B1(n13593), .B2(n14911), .A(n13592), .ZN(P2_U2878) );
  NAND2_X1 U16859 ( .A1(n13595), .A2(n13594), .ZN(n13596) );
  AND2_X1 U16860 ( .A1(n13733), .A2(n13596), .ZN(n19997) );
  INV_X1 U16861 ( .A(n19997), .ZN(n13597) );
  OAI222_X1 U16862 ( .A1(n13597), .A2(n20004), .B1(n20162), .B2(n20003), .C1(
        n20001), .C2(n11870), .ZN(P1_U2899) );
  OAI21_X1 U16863 ( .B1(n15394), .B2(n19866), .A(n13598), .ZN(n19121) );
  OR2_X1 U16864 ( .A1(n13600), .A2(n13599), .ZN(n13602) );
  NAND2_X1 U16865 ( .A1(n13602), .A2(n13601), .ZN(n19119) );
  XOR2_X1 U16866 ( .A(n19119), .B(n19854), .Z(n19122) );
  NAND2_X1 U16867 ( .A1(n19121), .A2(n19122), .ZN(n19120) );
  NAND2_X1 U16868 ( .A1(n19854), .A2(n19119), .ZN(n13607) );
  XNOR2_X1 U16869 ( .A(n13601), .B(n13606), .ZN(n14148) );
  INV_X1 U16870 ( .A(n14148), .ZN(n13610) );
  AOI21_X1 U16871 ( .B1(n19120), .B2(n13607), .A(n13610), .ZN(n19114) );
  OAI21_X1 U16872 ( .B1(n13609), .B2(n13608), .A(n13380), .ZN(n19113) );
  XNOR2_X1 U16873 ( .A(n19114), .B(n19113), .ZN(n13613) );
  AOI22_X1 U16874 ( .A1(n19127), .A2(n13610), .B1(n19126), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n13612) );
  NAND2_X1 U16875 ( .A1(n19102), .A2(n19260), .ZN(n13611) );
  OAI211_X1 U16876 ( .C1(n13613), .C2(n19112), .A(n13612), .B(n13611), .ZN(
        P2_U2915) );
  XNOR2_X1 U16877 ( .A(n13615), .B(n13758), .ZN(n13616) );
  XNOR2_X1 U16878 ( .A(n13614), .B(n13616), .ZN(n13635) );
  NOR2_X1 U16879 ( .A1(n13617), .A2(n13644), .ZN(n13620) );
  INV_X1 U16880 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14160) );
  OAI21_X1 U16881 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n13618), .A(
        n14131), .ZN(n14157) );
  OAI22_X1 U16882 ( .A1(n14160), .A2(n19212), .B1(n16262), .B2(n14157), .ZN(
        n13619) );
  AOI211_X1 U16883 ( .C1(n19030), .C2(P2_REIP_REG_3__SCAN_IN), .A(n13620), .B(
        n13619), .ZN(n13625) );
  NAND2_X1 U16884 ( .A1(n13622), .A2(n13623), .ZN(n13632) );
  NAND3_X1 U16885 ( .A1(n13621), .A2(n13632), .A3(n19204), .ZN(n13624) );
  OAI211_X1 U16886 ( .C1(n13635), .C2(n16263), .A(n13625), .B(n13624), .ZN(
        P2_U3011) );
  INV_X1 U16887 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n19797) );
  NAND2_X1 U16888 ( .A1(n15245), .A2(n13627), .ZN(n19218) );
  NAND2_X1 U16889 ( .A1(n19218), .A2(n13628), .ZN(n15318) );
  AOI22_X1 U16890 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15318), .B1(
        n13763), .B2(n13758), .ZN(n13629) );
  OAI21_X1 U16891 ( .B1(n15334), .B2(n19797), .A(n13629), .ZN(n13631) );
  NOR2_X1 U16892 ( .A1(n19119), .A2(n15346), .ZN(n13630) );
  AOI211_X1 U16893 ( .C1(n19220), .C2(n13626), .A(n13631), .B(n13630), .ZN(
        n13634) );
  NAND3_X1 U16894 ( .A1(n13621), .A2(n13632), .A3(n19233), .ZN(n13633) );
  OAI211_X1 U16895 ( .C1(n13635), .C2(n19225), .A(n13634), .B(n13633), .ZN(
        P2_U3043) );
  OR2_X1 U16896 ( .A1(n19854), .A2(n19420), .ZN(n19643) );
  OR2_X1 U16897 ( .A1(n19861), .A2(n19415), .ZN(n19675) );
  OAI21_X1 U16898 ( .B1(n19643), .B2(n19451), .A(n19675), .ZN(n13638) );
  INV_X1 U16899 ( .A(n10476), .ZN(n13636) );
  AOI21_X1 U16900 ( .B1(n13636), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n13637) );
  NAND2_X1 U16901 ( .A1(n13638), .A2(n13637), .ZN(n13639) );
  NAND2_X1 U16902 ( .A1(n13639), .A2(n19239), .ZN(n13640) );
  NAND2_X1 U16903 ( .A1(n13640), .A2(n19683), .ZN(n19757) );
  INV_X1 U16904 ( .A(n19239), .ZN(n19752) );
  OAI21_X1 U16905 ( .B1(n10476), .B2(n19752), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13641) );
  OAI21_X1 U16906 ( .B1(n19675), .B2(n19513), .A(n13641), .ZN(n19754) );
  NOR2_X2 U16907 ( .A1(n13642), .A2(n19424), .ZN(n19690) );
  NOR2_X2 U16908 ( .A1(n14666), .A2(n19278), .ZN(n19676) );
  INV_X1 U16909 ( .A(n19676), .ZN(n13822) );
  INV_X1 U16910 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n20118) );
  INV_X1 U16911 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n18223) );
  AOI22_X1 U16912 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19275), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19274), .ZN(n19693) );
  INV_X1 U16913 ( .A(n19693), .ZN(n19652) );
  AOI22_X1 U16914 ( .A1(n19756), .A2(n19677), .B1(n19740), .B2(n19652), .ZN(
        n13646) );
  OAI21_X1 U16915 ( .B1(n13822), .B2(n19239), .A(n13646), .ZN(n13647) );
  AOI21_X1 U16916 ( .B1(n19754), .B2(n19690), .A(n13647), .ZN(n13648) );
  OAI21_X1 U16917 ( .B1(n19724), .B2(n13649), .A(n13648), .ZN(P2_U3168) );
  INV_X1 U16918 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13656) );
  INV_X1 U16919 ( .A(n16199), .ZN(n13650) );
  NOR2_X2 U16920 ( .A1(n13650), .A2(n19424), .ZN(n19699) );
  INV_X1 U16921 ( .A(n19278), .ZN(n13651) );
  INV_X1 U16922 ( .A(n19697), .ZN(n13653) );
  INV_X1 U16923 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n20139) );
  INV_X1 U16924 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n18233) );
  AOI22_X1 U16925 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19275), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19274), .ZN(n19702) );
  INV_X1 U16926 ( .A(n19702), .ZN(n19620) );
  AOI22_X1 U16927 ( .A1(n19740), .A2(n19698), .B1(n19756), .B2(n19620), .ZN(
        n13652) );
  OAI21_X1 U16928 ( .B1(n13653), .B2(n19239), .A(n13652), .ZN(n13654) );
  AOI21_X1 U16929 ( .B1(n19754), .B2(n19699), .A(n13654), .ZN(n13655) );
  OAI21_X1 U16930 ( .B1(n19724), .B2(n13656), .A(n13655), .ZN(P2_U3170) );
  INV_X1 U16931 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n13668) );
  NOR2_X1 U16932 ( .A1(n13659), .A2(n13657), .ZN(n13662) );
  INV_X1 U16933 ( .A(n13775), .ZN(n13660) );
  OAI211_X1 U16934 ( .C1(n13662), .C2(n13661), .A(n13660), .B(n14894), .ZN(
        n13667) );
  OR2_X1 U16935 ( .A1(n13589), .A2(n13664), .ZN(n13665) );
  AND2_X1 U16936 ( .A1(n13663), .A2(n13665), .ZN(n16313) );
  NAND2_X1 U16937 ( .A1(n16313), .A2(n14901), .ZN(n13666) );
  OAI211_X1 U16938 ( .C1(n14901), .C2(n13668), .A(n13667), .B(n13666), .ZN(
        P2_U2877) );
  AND2_X1 U16939 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n11495), .ZN(n13670) );
  NAND2_X1 U16940 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20843), .ZN(n16105) );
  INV_X1 U16941 ( .A(n16105), .ZN(n13669) );
  AOI22_X1 U16942 ( .A1(n13671), .A2(n13670), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n13669), .ZN(n13672) );
  NAND2_X1 U16943 ( .A1(n16045), .A2(n13672), .ZN(n13673) );
  INV_X1 U16944 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13973) );
  INV_X1 U16945 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14179) );
  NAND3_X1 U16946 ( .A1(n15776), .A2(P1_STATE2_REG_2__SCAN_IN), .A3(n13677), 
        .ZN(n13678) );
  NAND2_X1 U16947 ( .A1(n19926), .A2(n13678), .ZN(n19980) );
  AND2_X1 U16948 ( .A1(n11464), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13679) );
  AND2_X1 U16949 ( .A1(n16106), .A2(n20643), .ZN(n15741) );
  NAND2_X1 U16950 ( .A1(n12355), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13683) );
  INV_X1 U16951 ( .A(n13683), .ZN(n13681) );
  NOR2_X1 U16952 ( .A1(n13687), .A2(n13681), .ZN(n13682) );
  NOR2_X1 U16953 ( .A1(n13683), .A2(n15741), .ZN(n13684) );
  AOI22_X1 U16954 ( .A1(n19942), .A2(P1_EBX_REG_3__SCAN_IN), .B1(n19974), .B2(
        n20063), .ZN(n13695) );
  NOR2_X1 U16955 ( .A1(n13685), .A2(n20742), .ZN(n13686) );
  AND2_X1 U16956 ( .A1(n15776), .A2(n13686), .ZN(n19962) );
  OAI221_X1 U16957 ( .B1(n19937), .B2(P1_REIP_REG_1__SCAN_IN), .C1(n19937), 
        .C2(P1_REIP_REG_2__SCAN_IN), .A(n15776), .ZN(n13689) );
  AOI22_X1 U16958 ( .A1(n19962), .A2(n20416), .B1(n13689), .B2(
        P1_REIP_REG_3__SCAN_IN), .ZN(n13694) );
  AOI22_X1 U16959 ( .A1(n13691), .A2(n15861), .B1(n19960), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13693) );
  NAND4_X1 U16960 ( .A1(n19964), .A2(P1_REIP_REG_2__SCAN_IN), .A3(n13563), 
        .A4(P1_REIP_REG_1__SCAN_IN), .ZN(n13692) );
  NAND4_X1 U16961 ( .A1(n13695), .A2(n13694), .A3(n13693), .A4(n13692), .ZN(
        n13696) );
  AOI21_X1 U16962 ( .B1(n13697), .B2(n19980), .A(n13696), .ZN(n13698) );
  INV_X1 U16963 ( .A(n13698), .ZN(P1_U2837) );
  NAND2_X1 U16964 ( .A1(n13775), .A2(n13699), .ZN(n13783) );
  OAI211_X1 U16965 ( .C1(n13775), .C2(n13699), .A(n13783), .B(n14894), .ZN(
        n13703) );
  AOI21_X1 U16966 ( .B1(n13701), .B2(n13663), .A(n13700), .ZN(n15296) );
  NAND2_X1 U16967 ( .A1(n14901), .A2(n15296), .ZN(n13702) );
  OAI211_X1 U16968 ( .C1(n14901), .C2(n13704), .A(n13703), .B(n13702), .ZN(
        P2_U2876) );
  AND2_X1 U16969 ( .A1(n13775), .A2(n13705), .ZN(n13708) );
  NAND2_X1 U16970 ( .A1(n13775), .A2(n13706), .ZN(n13776) );
  OAI211_X1 U16971 ( .C1(n13708), .C2(n13707), .A(n14894), .B(n13776), .ZN(
        n13715) );
  NAND2_X1 U16972 ( .A1(n13710), .A2(n13709), .ZN(n13713) );
  INV_X1 U16973 ( .A(n13711), .ZN(n13712) );
  NAND2_X1 U16974 ( .A1(n13713), .A2(n13712), .ZN(n18989) );
  OR2_X1 U16975 ( .A1(n13168), .A2(n18989), .ZN(n13714) );
  OAI211_X1 U16976 ( .C1(n14901), .C2(n10861), .A(n13715), .B(n13714), .ZN(
        P2_U2872) );
  NAND2_X1 U16977 ( .A1(n19854), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19452) );
  OR2_X1 U16978 ( .A1(n19452), .A2(n19650), .ZN(n13716) );
  NAND2_X1 U16979 ( .A1(n13716), .A2(n19856), .ZN(n13723) );
  NAND3_X1 U16980 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19861), .A3(
        n19877), .ZN(n13812) );
  NOR2_X1 U16981 ( .A1(n19886), .A2(n13812), .ZN(n19422) );
  OAI21_X1 U16982 ( .B1(n13718), .B2(n19422), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13717) );
  INV_X1 U16983 ( .A(n19410), .ZN(n13729) );
  INV_X1 U16984 ( .A(n19690), .ZN(n13728) );
  INV_X1 U16985 ( .A(n13812), .ZN(n13722) );
  OR2_X1 U16986 ( .A1(n13718), .A2(n19544), .ZN(n13719) );
  AOI21_X1 U16987 ( .B1(n13719), .B2(n19680), .A(n19422), .ZN(n13720) );
  NOR2_X1 U16988 ( .A1(n19424), .A2(n13720), .ZN(n13721) );
  INV_X1 U16989 ( .A(n19409), .ZN(n19396) );
  AOI22_X1 U16990 ( .A1(n19652), .A2(n19443), .B1(n19676), .B2(n19422), .ZN(
        n13725) );
  OAI21_X1 U16991 ( .B1(n19655), .B2(n19396), .A(n13725), .ZN(n13726) );
  AOI21_X1 U16992 ( .B1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B2(n19407), .A(
        n13726), .ZN(n13727) );
  OAI21_X1 U16993 ( .B1(n13729), .B2(n13728), .A(n13727), .ZN(P2_U3088) );
  AND2_X1 U16994 ( .A1(n16092), .A2(n13730), .ZN(n13731) );
  OR2_X1 U16995 ( .A1(n13731), .A2(n16074), .ZN(n19944) );
  XOR2_X1 U16996 ( .A(n13733), .B(n13732), .Z(n19950) );
  INV_X1 U16997 ( .A(n19950), .ZN(n13747) );
  INV_X1 U16998 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n13734) );
  OAI222_X1 U16999 ( .A1(n19944), .A2(n19986), .B1(n14389), .B2(n13747), .C1(
        n20000), .C2(n13734), .ZN(P1_U2866) );
  INV_X1 U17000 ( .A(n19980), .ZN(n13746) );
  NOR3_X1 U17001 ( .A1(n19937), .A2(P1_REIP_REG_2__SCAN_IN), .A3(n13735), .ZN(
        n13743) );
  INV_X1 U17002 ( .A(n13736), .ZN(n13737) );
  AOI22_X1 U17003 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n19960), .B1(
        n15861), .B2(n13737), .ZN(n13741) );
  NAND2_X1 U17004 ( .A1(n19974), .A2(n20075), .ZN(n13740) );
  OAI21_X1 U17005 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19937), .A(n15776), .ZN(
        n13738) );
  AOI22_X1 U17006 ( .A1(n19962), .A2(n20111), .B1(P1_REIP_REG_2__SCAN_IN), 
        .B2(n13738), .ZN(n13739) );
  NAND3_X1 U17007 ( .A1(n13741), .A2(n13740), .A3(n13739), .ZN(n13742) );
  AOI211_X1 U17008 ( .C1(n19942), .C2(P1_EBX_REG_2__SCAN_IN), .A(n13743), .B(
        n13742), .ZN(n13744) );
  OAI21_X1 U17009 ( .B1(n13746), .B2(n13745), .A(n13744), .ZN(P1_U2838) );
  OAI222_X1 U17010 ( .A1(n20001), .A2(n13748), .B1(n20168), .B2(n20003), .C1(
        n20004), .C2(n13747), .ZN(P1_U2898) );
  OR2_X1 U17011 ( .A1(n9803), .A2(n13750), .ZN(n13751) );
  AND2_X1 U17012 ( .A1(n13749), .A2(n13751), .ZN(n19991) );
  INV_X1 U17013 ( .A(n19991), .ZN(n13752) );
  INV_X1 U17014 ( .A(n14412), .ZN(n20181) );
  OAI222_X1 U17015 ( .A1(n13752), .A2(n20004), .B1(n20181), .B2(n20003), .C1(
        n20001), .C2(n11885), .ZN(P1_U2897) );
  XOR2_X1 U17016 ( .A(n13753), .B(n13754), .Z(n19208) );
  INV_X1 U17017 ( .A(n19208), .ZN(n13770) );
  XNOR2_X1 U17018 ( .A(n13755), .B(n13866), .ZN(n13756) );
  XNOR2_X1 U17019 ( .A(n13757), .B(n13756), .ZN(n19205) );
  AOI21_X1 U17020 ( .B1(n13758), .B2(n16294), .A(n15318), .ZN(n13862) );
  NOR2_X1 U17021 ( .A1(n13760), .A2(n13759), .ZN(n13761) );
  OR2_X1 U17022 ( .A1(n13762), .A2(n13761), .ZN(n14128) );
  INV_X1 U17023 ( .A(n14128), .ZN(n19206) );
  NAND2_X1 U17024 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13763), .ZN(
        n15316) );
  INV_X1 U17025 ( .A(n15316), .ZN(n15332) );
  INV_X1 U17026 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n19799) );
  NOR2_X1 U17027 ( .A1(n19799), .A2(n15334), .ZN(n13764) );
  AOI21_X1 U17028 ( .B1(n13866), .B2(n15332), .A(n13764), .ZN(n13765) );
  OAI21_X1 U17029 ( .B1(n15346), .B2(n14148), .A(n13765), .ZN(n13766) );
  AOI21_X1 U17030 ( .B1(n19206), .B2(n19220), .A(n13766), .ZN(n13767) );
  OAI21_X1 U17031 ( .B1(n13862), .B2(n13866), .A(n13767), .ZN(n13768) );
  AOI21_X1 U17032 ( .B1(n19205), .B2(n19233), .A(n13768), .ZN(n13769) );
  OAI21_X1 U17033 ( .B1(n13770), .B2(n19225), .A(n13769), .ZN(P2_U3042) );
  OR2_X1 U17034 ( .A1(n13771), .A2(n13711), .ZN(n13772) );
  NAND2_X1 U17035 ( .A1(n13772), .A2(n9799), .ZN(n15258) );
  INV_X1 U17036 ( .A(n13773), .ZN(n13777) );
  AND2_X1 U17037 ( .A1(n13775), .A2(n13774), .ZN(n13805) );
  AOI21_X1 U17038 ( .B1(n13777), .B2(n13776), .A(n13805), .ZN(n19080) );
  NAND2_X1 U17039 ( .A1(n19080), .A2(n14894), .ZN(n13779) );
  NAND2_X1 U17040 ( .A1(n14909), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n13778) );
  OAI211_X1 U17041 ( .C1(n15258), .C2(n14909), .A(n13779), .B(n13778), .ZN(
        P2_U2871) );
  OAI21_X1 U17042 ( .B1(n13781), .B2(n13700), .A(n13780), .ZN(n16298) );
  INV_X1 U17043 ( .A(n13783), .ZN(n13828) );
  OR2_X1 U17044 ( .A1(n13783), .A2(n13782), .ZN(n13881) );
  OAI211_X1 U17045 ( .C1(n13828), .C2(n13784), .A(n14894), .B(n13881), .ZN(
        n13786) );
  NAND2_X1 U17046 ( .A1(n14909), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13785) );
  OAI211_X1 U17047 ( .C1(n16298), .C2(n14909), .A(n13786), .B(n13785), .ZN(
        P2_U2875) );
  INV_X1 U17048 ( .A(n13787), .ZN(n13788) );
  AOI21_X1 U17049 ( .B1(n13789), .B2(n13749), .A(n13788), .ZN(n13850) );
  INV_X1 U17050 ( .A(n13850), .ZN(n13834) );
  INV_X1 U17051 ( .A(n13848), .ZN(n13798) );
  OR2_X1 U17052 ( .A1(n16076), .A2(n13791), .ZN(n13792) );
  NAND2_X1 U17053 ( .A1(n13790), .A2(n13792), .ZN(n16066) );
  NAND4_X1 U17054 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n19963)
         );
  INV_X1 U17055 ( .A(n19963), .ZN(n13793) );
  INV_X1 U17056 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n21092) );
  NAND4_X1 U17057 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .A4(n21092), .ZN(n13794) );
  OAI22_X1 U17058 ( .A1(n19945), .A2(n16066), .B1(n19954), .B2(n13794), .ZN(
        n13797) );
  NAND4_X1 U17059 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .A3(P1_REIP_REG_6__SCAN_IN), .A4(P1_REIP_REG_5__SCAN_IN), .ZN(n14026)
         );
  NOR2_X1 U17060 ( .A1(n19963), .A2(n14026), .ZN(n14103) );
  OAI21_X1 U17061 ( .B1(n14103), .B2(n19937), .A(n15776), .ZN(n19924) );
  INV_X1 U17062 ( .A(n19924), .ZN(n14028) );
  AOI22_X1 U17063 ( .A1(n19942), .A2(P1_EBX_REG_8__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19960), .ZN(n13795) );
  NAND2_X1 U17064 ( .A1(n15776), .A2(n19892), .ZN(n19969) );
  OAI211_X1 U17065 ( .C1(n14028), .C2(n21092), .A(n13795), .B(n19969), .ZN(
        n13796) );
  AOI211_X1 U17066 ( .C1(n15861), .C2(n13798), .A(n13797), .B(n13796), .ZN(
        n13799) );
  OAI21_X1 U17067 ( .B1(n13834), .B2(n19926), .A(n13799), .ZN(P1_U2832) );
  INV_X1 U17068 ( .A(DATAI_8_), .ZN(n13801) );
  NAND2_X1 U17069 ( .A1(n20116), .A2(BUF1_REG_8__SCAN_IN), .ZN(n13800) );
  OAI21_X1 U17070 ( .B1(n20116), .B2(n13801), .A(n13800), .ZN(n20011) );
  AOI22_X1 U17071 ( .A1(n15883), .A2(n20011), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n15884), .ZN(n13802) );
  OAI21_X1 U17072 ( .B1(n13834), .B2(n20004), .A(n13802), .ZN(P1_U2896) );
  INV_X1 U17073 ( .A(n13803), .ZN(n13840) );
  OAI21_X1 U17074 ( .B1(n13805), .B2(n13804), .A(n13840), .ZN(n13896) );
  NAND2_X1 U17075 ( .A1(n14909), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n13809) );
  AOI21_X1 U17076 ( .B1(n13807), .B2(n9799), .A(n13806), .ZN(n18956) );
  NAND2_X1 U17077 ( .A1(n18956), .A2(n14901), .ZN(n13808) );
  OAI211_X1 U17078 ( .C1(n13896), .C2(n14911), .A(n13809), .B(n13808), .ZN(
        P2_U2870) );
  NOR2_X1 U17079 ( .A1(n13811), .A2(n13810), .ZN(n19609) );
  NAND2_X1 U17080 ( .A1(n19609), .A2(n19861), .ZN(n13817) );
  OAI21_X1 U17081 ( .B1(n19390), .B2(n19409), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n13814) );
  NOR2_X1 U17082 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13812), .ZN(
        n19388) );
  NOR2_X1 U17083 ( .A1(n19680), .A2(n19388), .ZN(n13813) );
  AOI21_X1 U17084 ( .B1(n13817), .B2(n13814), .A(n13813), .ZN(n13816) );
  INV_X1 U17085 ( .A(n19388), .ZN(n13821) );
  NAND3_X1 U17086 ( .A1(n13815), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n13821), 
        .ZN(n13819) );
  NAND3_X1 U17087 ( .A1(n19683), .A2(n13816), .A3(n13819), .ZN(n19391) );
  INV_X1 U17088 ( .A(n19391), .ZN(n13826) );
  OAI21_X1 U17089 ( .B1(n13817), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19544), 
        .ZN(n13818) );
  AOI22_X1 U17090 ( .A1(n19390), .A2(n19677), .B1(n19409), .B2(n19652), .ZN(
        n13820) );
  OAI21_X1 U17091 ( .B1(n13822), .B2(n13821), .A(n13820), .ZN(n13823) );
  AOI21_X1 U17092 ( .B1(n19389), .B2(n19690), .A(n13823), .ZN(n13824) );
  OAI21_X1 U17093 ( .B1(n13826), .B2(n13825), .A(n13824), .ZN(P2_U3080) );
  XNOR2_X1 U17094 ( .A(n13880), .B(n13829), .ZN(n13833) );
  OAI21_X1 U17095 ( .B1(n13831), .B2(n13830), .A(n13709), .ZN(n16234) );
  MUX2_X1 U17096 ( .A(n16234), .B(n10661), .S(n14909), .Z(n13832) );
  OAI21_X1 U17097 ( .B1(n13833), .B2(n14911), .A(n13832), .ZN(P2_U2873) );
  INV_X1 U17098 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13835) );
  OAI222_X1 U17099 ( .A1(n16066), .A2(n19986), .B1(n20000), .B2(n13835), .C1(
        n14389), .C2(n13834), .ZN(P1_U2864) );
  OR2_X1 U17100 ( .A1(n13836), .A2(n13806), .ZN(n13837) );
  NAND2_X1 U17101 ( .A1(n13837), .A2(n9958), .ZN(n18949) );
  INV_X1 U17102 ( .A(n13838), .ZN(n13841) );
  AOI21_X1 U17103 ( .B1(n13841), .B2(n13840), .A(n13839), .ZN(n16201) );
  NAND2_X1 U17104 ( .A1(n16201), .A2(n14894), .ZN(n13843) );
  NAND2_X1 U17105 ( .A1(n13168), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n13842) );
  OAI211_X1 U17106 ( .C1(n18949), .C2(n14909), .A(n13843), .B(n13842), .ZN(
        P2_U2869) );
  XNOR2_X1 U17107 ( .A(n13845), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13846) );
  XNOR2_X1 U17108 ( .A(n13844), .B(n13846), .ZN(n16067) );
  AOI22_X1 U17109 ( .A1(n20039), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n20099), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n13847) );
  OAI21_X1 U17110 ( .B1(n20050), .B2(n13848), .A(n13847), .ZN(n13849) );
  AOI21_X1 U17111 ( .B1(n13850), .B2(n20045), .A(n13849), .ZN(n13851) );
  OAI21_X1 U17112 ( .B1(n16067), .B2(n19904), .A(n13851), .ZN(P1_U2991) );
  XNOR2_X1 U17113 ( .A(n13853), .B(n13852), .ZN(n13875) );
  NAND2_X1 U17114 ( .A1(n13855), .A2(n13854), .ZN(n13856) );
  XNOR2_X1 U17115 ( .A(n9849), .B(n13856), .ZN(n13873) );
  OAI21_X1 U17116 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n14130), .A(
        n14688), .ZN(n19047) );
  OAI22_X1 U17117 ( .A1(n19212), .A2(n10071), .B1(n16262), .B2(n19047), .ZN(
        n13860) );
  INV_X1 U17118 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n13857) );
  OAI22_X1 U17119 ( .A1(n13858), .A2(n13644), .B1(n15334), .B2(n13857), .ZN(
        n13859) );
  AOI211_X1 U17120 ( .C1(n13873), .C2(n19204), .A(n13860), .B(n13859), .ZN(
        n13861) );
  OAI21_X1 U17121 ( .B1(n13875), .B2(n16263), .A(n13861), .ZN(P2_U3009) );
  NOR2_X1 U17122 ( .A1(n13862), .A2(n13867), .ZN(n13872) );
  OAI21_X1 U17123 ( .B1(n13865), .B2(n13864), .A(n13863), .ZN(n19117) );
  AOI221_X1 U17124 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(n13867), .C2(n13866), .A(
        n15316), .ZN(n13869) );
  NOR2_X1 U17125 ( .A1(n18957), .A2(n13857), .ZN(n13868) );
  AOI211_X1 U17126 ( .C1(n19049), .C2(n19220), .A(n13869), .B(n13868), .ZN(
        n13870) );
  OAI21_X1 U17127 ( .B1(n19117), .B2(n15346), .A(n13870), .ZN(n13871) );
  AOI211_X1 U17128 ( .C1(n13873), .C2(n19233), .A(n13872), .B(n13871), .ZN(
        n13874) );
  OAI21_X1 U17129 ( .B1(n13875), .B2(n19225), .A(n13874), .ZN(P2_U3041) );
  NAND2_X1 U17130 ( .A1(n13787), .A2(n13876), .ZN(n13877) );
  NAND2_X1 U17131 ( .A1(n9843), .A2(n13877), .ZN(n19987) );
  MUX2_X1 U17132 ( .A(DATAI_9_), .B(BUF1_REG_9__SCAN_IN), .S(n20116), .Z(
        n20013) );
  AOI22_X1 U17133 ( .A1(n15883), .A2(n20013), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n15884), .ZN(n13878) );
  OAI21_X1 U17134 ( .B1(n19987), .B2(n20004), .A(n13878), .ZN(P1_U2895) );
  AOI21_X1 U17135 ( .B1(n13879), .B2(n13780), .A(n13830), .ZN(n15282) );
  NOR2_X1 U17136 ( .A1(n14901), .A2(n10657), .ZN(n13884) );
  AOI211_X1 U17137 ( .C1(n13882), .C2(n13881), .A(n14911), .B(n13880), .ZN(
        n13883) );
  AOI211_X1 U17138 ( .C1(n15282), .C2(n14901), .A(n13884), .B(n13883), .ZN(
        n13885) );
  INV_X1 U17139 ( .A(n13885), .ZN(P2_U2874) );
  OR2_X1 U17140 ( .A1(n13887), .A2(n13886), .ZN(n13889) );
  NAND2_X1 U17141 ( .A1(n13889), .A2(n13888), .ZN(n18971) );
  INV_X1 U17142 ( .A(n18971), .ZN(n13894) );
  INV_X1 U17143 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n19165) );
  OAI22_X1 U17144 ( .A1(n14973), .A2(n19248), .B1(n19110), .B2(n19165), .ZN(
        n13893) );
  INV_X1 U17145 ( .A(n19078), .ZN(n14977) );
  INV_X1 U17146 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n13891) );
  INV_X1 U17147 ( .A(n19077), .ZN(n14975) );
  INV_X1 U17148 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n13890) );
  OAI22_X1 U17149 ( .A1(n14977), .A2(n13891), .B1(n14975), .B2(n13890), .ZN(
        n13892) );
  AOI211_X1 U17150 ( .C1(n19127), .C2(n13894), .A(n13893), .B(n13892), .ZN(
        n13895) );
  OAI21_X1 U17151 ( .B1(n13896), .B2(n19112), .A(n13895), .ZN(P2_U2902) );
  XNOR2_X1 U17152 ( .A(n14460), .B(n16059), .ZN(n13898) );
  XNOR2_X1 U17153 ( .A(n13897), .B(n13898), .ZN(n16055) );
  NAND2_X1 U17154 ( .A1(n16055), .A2(n20046), .ZN(n13903) );
  INV_X1 U17155 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n13899) );
  OAI22_X1 U17156 ( .A1(n14518), .A2(n19921), .B1(n16045), .B2(n13899), .ZN(
        n13900) );
  AOI21_X1 U17157 ( .B1(n15919), .B2(n13901), .A(n13900), .ZN(n13902) );
  OAI211_X1 U17158 ( .C1(n20115), .C2(n19987), .A(n13903), .B(n13902), .ZN(
        P1_U2990) );
  AND2_X1 U17159 ( .A1(n14905), .A2(n13905), .ZN(n13906) );
  NOR2_X1 U17160 ( .A1(n13904), .A2(n13906), .ZN(n16195) );
  NAND2_X1 U17161 ( .A1(n16195), .A2(n14894), .ZN(n13908) );
  NAND2_X1 U17162 ( .A1(n14909), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n13907) );
  OAI211_X1 U17163 ( .C1(n18924), .C2(n14909), .A(n13908), .B(n13907), .ZN(
        P2_U2867) );
  AOI21_X1 U17164 ( .B1(n9876), .B2(n9843), .A(n13909), .ZN(n14563) );
  NAND2_X1 U17165 ( .A1(n16053), .A2(n13910), .ZN(n13911) );
  NAND2_X1 U17166 ( .A1(n15867), .A2(n13911), .ZN(n16044) );
  OAI22_X1 U17167 ( .A1(n19986), .A2(n16044), .B1(n13912), .B2(n20000), .ZN(
        n13913) );
  AOI21_X1 U17168 ( .B1(n14563), .B2(n19996), .A(n13913), .ZN(n13914) );
  INV_X1 U17169 ( .A(n13914), .ZN(P1_U2862) );
  INV_X1 U17170 ( .A(n14563), .ZN(n14297) );
  MUX2_X1 U17171 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n20116), .Z(
        n20015) );
  AOI22_X1 U17172 ( .A1(n15883), .A2(n20015), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n15884), .ZN(n13915) );
  OAI21_X1 U17173 ( .B1(n14297), .B2(n20004), .A(n13915), .ZN(P1_U2894) );
  AOI21_X1 U17174 ( .B1(n18685), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13936) );
  OR2_X1 U17175 ( .A1(n18684), .A2(n13936), .ZN(n18669) );
  NOR2_X1 U17176 ( .A1(n18837), .A2(n18669), .ZN(n13935) );
  NAND2_X1 U17177 ( .A1(n13916), .A2(n15627), .ZN(n17407) );
  INV_X1 U17178 ( .A(n18660), .ZN(n15631) );
  NAND2_X1 U17179 ( .A1(n15631), .A2(n18875), .ZN(n13933) );
  AOI211_X1 U17180 ( .C1(n15635), .C2(n15773), .A(n13918), .B(n13917), .ZN(
        n15626) );
  OAI211_X1 U17181 ( .C1(n15626), .C2(n13921), .A(n13920), .B(n13919), .ZN(
        n13922) );
  INV_X1 U17182 ( .A(n13922), .ZN(n15637) );
  INV_X1 U17183 ( .A(n13923), .ZN(n13928) );
  OAI21_X1 U17184 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18217), .A(
        n13924), .ZN(n15632) );
  OR2_X1 U17185 ( .A1(n13925), .A2(n15632), .ZN(n13927) );
  OAI211_X1 U17186 ( .C1(n13928), .C2(n13927), .A(n15633), .B(n13926), .ZN(
        n16380) );
  INV_X1 U17187 ( .A(n16380), .ZN(n18666) );
  INV_X1 U17188 ( .A(n15643), .ZN(n13930) );
  AOI21_X1 U17189 ( .B1(n18666), .B2(n15642), .A(n15771), .ZN(n13932) );
  OAI211_X1 U17190 ( .C1(n17407), .C2(n13933), .A(n15637), .B(n13932), .ZN(
        n18691) );
  NOR2_X1 U17191 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18824), .ZN(n18220) );
  INV_X1 U17192 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18211) );
  NAND3_X1 U17193 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18822)
         );
  NOR2_X1 U17194 ( .A1(n18211), .A2(n18822), .ZN(n13934) );
  AOI211_X1 U17195 ( .C1(n18868), .C2(n18691), .A(n18220), .B(n13934), .ZN(
        n18854) );
  MUX2_X1 U17196 ( .A(n13935), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n18854), .Z(P3_U3284) );
  NAND2_X1 U17197 ( .A1(n13936), .A2(n17012), .ZN(n18210) );
  NOR2_X1 U17198 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18210), .ZN(n13937) );
  INV_X1 U17199 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18727) );
  OAI21_X1 U17200 ( .B1(n13937), .B2(n18822), .A(n18515), .ZN(n18216) );
  INV_X1 U17201 ( .A(n18216), .ZN(n13938) );
  NAND2_X1 U17202 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n17515) );
  INV_X1 U17203 ( .A(n17515), .ZN(n17843) );
  OAI21_X1 U17204 ( .B1(n18834), .B2(n18888), .A(n18824), .ZN(n18867) );
  NOR2_X1 U17205 ( .A1(n17843), .A2(n18867), .ZN(n15499) );
  AOI21_X1 U17206 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n15499), .ZN(n15500) );
  NOR2_X1 U17207 ( .A1(n13938), .A2(n15500), .ZN(n13940) );
  NAND2_X1 U17208 ( .A1(n18824), .A2(n18888), .ZN(n16556) );
  NOR2_X1 U17209 ( .A1(n18824), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18265) );
  OR2_X1 U17210 ( .A1(n18265), .A2(n13938), .ZN(n15498) );
  OR2_X1 U17211 ( .A1(n18470), .A2(n15498), .ZN(n13939) );
  MUX2_X1 U17212 ( .A(n13940), .B(n13939), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  NAND2_X1 U17213 ( .A1(n14994), .A2(n14993), .ZN(n13942) );
  XNOR2_X1 U17214 ( .A(n13941), .B(n13942), .ZN(n13964) );
  AOI21_X1 U17215 ( .B1(n15167), .B2(n15292), .A(n15166), .ZN(n15154) );
  INV_X1 U17216 ( .A(n15154), .ZN(n13956) );
  NOR2_X1 U17217 ( .A1(n13944), .A2(n13945), .ZN(n13946) );
  OR2_X1 U17218 ( .A1(n13943), .A2(n13946), .ZN(n16158) );
  INV_X1 U17219 ( .A(n13947), .ZN(n13948) );
  XNOR2_X1 U17220 ( .A(n14950), .B(n13948), .ZN(n16159) );
  NAND2_X1 U17221 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15168), .ZN(
        n15152) );
  OR2_X1 U17222 ( .A1(n18957), .A2(n21016), .ZN(n13959) );
  OAI21_X1 U17223 ( .B1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n15152), .A(
        n13959), .ZN(n13949) );
  AOI21_X1 U17224 ( .B1(n19228), .B2(n16159), .A(n13949), .ZN(n13950) );
  OAI21_X1 U17225 ( .B1(n16158), .B2(n16299), .A(n13950), .ZN(n13955) );
  INV_X1 U17226 ( .A(n13951), .ZN(n13952) );
  NOR2_X1 U17227 ( .A1(n13952), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13960) );
  NOR3_X1 U17228 ( .A1(n13960), .A2(n13953), .A3(n16318), .ZN(n13954) );
  AOI211_X1 U17229 ( .C1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n13956), .A(
        n13955), .B(n13954), .ZN(n13957) );
  OAI21_X1 U17230 ( .B1(n19225), .B2(n13964), .A(n13957), .ZN(P2_U3021) );
  AOI21_X1 U17231 ( .B1(n14708), .B2(n16155), .A(n14681), .ZN(n14683) );
  NAND2_X1 U17232 ( .A1(n16247), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13958) );
  OAI211_X1 U17233 ( .C1(n16158), .C2(n13644), .A(n13959), .B(n13958), .ZN(
        n13962) );
  NOR3_X1 U17234 ( .A1(n13960), .A2(n13953), .A3(n16265), .ZN(n13961) );
  AOI211_X1 U17235 ( .C1(n19203), .C2(n14683), .A(n13962), .B(n13961), .ZN(
        n13963) );
  OAI21_X1 U17236 ( .B1(n16263), .B2(n13964), .A(n13963), .ZN(P2_U2989) );
  NAND2_X1 U17237 ( .A1(n13965), .A2(n14460), .ZN(n14478) );
  NAND2_X1 U17238 ( .A1(n14459), .A2(n14478), .ZN(n13969) );
  NAND2_X1 U17239 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14588) );
  NAND2_X1 U17240 ( .A1(n14460), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14449) );
  INV_X1 U17241 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14580) );
  NAND2_X1 U17242 ( .A1(n15893), .A2(n14580), .ZN(n14450) );
  NOR2_X1 U17243 ( .A1(n14450), .A2(n9881), .ZN(n13970) );
  OR2_X2 U17244 ( .A1(n14093), .A2(n10122), .ZN(n13971) );
  NAND2_X1 U17245 ( .A1(n15919), .A2(n14109), .ZN(n13972) );
  NAND2_X1 U17246 ( .A1(n20099), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n13976) );
  OAI211_X1 U17247 ( .C1(n14518), .C2(n13973), .A(n13972), .B(n13976), .ZN(
        n13974) );
  AOI21_X1 U17248 ( .B1(n14100), .B2(n20045), .A(n13974), .ZN(n13975) );
  OAI21_X1 U17249 ( .B1(n14001), .B2(n19904), .A(n13975), .ZN(P1_U2969) );
  INV_X1 U17250 ( .A(n13976), .ZN(n13999) );
  NAND2_X1 U17251 ( .A1(n20094), .A2(n20095), .ZN(n13977) );
  NAND3_X1 U17252 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16048) );
  NOR3_X1 U17253 ( .A1(n14557), .A2(n16059), .A3(n16048), .ZN(n16026) );
  NAND2_X1 U17254 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16026), .ZN(
        n16023) );
  NOR2_X1 U17255 ( .A1(n11742), .A2(n16023), .ZN(n13979) );
  NOR2_X1 U17256 ( .A1(n20062), .A2(n20069), .ZN(n20055) );
  NAND2_X1 U17257 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20071) );
  INV_X1 U17258 ( .A(n20071), .ZN(n16061) );
  AND3_X1 U17259 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n20055), .A3(
        n16061), .ZN(n16042) );
  NAND2_X1 U17260 ( .A1(n13979), .A2(n16042), .ZN(n15973) );
  INV_X1 U17261 ( .A(n15973), .ZN(n13978) );
  NAND2_X1 U17262 ( .A1(n20081), .A2(n13978), .ZN(n13982) );
  OAI21_X1 U17263 ( .B1(n20095), .B2(n20090), .A(n20082), .ZN(n20051) );
  AND3_X1 U17264 ( .A1(n20051), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        n20055), .ZN(n16022) );
  NAND2_X1 U17265 ( .A1(n16022), .A2(n13979), .ZN(n15972) );
  INV_X1 U17266 ( .A(n15972), .ZN(n13980) );
  NAND2_X1 U17267 ( .A1(n16024), .A2(n13980), .ZN(n13981) );
  NAND2_X1 U17268 ( .A1(n13982), .A2(n13981), .ZN(n16016) );
  AND2_X1 U17269 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n13986) );
  NAND2_X1 U17270 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15991) );
  NOR2_X1 U17271 ( .A1(n15984), .A2(n15991), .ZN(n15976) );
  INV_X1 U17272 ( .A(n15976), .ZN(n13983) );
  NOR2_X1 U17273 ( .A1(n14603), .A2(n14606), .ZN(n13984) );
  NAND3_X1 U17274 ( .A1(n14600), .A2(n9998), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14568) );
  NAND2_X1 U17275 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14604) );
  INV_X1 U17276 ( .A(n14604), .ZN(n13993) );
  NOR2_X1 U17277 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n13994), .ZN(
        n13985) );
  AND2_X1 U17278 ( .A1(n13986), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13987) );
  NAND2_X1 U17279 ( .A1(n15976), .A2(n13987), .ZN(n13988) );
  OAI21_X1 U17280 ( .B1(n15973), .B2(n13988), .A(n20054), .ZN(n13990) );
  OAI21_X1 U17281 ( .B1(n15972), .B2(n13988), .A(n16024), .ZN(n13989) );
  NAND3_X1 U17282 ( .A1(n20052), .A2(n13990), .A3(n13989), .ZN(n15966) );
  NAND2_X1 U17283 ( .A1(n20093), .A2(n20052), .ZN(n16065) );
  OAI21_X1 U17284 ( .B1(n15966), .B2(n14642), .A(n16065), .ZN(n15956) );
  OAI221_X1 U17285 ( .B1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n20093), 
        .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n20093), .A(n15956), .ZN(
        n15947) );
  AOI21_X1 U17286 ( .B1(n16024), .B2(n13967), .A(n15947), .ZN(n14624) );
  OAI21_X1 U17287 ( .B1(n13991), .B2(n16024), .A(n14603), .ZN(n13992) );
  OAI211_X1 U17288 ( .C1(n13994), .C2(n13993), .A(n14624), .B(n13992), .ZN(
        n14616) );
  OR2_X1 U17289 ( .A1(n14616), .A2(n15975), .ZN(n14569) );
  OR3_X1 U17290 ( .A1(n14616), .A2(n13995), .A3(n14606), .ZN(n13996) );
  AOI21_X1 U17291 ( .B1(n14588), .B2(n14569), .A(n14595), .ZN(n14581) );
  OAI211_X1 U17292 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n20093), .A(
        n14581), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14570) );
  INV_X1 U17293 ( .A(n14570), .ZN(n13997) );
  AOI21_X1 U17294 ( .B1(n14568), .B2(n14567), .A(n13997), .ZN(n13998) );
  AOI211_X1 U17295 ( .C1(n14114), .C2(n20076), .A(n13999), .B(n13998), .ZN(
        n14000) );
  OAI21_X1 U17296 ( .B1(n14001), .B2(n20088), .A(n14000), .ZN(P1_U3001) );
  OR2_X1 U17297 ( .A1(n13909), .A2(n14003), .ZN(n14004) );
  NAND2_X1 U17298 ( .A1(n14002), .A2(n14004), .ZN(n15875) );
  INV_X1 U17299 ( .A(n15874), .ZN(n14005) );
  OAI21_X1 U17300 ( .B1(n15875), .B2(n14005), .A(n14002), .ZN(n14386) );
  AND2_X1 U17301 ( .A1(n14386), .A2(n14385), .ZN(n14388) );
  NAND2_X1 U17302 ( .A1(n14006), .A2(n14007), .ZN(n14376) );
  OAI22_X1 U17303 ( .A1(n14554), .A2(n14011), .B1(n14010), .B2(n14460), .ZN(
        n14012) );
  INV_X1 U17304 ( .A(n14012), .ZN(n15915) );
  INV_X1 U17305 ( .A(n14543), .ZN(n14013) );
  AOI21_X1 U17306 ( .B1(n14014), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n14013), .ZN(n15914) );
  NAND2_X1 U17307 ( .A1(n15915), .A2(n15914), .ZN(n15913) );
  NAND2_X1 U17308 ( .A1(n15913), .A2(n14543), .ZN(n14015) );
  XOR2_X1 U17309 ( .A(n14016), .B(n14015), .Z(n16014) );
  NAND2_X1 U17310 ( .A1(n16014), .A2(n20046), .ZN(n14020) );
  INV_X1 U17311 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n14017) );
  OAI22_X1 U17312 ( .A1(n14518), .A2(n14033), .B1(n16045), .B2(n14017), .ZN(
        n14018) );
  AOI21_X1 U17313 ( .B1(n15919), .B2(n14030), .A(n14018), .ZN(n14019) );
  OAI211_X1 U17314 ( .C1(n20115), .C2(n14039), .A(n14020), .B(n14019), .ZN(
        P1_U2986) );
  MUX2_X1 U17315 ( .A(DATAI_13_), .B(BUF1_REG_13__SCAN_IN), .S(n20116), .Z(
        n20019) );
  AOI22_X1 U17316 ( .A1(n15883), .A2(n20019), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n15884), .ZN(n14021) );
  OAI21_X1 U17317 ( .B1(n14039), .B2(n20004), .A(n14021), .ZN(P1_U2891) );
  NAND2_X1 U17318 ( .A1(n14022), .A2(n14023), .ZN(n14024) );
  AND2_X1 U17319 ( .A1(n14380), .A2(n14024), .ZN(n16013) );
  AOI22_X1 U17320 ( .A1(n19995), .A2(n16013), .B1(n14381), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14025) );
  OAI21_X1 U17321 ( .B1(n14039), .B2(n14389), .A(n14025), .ZN(P1_U2859) );
  INV_X1 U17322 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n20772) );
  INV_X1 U17323 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20771) );
  NOR2_X1 U17324 ( .A1(n20772), .A2(n20771), .ZN(n14101) );
  INV_X1 U17325 ( .A(n14101), .ZN(n14027) );
  INV_X1 U17326 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20768) );
  NOR2_X1 U17327 ( .A1(n20768), .A2(n13899), .ZN(n14102) );
  NAND2_X1 U17328 ( .A1(n14102), .A2(n19923), .ZN(n15855) );
  OAI21_X1 U17329 ( .B1(n14102), .B2(n14281), .A(n14028), .ZN(n15872) );
  NOR2_X1 U17330 ( .A1(n19937), .A2(n14101), .ZN(n14029) );
  NOR2_X1 U17331 ( .A1(n15872), .A2(n14029), .ZN(n15865) );
  INV_X1 U17332 ( .A(n14030), .ZN(n14032) );
  OAI22_X1 U17333 ( .A1(n14032), .A2(n19983), .B1(n19977), .B2(n14031), .ZN(
        n14035) );
  OAI21_X1 U17334 ( .B1(n19931), .B2(n14033), .A(n19969), .ZN(n14034) );
  AOI211_X1 U17335 ( .C1(n16013), .C2(n19974), .A(n14035), .B(n14034), .ZN(
        n14036) );
  OAI21_X1 U17336 ( .B1(n15865), .B2(n14017), .A(n14036), .ZN(n14037) );
  AOI21_X1 U17337 ( .B1(n14017), .B2(n15844), .A(n14037), .ZN(n14038) );
  OAI21_X1 U17338 ( .B1(n14039), .B2(n19926), .A(n14038), .ZN(P1_U2827) );
  XNOR2_X1 U17339 ( .A(n14040), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15149) );
  INV_X1 U17340 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14044) );
  INV_X1 U17341 ( .A(n14041), .ZN(n14043) );
  AOI21_X1 U17342 ( .B1(n14044), .B2(n14043), .A(n14042), .ZN(n14680) );
  INV_X1 U17343 ( .A(n14680), .ZN(n14054) );
  NAND2_X1 U17344 ( .A1(n14045), .A2(n14046), .ZN(n14047) );
  NAND2_X1 U17345 ( .A1(n9815), .A2(n14047), .ZN(n16133) );
  NOR2_X1 U17346 ( .A1(n18957), .A2(n19831), .ZN(n15140) );
  AOI21_X1 U17347 ( .B1(n16247), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15140), .ZN(n14048) );
  OAI21_X1 U17348 ( .B1(n16133), .B2(n13644), .A(n14048), .ZN(n14049) );
  INV_X1 U17349 ( .A(n14049), .ZN(n14053) );
  INV_X1 U17350 ( .A(n14050), .ZN(n14997) );
  NOR2_X1 U17351 ( .A1(n14997), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15138) );
  NOR3_X1 U17352 ( .A1(n15138), .A2(n15137), .A3(n16265), .ZN(n14051) );
  INV_X1 U17353 ( .A(n14051), .ZN(n14052) );
  OAI211_X1 U17354 ( .C1(n16262), .C2(n14054), .A(n14053), .B(n14052), .ZN(
        n14055) );
  INV_X1 U17355 ( .A(n14055), .ZN(n14056) );
  OAI21_X1 U17356 ( .B1(n15149), .B2(n16263), .A(n14056), .ZN(P2_U2987) );
  NOR2_X1 U17357 ( .A1(n14840), .A2(n13644), .ZN(n14062) );
  NAND2_X1 U17358 ( .A1(n14677), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14058) );
  AOI21_X1 U17359 ( .B1(n16247), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14059), .ZN(n14060) );
  AOI21_X1 U17360 ( .B1(n14064), .B2(n19204), .A(n14063), .ZN(n14065) );
  OAI21_X1 U17361 ( .B1(n14066), .B2(n16263), .A(n14065), .ZN(P2_U2983) );
  NOR3_X1 U17362 ( .A1(n14068), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n14067), .ZN(n14077) );
  NAND2_X1 U17363 ( .A1(n14069), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14072) );
  AOI21_X1 U17364 ( .B1(n14717), .B2(n19220), .A(n14073), .ZN(n14075) );
  NAND2_X1 U17365 ( .A1(n14712), .A2(n19228), .ZN(n14074) );
  OAI21_X1 U17366 ( .B1(n14080), .B2(n19225), .A(n14079), .ZN(P2_U3016) );
  INV_X1 U17367 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n20176) );
  NOR2_X1 U17368 ( .A1(n14088), .A2(n20114), .ZN(n14081) );
  NAND2_X1 U17369 ( .A1(n20001), .A2(n14081), .ZN(n14410) );
  AOI22_X1 U17370 ( .A1(n14084), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n14083), .ZN(n14085) );
  INV_X1 U17371 ( .A(n14085), .ZN(n14086) );
  XNOR2_X2 U17372 ( .A(n9797), .B(n14086), .ZN(n14178) );
  NAND3_X1 U17373 ( .A1(n14178), .A2(n14087), .A3(n20001), .ZN(n14091) );
  NOR3_X1 U17374 ( .A1(n15884), .A2(n20116), .A3(n14088), .ZN(n14089) );
  AOI22_X1 U17375 ( .A1(n14441), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15884), .ZN(n14090) );
  OAI211_X1 U17376 ( .C1(n20176), .C2(n14410), .A(n14091), .B(n14090), .ZN(
        P1_U2873) );
  XNOR2_X1 U17377 ( .A(n14095), .B(n14094), .ZN(n14576) );
  NAND2_X1 U17378 ( .A1(n20099), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n14571) );
  NAND2_X1 U17379 ( .A1(n20039), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14096) );
  OAI211_X1 U17380 ( .C1(n20050), .C2(n14097), .A(n14571), .B(n14096), .ZN(
        n14098) );
  OAI21_X1 U17381 ( .B1(n14576), .B2(n19904), .A(n14099), .ZN(P1_U2968) );
  INV_X1 U17382 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20791) );
  INV_X1 U17383 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20788) );
  NAND4_X1 U17384 ( .A1(n14102), .A2(n14101), .A3(P1_REIP_REG_14__SCAN_IN), 
        .A4(P1_REIP_REG_13__SCAN_IN), .ZN(n14278) );
  INV_X1 U17385 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20780) );
  NAND2_X1 U17386 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n15830) );
  NOR2_X1 U17387 ( .A1(n20780), .A2(n15830), .ZN(n15813) );
  NAND2_X1 U17388 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n15813), .ZN(n15799) );
  NAND3_X1 U17389 ( .A1(n14103), .A2(P1_REIP_REG_20__SCAN_IN), .A3(
        P1_REIP_REG_19__SCAN_IN), .ZN(n14104) );
  NOR3_X1 U17390 ( .A1(n14278), .A2(n15799), .A3(n14104), .ZN(n15787) );
  NAND2_X1 U17391 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n15787), .ZN(n15778) );
  NOR2_X1 U17392 ( .A1(n20788), .A2(n15778), .ZN(n14267) );
  NAND2_X1 U17393 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n14267), .ZN(n14241) );
  NOR2_X1 U17394 ( .A1(n20791), .A2(n14241), .ZN(n14244) );
  AND2_X1 U17395 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n14244), .ZN(n14105) );
  NAND2_X1 U17396 ( .A1(n19964), .A2(n14105), .ZN(n14227) );
  INV_X1 U17397 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20797) );
  INV_X1 U17398 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20795) );
  NOR3_X1 U17399 ( .A1(n14227), .A2(n20797), .A3(n20795), .ZN(n14202) );
  NAND2_X1 U17400 ( .A1(n14202), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14194) );
  INV_X1 U17401 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20799) );
  NOR2_X1 U17402 ( .A1(n14194), .A2(n20799), .ZN(n14108) );
  AND2_X1 U17403 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n14107) );
  INV_X1 U17404 ( .A(n14281), .ZN(n14309) );
  NAND2_X1 U17405 ( .A1(n15776), .A2(n14105), .ZN(n14226) );
  NOR2_X1 U17406 ( .A1(n14226), .A2(n20795), .ZN(n14213) );
  NAND3_X1 U17407 ( .A1(n14213), .A2(P1_REIP_REG_27__SCAN_IN), .A3(
        P1_REIP_REG_28__SCAN_IN), .ZN(n14106) );
  NAND2_X1 U17408 ( .A1(n14309), .A2(n14106), .ZN(n14200) );
  OAI21_X1 U17409 ( .B1(n14281), .B2(n14107), .A(n14200), .ZN(n14183) );
  OAI21_X1 U17410 ( .B1(n14108), .B2(P1_REIP_REG_30__SCAN_IN), .A(n14183), 
        .ZN(n14111) );
  AOI22_X1 U17411 ( .A1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19960), .B1(
        n15861), .B2(n14109), .ZN(n14110) );
  OAI211_X1 U17412 ( .C1(n19977), .C2(n14112), .A(n14111), .B(n14110), .ZN(
        n14113) );
  AOI21_X1 U17413 ( .B1(n14114), .B2(n19974), .A(n14113), .ZN(n14115) );
  OAI21_X1 U17414 ( .B1(n14118), .B2(n19926), .A(n14115), .ZN(P1_U2810) );
  AOI22_X1 U17415 ( .A1(n14438), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n15884), .ZN(n14117) );
  MUX2_X1 U17416 ( .A(DATAI_14_), .B(BUF1_REG_14__SCAN_IN), .S(n20116), .Z(
        n20021) );
  AOI22_X1 U17417 ( .A1(n14441), .A2(DATAI_30_), .B1(n14440), .B2(n20021), 
        .ZN(n14116) );
  OAI211_X1 U17418 ( .C1(n14118), .C2(n20004), .A(n14117), .B(n14116), .ZN(
        P1_U2874) );
  NOR2_X1 U17419 ( .A1(n16265), .A2(n14119), .ZN(n14120) );
  AOI211_X1 U17420 ( .C1(n14122), .C2(n11305), .A(n14121), .B(n14120), .ZN(
        n14125) );
  OAI21_X1 U17421 ( .B1(n16247), .B2(n14123), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14124) );
  OAI211_X1 U17422 ( .C1(n13644), .C2(n14126), .A(n14125), .B(n14124), .ZN(
        P2_U3014) );
  MUX2_X1 U17423 ( .A(n14128), .B(n14127), .S(n13168), .Z(n14129) );
  OAI21_X1 U17424 ( .B1(n19113), .B2(n14911), .A(n14129), .ZN(P2_U2883) );
  AOI21_X1 U17425 ( .B1(n19211), .B2(n14131), .A(n14130), .ZN(n19202) );
  INV_X1 U17426 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n18894) );
  AOI22_X1 U17427 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18894), .ZN(n19072) );
  AOI22_X1 U17428 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n14833), .B2(n18894), .ZN(
        n14830) );
  NAND2_X1 U17429 ( .A1(n19072), .A2(n14830), .ZN(n14829) );
  NOR2_X1 U17430 ( .A1(n14820), .A2(n14829), .ZN(n14156) );
  NAND2_X1 U17431 ( .A1(n14156), .A2(n14157), .ZN(n14689) );
  AND2_X1 U17432 ( .A1(n19032), .A2(n14689), .ZN(n14134) );
  NOR4_X1 U17433 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .A4(n10329), .ZN(n18939) );
  AOI21_X1 U17434 ( .B1(n19202), .B2(n14134), .A(n19771), .ZN(n14133) );
  OAI21_X1 U17435 ( .B1(n19202), .B2(n14134), .A(n14133), .ZN(n14154) );
  NAND2_X1 U17436 ( .A1(n19420), .A2(n19765), .ZN(n14142) );
  INV_X1 U17437 ( .A(n14142), .ZN(n14135) );
  NAND2_X1 U17438 ( .A1(n10257), .A2(n14135), .ZN(n14136) );
  NOR2_X2 U17439 ( .A1(n14137), .A2(n14136), .ZN(n19066) );
  NOR3_X1 U17440 ( .A1(n18894), .A2(n19680), .A3(n14670), .ZN(n16359) );
  NAND2_X1 U17441 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n14142), .ZN(n14138) );
  NOR2_X1 U17442 ( .A1(n10279), .A2(n14138), .ZN(n14139) );
  INV_X1 U17443 ( .A(n15359), .ZN(n14140) );
  NOR2_X1 U17444 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n14140), .ZN(n16365) );
  INV_X1 U17445 ( .A(n16365), .ZN(n14145) );
  INV_X1 U17446 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n14141) );
  NAND3_X1 U17447 ( .A1(n14143), .A2(n14142), .A3(n14141), .ZN(n14144) );
  NAND2_X1 U17448 ( .A1(n19136), .A2(n14144), .ZN(n14146) );
  AOI22_X1 U17449 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19024), .B1(
        P2_EBX_REG_4__SCAN_IN), .B2(n19054), .ZN(n14147) );
  OAI211_X1 U17450 ( .C1(n19063), .C2(n14148), .A(n14147), .B(n18957), .ZN(
        n14149) );
  AOI21_X1 U17451 ( .B1(n14150), .B2(n19060), .A(n14149), .ZN(n14151) );
  OAI21_X1 U17452 ( .B1(n9807), .B2(n19799), .A(n14151), .ZN(n14152) );
  AOI21_X1 U17453 ( .B1(n19066), .B2(n19206), .A(n14152), .ZN(n14153) );
  OAI211_X1 U17454 ( .C1(n19068), .C2(n19113), .A(n14154), .B(n14153), .ZN(
        P2_U2851) );
  MUX2_X1 U17455 ( .A(n13617), .B(n10552), .S(n14909), .Z(n14155) );
  OAI21_X1 U17456 ( .B1(n19854), .B2(n14911), .A(n14155), .ZN(P2_U2884) );
  NOR2_X1 U17457 ( .A1(n14704), .A2(n14156), .ZN(n14158) );
  XNOR2_X1 U17458 ( .A(n14158), .B(n14157), .ZN(n14159) );
  NAND2_X1 U17459 ( .A1(n14159), .A2(n18939), .ZN(n14167) );
  OAI22_X1 U17460 ( .A1(n19797), .A2(n9807), .B1(n10552), .B2(n19028), .ZN(
        n14161) );
  AOI21_X1 U17461 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n19024), .A(
        n14161), .ZN(n14162) );
  OAI21_X1 U17462 ( .B1(n19042), .B2(n14163), .A(n14162), .ZN(n14165) );
  NOR2_X1 U17463 ( .A1(n19119), .A2(n19063), .ZN(n14164) );
  AOI211_X1 U17464 ( .C1(n19066), .C2(n10351), .A(n14165), .B(n14164), .ZN(
        n14166) );
  OAI211_X1 U17465 ( .C1(n19068), .C2(n19854), .A(n14167), .B(n14166), .ZN(
        P2_U2852) );
  NOR2_X1 U17466 ( .A1(n14168), .A2(n13168), .ZN(n14169) );
  AOI21_X1 U17467 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n14909), .A(n14169), .ZN(
        n14170) );
  OAI21_X1 U17468 ( .B1(n14171), .B2(n14911), .A(n14170), .ZN(P2_U2857) );
  AOI22_X1 U17469 ( .A1(n14176), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n14175), .ZN(n14177) );
  NAND2_X1 U17470 ( .A1(n14178), .A2(n19949), .ZN(n14185) );
  INV_X1 U17471 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14315) );
  OAI22_X1 U17472 ( .A1(n14179), .A2(n19931), .B1(n19977), .B2(n14315), .ZN(
        n14182) );
  INV_X1 U17473 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14180) );
  NOR4_X1 U17474 ( .A1(n14194), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14180), 
        .A4(n20799), .ZN(n14181) );
  AOI211_X1 U17475 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n14183), .A(n14182), 
        .B(n14181), .ZN(n14184) );
  OAI211_X1 U17476 ( .C1(n14566), .C2(n19945), .A(n14185), .B(n14184), .ZN(
        P1_U2809) );
  AOI21_X1 U17477 ( .B1(n14187), .B2(n12313), .A(n14186), .ZN(n14456) );
  INV_X1 U17478 ( .A(n14456), .ZN(n14393) );
  AOI21_X1 U17479 ( .B1(n14189), .B2(n14199), .A(n14188), .ZN(n14583) );
  OAI22_X1 U17480 ( .A1(n14190), .A2(n19931), .B1(n19983), .B2(n14454), .ZN(
        n14192) );
  NOR2_X1 U17481 ( .A1(n14200), .A2(n20799), .ZN(n14191) );
  AOI211_X1 U17482 ( .C1(P1_EBX_REG_29__SCAN_IN), .C2(n19942), .A(n14192), .B(
        n14191), .ZN(n14193) );
  OAI21_X1 U17483 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(n14194), .A(n14193), 
        .ZN(n14195) );
  AOI21_X1 U17484 ( .B1(n14583), .B2(n19974), .A(n14195), .ZN(n14196) );
  OAI21_X1 U17485 ( .B1(n14393), .B2(n19926), .A(n14196), .ZN(P1_U2811) );
  OR2_X1 U17486 ( .A1(n14208), .A2(n14197), .ZN(n14198) );
  INV_X1 U17487 ( .A(n14200), .ZN(n14201) );
  OAI21_X1 U17488 ( .B1(n14202), .B2(P1_REIP_REG_28__SCAN_IN), .A(n14201), 
        .ZN(n14205) );
  AOI22_X1 U17489 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19960), .B1(
        n15861), .B2(n14203), .ZN(n14204) );
  OAI211_X1 U17490 ( .C1(n19977), .C2(n14318), .A(n14205), .B(n14204), .ZN(
        n14206) );
  AOI21_X1 U17491 ( .B1(n14589), .B2(n19974), .A(n14206), .ZN(n14207) );
  OAI21_X1 U17492 ( .B1(n14396), .B2(n19926), .A(n14207), .ZN(P1_U2812) );
  INV_X1 U17493 ( .A(n14208), .ZN(n14209) );
  OAI21_X1 U17494 ( .B1(n14210), .B2(n14224), .A(n14209), .ZN(n14597) );
  AOI21_X1 U17495 ( .B1(n14212), .B2(n14211), .A(n12277), .ZN(n14466) );
  NAND2_X1 U17496 ( .A1(n14466), .A2(n19949), .ZN(n14220) );
  NOR3_X1 U17497 ( .A1(n14227), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n20795), 
        .ZN(n14218) );
  NOR3_X1 U17498 ( .A1(n14281), .A2(n14213), .A3(n20797), .ZN(n14217) );
  NOR2_X1 U17499 ( .A1(n19977), .A2(n14319), .ZN(n14216) );
  OAI22_X1 U17500 ( .A1(n14214), .A2(n19931), .B1(n19983), .B2(n14464), .ZN(
        n14215) );
  NOR4_X1 U17501 ( .A1(n14218), .A2(n14217), .A3(n14216), .A4(n14215), .ZN(
        n14219) );
  OAI211_X1 U17502 ( .C1(n19945), .C2(n14597), .A(n14220), .B(n14219), .ZN(
        P1_U2813) );
  OAI21_X1 U17503 ( .B1(n14221), .B2(n14222), .A(n14211), .ZN(n14472) );
  AND2_X1 U17504 ( .A1(n14238), .A2(n14223), .ZN(n14225) );
  OR2_X1 U17505 ( .A1(n14225), .A2(n14224), .ZN(n14609) );
  INV_X1 U17506 ( .A(n14609), .ZN(n14233) );
  NAND3_X1 U17507 ( .A1(n14309), .A2(P1_REIP_REG_26__SCAN_IN), .A3(n14226), 
        .ZN(n14231) );
  OR2_X1 U17508 ( .A1(n14227), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14230) );
  AOI22_X1 U17509 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19960), .B1(
        n15861), .B2(n14475), .ZN(n14229) );
  NAND2_X1 U17510 ( .A1(n19942), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n14228) );
  NAND4_X1 U17511 ( .A1(n14231), .A2(n14230), .A3(n14229), .A4(n14228), .ZN(
        n14232) );
  AOI21_X1 U17512 ( .B1(n14233), .B2(n19974), .A(n14232), .ZN(n14234) );
  OAI21_X1 U17513 ( .B1(n14472), .B2(n19926), .A(n14234), .ZN(P1_U2814) );
  NAND2_X1 U17514 ( .A1(n14235), .A2(n14236), .ZN(n14237) );
  NAND2_X1 U17515 ( .A1(n14238), .A2(n14237), .ZN(n14619) );
  AOI21_X1 U17516 ( .B1(n14240), .B2(n14239), .A(n14221), .ZN(n14485) );
  NAND2_X1 U17517 ( .A1(n14485), .A2(n19949), .ZN(n14251) );
  INV_X1 U17518 ( .A(n14241), .ZN(n14253) );
  AND2_X1 U17519 ( .A1(n15776), .A2(n14253), .ZN(n14242) );
  NOR2_X1 U17520 ( .A1(n14281), .A2(n14242), .ZN(n14266) );
  NAND2_X1 U17521 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n14243) );
  OAI21_X1 U17522 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(n14244), .A(n14243), 
        .ZN(n14248) );
  NAND2_X1 U17523 ( .A1(n19942), .A2(P1_EBX_REG_25__SCAN_IN), .ZN(n14247) );
  INV_X1 U17524 ( .A(n14483), .ZN(n14245) );
  AOI22_X1 U17525 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19960), .B1(
        n15861), .B2(n14245), .ZN(n14246) );
  OAI211_X1 U17526 ( .C1(n14248), .C2(n19937), .A(n14247), .B(n14246), .ZN(
        n14249) );
  AOI21_X1 U17527 ( .B1(n14266), .B2(P1_REIP_REG_25__SCAN_IN), .A(n14249), 
        .ZN(n14250) );
  OAI211_X1 U17528 ( .C1(n19945), .C2(n14619), .A(n14251), .B(n14250), .ZN(
        P1_U2815) );
  OAI21_X1 U17529 ( .B1(n14263), .B2(n14252), .A(n14239), .ZN(n14492) );
  NAND3_X1 U17530 ( .A1(n19964), .A2(n20791), .A3(n14253), .ZN(n14255) );
  AOI22_X1 U17531 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19960), .B1(
        n15861), .B2(n14495), .ZN(n14254) );
  OAI211_X1 U17532 ( .C1(n14322), .C2(n19977), .A(n14255), .B(n14254), .ZN(
        n14258) );
  OAI21_X1 U17533 ( .B1(n14261), .B2(n14256), .A(n14235), .ZN(n14623) );
  NOR2_X1 U17534 ( .A1(n14623), .A2(n19945), .ZN(n14257) );
  AOI211_X1 U17535 ( .C1(n14266), .C2(P1_REIP_REG_24__SCAN_IN), .A(n14258), 
        .B(n14257), .ZN(n14259) );
  OAI21_X1 U17536 ( .B1(n14492), .B2(n19926), .A(n14259), .ZN(P1_U2816) );
  AND2_X1 U17537 ( .A1(n14327), .A2(n14260), .ZN(n14262) );
  OR2_X1 U17538 ( .A1(n14262), .A2(n14261), .ZN(n15953) );
  AOI21_X1 U17539 ( .B1(n14264), .B2(n14331), .A(n14263), .ZN(n14501) );
  NAND2_X1 U17540 ( .A1(n14501), .A2(n19949), .ZN(n14273) );
  OAI22_X1 U17541 ( .A1(n14265), .A2(n19931), .B1(n19983), .B2(n14499), .ZN(
        n14271) );
  INV_X1 U17542 ( .A(n14266), .ZN(n14269) );
  AOI21_X1 U17543 ( .B1(n19964), .B2(n14267), .A(P1_REIP_REG_23__SCAN_IN), 
        .ZN(n14268) );
  NOR2_X1 U17544 ( .A1(n14269), .A2(n14268), .ZN(n14270) );
  AOI211_X1 U17545 ( .C1(P1_EBX_REG_23__SCAN_IN), .C2(n19942), .A(n14271), .B(
        n14270), .ZN(n14272) );
  OAI211_X1 U17546 ( .C1(n15953), .C2(n19945), .A(n14273), .B(n14272), .ZN(
        P1_U2817) );
  AND2_X1 U17547 ( .A1(n14006), .A2(n14274), .ZN(n14359) );
  OR2_X1 U17548 ( .A1(n14359), .A2(n14275), .ZN(n14277) );
  NAND2_X1 U17549 ( .A1(n14006), .A2(n14276), .ZN(n14350) );
  NAND3_X1 U17550 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(n15844), .ZN(n15843) );
  OAI21_X1 U17551 ( .B1(n15830), .B2(n15843), .A(n20780), .ZN(n14289) );
  INV_X1 U17552 ( .A(n14278), .ZN(n14279) );
  NOR2_X1 U17553 ( .A1(n14281), .A2(n14279), .ZN(n14280) );
  OR2_X1 U17554 ( .A1(n19924), .A2(n14280), .ZN(n15837) );
  INV_X1 U17555 ( .A(n15837), .ZN(n15854) );
  OAI21_X1 U17556 ( .B1(n15813), .B2(n14281), .A(n15854), .ZN(n15818) );
  NAND2_X1 U17557 ( .A1(n15861), .A2(n15901), .ZN(n14283) );
  NAND2_X1 U17558 ( .A1(n19960), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14282) );
  NAND3_X1 U17559 ( .A1(n14283), .A2(n14282), .A3(n19969), .ZN(n14288) );
  OAI21_X1 U17560 ( .B1(n14284), .B2(n14285), .A(n14353), .ZN(n15983) );
  INV_X1 U17561 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14286) );
  OAI22_X1 U17562 ( .A1(n19945), .A2(n15983), .B1(n14286), .B2(n19977), .ZN(
        n14287) );
  AOI211_X1 U17563 ( .C1(n14289), .C2(n15818), .A(n14288), .B(n14287), .ZN(
        n14290) );
  OAI21_X1 U17564 ( .B1(n14437), .B2(n19926), .A(n14290), .ZN(P1_U2823) );
  NAND3_X1 U17565 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n19923), .A3(n20768), 
        .ZN(n14294) );
  INV_X1 U17566 ( .A(n19969), .ZN(n19947) );
  AOI21_X1 U17567 ( .B1(n19960), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n19947), .ZN(n14291) );
  OAI21_X1 U17568 ( .B1(n19983), .B2(n14561), .A(n14291), .ZN(n14292) );
  AOI21_X1 U17569 ( .B1(n19942), .B2(P1_EBX_REG_10__SCAN_IN), .A(n14292), .ZN(
        n14293) );
  OAI211_X1 U17570 ( .C1(n19945), .C2(n16044), .A(n14294), .B(n14293), .ZN(
        n14295) );
  AOI21_X1 U17571 ( .B1(n15872), .B2(P1_REIP_REG_10__SCAN_IN), .A(n14295), 
        .ZN(n14296) );
  OAI21_X1 U17572 ( .B1(n14297), .B2(n19926), .A(n14296), .ZN(P1_U2830) );
  MUX2_X1 U17573 ( .A(n19983), .B(n19931), .S(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n14305) );
  INV_X1 U17574 ( .A(n14298), .ZN(n14299) );
  AOI22_X1 U17575 ( .A1(n14299), .A2(n19980), .B1(n19964), .B2(n13735), .ZN(
        n14304) );
  INV_X1 U17576 ( .A(n15776), .ZN(n19935) );
  AOI22_X1 U17577 ( .A1(n19962), .A2(n20645), .B1(n19935), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n14303) );
  AOI22_X1 U17578 ( .A1(n19942), .A2(P1_EBX_REG_1__SCAN_IN), .B1(n19974), .B2(
        n14301), .ZN(n14302) );
  NAND4_X1 U17579 ( .A1(n14305), .A2(n14304), .A3(n14303), .A4(n14302), .ZN(
        P1_U2839) );
  OAI22_X1 U17580 ( .A1(n19945), .A2(n14307), .B1(n14306), .B2(n19977), .ZN(
        n14308) );
  AOI21_X1 U17581 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(n14309), .A(n14308), .ZN(
        n14314) );
  INV_X1 U17582 ( .A(n20005), .ZN(n14310) );
  NAND2_X1 U17583 ( .A1(n19980), .A2(n14310), .ZN(n14313) );
  NAND2_X1 U17584 ( .A1(n19962), .A2(n11849), .ZN(n14312) );
  OAI21_X1 U17585 ( .B1(n19960), .B2(n15861), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14311) );
  NAND4_X1 U17586 ( .A1(n14314), .A2(n14313), .A3(n14312), .A4(n14311), .ZN(
        P1_U2840) );
  OAI22_X1 U17587 ( .A1(n14566), .A2(n19986), .B1(n14315), .B2(n20000), .ZN(
        P1_U2841) );
  AOI22_X1 U17588 ( .A1(n14583), .A2(n19995), .B1(n14381), .B2(
        P1_EBX_REG_29__SCAN_IN), .ZN(n14316) );
  OAI21_X1 U17589 ( .B1(n14393), .B2(n14389), .A(n14316), .ZN(P1_U2843) );
  INV_X1 U17590 ( .A(n14589), .ZN(n14317) );
  OAI222_X1 U17591 ( .A1(n14318), .A2(n20000), .B1(n19986), .B2(n14317), .C1(
        n14396), .C2(n14389), .ZN(P1_U2844) );
  INV_X1 U17592 ( .A(n14466), .ZN(n14401) );
  OAI222_X1 U17593 ( .A1(n14319), .A2(n20000), .B1(n19986), .B2(n14597), .C1(
        n14401), .C2(n14389), .ZN(P1_U2845) );
  OAI222_X1 U17594 ( .A1(n14320), .A2(n20000), .B1(n19986), .B2(n14609), .C1(
        n14472), .C2(n14389), .ZN(P1_U2846) );
  INV_X1 U17595 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14321) );
  INV_X1 U17596 ( .A(n14485), .ZN(n14406) );
  OAI222_X1 U17597 ( .A1(n14321), .A2(n20000), .B1(n19986), .B2(n14619), .C1(
        n14406), .C2(n14389), .ZN(P1_U2847) );
  OAI222_X1 U17598 ( .A1(n14322), .A2(n20000), .B1(n19986), .B2(n14623), .C1(
        n14492), .C2(n14389), .ZN(P1_U2848) );
  INV_X1 U17599 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14323) );
  INV_X1 U17600 ( .A(n14501), .ZN(n14415) );
  OAI222_X1 U17601 ( .A1(n15953), .A2(n19986), .B1(n14323), .B2(n20000), .C1(
        n14389), .C2(n14415), .ZN(P1_U2849) );
  NAND2_X1 U17602 ( .A1(n14324), .A2(n14325), .ZN(n14326) );
  NAND2_X1 U17603 ( .A1(n14327), .A2(n14326), .ZN(n15962) );
  INV_X1 U17604 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n20858) );
  NAND2_X1 U17605 ( .A1(n14328), .A2(n14329), .ZN(n14330) );
  OAI222_X1 U17606 ( .A1(n15962), .A2(n19986), .B1(n20000), .B2(n20858), .C1(
        n14389), .C2(n14509), .ZN(P1_U2850) );
  INV_X1 U17607 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14337) );
  NAND2_X1 U17608 ( .A1(n14340), .A2(n14332), .ZN(n14333) );
  NAND2_X1 U17609 ( .A1(n14324), .A2(n14333), .ZN(n15792) );
  OR2_X1 U17610 ( .A1(n14334), .A2(n14335), .ZN(n14336) );
  OAI222_X1 U17611 ( .A1(n14337), .A2(n20000), .B1(n19986), .B2(n15792), .C1(
        n14422), .C2(n14389), .ZN(P1_U2851) );
  OR2_X1 U17612 ( .A1(n14347), .A2(n14338), .ZN(n14339) );
  NAND2_X1 U17613 ( .A1(n14340), .A2(n14339), .ZN(n15800) );
  INV_X1 U17614 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14344) );
  INV_X1 U17615 ( .A(n14334), .ZN(n14342) );
  OAI21_X1 U17616 ( .B1(n14343), .B2(n14341), .A(n14342), .ZN(n15801) );
  OAI222_X1 U17617 ( .A1(n15800), .A2(n19986), .B1(n20000), .B2(n14344), .C1(
        n14389), .C2(n15801), .ZN(P1_U2852) );
  AOI21_X1 U17618 ( .B1(n14346), .B2(n14345), .A(n14341), .ZN(n15889) );
  INV_X1 U17619 ( .A(n15889), .ZN(n14429) );
  AOI21_X1 U17620 ( .B1(n14348), .B2(n14355), .A(n14347), .ZN(n15964) );
  AOI22_X1 U17621 ( .A1(n15964), .A2(n19995), .B1(n14381), .B2(
        P1_EBX_REG_19__SCAN_IN), .ZN(n14349) );
  OAI21_X1 U17622 ( .B1(n14429), .B2(n14389), .A(n14349), .ZN(P1_U2853) );
  XOR2_X1 U17623 ( .A(n14351), .B(n14350), .Z(n15825) );
  INV_X1 U17624 ( .A(n15825), .ZN(n14433) );
  NAND2_X1 U17625 ( .A1(n14353), .A2(n14352), .ZN(n14354) );
  NAND2_X1 U17626 ( .A1(n14355), .A2(n14354), .ZN(n15977) );
  OAI22_X1 U17627 ( .A1(n15977), .A2(n19986), .B1(n15821), .B2(n20000), .ZN(
        n14356) );
  INV_X1 U17628 ( .A(n14356), .ZN(n14357) );
  OAI21_X1 U17629 ( .B1(n14433), .B2(n14389), .A(n14357), .ZN(P1_U2854) );
  OAI222_X1 U17630 ( .A1(n14437), .A2(n14389), .B1(n20000), .B2(n14286), .C1(
        n19986), .C2(n15983), .ZN(P1_U2855) );
  NAND2_X1 U17631 ( .A1(n14006), .A2(n14358), .ZN(n14367) );
  AOI21_X1 U17632 ( .B1(n14360), .B2(n14367), .A(n14359), .ZN(n14540) );
  INV_X1 U17633 ( .A(n14540), .ZN(n15832) );
  NOR2_X1 U17634 ( .A1(n14372), .A2(n14361), .ZN(n14362) );
  OR2_X1 U17635 ( .A1(n14284), .A2(n14362), .ZN(n15994) );
  OAI22_X1 U17636 ( .A1(n15994), .A2(n19986), .B1(n14363), .B2(n20000), .ZN(
        n14364) );
  INV_X1 U17637 ( .A(n14364), .ZN(n14365) );
  OAI21_X1 U17638 ( .B1(n15832), .B2(n14389), .A(n14365), .ZN(P1_U2856) );
  NAND2_X1 U17639 ( .A1(n14006), .A2(n14366), .ZN(n14378) );
  INV_X1 U17640 ( .A(n14367), .ZN(n14368) );
  AOI21_X1 U17641 ( .B1(n14369), .B2(n14378), .A(n14368), .ZN(n15910) );
  INV_X1 U17642 ( .A(n15910), .ZN(n14446) );
  INV_X1 U17643 ( .A(n14380), .ZN(n14371) );
  AOI21_X1 U17644 ( .B1(n14371), .B2(n14379), .A(n14370), .ZN(n14373) );
  NOR2_X1 U17645 ( .A1(n14373), .A2(n14372), .ZN(n16003) );
  AOI22_X1 U17646 ( .A1(n16003), .A2(n19995), .B1(n14381), .B2(
        P1_EBX_REG_15__SCAN_IN), .ZN(n14374) );
  OAI21_X1 U17647 ( .B1(n14446), .B2(n14389), .A(n14374), .ZN(P1_U2857) );
  NAND2_X1 U17648 ( .A1(n14376), .A2(n14375), .ZN(n14377) );
  XNOR2_X1 U17649 ( .A(n14380), .B(n14379), .ZN(n16007) );
  AOI22_X1 U17650 ( .A1(n19995), .A2(n16007), .B1(n14381), .B2(
        P1_EBX_REG_14__SCAN_IN), .ZN(n14382) );
  OAI21_X1 U17651 ( .B1(n14448), .B2(n14389), .A(n14382), .ZN(P1_U2858) );
  OR2_X1 U17652 ( .A1(n15866), .A2(n14383), .ZN(n14384) );
  NAND2_X1 U17653 ( .A1(n14022), .A2(n14384), .ZN(n16029) );
  INV_X1 U17654 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n21094) );
  NOR2_X1 U17655 ( .A1(n14386), .A2(n14385), .ZN(n14387) );
  OAI222_X1 U17656 ( .A1(n16029), .A2(n19986), .B1(n20000), .B2(n21094), .C1(
        n14389), .C2(n15881), .ZN(P1_U2860) );
  INV_X1 U17657 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n19264) );
  OAI22_X1 U17658 ( .A1(n14410), .A2(n19264), .B1(n13500), .B2(n20001), .ZN(
        n14390) );
  INV_X1 U17659 ( .A(n14390), .ZN(n14392) );
  AOI22_X1 U17660 ( .A1(n14441), .A2(DATAI_29_), .B1(n14440), .B2(n20019), 
        .ZN(n14391) );
  OAI211_X1 U17661 ( .C1(n14393), .C2(n20004), .A(n14392), .B(n14391), .ZN(
        P1_U2875) );
  AOI22_X1 U17662 ( .A1(n14438), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n15884), .ZN(n14395) );
  MUX2_X1 U17663 ( .A(DATAI_12_), .B(BUF1_REG_12__SCAN_IN), .S(n20116), .Z(
        n20017) );
  AOI22_X1 U17664 ( .A1(n14441), .A2(DATAI_28_), .B1(n14440), .B2(n20017), 
        .ZN(n14394) );
  OAI211_X1 U17665 ( .C1(n14396), .C2(n20004), .A(n14395), .B(n14394), .ZN(
        P1_U2876) );
  INV_X1 U17666 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n21078) );
  OAI22_X1 U17667 ( .A1(n14410), .A2(n21078), .B1(n14397), .B2(n20001), .ZN(
        n14398) );
  INV_X1 U17668 ( .A(n14398), .ZN(n14400) );
  AOI22_X1 U17669 ( .A1(n14441), .A2(DATAI_27_), .B1(n14440), .B2(n15882), 
        .ZN(n14399) );
  OAI211_X1 U17670 ( .C1(n14401), .C2(n20004), .A(n14400), .B(n14399), .ZN(
        P1_U2877) );
  AOI22_X1 U17671 ( .A1(n14438), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n15884), .ZN(n14403) );
  AOI22_X1 U17672 ( .A1(n14441), .A2(DATAI_26_), .B1(n14440), .B2(n20015), 
        .ZN(n14402) );
  OAI211_X1 U17673 ( .C1(n14472), .C2(n20004), .A(n14403), .B(n14402), .ZN(
        P1_U2878) );
  AOI22_X1 U17674 ( .A1(n14438), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n15884), .ZN(n14405) );
  AOI22_X1 U17675 ( .A1(n14441), .A2(DATAI_25_), .B1(n14440), .B2(n20013), 
        .ZN(n14404) );
  OAI211_X1 U17676 ( .C1(n14406), .C2(n20004), .A(n14405), .B(n14404), .ZN(
        P1_U2879) );
  AOI22_X1 U17677 ( .A1(n14438), .A2(BUF1_REG_24__SCAN_IN), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(n15884), .ZN(n14408) );
  AOI22_X1 U17678 ( .A1(n14441), .A2(DATAI_24_), .B1(n14440), .B2(n20011), 
        .ZN(n14407) );
  OAI211_X1 U17679 ( .C1(n14492), .C2(n20004), .A(n14408), .B(n14407), .ZN(
        P1_U2880) );
  INV_X1 U17680 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16478) );
  OAI22_X1 U17681 ( .A1(n14410), .A2(n16478), .B1(n14409), .B2(n20001), .ZN(
        n14411) );
  INV_X1 U17682 ( .A(n14411), .ZN(n14414) );
  AOI22_X1 U17683 ( .A1(n14441), .A2(DATAI_23_), .B1(n14440), .B2(n14412), 
        .ZN(n14413) );
  OAI211_X1 U17684 ( .C1(n14415), .C2(n20004), .A(n14414), .B(n14413), .ZN(
        P1_U2881) );
  AOI22_X1 U17685 ( .A1(n14438), .A2(BUF1_REG_22__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n15884), .ZN(n14418) );
  AOI22_X1 U17686 ( .A1(n14441), .A2(DATAI_22_), .B1(n14440), .B2(n14416), 
        .ZN(n14417) );
  OAI211_X1 U17687 ( .C1(n14509), .C2(n20004), .A(n14418), .B(n14417), .ZN(
        P1_U2882) );
  AOI22_X1 U17688 ( .A1(n14438), .A2(BUF1_REG_21__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n15884), .ZN(n14421) );
  AOI22_X1 U17689 ( .A1(n14441), .A2(DATAI_21_), .B1(n14440), .B2(n14419), 
        .ZN(n14420) );
  OAI211_X1 U17690 ( .C1(n14422), .C2(n20004), .A(n14421), .B(n14420), .ZN(
        P1_U2883) );
  AOI22_X1 U17691 ( .A1(n14438), .A2(BUF1_REG_20__SCAN_IN), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(n15884), .ZN(n14425) );
  AOI22_X1 U17692 ( .A1(n14441), .A2(DATAI_20_), .B1(n14440), .B2(n14423), 
        .ZN(n14424) );
  OAI211_X1 U17693 ( .C1(n15801), .C2(n20004), .A(n14425), .B(n14424), .ZN(
        P1_U2884) );
  AOI22_X1 U17694 ( .A1(n14438), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n15884), .ZN(n14428) );
  AOI22_X1 U17695 ( .A1(n14441), .A2(DATAI_19_), .B1(n14440), .B2(n14426), 
        .ZN(n14427) );
  OAI211_X1 U17696 ( .C1(n14429), .C2(n20004), .A(n14428), .B(n14427), .ZN(
        P1_U2885) );
  AOI22_X1 U17697 ( .A1(n14438), .A2(BUF1_REG_18__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n15884), .ZN(n14432) );
  AOI22_X1 U17698 ( .A1(n14441), .A2(DATAI_18_), .B1(n14440), .B2(n14430), 
        .ZN(n14431) );
  OAI211_X1 U17699 ( .C1(n14433), .C2(n20004), .A(n14432), .B(n14431), .ZN(
        P1_U2886) );
  AOI22_X1 U17700 ( .A1(n14438), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n15884), .ZN(n14436) );
  AOI22_X1 U17701 ( .A1(n14441), .A2(DATAI_17_), .B1(n14440), .B2(n14434), 
        .ZN(n14435) );
  OAI211_X1 U17702 ( .C1(n14437), .C2(n20004), .A(n14436), .B(n14435), .ZN(
        P1_U2887) );
  AOI22_X1 U17703 ( .A1(n14438), .A2(BUF1_REG_16__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n15884), .ZN(n14443) );
  AOI22_X1 U17704 ( .A1(n14441), .A2(DATAI_16_), .B1(n14440), .B2(n14439), 
        .ZN(n14442) );
  OAI211_X1 U17705 ( .C1(n15832), .C2(n20004), .A(n14443), .B(n14442), .ZN(
        P1_U2888) );
  OAI222_X1 U17706 ( .A1(n14446), .A2(n20004), .B1(n20003), .B2(n14445), .C1(
        n20001), .C2(n14444), .ZN(P1_U2889) );
  AOI22_X1 U17707 ( .A1(n15883), .A2(n20021), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n15884), .ZN(n14447) );
  OAI21_X1 U17708 ( .B1(n14448), .B2(n20004), .A(n14447), .ZN(P1_U2890) );
  NAND2_X1 U17709 ( .A1(n14450), .A2(n14449), .ZN(n14452) );
  XOR2_X1 U17710 ( .A(n14452), .B(n14451), .Z(n14585) );
  NOR2_X1 U17711 ( .A1(n16045), .A2(n20799), .ZN(n14577) );
  AOI21_X1 U17712 ( .B1(n20039), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14577), .ZN(n14453) );
  OAI21_X1 U17713 ( .B1(n20050), .B2(n14454), .A(n14453), .ZN(n14455) );
  AOI21_X1 U17714 ( .B1(n14456), .B2(n20045), .A(n14455), .ZN(n14457) );
  OAI21_X1 U17715 ( .B1(n19904), .B2(n14585), .A(n14457), .ZN(P1_U2970) );
  INV_X1 U17716 ( .A(n13965), .ZN(n14458) );
  AND2_X1 U17717 ( .A1(n14459), .A2(n14458), .ZN(n14461) );
  MUX2_X1 U17718 ( .A(n14461), .B(n14092), .S(n15893), .Z(n14462) );
  XNOR2_X1 U17719 ( .A(n14462), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14602) );
  NOR2_X1 U17720 ( .A1(n16045), .A2(n20797), .ZN(n14594) );
  AOI21_X1 U17721 ( .B1(n20039), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n14594), .ZN(n14463) );
  OAI21_X1 U17722 ( .B1(n20050), .B2(n14464), .A(n14463), .ZN(n14465) );
  AOI21_X1 U17723 ( .B1(n14466), .B2(n20045), .A(n14465), .ZN(n14467) );
  OAI21_X1 U17724 ( .B1(n19904), .B2(n14602), .A(n14467), .ZN(P1_U2972) );
  OAI21_X1 U17725 ( .B1(n14487), .B2(n14603), .A(n14460), .ZN(n14468) );
  NAND2_X1 U17726 ( .A1(n14469), .A2(n14468), .ZN(n14470) );
  XNOR2_X1 U17727 ( .A(n14470), .B(n14606), .ZN(n14614) );
  NAND2_X1 U17728 ( .A1(n20099), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14608) );
  OAI21_X1 U17729 ( .B1(n14518), .B2(n14471), .A(n14608), .ZN(n14474) );
  NOR2_X1 U17730 ( .A1(n14472), .A2(n20115), .ZN(n14473) );
  AOI211_X1 U17731 ( .C1(n15919), .C2(n14475), .A(n14474), .B(n14473), .ZN(
        n14476) );
  OAI21_X1 U17732 ( .B1(n19904), .B2(n14614), .A(n14476), .ZN(P1_U2973) );
  MUX2_X1 U17733 ( .A(n21048), .B(n14477), .S(n15893), .Z(n14480) );
  NAND2_X1 U17734 ( .A1(n14478), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14489) );
  AND2_X1 U17735 ( .A1(n14489), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14479) );
  NOR2_X1 U17736 ( .A1(n14480), .A2(n14479), .ZN(n14481) );
  XNOR2_X1 U17737 ( .A(n14481), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14622) );
  INV_X1 U17738 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20793) );
  NOR2_X1 U17739 ( .A1(n16045), .A2(n20793), .ZN(n14615) );
  AOI21_X1 U17740 ( .B1(n20039), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n14615), .ZN(n14482) );
  OAI21_X1 U17741 ( .B1(n20050), .B2(n14483), .A(n14482), .ZN(n14484) );
  AOI21_X1 U17742 ( .B1(n14485), .B2(n20045), .A(n14484), .ZN(n14486) );
  OAI21_X1 U17743 ( .B1(n19904), .B2(n14622), .A(n14486), .ZN(P1_U2974) );
  NAND2_X1 U17744 ( .A1(n14487), .A2(n14489), .ZN(n14488) );
  MUX2_X1 U17745 ( .A(n14489), .B(n14488), .S(n15893), .Z(n14490) );
  XNOR2_X1 U17746 ( .A(n14490), .B(n21048), .ZN(n14633) );
  NAND2_X1 U17747 ( .A1(n20099), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14626) );
  OAI21_X1 U17748 ( .B1(n14518), .B2(n14491), .A(n14626), .ZN(n14494) );
  NOR2_X1 U17749 ( .A1(n14492), .A2(n20115), .ZN(n14493) );
  AOI211_X1 U17750 ( .C1(n15919), .C2(n14495), .A(n14494), .B(n14493), .ZN(
        n14496) );
  OAI21_X1 U17751 ( .B1(n19904), .B2(n14633), .A(n14496), .ZN(P1_U2975) );
  XNOR2_X1 U17752 ( .A(n14460), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14497) );
  XNOR2_X1 U17753 ( .A(n13966), .B(n14497), .ZN(n15948) );
  AOI22_X1 U17754 ( .A1(n20039), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B1(
        n20099), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n14498) );
  OAI21_X1 U17755 ( .B1(n20050), .B2(n14499), .A(n14498), .ZN(n14500) );
  AOI21_X1 U17756 ( .B1(n14501), .B2(n20045), .A(n14500), .ZN(n14502) );
  OAI21_X1 U17757 ( .B1(n15948), .B2(n19904), .A(n14502), .ZN(P1_U2976) );
  OAI22_X1 U17758 ( .A1(n14518), .A2(n15779), .B1(n16045), .B2(n20788), .ZN(
        n14503) );
  AOI21_X1 U17759 ( .B1(n15783), .B2(n15919), .A(n14503), .ZN(n14508) );
  NAND2_X1 U17760 ( .A1(n14505), .A2(n14504), .ZN(n14506) );
  XNOR2_X1 U17761 ( .A(n14506), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15958) );
  NAND2_X1 U17762 ( .A1(n15958), .A2(n20046), .ZN(n14507) );
  OAI211_X1 U17763 ( .C1(n14509), .C2(n20115), .A(n14508), .B(n14507), .ZN(
        P1_U2977) );
  INV_X1 U17764 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15967) );
  OR3_X1 U17765 ( .A1(n14510), .A2(n15893), .A3(n15967), .ZN(n14512) );
  OAI21_X1 U17766 ( .B1(n14460), .B2(n14511), .A(n14512), .ZN(n14522) );
  NAND2_X1 U17767 ( .A1(n14522), .A2(n14521), .ZN(n14520) );
  OAI22_X1 U17768 ( .A1(n14520), .A2(n14460), .B1(n14521), .B2(n14512), .ZN(
        n14513) );
  XNOR2_X1 U17769 ( .A(n14513), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14639) );
  INV_X1 U17770 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n14514) );
  OR2_X1 U17771 ( .A1(n16045), .A2(n14514), .ZN(n14634) );
  NAND2_X1 U17772 ( .A1(n20039), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14515) );
  OAI211_X1 U17773 ( .C1(n20050), .C2(n15797), .A(n14634), .B(n14515), .ZN(
        n14516) );
  AOI21_X1 U17774 ( .B1(n15794), .B2(n20045), .A(n14516), .ZN(n14517) );
  OAI21_X1 U17775 ( .B1(n14639), .B2(n19904), .A(n14517), .ZN(P1_U2978) );
  NAND2_X1 U17776 ( .A1(n20099), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n14643) );
  OAI21_X1 U17777 ( .B1(n14518), .B2(n15807), .A(n14643), .ZN(n14519) );
  AOI21_X1 U17778 ( .B1(n15798), .B2(n15919), .A(n14519), .ZN(n14524) );
  OAI21_X1 U17779 ( .B1(n14522), .B2(n14521), .A(n14520), .ZN(n14640) );
  NAND2_X1 U17780 ( .A1(n14640), .A2(n20046), .ZN(n14523) );
  OAI211_X1 U17781 ( .C1(n15801), .C2(n20115), .A(n14524), .B(n14523), .ZN(
        P1_U2979) );
  OAI21_X1 U17782 ( .B1(n14526), .B2(n14525), .A(n14510), .ZN(n15978) );
  INV_X1 U17783 ( .A(n15824), .ZN(n14528) );
  AOI22_X1 U17784 ( .A1(n20039), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n20099), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n14527) );
  OAI21_X1 U17785 ( .B1(n20050), .B2(n14528), .A(n14527), .ZN(n14529) );
  AOI21_X1 U17786 ( .B1(n15825), .B2(n20045), .A(n14529), .ZN(n14530) );
  OAI21_X1 U17787 ( .B1(n19904), .B2(n15978), .A(n14530), .ZN(P1_U2981) );
  OAI21_X1 U17788 ( .B1(n14554), .B2(n14532), .A(n14531), .ZN(n15908) );
  NAND2_X1 U17789 ( .A1(n14533), .A2(n14534), .ZN(n15907) );
  OR2_X1 U17790 ( .A1(n15908), .A2(n15907), .ZN(n15905) );
  NAND2_X1 U17791 ( .A1(n15905), .A2(n14534), .ZN(n14535) );
  XOR2_X1 U17792 ( .A(n14536), .B(n14535), .Z(n15992) );
  INV_X1 U17793 ( .A(n15835), .ZN(n14538) );
  AOI22_X1 U17794 ( .A1(n20039), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n20099), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n14537) );
  OAI21_X1 U17795 ( .B1(n20050), .B2(n14538), .A(n14537), .ZN(n14539) );
  AOI21_X1 U17796 ( .B1(n14540), .B2(n20045), .A(n14539), .ZN(n14541) );
  OAI21_X1 U17797 ( .B1(n15992), .B2(n19904), .A(n14541), .ZN(P1_U2983) );
  NOR2_X1 U17798 ( .A1(n11747), .A2(n14542), .ZN(n15897) );
  NAND2_X1 U17799 ( .A1(n14544), .A2(n14543), .ZN(n14546) );
  OAI21_X1 U17800 ( .B1(n15897), .B2(n14546), .A(n14545), .ZN(n14548) );
  XNOR2_X1 U17801 ( .A(n14460), .B(n16008), .ZN(n14547) );
  XNOR2_X1 U17802 ( .A(n14548), .B(n14547), .ZN(n16006) );
  INV_X1 U17803 ( .A(n16006), .ZN(n14552) );
  AOI22_X1 U17804 ( .A1(n20039), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n20099), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n14549) );
  OAI21_X1 U17805 ( .B1(n20050), .B2(n15848), .A(n14549), .ZN(n14550) );
  AOI21_X1 U17806 ( .B1(n15850), .B2(n20045), .A(n14550), .ZN(n14551) );
  OAI21_X1 U17807 ( .B1(n14552), .B2(n19904), .A(n14551), .ZN(P1_U2985) );
  NAND2_X1 U17808 ( .A1(n14553), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14556) );
  XNOR2_X1 U17809 ( .A(n14554), .B(n14557), .ZN(n14555) );
  MUX2_X1 U17810 ( .A(n14556), .B(n14555), .S(n14460), .Z(n14559) );
  INV_X1 U17811 ( .A(n14553), .ZN(n14558) );
  NAND3_X1 U17812 ( .A1(n14558), .A2(n15893), .A3(n14557), .ZN(n15922) );
  NAND2_X1 U17813 ( .A1(n14559), .A2(n15922), .ZN(n16047) );
  INV_X1 U17814 ( .A(n16047), .ZN(n14565) );
  AOI22_X1 U17815 ( .A1(n20039), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n20099), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14560) );
  OAI21_X1 U17816 ( .B1(n20050), .B2(n14561), .A(n14560), .ZN(n14562) );
  AOI21_X1 U17817 ( .B1(n14563), .B2(n20045), .A(n14562), .ZN(n14564) );
  OAI21_X1 U17818 ( .B1(n14565), .B2(n19904), .A(n14564), .ZN(P1_U2989) );
  NOR3_X1 U17819 ( .A1(n14568), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14567), .ZN(n14574) );
  NAND3_X1 U17820 ( .A1(n14570), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14569), .ZN(n14572) );
  NAND2_X1 U17821 ( .A1(n14572), .A2(n14571), .ZN(n14573) );
  OAI21_X1 U17822 ( .B1(n14576), .B2(n20088), .A(n14575), .ZN(P1_U3000) );
  NAND3_X1 U17823 ( .A1(n14600), .A2(n9998), .A3(n14580), .ZN(n14579) );
  INV_X1 U17824 ( .A(n14577), .ZN(n14578) );
  OAI211_X1 U17825 ( .C1(n14581), .C2(n14580), .A(n14579), .B(n14578), .ZN(
        n14582) );
  AOI21_X1 U17826 ( .B1(n14583), .B2(n20076), .A(n14582), .ZN(n14584) );
  OAI21_X1 U17827 ( .B1(n14585), .B2(n20088), .A(n14584), .ZN(P1_U3002) );
  NAND2_X1 U17828 ( .A1(n14586), .A2(n20079), .ZN(n14593) );
  AOI21_X1 U17829 ( .B1(n14595), .B2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14587), .ZN(n14592) );
  NAND3_X1 U17830 ( .A1(n14600), .A2(n14588), .A3(n9881), .ZN(n14591) );
  NAND2_X1 U17831 ( .A1(n14589), .A2(n20076), .ZN(n14590) );
  NAND4_X1 U17832 ( .A1(n14593), .A2(n14592), .A3(n14591), .A4(n14590), .ZN(
        P1_U3003) );
  AOI21_X1 U17833 ( .B1(n14595), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n14594), .ZN(n14596) );
  OAI21_X1 U17834 ( .B1(n14597), .B2(n20102), .A(n14596), .ZN(n14598) );
  AOI21_X1 U17835 ( .B1(n14600), .B2(n14599), .A(n14598), .ZN(n14601) );
  OAI21_X1 U17836 ( .B1(n14602), .B2(n20088), .A(n14601), .ZN(P1_U3004) );
  NOR2_X1 U17837 ( .A1(n14603), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14612) );
  NOR2_X1 U17838 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n14604), .ZN(
        n14605) );
  NAND2_X1 U17839 ( .A1(n14630), .A2(n14605), .ZN(n14617) );
  INV_X1 U17840 ( .A(n14616), .ZN(n14607) );
  AOI21_X1 U17841 ( .B1(n14617), .B2(n14607), .A(n14606), .ZN(n14611) );
  OAI21_X1 U17842 ( .B1(n14609), .B2(n20102), .A(n14608), .ZN(n14610) );
  AOI211_X1 U17843 ( .C1(n14630), .C2(n14612), .A(n14611), .B(n14610), .ZN(
        n14613) );
  OAI21_X1 U17844 ( .B1(n14614), .B2(n20088), .A(n14613), .ZN(P1_U3005) );
  AOI21_X1 U17845 ( .B1(n14616), .B2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n14615), .ZN(n14618) );
  OAI211_X1 U17846 ( .C1(n14619), .C2(n20102), .A(n14618), .B(n14617), .ZN(
        n14620) );
  INV_X1 U17847 ( .A(n14620), .ZN(n14621) );
  OAI21_X1 U17848 ( .B1(n14622), .B2(n20088), .A(n14621), .ZN(P1_U3006) );
  INV_X1 U17849 ( .A(n14623), .ZN(n14629) );
  INV_X1 U17850 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15954) );
  NOR2_X1 U17851 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n15954), .ZN(
        n15949) );
  INV_X1 U17852 ( .A(n14624), .ZN(n14625) );
  AOI21_X1 U17853 ( .B1(n20081), .B2(n15949), .A(n14625), .ZN(n14627) );
  OAI21_X1 U17854 ( .B1(n14627), .B2(n21048), .A(n14626), .ZN(n14628) );
  AOI21_X1 U17855 ( .B1(n14629), .B2(n20076), .A(n14628), .ZN(n14632) );
  NAND3_X1 U17856 ( .A1(n14630), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n21048), .ZN(n14631) );
  OAI211_X1 U17857 ( .C1(n14633), .C2(n20088), .A(n14632), .B(n14631), .ZN(
        P1_U3007) );
  INV_X1 U17858 ( .A(n15956), .ZN(n14637) );
  NOR2_X1 U17859 ( .A1(n15957), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14636) );
  OAI21_X1 U17860 ( .B1(n15792), .B2(n20102), .A(n14634), .ZN(n14635) );
  AOI211_X1 U17861 ( .C1(n14637), .C2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n14636), .B(n14635), .ZN(n14638) );
  OAI21_X1 U17862 ( .B1(n14639), .B2(n20088), .A(n14638), .ZN(P1_U3010) );
  INV_X1 U17863 ( .A(n14640), .ZN(n14647) );
  INV_X1 U17864 ( .A(n14641), .ZN(n15968) );
  OAI211_X1 U17865 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(n15968), .B(n14642), .ZN(
        n14644) );
  OAI211_X1 U17866 ( .C1(n20102), .C2(n15800), .A(n14644), .B(n14643), .ZN(
        n14645) );
  AOI21_X1 U17867 ( .B1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n15966), .A(
        n14645), .ZN(n14646) );
  OAI21_X1 U17868 ( .B1(n14647), .B2(n20088), .A(n14646), .ZN(P1_U3011) );
  XNOR2_X1 U17869 ( .A(n20214), .B(P1_STATEBS16_REG_SCAN_IN), .ZN(n14649) );
  OAI22_X1 U17870 ( .A1(n14649), .A2(n20836), .B1(n20642), .B2(n14648), .ZN(
        n14650) );
  MUX2_X1 U17871 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n14650), .S(
        n20104), .Z(P1_U3477) );
  NOR2_X1 U17872 ( .A1(n14651), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14654) );
  NOR3_X1 U17873 ( .A1(n14652), .A2(n13411), .A3(n13393), .ZN(n14653) );
  AOI211_X1 U17874 ( .C1(n20645), .C2(n14655), .A(n14654), .B(n14653), .ZN(
        n15718) );
  AOI22_X1 U17875 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n20090), .B2(n14094), .ZN(
        n14662) );
  INV_X1 U17876 ( .A(n14662), .ZN(n14657) );
  NOR2_X1 U17877 ( .A1(n20739), .A2(n20095), .ZN(n14661) );
  NOR3_X1 U17878 ( .A1(n13411), .A2(n13393), .A3(n20821), .ZN(n14656) );
  AOI21_X1 U17879 ( .B1(n14657), .B2(n14661), .A(n14656), .ZN(n14658) );
  OAI21_X1 U17880 ( .B1(n15718), .B2(n20822), .A(n14658), .ZN(n14659) );
  MUX2_X1 U17881 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14659), .S(
        n20824), .Z(P1_U3473) );
  INV_X1 U17882 ( .A(n20821), .ZN(n15750) );
  AOI22_X1 U17883 ( .A1(n14662), .A2(n14661), .B1(n14660), .B2(n15750), .ZN(
        n14663) );
  OAI21_X1 U17884 ( .B1(n14664), .B2(n20822), .A(n14663), .ZN(n14665) );
  MUX2_X1 U17885 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14665), .S(
        n20824), .Z(P1_U3472) );
  NAND2_X1 U17886 ( .A1(n14666), .A2(n14667), .ZN(n14669) );
  OAI21_X1 U17887 ( .B1(n14667), .B2(n19420), .A(n10274), .ZN(n14668) );
  MUX2_X1 U17888 ( .A(n14669), .B(n14668), .S(n9788), .Z(n14672) );
  INV_X1 U17889 ( .A(n14670), .ZN(n16367) );
  OAI22_X1 U17890 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16367), .B1(n19785), 
        .B2(n19544), .ZN(n14671) );
  OAI21_X1 U17891 ( .B1(n14672), .B2(n18894), .A(n14671), .ZN(n14675) );
  NOR2_X1 U17892 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n15363), .ZN(n19199) );
  CLKBUF_X2 U17893 ( .A(n19199), .Z(n19178) );
  AOI21_X1 U17894 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n16363), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n14673) );
  AOI211_X1 U17895 ( .C1(n19178), .C2(n19765), .A(n14673), .B(n18895), .ZN(
        n14674) );
  MUX2_X1 U17896 ( .A(n14675), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n14674), 
        .Z(P2_U3610) );
  INV_X1 U17897 ( .A(n14676), .ZN(n14720) );
  AOI21_X1 U17898 ( .B1(n14679), .B2(n14678), .A(n14677), .ZN(n14988) );
  INV_X1 U17899 ( .A(n14988), .ZN(n16128) );
  NOR2_X1 U17900 ( .A1(n14681), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14682) );
  OR2_X1 U17901 ( .A1(n14041), .A2(n14682), .ZN(n16150) );
  INV_X1 U17902 ( .A(n14683), .ZN(n16163) );
  AOI21_X1 U17903 ( .B1(n15029), .B2(n14684), .A(n14705), .ZN(n15032) );
  OAI21_X1 U17904 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n14685), .A(
        n14703), .ZN(n18945) );
  INV_X1 U17905 ( .A(n18945), .ZN(n14702) );
  AOI21_X1 U17906 ( .B1(n18975), .B2(n14698), .A(n14701), .ZN(n18974) );
  OAI21_X1 U17907 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n14696), .A(
        n14686), .ZN(n16237) );
  INV_X1 U17908 ( .A(n16237), .ZN(n14750) );
  OAI21_X1 U17909 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n9845), .A(
        n14697), .ZN(n16246) );
  INV_X1 U17910 ( .A(n16246), .ZN(n14778) );
  OAI21_X1 U17911 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n14692), .A(
        n14695), .ZN(n16261) );
  INV_X1 U17912 ( .A(n16261), .ZN(n14795) );
  AOI21_X1 U17913 ( .B1(n16282), .B2(n14690), .A(n14687), .ZN(n16272) );
  AOI21_X1 U17914 ( .B1(n19041), .B2(n14688), .A(n14691), .ZN(n19034) );
  NOR2_X1 U17915 ( .A1(n19202), .A2(n14689), .ZN(n19046) );
  NAND2_X1 U17916 ( .A1(n19046), .A2(n19047), .ZN(n19031) );
  NOR2_X1 U17917 ( .A1(n19034), .A2(n19031), .ZN(n19016) );
  OAI21_X1 U17918 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n14691), .A(
        n14690), .ZN(n19018) );
  NAND2_X1 U17919 ( .A1(n19016), .A2(n19018), .ZN(n14805) );
  NOR2_X1 U17920 ( .A1(n16272), .A2(n14805), .ZN(n19006) );
  AOI21_X1 U17921 ( .B1(n16271), .B2(n14693), .A(n14692), .ZN(n19007) );
  INV_X1 U17922 ( .A(n19007), .ZN(n14694) );
  NAND2_X1 U17923 ( .A1(n19006), .A2(n14694), .ZN(n14793) );
  NOR2_X1 U17924 ( .A1(n14795), .A2(n14793), .ZN(n18995) );
  AOI21_X1 U17925 ( .B1(n15100), .B2(n14695), .A(n9845), .ZN(n18997) );
  INV_X1 U17926 ( .A(n18997), .ZN(n15099) );
  NAND2_X1 U17927 ( .A1(n18995), .A2(n15099), .ZN(n14776) );
  NOR2_X1 U17928 ( .A1(n14778), .A2(n14776), .ZN(n14765) );
  AOI21_X1 U17929 ( .B1(n15084), .B2(n14697), .A(n14696), .ZN(n15087) );
  INV_X1 U17930 ( .A(n15087), .ZN(n14764) );
  NAND2_X1 U17931 ( .A1(n14765), .A2(n14764), .ZN(n14749) );
  NOR2_X1 U17932 ( .A1(n14750), .A2(n14749), .ZN(n18986) );
  OAI21_X1 U17933 ( .B1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n14699), .A(
        n14698), .ZN(n18988) );
  NAND2_X1 U17934 ( .A1(n18986), .A2(n18988), .ZN(n18972) );
  NOR2_X1 U17935 ( .A1(n18974), .A2(n18972), .ZN(n18968) );
  OAI21_X1 U17936 ( .B1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n14701), .A(
        n14700), .ZN(n18967) );
  NAND2_X1 U17937 ( .A1(n18968), .A2(n18967), .ZN(n18944) );
  NOR2_X1 U17938 ( .A1(n14702), .A2(n18944), .ZN(n18935) );
  AOI21_X1 U17939 ( .B1(n21034), .B2(n14703), .A(n9844), .ZN(n15045) );
  INV_X1 U17940 ( .A(n15045), .ZN(n18936) );
  NAND2_X1 U17941 ( .A1(n18935), .A2(n18936), .ZN(n18920) );
  NOR2_X1 U17942 ( .A1(n18923), .A2(n18920), .ZN(n14732) );
  OAI21_X1 U17943 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n14705), .A(
        n14706), .ZN(n16223) );
  NAND2_X1 U17944 ( .A1(n15712), .A2(n16223), .ZN(n15711) );
  NAND2_X1 U17945 ( .A1(n14707), .A2(n15711), .ZN(n16183) );
  AOI21_X1 U17946 ( .B1(n15010), .B2(n14706), .A(n14709), .ZN(n15013) );
  INV_X1 U17947 ( .A(n15013), .ZN(n16184) );
  NAND2_X1 U17948 ( .A1(n16183), .A2(n16184), .ZN(n16182) );
  NAND2_X1 U17949 ( .A1(n14707), .A2(n16182), .ZN(n16174) );
  OAI21_X1 U17950 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n14709), .A(
        n14708), .ZN(n16213) );
  NAND2_X1 U17951 ( .A1(n16174), .A2(n16213), .ZN(n16173) );
  NAND2_X1 U17952 ( .A1(n19032), .A2(n16173), .ZN(n16162) );
  NAND2_X1 U17953 ( .A1(n16163), .A2(n16162), .ZN(n16161) );
  NAND2_X1 U17954 ( .A1(n19032), .A2(n16161), .ZN(n16149) );
  NAND2_X1 U17955 ( .A1(n16150), .A2(n16149), .ZN(n16148) );
  NAND2_X1 U17956 ( .A1(n19032), .A2(n16148), .ZN(n16140) );
  NAND2_X1 U17957 ( .A1(n14054), .A2(n16140), .ZN(n16139) );
  NAND2_X1 U17958 ( .A1(n19032), .A2(n16139), .ZN(n14723) );
  NAND2_X1 U17959 ( .A1(n14722), .A2(n14723), .ZN(n14721) );
  NAND2_X1 U17960 ( .A1(n19032), .A2(n14721), .ZN(n16127) );
  NAND2_X1 U17961 ( .A1(n16128), .A2(n16127), .ZN(n16126) );
  NAND2_X1 U17962 ( .A1(n19032), .A2(n16126), .ZN(n14711) );
  NAND2_X1 U17963 ( .A1(n14711), .A2(n14710), .ZN(n16120) );
  OAI211_X1 U17964 ( .C1(n14711), .C2(n14710), .A(n16120), .B(n18939), .ZN(
        n14719) );
  INV_X1 U17965 ( .A(n14712), .ZN(n14713) );
  OAI22_X1 U17966 ( .A1(n14713), .A2(n19063), .B1(n10946), .B2(n19028), .ZN(
        n14716) );
  INV_X1 U17967 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14714) );
  OAI22_X1 U17968 ( .A1(n14714), .A2(n19057), .B1(n19836), .B2(n9807), .ZN(
        n14715) );
  AOI211_X1 U17969 ( .C1(n14717), .C2(n19066), .A(n14716), .B(n14715), .ZN(
        n14718) );
  OAI211_X1 U17970 ( .C1(n14720), .C2(n19042), .A(n14719), .B(n14718), .ZN(
        P2_U2825) );
  OAI211_X1 U17971 ( .C1(n14723), .C2(n14722), .A(n19050), .B(n14721), .ZN(
        n14730) );
  INV_X1 U17972 ( .A(n14852), .ZN(n14728) );
  OAI22_X1 U17973 ( .A1(n12478), .A2(n9807), .B1(n10904), .B2(n19028), .ZN(
        n14727) );
  INV_X1 U17974 ( .A(n14922), .ZN(n14725) );
  INV_X1 U17975 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14724) );
  OAI22_X1 U17976 ( .A1(n14725), .A2(n19063), .B1(n14724), .B2(n19057), .ZN(
        n14726) );
  AOI211_X1 U17977 ( .C1(n14728), .C2(n19066), .A(n14727), .B(n14726), .ZN(
        n14729) );
  OAI211_X1 U17978 ( .C1(n19042), .C2(n14731), .A(n14730), .B(n14729), .ZN(
        P2_U2827) );
  OAI22_X1 U17979 ( .A1(n19823), .A2(n9807), .B1(n14903), .B2(n19028), .ZN(
        n14737) );
  NAND2_X1 U17980 ( .A1(n19050), .A2(n19032), .ZN(n19071) );
  OR2_X1 U17981 ( .A1(n14732), .A2(n19071), .ZN(n18919) );
  INV_X1 U17982 ( .A(n18919), .ZN(n14735) );
  NOR2_X1 U17983 ( .A1(n14733), .A2(n19771), .ZN(n14734) );
  MUX2_X1 U17984 ( .A(n14735), .B(n14734), .S(n15032), .Z(n14736) );
  AOI211_X1 U17985 ( .C1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(n19003), .A(
        n14737), .B(n14736), .ZN(n14747) );
  NAND2_X1 U17986 ( .A1(n11292), .A2(n14739), .ZN(n14740) );
  NAND2_X1 U17987 ( .A1(n14738), .A2(n14740), .ZN(n15204) );
  OR2_X1 U17988 ( .A1(n14741), .A2(n12497), .ZN(n14744) );
  INV_X1 U17989 ( .A(n15194), .ZN(n14743) );
  NAND2_X1 U17990 ( .A1(n14744), .A2(n14743), .ZN(n15207) );
  OAI22_X1 U17991 ( .A1(n15204), .A2(n19036), .B1(n19063), .B2(n15207), .ZN(
        n14745) );
  INV_X1 U17992 ( .A(n14745), .ZN(n14746) );
  OAI211_X1 U17993 ( .C1(n14748), .C2(n19042), .A(n14747), .B(n14746), .ZN(
        P2_U2834) );
  NAND2_X1 U17994 ( .A1(n19032), .A2(n14749), .ZN(n14762) );
  XNOR2_X1 U17995 ( .A(n14750), .B(n14762), .ZN(n14751) );
  NAND2_X1 U17996 ( .A1(n14751), .A2(n19050), .ZN(n14760) );
  AOI21_X1 U17997 ( .B1(n14754), .B2(n14753), .A(n14752), .ZN(n19087) );
  INV_X1 U17998 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n19813) );
  OAI21_X1 U17999 ( .B1(n19813), .B2(n9807), .A(n18957), .ZN(n14755) );
  AOI21_X1 U18000 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19024), .A(
        n14755), .ZN(n14756) );
  OAI21_X1 U18001 ( .B1(n16234), .B2(n19036), .A(n14756), .ZN(n14758) );
  NOR2_X1 U18002 ( .A1(n19028), .A2(n10661), .ZN(n14757) );
  AOI211_X1 U18003 ( .C1(n18980), .C2(n19087), .A(n14758), .B(n14757), .ZN(
        n14759) );
  OAI211_X1 U18004 ( .C1(n19042), .C2(n14761), .A(n14760), .B(n14759), .ZN(
        P2_U2841) );
  INV_X1 U18005 ( .A(n14762), .ZN(n14763) );
  OAI211_X1 U18006 ( .C1(n14765), .C2(n14764), .A(n19050), .B(n14763), .ZN(
        n14775) );
  OAI22_X1 U18007 ( .A1(n15084), .A2(n19057), .B1(n10657), .B2(n19028), .ZN(
        n14773) );
  XNOR2_X1 U18008 ( .A(n14766), .B(n14767), .ZN(n19092) );
  AOI22_X1 U18009 ( .A1(n19055), .A2(n15087), .B1(n19060), .B2(n14768), .ZN(
        n14769) );
  OAI211_X1 U18010 ( .C1(n10855), .C2(n9807), .A(n14769), .B(n18957), .ZN(
        n14770) );
  AOI21_X1 U18011 ( .B1(n15282), .B2(n19066), .A(n14770), .ZN(n14771) );
  OAI21_X1 U18012 ( .B1(n19092), .B2(n19063), .A(n14771), .ZN(n14772) );
  NOR2_X1 U18013 ( .A1(n14773), .A2(n14772), .ZN(n14774) );
  NAND2_X1 U18014 ( .A1(n14775), .A2(n14774), .ZN(P2_U2842) );
  INV_X1 U18015 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n14789) );
  NAND2_X1 U18016 ( .A1(n19032), .A2(n14776), .ZN(n14777) );
  XNOR2_X1 U18017 ( .A(n14778), .B(n14777), .ZN(n14779) );
  NAND2_X1 U18018 ( .A1(n14779), .A2(n19050), .ZN(n14788) );
  AOI21_X1 U18019 ( .B1(n14781), .B2(n14780), .A(n14766), .ZN(n19093) );
  NAND2_X1 U18020 ( .A1(n18980), .A2(n19093), .ZN(n14783) );
  AOI21_X1 U18021 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19024), .A(
        n19030), .ZN(n14782) );
  OAI211_X1 U18022 ( .C1(n16298), .C2(n19036), .A(n14783), .B(n14782), .ZN(
        n14786) );
  NOR2_X1 U18023 ( .A1(n14784), .A2(n19042), .ZN(n14785) );
  AOI211_X1 U18024 ( .C1(n19054), .C2(P2_EBX_REG_12__SCAN_IN), .A(n14786), .B(
        n14785), .ZN(n14787) );
  OAI211_X1 U18025 ( .C1(n9807), .C2(n14789), .A(n14788), .B(n14787), .ZN(
        P2_U2843) );
  AOI21_X1 U18026 ( .B1(n15309), .B2(n14792), .A(n14791), .ZN(n16312) );
  INV_X1 U18027 ( .A(n16312), .ZN(n19101) );
  NAND2_X1 U18028 ( .A1(n19032), .A2(n14793), .ZN(n14794) );
  XNOR2_X1 U18029 ( .A(n14795), .B(n14794), .ZN(n14796) );
  NAND2_X1 U18030 ( .A1(n14796), .A2(n19050), .ZN(n14804) );
  AOI21_X1 U18031 ( .B1(n19024), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n19030), .ZN(n14798) );
  NAND2_X1 U18032 ( .A1(n19054), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n14797) );
  OAI211_X1 U18033 ( .C1(n14799), .C2(n19042), .A(n14798), .B(n14797), .ZN(
        n14802) );
  INV_X1 U18034 ( .A(n16313), .ZN(n14800) );
  NOR2_X1 U18035 ( .A1(n14800), .A2(n19036), .ZN(n14801) );
  AOI211_X1 U18036 ( .C1(n9882), .C2(P2_REIP_REG_10__SCAN_IN), .A(n14802), .B(
        n14801), .ZN(n14803) );
  OAI211_X1 U18037 ( .C1(n19063), .C2(n19101), .A(n14804), .B(n14803), .ZN(
        P2_U2845) );
  NAND2_X1 U18038 ( .A1(n19032), .A2(n14805), .ZN(n14806) );
  XNOR2_X1 U18039 ( .A(n16272), .B(n14806), .ZN(n14807) );
  NAND2_X1 U18040 ( .A1(n14807), .A2(n19050), .ZN(n14817) );
  AOI21_X1 U18041 ( .B1(n14810), .B2(n14808), .A(n14809), .ZN(n16319) );
  INV_X1 U18042 ( .A(n16319), .ZN(n19107) );
  NAND2_X1 U18043 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19024), .ZN(
        n14811) );
  OAI211_X1 U18044 ( .C1(n19063), .C2(n19107), .A(n18957), .B(n14811), .ZN(
        n14812) );
  AOI21_X1 U18045 ( .B1(P2_EBX_REG_8__SCAN_IN), .B2(n19054), .A(n14812), .ZN(
        n14813) );
  OAI21_X1 U18046 ( .B1(n14814), .B2(n19042), .A(n14813), .ZN(n14815) );
  AOI21_X1 U18047 ( .B1(n9882), .B2(P2_REIP_REG_8__SCAN_IN), .A(n14815), .ZN(
        n14816) );
  OAI211_X1 U18048 ( .C1(n14818), .C2(n19036), .A(n14817), .B(n14816), .ZN(
        P2_U2847) );
  NAND2_X1 U18049 ( .A1(n19032), .A2(n14829), .ZN(n14819) );
  XNOR2_X1 U18050 ( .A(n14820), .B(n14819), .ZN(n14821) );
  NAND2_X1 U18051 ( .A1(n14821), .A2(n19050), .ZN(n14828) );
  NAND2_X1 U18052 ( .A1(n13265), .A2(n19066), .ZN(n14824) );
  OAI22_X1 U18053 ( .A1(n19795), .A2(n9807), .B1(n10325), .B2(n19028), .ZN(
        n14822) );
  AOI21_X1 U18054 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19003), .A(
        n14822), .ZN(n14823) );
  OAI211_X1 U18055 ( .C1(n19042), .C2(n14825), .A(n14824), .B(n14823), .ZN(
        n14826) );
  AOI21_X1 U18056 ( .B1(n19866), .B2(n18980), .A(n14826), .ZN(n14827) );
  OAI211_X1 U18057 ( .C1(n19068), .C2(n19864), .A(n14828), .B(n14827), .ZN(
        P2_U2853) );
  OAI211_X1 U18058 ( .C1(n19072), .C2(n14830), .A(n19032), .B(n14829), .ZN(
        n15369) );
  NAND2_X1 U18059 ( .A1(n18980), .A2(n19875), .ZN(n14835) );
  AOI22_X1 U18060 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n9882), .B1(
        P2_EBX_REG_1__SCAN_IN), .B2(n19054), .ZN(n14831) );
  OAI21_X1 U18061 ( .B1(n19057), .B2(n14833), .A(n14831), .ZN(n14832) );
  AOI21_X1 U18062 ( .B1(n19055), .B2(n14833), .A(n14832), .ZN(n14834) );
  OAI211_X1 U18063 ( .C1(n19042), .C2(n14836), .A(n14835), .B(n14834), .ZN(
        n14838) );
  NOR2_X1 U18064 ( .A1(n19871), .A2(n19068), .ZN(n14837) );
  AOI211_X1 U18065 ( .C1(n19066), .C2(n9792), .A(n14838), .B(n14837), .ZN(
        n14839) );
  OAI21_X1 U18066 ( .B1(n15369), .B2(n19771), .A(n14839), .ZN(P2_U2854) );
  INV_X1 U18067 ( .A(n14840), .ZN(n16117) );
  MUX2_X1 U18068 ( .A(P2_EBX_REG_31__SCAN_IN), .B(n16117), .S(n14901), .Z(
        P2_U2856) );
  NOR2_X1 U18069 ( .A1(n14842), .A2(n14841), .ZN(n14843) );
  NAND2_X1 U18070 ( .A1(n14845), .A2(n14844), .ZN(n14912) );
  NAND3_X1 U18071 ( .A1(n9821), .A2(n14894), .A3(n14912), .ZN(n14847) );
  NAND2_X1 U18072 ( .A1(n14909), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14846) );
  OAI211_X1 U18073 ( .C1(n14909), .C2(n16124), .A(n14847), .B(n14846), .ZN(
        P2_U2858) );
  NAND2_X1 U18074 ( .A1(n14848), .A2(n14849), .ZN(n14851) );
  XNOR2_X1 U18075 ( .A(n14851), .B(n14850), .ZN(n14925) );
  NOR2_X1 U18076 ( .A1(n14852), .A2(n14909), .ZN(n14853) );
  AOI21_X1 U18077 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n13168), .A(n14853), .ZN(
        n14854) );
  OAI21_X1 U18078 ( .B1(n14925), .B2(n14911), .A(n14854), .ZN(P2_U2859) );
  AOI21_X1 U18079 ( .B1(n14857), .B2(n14856), .A(n14855), .ZN(n14858) );
  INV_X1 U18080 ( .A(n14858), .ZN(n14932) );
  NOR2_X1 U18081 ( .A1(n16133), .A2(n13168), .ZN(n14859) );
  AOI21_X1 U18082 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n14909), .A(n14859), .ZN(
        n14860) );
  OAI21_X1 U18083 ( .B1(n14932), .B2(n14911), .A(n14860), .ZN(P2_U2860) );
  OR2_X1 U18084 ( .A1(n13943), .A2(n14861), .ZN(n14862) );
  NAND2_X1 U18085 ( .A1(n14045), .A2(n14862), .ZN(n14999) );
  AOI21_X1 U18086 ( .B1(n14866), .B2(n14865), .A(n14864), .ZN(n14939) );
  NAND2_X1 U18087 ( .A1(n14939), .A2(n14894), .ZN(n14868) );
  NAND2_X1 U18088 ( .A1(n13168), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n14867) );
  OAI211_X1 U18089 ( .C1(n13168), .C2(n14999), .A(n14868), .B(n14867), .ZN(
        P2_U2861) );
  OAI21_X1 U18090 ( .B1(n14871), .B2(n14870), .A(n14869), .ZN(n14947) );
  MUX2_X1 U18091 ( .A(n16158), .B(n14872), .S(n14909), .Z(n14873) );
  OAI21_X1 U18092 ( .B1(n14947), .B2(n14911), .A(n14873), .ZN(P2_U2862) );
  AOI21_X1 U18093 ( .B1(n9854), .B2(n14875), .A(n14874), .ZN(n14876) );
  XOR2_X1 U18094 ( .A(n14877), .B(n14876), .Z(n14955) );
  NOR2_X1 U18095 ( .A1(n14886), .A2(n14878), .ZN(n14879) );
  OR2_X1 U18096 ( .A1(n13944), .A2(n14879), .ZN(n16169) );
  NOR2_X1 U18097 ( .A1(n16169), .A2(n13168), .ZN(n14880) );
  AOI21_X1 U18098 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n14909), .A(n14880), .ZN(
        n14881) );
  OAI21_X1 U18099 ( .B1(n14955), .B2(n14911), .A(n14881), .ZN(P2_U2863) );
  AOI21_X1 U18100 ( .B1(n14884), .B2(n14883), .A(n14882), .ZN(n14885) );
  INV_X1 U18101 ( .A(n14885), .ZN(n14962) );
  INV_X1 U18102 ( .A(n14886), .ZN(n14889) );
  NAND2_X1 U18103 ( .A1(n14897), .A2(n14887), .ZN(n14888) );
  NAND2_X1 U18104 ( .A1(n14889), .A2(n14888), .ZN(n16179) );
  MUX2_X1 U18105 ( .A(n10888), .B(n16179), .S(n14901), .Z(n14890) );
  OAI21_X1 U18106 ( .B1(n14962), .B2(n14911), .A(n14890), .ZN(P2_U2864) );
  INV_X1 U18107 ( .A(n14891), .ZN(n14893) );
  AOI21_X1 U18108 ( .B1(n14893), .B2(n9842), .A(n14892), .ZN(n16191) );
  NAND2_X1 U18109 ( .A1(n16191), .A2(n14894), .ZN(n14899) );
  NAND2_X1 U18110 ( .A1(n14738), .A2(n14895), .ZN(n14896) );
  NAND2_X1 U18111 ( .A1(n14897), .A2(n14896), .ZN(n15196) );
  NAND2_X1 U18112 ( .A1(n14901), .A2(n16217), .ZN(n14898) );
  OAI211_X1 U18113 ( .C1(n14901), .C2(n14900), .A(n14899), .B(n14898), .ZN(
        P2_U2865) );
  OAI21_X1 U18114 ( .B1(n13904), .B2(n14902), .A(n9842), .ZN(n14969) );
  MUX2_X1 U18115 ( .A(n15204), .B(n14903), .S(n14909), .Z(n14904) );
  OAI21_X1 U18116 ( .B1(n14969), .B2(n14911), .A(n14904), .ZN(P2_U2866) );
  OAI21_X1 U18117 ( .B1(n13839), .B2(n14906), .A(n14905), .ZN(n14982) );
  AOI21_X1 U18118 ( .B1(n14907), .B2(n9958), .A(n11293), .ZN(n18938) );
  INV_X1 U18119 ( .A(n18938), .ZN(n15042) );
  NOR2_X1 U18120 ( .A1(n14909), .A2(n15042), .ZN(n14908) );
  AOI21_X1 U18121 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n14909), .A(n14908), .ZN(
        n14910) );
  OAI21_X1 U18122 ( .B1(n14982), .B2(n14911), .A(n14910), .ZN(P2_U2868) );
  NAND3_X1 U18123 ( .A1(n9821), .A2(n19131), .A3(n14912), .ZN(n14919) );
  OR2_X1 U18124 ( .A1(n14914), .A2(n14913), .ZN(n14915) );
  INV_X1 U18125 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n19143) );
  OAI22_X1 U18126 ( .A1(n14973), .A2(n19091), .B1(n19110), .B2(n19143), .ZN(
        n14916) );
  AOI21_X1 U18127 ( .B1(n19127), .B2(n16122), .A(n14916), .ZN(n14918) );
  AOI22_X1 U18128 ( .A1(n19078), .A2(BUF1_REG_29__SCAN_IN), .B1(n19077), .B2(
        BUF2_REG_29__SCAN_IN), .ZN(n14917) );
  NAND3_X1 U18129 ( .A1(n14919), .A2(n14918), .A3(n14917), .ZN(P2_U2890) );
  INV_X1 U18130 ( .A(n19094), .ZN(n14920) );
  OAI22_X1 U18131 ( .A1(n14973), .A2(n14920), .B1(n19110), .B2(n20973), .ZN(
        n14921) );
  AOI21_X1 U18132 ( .B1(n19127), .B2(n14922), .A(n14921), .ZN(n14924) );
  AOI22_X1 U18133 ( .A1(n19078), .A2(BUF1_REG_28__SCAN_IN), .B1(n19077), .B2(
        BUF2_REG_28__SCAN_IN), .ZN(n14923) );
  OAI211_X1 U18134 ( .C1(n14925), .C2(n19112), .A(n14924), .B(n14923), .ZN(
        P2_U2891) );
  NAND2_X1 U18135 ( .A1(n14933), .A2(n14926), .ZN(n14927) );
  NAND2_X1 U18136 ( .A1(n14928), .A2(n14927), .ZN(n16143) );
  INV_X1 U18137 ( .A(n16143), .ZN(n15141) );
  INV_X1 U18138 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n19146) );
  OAI22_X1 U18139 ( .A1(n14973), .A2(n19097), .B1(n19110), .B2(n19146), .ZN(
        n14929) );
  AOI21_X1 U18140 ( .B1(n19127), .B2(n15141), .A(n14929), .ZN(n14931) );
  AOI22_X1 U18141 ( .A1(n19078), .A2(BUF1_REG_27__SCAN_IN), .B1(n19077), .B2(
        BUF2_REG_27__SCAN_IN), .ZN(n14930) );
  OAI211_X1 U18142 ( .C1(n14932), .C2(n19112), .A(n14931), .B(n14930), .ZN(
        P2_U2892) );
  OAI21_X1 U18143 ( .B1(n14935), .B2(n14934), .A(n14933), .ZN(n16145) );
  AOI22_X1 U18144 ( .A1(n19078), .A2(BUF1_REG_26__SCAN_IN), .B1(n19077), .B2(
        BUF2_REG_26__SCAN_IN), .ZN(n14937) );
  INV_X1 U18145 ( .A(n14973), .ZN(n19076) );
  AOI22_X1 U18146 ( .A1(n19076), .A2(n19099), .B1(P2_EAX_REG_26__SCAN_IN), 
        .B2(n19126), .ZN(n14936) );
  OAI211_X1 U18147 ( .C1(n19084), .C2(n16145), .A(n14937), .B(n14936), .ZN(
        n14938) );
  AOI21_X1 U18148 ( .B1(n14939), .B2(n19131), .A(n14938), .ZN(n14940) );
  INV_X1 U18149 ( .A(n14940), .ZN(P2_U2893) );
  INV_X1 U18150 ( .A(n19103), .ZN(n14941) );
  INV_X1 U18151 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n19149) );
  OAI22_X1 U18152 ( .A1(n14973), .A2(n14941), .B1(n19110), .B2(n19149), .ZN(
        n14945) );
  INV_X1 U18153 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n14943) );
  INV_X1 U18154 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n14942) );
  OAI22_X1 U18155 ( .A1(n14977), .A2(n14943), .B1(n14975), .B2(n14942), .ZN(
        n14944) );
  AOI211_X1 U18156 ( .C1(n19127), .C2(n16159), .A(n14945), .B(n14944), .ZN(
        n14946) );
  OAI21_X1 U18157 ( .B1(n14947), .B2(n19112), .A(n14946), .ZN(P2_U2894) );
  AND2_X1 U18158 ( .A1(n14949), .A2(n14948), .ZN(n14951) );
  OR2_X1 U18159 ( .A1(n14951), .A2(n14950), .ZN(n16177) );
  INV_X1 U18160 ( .A(n16177), .ZN(n15169) );
  INV_X1 U18161 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n19151) );
  OAI22_X1 U18162 ( .A1(n14973), .A2(n19106), .B1(n19110), .B2(n19151), .ZN(
        n14952) );
  AOI21_X1 U18163 ( .B1(n19127), .B2(n15169), .A(n14952), .ZN(n14954) );
  AOI22_X1 U18164 ( .A1(n19078), .A2(BUF1_REG_24__SCAN_IN), .B1(n19077), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n14953) );
  OAI211_X1 U18165 ( .C1(n14955), .C2(n19112), .A(n14954), .B(n14953), .ZN(
        P2_U2895) );
  XNOR2_X1 U18166 ( .A(n14956), .B(n14957), .ZN(n15176) );
  INV_X1 U18167 ( .A(n15176), .ZN(n16180) );
  INV_X1 U18168 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n19153) );
  OAI22_X1 U18169 ( .A1(n14973), .A2(n19281), .B1(n19110), .B2(n19153), .ZN(
        n14960) );
  INV_X1 U18170 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n14958) );
  OAI22_X1 U18171 ( .A1(n14977), .A2(n16478), .B1(n14975), .B2(n14958), .ZN(
        n14959) );
  AOI211_X1 U18172 ( .C1(n19127), .C2(n16180), .A(n14960), .B(n14959), .ZN(
        n14961) );
  OAI21_X1 U18173 ( .B1(n14962), .B2(n19112), .A(n14961), .ZN(P2_U2896) );
  INV_X1 U18174 ( .A(n15207), .ZN(n14967) );
  INV_X1 U18175 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n19157) );
  OAI22_X1 U18176 ( .A1(n14973), .A2(n19266), .B1(n19110), .B2(n19157), .ZN(
        n14966) );
  INV_X1 U18177 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n14964) );
  INV_X1 U18178 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n14963) );
  OAI22_X1 U18179 ( .A1(n14977), .A2(n14964), .B1(n14975), .B2(n14963), .ZN(
        n14965) );
  AOI211_X1 U18180 ( .C1(n19127), .C2(n14967), .A(n14966), .B(n14965), .ZN(
        n14968) );
  OAI21_X1 U18181 ( .B1(n14969), .B2(n19112), .A(n14968), .ZN(P2_U2898) );
  OR2_X1 U18182 ( .A1(n14971), .A2(n14970), .ZN(n14972) );
  NAND2_X1 U18183 ( .A1(n14972), .A2(n9798), .ZN(n18943) );
  INV_X1 U18184 ( .A(n18943), .ZN(n14980) );
  INV_X1 U18185 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n19161) );
  OAI22_X1 U18186 ( .A1(n14973), .A2(n19254), .B1(n19110), .B2(n19161), .ZN(
        n14979) );
  INV_X1 U18187 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n14976) );
  INV_X1 U18188 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n14974) );
  OAI22_X1 U18189 ( .A1(n14977), .A2(n14976), .B1(n14975), .B2(n14974), .ZN(
        n14978) );
  AOI211_X1 U18190 ( .C1(n19127), .C2(n14980), .A(n14979), .B(n14978), .ZN(
        n14981) );
  OAI21_X1 U18191 ( .B1(n14982), .B2(n19112), .A(n14981), .ZN(P2_U2900) );
  NAND2_X1 U18192 ( .A1(n14984), .A2(n14983), .ZN(n14986) );
  XOR2_X1 U18193 ( .A(n14986), .B(n14985), .Z(n15136) );
  AOI21_X1 U18194 ( .B1(n15137), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14987) );
  NOR2_X1 U18195 ( .A1(n14987), .A2(n10979), .ZN(n15126) );
  NAND2_X1 U18196 ( .A1(n14988), .A2(n19203), .ZN(n14990) );
  NOR2_X1 U18197 ( .A1(n15334), .A2(n19833), .ZN(n15129) );
  AOI21_X1 U18198 ( .B1(n16247), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15129), .ZN(n14989) );
  OAI211_X1 U18199 ( .C1(n13644), .C2(n16124), .A(n14990), .B(n14989), .ZN(
        n14991) );
  AOI21_X1 U18200 ( .B1(n15126), .B2(n19204), .A(n14991), .ZN(n14992) );
  OAI21_X1 U18201 ( .B1(n15136), .B2(n16263), .A(n14992), .ZN(P2_U2985) );
  OAI21_X1 U18202 ( .B1(n13941), .B2(n10732), .A(n14994), .ZN(n14995) );
  XOR2_X1 U18203 ( .A(n14996), .B(n14995), .Z(n15160) );
  INV_X1 U18204 ( .A(n13953), .ZN(n14998) );
  AOI21_X1 U18205 ( .B1(n15153), .B2(n14998), .A(n14997), .ZN(n15158) );
  INV_X1 U18206 ( .A(n14999), .ZN(n16147) );
  INV_X1 U18207 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15001) );
  OAI22_X1 U18208 ( .A1(n19212), .A2(n15001), .B1(n15000), .B2(n18957), .ZN(
        n15002) );
  AOI21_X1 U18209 ( .B1(n16147), .B2(n19207), .A(n15002), .ZN(n15003) );
  OAI21_X1 U18210 ( .B1(n16150), .B2(n16262), .A(n15003), .ZN(n15004) );
  AOI21_X1 U18211 ( .B1(n15158), .B2(n19204), .A(n15004), .ZN(n15005) );
  OAI21_X1 U18212 ( .B1(n15160), .B2(n16263), .A(n15005), .ZN(P2_U2988) );
  INV_X1 U18213 ( .A(n16215), .ZN(n15009) );
  INV_X1 U18214 ( .A(n15007), .ZN(n15008) );
  OAI21_X1 U18215 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15009), .A(
        n15008), .ZN(n15185) );
  OAI22_X1 U18216 ( .A1(n19212), .A2(n15010), .B1(n19825), .B2(n15334), .ZN(
        n15012) );
  NOR2_X1 U18217 ( .A1(n16179), .A2(n13644), .ZN(n15011) );
  AOI211_X1 U18218 ( .C1(n15013), .C2(n19203), .A(n15012), .B(n15011), .ZN(
        n15018) );
  OR2_X1 U18219 ( .A1(n15015), .A2(n15014), .ZN(n15174) );
  NAND3_X1 U18220 ( .A1(n15174), .A2(n15016), .A3(n11305), .ZN(n15017) );
  OAI211_X1 U18221 ( .C1(n15185), .C2(n16265), .A(n15018), .B(n15017), .ZN(
        P2_U2991) );
  INV_X1 U18222 ( .A(n15019), .ZN(n15021) );
  NAND2_X1 U18223 ( .A1(n11284), .A2(n15020), .ZN(n15190) );
  OAI21_X1 U18224 ( .B1(n15021), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15190), .ZN(n15215) );
  NAND2_X1 U18225 ( .A1(n15023), .A2(n15022), .ZN(n15028) );
  OAI21_X1 U18226 ( .B1(n15026), .B2(n15025), .A(n15024), .ZN(n15027) );
  XNOR2_X1 U18227 ( .A(n15028), .B(n15027), .ZN(n15202) );
  NAND2_X1 U18228 ( .A1(n15202), .A2(n11305), .ZN(n15034) );
  OAI22_X1 U18229 ( .A1(n19212), .A2(n15029), .B1(n19823), .B2(n15334), .ZN(
        n15031) );
  NOR2_X1 U18230 ( .A1(n13644), .A2(n15204), .ZN(n15030) );
  AOI211_X1 U18231 ( .C1(n15032), .C2(n19203), .A(n15031), .B(n15030), .ZN(
        n15033) );
  OAI211_X1 U18232 ( .C1(n16265), .C2(n15215), .A(n15034), .B(n15033), .ZN(
        P2_U2993) );
  OAI21_X1 U18233 ( .B1(n15225), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15035), .ZN(n15223) );
  NAND2_X1 U18234 ( .A1(n15037), .A2(n15036), .ZN(n15041) );
  INV_X1 U18235 ( .A(n15038), .ZN(n15229) );
  INV_X1 U18236 ( .A(n15227), .ZN(n15039) );
  AOI21_X1 U18237 ( .B1(n15226), .B2(n15229), .A(n15039), .ZN(n15040) );
  XNOR2_X1 U18238 ( .A(n15041), .B(n15040), .ZN(n15216) );
  NAND2_X1 U18239 ( .A1(n15216), .A2(n11305), .ZN(n15047) );
  OAI22_X1 U18240 ( .A1(n19212), .A2(n21034), .B1(n10873), .B2(n18957), .ZN(
        n15044) );
  NOR2_X1 U18241 ( .A1(n13644), .A2(n15042), .ZN(n15043) );
  AOI211_X1 U18242 ( .C1(n15045), .C2(n19203), .A(n15044), .B(n15043), .ZN(
        n15046) );
  OAI211_X1 U18243 ( .C1(n16265), .C2(n15223), .A(n15047), .B(n15046), .ZN(
        P2_U2995) );
  NAND2_X1 U18244 ( .A1(n15048), .A2(n15049), .ZN(n15053) );
  NAND2_X1 U18245 ( .A1(n15051), .A2(n15050), .ZN(n15052) );
  XOR2_X1 U18246 ( .A(n15053), .B(n15052), .Z(n15255) );
  NOR2_X1 U18247 ( .A1(n19818), .A2(n15334), .ZN(n15055) );
  OAI22_X1 U18248 ( .A1(n19212), .A2(n10866), .B1(n16262), .B2(n18967), .ZN(
        n15054) );
  AOI211_X1 U18249 ( .C1(n19207), .C2(n18956), .A(n15055), .B(n15054), .ZN(
        n15058) );
  XOR2_X1 U18250 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B(n15247), .Z(
        n15056) );
  NAND2_X1 U18251 ( .A1(n15056), .A2(n19204), .ZN(n15057) );
  OAI211_X1 U18252 ( .C1(n15255), .C2(n16263), .A(n15058), .B(n15057), .ZN(
        P2_U2997) );
  OAI21_X1 U18253 ( .B1(n15060), .B2(n15059), .A(n15048), .ZN(n15266) );
  OR2_X1 U18254 ( .A1(n15266), .A2(n16263), .ZN(n15068) );
  INV_X1 U18255 ( .A(n15258), .ZN(n18979) );
  INV_X1 U18256 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19816) );
  NOR2_X1 U18257 ( .A1(n19816), .A2(n15334), .ZN(n15061) );
  AOI21_X1 U18258 ( .B1(n19207), .B2(n18979), .A(n15061), .ZN(n15067) );
  AOI21_X1 U18259 ( .B1(n11284), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15062) );
  OR3_X1 U18260 ( .A1(n15247), .A2(n15062), .A3(n16265), .ZN(n15066) );
  INV_X1 U18261 ( .A(n18974), .ZN(n15063) );
  OAI22_X1 U18262 ( .A1(n19212), .A2(n18975), .B1(n16262), .B2(n15063), .ZN(
        n15064) );
  INV_X1 U18263 ( .A(n15064), .ZN(n15065) );
  NAND4_X1 U18264 ( .A1(n15068), .A2(n15067), .A3(n15066), .A4(n15065), .ZN(
        P2_U2998) );
  NAND2_X1 U18265 ( .A1(n15070), .A2(n9916), .ZN(n15071) );
  XNOR2_X1 U18266 ( .A(n15072), .B(n15071), .ZN(n15278) );
  INV_X1 U18267 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15271) );
  XNOR2_X1 U18268 ( .A(n11284), .B(n15271), .ZN(n15276) );
  INV_X1 U18269 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18994) );
  OAI22_X1 U18270 ( .A1(n19212), .A2(n18994), .B1(n16262), .B2(n18988), .ZN(
        n15075) );
  INV_X1 U18271 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n15073) );
  OAI22_X1 U18272 ( .A1(n13644), .A2(n18989), .B1(n15334), .B2(n15073), .ZN(
        n15074) );
  AOI211_X1 U18273 ( .C1(n15276), .C2(n19204), .A(n15075), .B(n15074), .ZN(
        n15076) );
  OAI21_X1 U18274 ( .B1(n15278), .B2(n16263), .A(n15076), .ZN(P2_U2999) );
  NOR2_X1 U18275 ( .A1(n15077), .A2(n16239), .ZN(n15082) );
  INV_X1 U18276 ( .A(n15078), .ZN(n15080) );
  NOR2_X1 U18277 ( .A1(n15080), .A2(n15079), .ZN(n15081) );
  XNOR2_X1 U18278 ( .A(n15082), .B(n15081), .ZN(n15286) );
  INV_X1 U18279 ( .A(n15282), .ZN(n15083) );
  NOR2_X1 U18280 ( .A1(n13644), .A2(n15083), .ZN(n15086) );
  OAI22_X1 U18281 ( .A1(n19212), .A2(n15084), .B1(n10855), .B2(n15334), .ZN(
        n15085) );
  AOI211_X1 U18282 ( .C1(n19203), .C2(n15087), .A(n15086), .B(n15085), .ZN(
        n15091) );
  NAND2_X1 U18283 ( .A1(n15089), .A2(n15279), .ZN(n15283) );
  NAND3_X1 U18284 ( .A1(n15088), .A2(n19204), .A3(n15283), .ZN(n15090) );
  OAI211_X1 U18285 ( .C1(n15286), .C2(n16263), .A(n15091), .B(n15090), .ZN(
        P2_U3001) );
  NAND3_X1 U18286 ( .A1(n15092), .A2(n16252), .A3(n16253), .ZN(n15097) );
  INV_X1 U18287 ( .A(n15093), .ZN(n15094) );
  NOR2_X1 U18288 ( .A1(n15095), .A2(n15094), .ZN(n15096) );
  XNOR2_X1 U18289 ( .A(n15097), .B(n15096), .ZN(n15302) );
  INV_X1 U18290 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15293) );
  NAND2_X1 U18291 ( .A1(n15098), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16249) );
  OR2_X1 U18292 ( .A1(n16249), .A2(n16248), .ZN(n16251) );
  NAND2_X1 U18293 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15290) );
  NOR2_X1 U18294 ( .A1(n16249), .A2(n15290), .ZN(n16242) );
  AOI21_X1 U18295 ( .B1(n15293), .B2(n16251), .A(n16242), .ZN(n15300) );
  OAI22_X1 U18296 ( .A1(n19212), .A2(n15100), .B1(n16262), .B2(n15099), .ZN(
        n15103) );
  INV_X1 U18297 ( .A(n15296), .ZN(n19000) );
  OAI22_X1 U18298 ( .A1(n13644), .A2(n19000), .B1(n15334), .B2(n15101), .ZN(
        n15102) );
  AOI211_X1 U18299 ( .C1(n15300), .C2(n19204), .A(n15103), .B(n15102), .ZN(
        n15104) );
  OAI21_X1 U18300 ( .B1(n15302), .B2(n16263), .A(n15104), .ZN(P2_U3003) );
  NAND2_X1 U18301 ( .A1(n15106), .A2(n15105), .ZN(n15107) );
  XNOR2_X1 U18302 ( .A(n15107), .B(n16326), .ZN(n15330) );
  NOR2_X1 U18303 ( .A1(n15109), .A2(n15108), .ZN(n15113) );
  NAND2_X1 U18304 ( .A1(n15110), .A2(n15111), .ZN(n15112) );
  XOR2_X1 U18305 ( .A(n15113), .B(n15112), .Z(n15327) );
  INV_X1 U18306 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15114) );
  OAI22_X1 U18307 ( .A1(n19212), .A2(n15114), .B1(n16262), .B2(n19018), .ZN(
        n15116) );
  OAI22_X1 U18308 ( .A1(n19021), .A2(n13644), .B1(n15334), .B2(n19803), .ZN(
        n15115) );
  AOI211_X1 U18309 ( .C1(n15327), .C2(n11305), .A(n15116), .B(n15115), .ZN(
        n15117) );
  OAI21_X1 U18310 ( .B1(n16265), .B2(n15330), .A(n15117), .ZN(P2_U3007) );
  XNOR2_X1 U18311 ( .A(n15118), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15341) );
  XOR2_X1 U18312 ( .A(n15119), .B(n15120), .Z(n15339) );
  OAI22_X1 U18313 ( .A1(n19212), .A2(n19041), .B1(n19801), .B2(n18957), .ZN(
        n15121) );
  INV_X1 U18314 ( .A(n15121), .ZN(n15123) );
  NAND2_X1 U18315 ( .A1(n19203), .A2(n19034), .ZN(n15122) );
  OAI211_X1 U18316 ( .C1(n19035), .C2(n13644), .A(n15123), .B(n15122), .ZN(
        n15124) );
  AOI21_X1 U18317 ( .B1(n15339), .B2(n11305), .A(n15124), .ZN(n15125) );
  OAI21_X1 U18318 ( .B1(n15341), .B2(n16265), .A(n15125), .ZN(P2_U3008) );
  NAND2_X1 U18319 ( .A1(n15126), .A2(n19233), .ZN(n15135) );
  OAI21_X1 U18320 ( .B1(n15144), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15127) );
  OAI211_X1 U18321 ( .C1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(n15128), .B(n15127), .ZN(
        n15131) );
  AOI21_X1 U18322 ( .B1(n19228), .B2(n16122), .A(n15129), .ZN(n15130) );
  OAI211_X1 U18323 ( .C1(n16299), .C2(n16124), .A(n15131), .B(n15130), .ZN(
        n15132) );
  AOI21_X1 U18324 ( .B1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15133), .A(
        n15132), .ZN(n15134) );
  OAI211_X1 U18325 ( .C1(n15136), .C2(n19225), .A(n15135), .B(n15134), .ZN(
        P2_U3017) );
  NOR3_X1 U18326 ( .A1(n15138), .A2(n15137), .A3(n16318), .ZN(n15147) );
  NOR2_X1 U18327 ( .A1(n16133), .A2(n16299), .ZN(n15139) );
  AOI211_X1 U18328 ( .C1(n15141), .C2(n19228), .A(n15140), .B(n15139), .ZN(
        n15142) );
  OAI211_X1 U18329 ( .C1(n15145), .C2(n15144), .A(n15143), .B(n15142), .ZN(
        n15146) );
  NOR2_X1 U18330 ( .A1(n15147), .A2(n15146), .ZN(n15148) );
  OAI21_X1 U18331 ( .B1(n15149), .B2(n19225), .A(n15148), .ZN(P2_U3019) );
  OAI21_X1 U18332 ( .B1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n15150), .ZN(n15151) );
  OAI22_X1 U18333 ( .A1(n15154), .A2(n15153), .B1(n15152), .B2(n15151), .ZN(
        n15157) );
  AOI22_X1 U18334 ( .A1(n16147), .A2(n19220), .B1(n19030), .B2(
        P2_REIP_REG_26__SCAN_IN), .ZN(n15155) );
  OAI21_X1 U18335 ( .B1(n15346), .B2(n16145), .A(n15155), .ZN(n15156) );
  AOI211_X1 U18336 ( .C1(n15158), .C2(n19233), .A(n15157), .B(n15156), .ZN(
        n15159) );
  OAI21_X1 U18337 ( .B1(n15160), .B2(n19225), .A(n15159), .ZN(P2_U3020) );
  NAND2_X1 U18338 ( .A1(n9851), .A2(n15162), .ZN(n15163) );
  XNOR2_X1 U18339 ( .A(n15161), .B(n15163), .ZN(n16205) );
  OR2_X1 U18340 ( .A1(n15007), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15164) );
  NAND2_X1 U18341 ( .A1(n13951), .A2(n15164), .ZN(n16209) );
  NOR2_X1 U18342 ( .A1(n11240), .A2(n15334), .ZN(n15165) );
  AOI221_X1 U18343 ( .B1(n15168), .B2(n15167), .C1(n15166), .C2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(n15165), .ZN(n15171) );
  INV_X1 U18344 ( .A(n16169), .ZN(n16206) );
  AOI22_X1 U18345 ( .A1(n16206), .A2(n19220), .B1(n19228), .B2(n15169), .ZN(
        n15170) );
  OAI211_X1 U18346 ( .C1(n16209), .C2(n16318), .A(n15171), .B(n15170), .ZN(
        n15172) );
  AOI21_X1 U18347 ( .B1(n16323), .B2(n16205), .A(n15172), .ZN(n15173) );
  INV_X1 U18348 ( .A(n15173), .ZN(P2_U3022) );
  AND3_X1 U18349 ( .A1(n15016), .A2(n15174), .A3(n16323), .ZN(n15183) );
  AOI211_X1 U18350 ( .C1(n15180), .C2(n15192), .A(n15175), .B(n15193), .ZN(
        n15182) );
  NOR2_X1 U18351 ( .A1(n16179), .A2(n16299), .ZN(n15178) );
  OAI22_X1 U18352 ( .A1(n15346), .A2(n15176), .B1(n19825), .B2(n18957), .ZN(
        n15177) );
  NOR2_X1 U18353 ( .A1(n15178), .A2(n15177), .ZN(n15179) );
  OAI21_X1 U18354 ( .B1(n15203), .B2(n15180), .A(n15179), .ZN(n15181) );
  NOR3_X1 U18355 ( .A1(n15183), .A2(n15182), .A3(n15181), .ZN(n15184) );
  OAI21_X1 U18356 ( .B1(n15185), .B2(n16318), .A(n15184), .ZN(P2_U3023) );
  NAND2_X1 U18357 ( .A1(n15188), .A2(n15187), .ZN(n15189) );
  XNOR2_X1 U18358 ( .A(n15186), .B(n15189), .ZN(n16216) );
  INV_X1 U18359 ( .A(n16216), .ZN(n15201) );
  NAND2_X1 U18360 ( .A1(n15190), .A2(n15192), .ZN(n16214) );
  NAND3_X1 U18361 ( .A1(n16215), .A2(n19233), .A3(n16214), .ZN(n15200) );
  NAND2_X1 U18362 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19030), .ZN(n15191) );
  OAI221_X1 U18363 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n15193), 
        .C1(n15192), .C2(n15203), .A(n15191), .ZN(n15198) );
  OAI21_X1 U18364 ( .B1(n15195), .B2(n15194), .A(n14956), .ZN(n15710) );
  OAI22_X1 U18365 ( .A1(n16299), .A2(n15196), .B1(n15346), .B2(n15710), .ZN(
        n15197) );
  NOR2_X1 U18366 ( .A1(n15198), .A2(n15197), .ZN(n15199) );
  OAI211_X1 U18367 ( .C1(n15201), .C2(n19225), .A(n15200), .B(n15199), .ZN(
        P2_U3024) );
  NAND2_X1 U18368 ( .A1(n15202), .A2(n16323), .ZN(n15214) );
  INV_X1 U18369 ( .A(n15203), .ZN(n15212) );
  INV_X1 U18370 ( .A(n15204), .ZN(n15205) );
  AOI22_X1 U18371 ( .A1(n19220), .A2(n15205), .B1(P2_REIP_REG_21__SCAN_IN), 
        .B2(n19030), .ZN(n15206) );
  OAI21_X1 U18372 ( .B1(n15346), .B2(n15207), .A(n15206), .ZN(n15211) );
  INV_X1 U18373 ( .A(n15220), .ZN(n15208) );
  NOR3_X1 U18374 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n15209), .A3(
        n15208), .ZN(n15210) );
  AOI211_X1 U18375 ( .C1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15212), .A(
        n15211), .B(n15210), .ZN(n15213) );
  OAI211_X1 U18376 ( .C1(n15215), .C2(n16318), .A(n15214), .B(n15213), .ZN(
        P2_U3025) );
  NAND2_X1 U18377 ( .A1(n15216), .A2(n16323), .ZN(n15222) );
  INV_X1 U18378 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21008) );
  OAI22_X1 U18379 ( .A1(n15346), .A2(n18943), .B1(n10873), .B2(n18957), .ZN(
        n15217) );
  AOI21_X1 U18380 ( .B1(n19220), .B2(n18938), .A(n15217), .ZN(n15218) );
  OAI21_X1 U18381 ( .B1(n15231), .B2(n21008), .A(n15218), .ZN(n15219) );
  AOI21_X1 U18382 ( .B1(n15220), .B2(n21008), .A(n15219), .ZN(n15221) );
  OAI211_X1 U18383 ( .C1(n15223), .C2(n16318), .A(n15222), .B(n15221), .ZN(
        P2_U3027) );
  AOI21_X1 U18384 ( .B1(n15247), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15224) );
  OR2_X1 U18385 ( .A1(n15225), .A2(n15224), .ZN(n16224) );
  NAND2_X1 U18386 ( .A1(n15227), .A2(n15226), .ZN(n15228) );
  XNOR2_X1 U18387 ( .A(n15229), .B(n15228), .ZN(n16225) );
  OR2_X1 U18388 ( .A1(n16225), .A2(n19225), .ZN(n15240) );
  NAND2_X1 U18389 ( .A1(P2_REIP_REG_18__SCAN_IN), .A2(n19030), .ZN(n15230) );
  OAI221_X1 U18390 ( .B1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n15233), 
        .C1(n15232), .C2(n15231), .A(n15230), .ZN(n15238) );
  NAND2_X1 U18391 ( .A1(n15234), .A2(n13888), .ZN(n15236) );
  INV_X1 U18392 ( .A(n14970), .ZN(n15235) );
  NAND2_X1 U18393 ( .A1(n15236), .A2(n15235), .ZN(n16200) );
  OAI22_X1 U18394 ( .A1(n16299), .A2(n18949), .B1(n15346), .B2(n16200), .ZN(
        n15237) );
  NOR2_X1 U18395 ( .A1(n15238), .A2(n15237), .ZN(n15239) );
  OAI211_X1 U18396 ( .C1(n16224), .C2(n16318), .A(n15240), .B(n15239), .ZN(
        P2_U3028) );
  OAI22_X1 U18397 ( .A1(n15346), .A2(n18971), .B1(n19818), .B2(n18957), .ZN(
        n15244) );
  AOI22_X1 U18398 ( .A1(n15247), .A2(n19233), .B1(n15241), .B2(n15272), .ZN(
        n15242) );
  NOR2_X1 U18399 ( .A1(n15242), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15243) );
  AOI211_X1 U18400 ( .C1(n18956), .C2(n19220), .A(n15244), .B(n15243), .ZN(
        n15254) );
  NOR2_X1 U18401 ( .A1(n19233), .A2(n15245), .ZN(n15246) );
  OR2_X1 U18402 ( .A1(n15247), .A2(n15246), .ZN(n15250) );
  NOR2_X1 U18403 ( .A1(n19213), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15248) );
  NOR2_X1 U18404 ( .A1(n15270), .A2(n15248), .ZN(n15249) );
  NAND2_X1 U18405 ( .A1(n15250), .A2(n15249), .ZN(n15264) );
  AOI21_X1 U18406 ( .B1(n10865), .B2(n16294), .A(n15264), .ZN(n15252) );
  OR2_X1 U18407 ( .A1(n15252), .A2(n15251), .ZN(n15253) );
  OAI211_X1 U18408 ( .C1(n15255), .C2(n19225), .A(n15254), .B(n15253), .ZN(
        P2_U3029) );
  AOI21_X1 U18409 ( .B1(n11284), .B2(n19233), .A(n15272), .ZN(n15262) );
  NAND2_X1 U18410 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n10865), .ZN(
        n15261) );
  AOI21_X1 U18411 ( .B1(n15256), .B2(n15257), .A(n13886), .ZN(n19079) );
  OAI22_X1 U18412 ( .A1(n16299), .A2(n15258), .B1(n15334), .B2(n19816), .ZN(
        n15259) );
  AOI21_X1 U18413 ( .B1(n19079), .B2(n19228), .A(n15259), .ZN(n15260) );
  OAI21_X1 U18414 ( .B1(n15262), .B2(n15261), .A(n15260), .ZN(n15263) );
  AOI21_X1 U18415 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15264), .A(
        n15263), .ZN(n15265) );
  OAI21_X1 U18416 ( .B1(n15266), .B2(n19225), .A(n15265), .ZN(P2_U3030) );
  OAI21_X1 U18417 ( .B1(n14752), .B2(n15267), .A(n15256), .ZN(n19086) );
  NOR2_X1 U18418 ( .A1(n16299), .A2(n18989), .ZN(n15269) );
  NOR2_X1 U18419 ( .A1(n15073), .A2(n15334), .ZN(n15268) );
  AOI211_X1 U18420 ( .C1(n15270), .C2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15269), .B(n15268), .ZN(n15274) );
  NAND2_X1 U18421 ( .A1(n15272), .A2(n15271), .ZN(n15273) );
  OAI211_X1 U18422 ( .C1(n19086), .C2(n15346), .A(n15274), .B(n15273), .ZN(
        n15275) );
  AOI21_X1 U18423 ( .B1(n15276), .B2(n19233), .A(n15275), .ZN(n15277) );
  OAI21_X1 U18424 ( .B1(n15278), .B2(n19225), .A(n15277), .ZN(P2_U3031) );
  OAI22_X1 U18425 ( .A1(n15346), .A2(n19092), .B1(n10855), .B2(n18957), .ZN(
        n15281) );
  NOR3_X1 U18426 ( .A1(n15289), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        n16295), .ZN(n16296) );
  AOI211_X1 U18427 ( .C1(n16295), .C2(n16294), .A(n16296), .B(n16293), .ZN(
        n16284) );
  OR3_X1 U18428 ( .A1(n16295), .A2(n15289), .A3(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16283) );
  OAI22_X1 U18429 ( .A1(n16284), .A2(n15279), .B1(n16305), .B2(n16283), .ZN(
        n15280) );
  AOI211_X1 U18430 ( .C1(n15282), .C2(n19220), .A(n15281), .B(n15280), .ZN(
        n15285) );
  NAND3_X1 U18431 ( .A1(n15088), .A2(n19233), .A3(n15283), .ZN(n15284) );
  OAI211_X1 U18432 ( .C1(n15286), .C2(n19225), .A(n15285), .B(n15284), .ZN(
        P2_U3033) );
  OR2_X1 U18433 ( .A1(n15287), .A2(n14791), .ZN(n15288) );
  NAND2_X1 U18434 ( .A1(n15288), .A2(n14780), .ZN(n19098) );
  AOI211_X1 U18435 ( .C1(n16248), .C2(n15293), .A(n15308), .B(n15289), .ZN(
        n15291) );
  NAND2_X1 U18436 ( .A1(n15291), .A2(n15290), .ZN(n15298) );
  NOR2_X1 U18437 ( .A1(n15101), .A2(n15334), .ZN(n15295) );
  OAI21_X1 U18438 ( .B1(n16293), .B2(n15308), .A(n15292), .ZN(n16309) );
  NOR2_X1 U18439 ( .A1(n15293), .A2(n16309), .ZN(n15294) );
  AOI211_X1 U18440 ( .C1(n19220), .C2(n15296), .A(n15295), .B(n15294), .ZN(
        n15297) );
  OAI211_X1 U18441 ( .C1(n15346), .C2(n19098), .A(n15298), .B(n15297), .ZN(
        n15299) );
  AOI21_X1 U18442 ( .B1(n15300), .B2(n19233), .A(n15299), .ZN(n15301) );
  OAI21_X1 U18443 ( .B1(n15302), .B2(n19225), .A(n15301), .ZN(P2_U3035) );
  OAI21_X1 U18444 ( .B1(n15098), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n16249), .ZN(n16266) );
  INV_X1 U18445 ( .A(n16252), .ZN(n15306) );
  AND2_X1 U18446 ( .A1(n16252), .A2(n15304), .ZN(n15305) );
  OAI22_X1 U18447 ( .A1(n15303), .A2(n15306), .B1(n9826), .B2(n15305), .ZN(
        n16264) );
  INV_X1 U18448 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n19807) );
  NOR2_X1 U18449 ( .A1(n19807), .A2(n18957), .ZN(n15307) );
  AOI221_X1 U18450 ( .B1(n16307), .B2(n15308), .C1(n16293), .C2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n15307), .ZN(n15313) );
  OAI21_X1 U18451 ( .B1(n14809), .B2(n15310), .A(n15309), .ZN(n19105) );
  INV_X1 U18452 ( .A(n19105), .ZN(n15311) );
  INV_X1 U18453 ( .A(n19011), .ZN(n16268) );
  AOI22_X1 U18454 ( .A1(n15311), .A2(n19228), .B1(n19220), .B2(n16268), .ZN(
        n15312) );
  OAI211_X1 U18455 ( .C1(n16264), .C2(n19225), .A(n15313), .B(n15312), .ZN(
        n15314) );
  INV_X1 U18456 ( .A(n15314), .ZN(n15315) );
  OAI21_X1 U18457 ( .B1(n16318), .B2(n16266), .A(n15315), .ZN(P2_U3037) );
  NOR2_X1 U18458 ( .A1(n15317), .A2(n15316), .ZN(n16325) );
  INV_X1 U18459 ( .A(n15318), .ZN(n15319) );
  OAI21_X1 U18460 ( .B1(n15321), .B2(n15320), .A(n15319), .ZN(n16320) );
  AOI22_X1 U18461 ( .A1(n16320), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B1(
        n19030), .B2(P2_REIP_REG_7__SCAN_IN), .ZN(n15322) );
  OAI21_X1 U18462 ( .B1(n19021), .B2(n16299), .A(n15322), .ZN(n15326) );
  OAI21_X1 U18463 ( .B1(n15324), .B2(n15323), .A(n14808), .ZN(n19108) );
  NOR2_X1 U18464 ( .A1(n19108), .A2(n15346), .ZN(n15325) );
  AOI211_X1 U18465 ( .C1(n16325), .C2(n16326), .A(n15326), .B(n15325), .ZN(
        n15329) );
  NAND2_X1 U18466 ( .A1(n15327), .A2(n16323), .ZN(n15328) );
  OAI211_X1 U18467 ( .C1(n15330), .C2(n16318), .A(n15329), .B(n15328), .ZN(
        P2_U3039) );
  XNOR2_X1 U18468 ( .A(n9868), .B(n15331), .ZN(n19109) );
  NAND4_X1 U18469 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n15332), .A4(n20863), .ZN(
        n15333) );
  OAI21_X1 U18470 ( .B1(n15334), .B2(n19801), .A(n15333), .ZN(n15336) );
  NOR2_X1 U18471 ( .A1(n19035), .A2(n16299), .ZN(n15335) );
  AOI211_X1 U18472 ( .C1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n16320), .A(
        n15336), .B(n15335), .ZN(n15337) );
  OAI21_X1 U18473 ( .B1(n19109), .B2(n15346), .A(n15337), .ZN(n15338) );
  AOI21_X1 U18474 ( .B1(n15339), .B2(n16323), .A(n15338), .ZN(n15340) );
  OAI21_X1 U18475 ( .B1(n15341), .B2(n16318), .A(n15340), .ZN(P2_U3040) );
  AOI22_X1 U18476 ( .A1(n16323), .A2(n15343), .B1(n19233), .B2(n15342), .ZN(
        n15351) );
  INV_X1 U18477 ( .A(n19875), .ZN(n15345) );
  OAI21_X1 U18478 ( .B1(n15346), .B2(n15345), .A(n15344), .ZN(n15347) );
  AOI21_X1 U18479 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n19216), .A(
        n15347), .ZN(n15350) );
  NAND2_X1 U18480 ( .A1(n19220), .A2(n9791), .ZN(n15349) );
  OAI211_X1 U18481 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n16294), .B(n19217), .ZN(n15348) );
  NAND4_X1 U18482 ( .A1(n15351), .A2(n15350), .A3(n15349), .A4(n15348), .ZN(
        P2_U3045) );
  INV_X1 U18483 ( .A(n16368), .ZN(n15416) );
  INV_X1 U18484 ( .A(n19764), .ZN(n19851) );
  INV_X1 U18485 ( .A(n15400), .ZN(n15377) );
  INV_X1 U18486 ( .A(n11254), .ZN(n15353) );
  NAND2_X1 U18487 ( .A1(n15353), .A2(n15352), .ZN(n15371) );
  MUX2_X1 U18488 ( .A(n15371), .B(n11010), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n15354) );
  AOI21_X1 U18489 ( .B1(n13216), .B2(n15377), .A(n15354), .ZN(n16332) );
  OAI22_X1 U18490 ( .A1(n19032), .A2(n13219), .B1(n19072), .B2(n14704), .ZN(
        n15367) );
  OAI222_X1 U18491 ( .A1(n15416), .A2(n15355), .B1(n19851), .B2(n16332), .C1(
        n10329), .C2(n15367), .ZN(n15365) );
  NAND3_X1 U18492 ( .A1(n15358), .A2(n15357), .A3(n15356), .ZN(n15362) );
  NAND2_X1 U18493 ( .A1(n16348), .A2(n15359), .ZN(n15360) );
  NOR2_X1 U18494 ( .A1(n19138), .A2(n15360), .ZN(n15361) );
  NOR2_X1 U18495 ( .A1(n18894), .A2(n15363), .ZN(n16377) );
  AOI22_X1 U18496 ( .A1(n16377), .A2(P2_FLUSH_REG_SCAN_IN), .B1(
        P2_STATE2_REG_3__SCAN_IN), .B2(n18894), .ZN(n15364) );
  OAI21_X1 U18497 ( .B1(n16354), .B2(n16375), .A(n15364), .ZN(n15506) );
  MUX2_X1 U18498 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n15365), .S(
        n15506), .Z(P2_U3601) );
  INV_X1 U18499 ( .A(n15367), .ZN(n15368) );
  NOR2_X1 U18500 ( .A1(n15368), .A2(n10329), .ZN(n15396) );
  INV_X1 U18501 ( .A(n15396), .ZN(n15375) );
  OAI21_X1 U18502 ( .B1(n19032), .B2(n15370), .A(n15369), .ZN(n15395) );
  INV_X1 U18503 ( .A(n11010), .ZN(n15373) );
  OAI21_X1 U18504 ( .B1(n10387), .B2(n10385), .A(n15371), .ZN(n15372) );
  OAI21_X1 U18505 ( .B1(n15373), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n15372), .ZN(n15374) );
  AOI21_X1 U18506 ( .B1(n9792), .B2(n15377), .A(n15374), .ZN(n16335) );
  OAI222_X1 U18507 ( .A1(n15416), .A2(n19871), .B1(n15375), .B2(n15395), .C1(
        n19851), .C2(n16335), .ZN(n15376) );
  INV_X1 U18508 ( .A(n15506), .ZN(n15398) );
  MUX2_X1 U18509 ( .A(n15376), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n15398), .Z(P2_U3600) );
  NAND2_X1 U18510 ( .A1(n13265), .A2(n15377), .ZN(n15393) );
  NOR2_X1 U18511 ( .A1(n15379), .A2(n15378), .ZN(n15404) );
  INV_X1 U18512 ( .A(n10388), .ZN(n15380) );
  NAND2_X1 U18513 ( .A1(n15380), .A2(n9780), .ZN(n15401) );
  AND2_X1 U18514 ( .A1(n15381), .A2(n15401), .ZN(n15390) );
  INV_X1 U18515 ( .A(n15382), .ZN(n15383) );
  OAI21_X1 U18516 ( .B1(n16336), .B2(n15384), .A(n15383), .ZN(n15385) );
  NAND2_X1 U18517 ( .A1(n11010), .A2(n15385), .ZN(n15389) );
  NAND2_X1 U18518 ( .A1(n10297), .A2(n11001), .ZN(n15386) );
  NAND2_X1 U18519 ( .A1(n15386), .A2(n15381), .ZN(n15406) );
  INV_X1 U18520 ( .A(n15406), .ZN(n15387) );
  NAND2_X1 U18521 ( .A1(n15387), .A2(n15401), .ZN(n15388) );
  OAI211_X1 U18522 ( .C1(n15404), .C2(n15390), .A(n15389), .B(n15388), .ZN(
        n15391) );
  INV_X1 U18523 ( .A(n15391), .ZN(n15392) );
  NAND2_X1 U18524 ( .A1(n15393), .A2(n15392), .ZN(n16337) );
  AOI222_X1 U18525 ( .A1(n16337), .A2(n19764), .B1(n15396), .B2(n15395), .C1(
        n16368), .C2(n15394), .ZN(n15399) );
  NAND2_X1 U18526 ( .A1(n15398), .A2(n16336), .ZN(n15397) );
  OAI21_X1 U18527 ( .B1(n15399), .B2(n15398), .A(n15397), .ZN(P2_U3599) );
  OR2_X1 U18528 ( .A1(n13617), .A2(n15400), .ZN(n15414) );
  XNOR2_X1 U18529 ( .A(n15401), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n15403) );
  OAI21_X1 U18530 ( .B1(n15404), .B2(n15403), .A(n15402), .ZN(n15412) );
  NAND2_X1 U18531 ( .A1(n16336), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15407) );
  NAND2_X1 U18532 ( .A1(n11010), .A2(n15407), .ZN(n15405) );
  NAND2_X1 U18533 ( .A1(n15406), .A2(n15405), .ZN(n15410) );
  AND2_X1 U18534 ( .A1(n11010), .A2(n9776), .ZN(n15409) );
  MUX2_X1 U18535 ( .A(n15410), .B(n15409), .S(n15408), .Z(n15411) );
  NOR2_X1 U18536 ( .A1(n15412), .A2(n15411), .ZN(n15413) );
  NAND2_X1 U18537 ( .A1(n15414), .A2(n15413), .ZN(n16340) );
  INV_X1 U18538 ( .A(n16340), .ZN(n15415) );
  OAI22_X1 U18539 ( .A1(n19854), .A2(n15416), .B1(n15415), .B2(n19851), .ZN(
        n15417) );
  MUX2_X1 U18540 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n15417), .S(
        n15506), .Z(P2_U3596) );
  INV_X1 U18541 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16639) );
  INV_X1 U18542 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16661) );
  INV_X1 U18543 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16681) );
  INV_X1 U18544 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17037) );
  INV_X1 U18545 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n16715) );
  INV_X1 U18546 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16796) );
  INV_X1 U18547 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n21019) );
  NAND3_X1 U18548 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17235) );
  NAND4_X1 U18549 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .A3(P3_EBX_REG_4__SCAN_IN), .A4(P3_EBX_REG_3__SCAN_IN), .ZN(n15420) );
  NOR2_X1 U18550 ( .A1(n17235), .A2(n15420), .ZN(n17236) );
  NOR3_X2 U18551 ( .A1(n16715), .A2(n17062), .A3(n17065), .ZN(n17025) );
  NAND2_X1 U18552 ( .A1(n9796), .A2(n17025), .ZN(n17038) );
  NAND2_X1 U18553 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17010), .ZN(n17005) );
  NOR2_X2 U18554 ( .A1(n16681), .A2(n17005), .ZN(n17009) );
  NAND2_X1 U18555 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17009), .ZN(n16996) );
  NOR2_X2 U18556 ( .A1(n16661), .A2(n16996), .ZN(n16999) );
  NAND2_X1 U18557 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16999), .ZN(n16987) );
  NOR2_X2 U18558 ( .A1(n16639), .A2(n16987), .ZN(n16990) );
  NAND2_X1 U18559 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16990), .ZN(n16986) );
  INV_X1 U18560 ( .A(n16986), .ZN(n15497) );
  INV_X1 U18561 ( .A(n9796), .ZN(n17247) );
  INV_X2 U18562 ( .A(n17254), .ZN(n17251) );
  AOI21_X1 U18563 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n17251), .A(n16990), .ZN(
        n15496) );
  AOI22_X1 U18564 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(n9763), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15424) );
  AOI22_X1 U18565 ( .A1(n9758), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15423) );
  AOI22_X1 U18566 ( .A1(n17209), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15422) );
  AOI22_X1 U18567 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15421) );
  NAND4_X1 U18568 ( .A1(n15424), .A2(n15423), .A3(n15422), .A4(n15421), .ZN(
        n15430) );
  AOI22_X1 U18569 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15428) );
  AOI22_X1 U18570 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n15550), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15427) );
  AOI22_X1 U18571 ( .A1(n17207), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15426) );
  AOI22_X1 U18572 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15425) );
  NAND4_X1 U18573 ( .A1(n15428), .A2(n15427), .A3(n15426), .A4(n15425), .ZN(
        n15429) );
  NOR2_X1 U18574 ( .A1(n15430), .A2(n15429), .ZN(n16988) );
  AOI22_X1 U18575 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15434) );
  AOI22_X1 U18576 ( .A1(n9758), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15433) );
  AOI22_X1 U18577 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15432) );
  AOI22_X1 U18578 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15431) );
  NAND4_X1 U18579 ( .A1(n15434), .A2(n15433), .A3(n15432), .A4(n15431), .ZN(
        n15441) );
  AOI22_X1 U18580 ( .A1(n9763), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15550), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15439) );
  AOI22_X1 U18581 ( .A1(n17207), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15438) );
  AOI22_X1 U18582 ( .A1(n17209), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15437) );
  AOI22_X1 U18583 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17205), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15436) );
  NAND4_X1 U18584 ( .A1(n15439), .A2(n15438), .A3(n15437), .A4(n15436), .ZN(
        n15440) );
  NOR2_X1 U18585 ( .A1(n15441), .A2(n15440), .ZN(n16997) );
  AOI22_X1 U18586 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15445) );
  AOI22_X1 U18587 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15444) );
  AOI22_X1 U18588 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17205), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15443) );
  AOI22_X1 U18589 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15442) );
  NAND4_X1 U18590 ( .A1(n15445), .A2(n15444), .A3(n15443), .A4(n15442), .ZN(
        n15451) );
  AOI22_X1 U18591 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15449) );
  AOI22_X1 U18592 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15448) );
  AOI22_X1 U18593 ( .A1(n17209), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n15550), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15447) );
  AOI22_X1 U18594 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n15446) );
  NAND4_X1 U18595 ( .A1(n15449), .A2(n15448), .A3(n15447), .A4(n15446), .ZN(
        n15450) );
  NOR2_X1 U18596 ( .A1(n15451), .A2(n15450), .ZN(n17007) );
  AOI22_X1 U18597 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15455) );
  AOI22_X1 U18598 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17205), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15454) );
  AOI22_X1 U18599 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15453) );
  AOI22_X1 U18600 ( .A1(n17209), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15452) );
  NAND4_X1 U18601 ( .A1(n15455), .A2(n15454), .A3(n15453), .A4(n15452), .ZN(
        n15461) );
  AOI22_X1 U18602 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15459) );
  AOI22_X1 U18603 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n15458) );
  AOI22_X1 U18604 ( .A1(n17207), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17224), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15457) );
  AOI22_X1 U18605 ( .A1(n9763), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n15550), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15456) );
  NAND4_X1 U18606 ( .A1(n15459), .A2(n15458), .A3(n15457), .A4(n15456), .ZN(
        n15460) );
  NOR2_X1 U18607 ( .A1(n15461), .A2(n15460), .ZN(n17006) );
  NOR2_X1 U18608 ( .A1(n17007), .A2(n17006), .ZN(n17002) );
  AOI22_X1 U18609 ( .A1(n17208), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n15550), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n15472) );
  AOI22_X1 U18610 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n15471) );
  AOI22_X1 U18611 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15462) );
  OAI21_X1 U18612 ( .B1(n15474), .B2(n18230), .A(n15462), .ZN(n15469) );
  AOI22_X1 U18613 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17205), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n15467) );
  AOI22_X1 U18614 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15466) );
  AOI22_X1 U18615 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n15465) );
  AOI22_X1 U18616 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15464) );
  NAND4_X1 U18617 ( .A1(n15467), .A2(n15466), .A3(n15465), .A4(n15464), .ZN(
        n15468) );
  AOI211_X1 U18618 ( .C1(n17214), .C2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n15469), .B(n15468), .ZN(n15470) );
  NAND3_X1 U18619 ( .A1(n15472), .A2(n15471), .A3(n15470), .ZN(n17001) );
  NAND2_X1 U18620 ( .A1(n17002), .A2(n17001), .ZN(n17000) );
  NOR2_X1 U18621 ( .A1(n16997), .A2(n17000), .ZN(n16993) );
  AOI22_X1 U18622 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9758), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15483) );
  AOI22_X1 U18623 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15482) );
  INV_X1 U18624 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n20907) );
  AOI22_X1 U18625 ( .A1(n9763), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15473) );
  OAI21_X1 U18626 ( .B1(n15474), .B2(n20907), .A(n15473), .ZN(n15480) );
  AOI22_X1 U18627 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15478) );
  AOI22_X1 U18628 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15477) );
  AOI22_X1 U18629 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n15550), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15476) );
  AOI22_X1 U18630 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15475) );
  NAND4_X1 U18631 ( .A1(n15478), .A2(n15477), .A3(n15476), .A4(n15475), .ZN(
        n15479) );
  AOI211_X1 U18632 ( .C1(n17176), .C2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A(
        n15480), .B(n15479), .ZN(n15481) );
  NAND3_X1 U18633 ( .A1(n15483), .A2(n15482), .A3(n15481), .ZN(n16992) );
  NAND2_X1 U18634 ( .A1(n16993), .A2(n16992), .ZN(n16991) );
  NOR2_X1 U18635 ( .A1(n16988), .A2(n16991), .ZN(n15495) );
  AOI22_X1 U18636 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n15550), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15493) );
  AOI22_X1 U18637 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17224), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15492) );
  AOI22_X1 U18638 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n15559), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15484) );
  OAI21_X1 U18639 ( .B1(n15594), .B2(n20954), .A(n15484), .ZN(n15490) );
  AOI22_X1 U18640 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17205), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15488) );
  AOI22_X1 U18641 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15487) );
  AOI22_X1 U18642 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n15600), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15486) );
  AOI22_X1 U18643 ( .A1(n9763), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15485) );
  NAND4_X1 U18644 ( .A1(n15488), .A2(n15487), .A3(n15486), .A4(n15485), .ZN(
        n15489) );
  AOI211_X1 U18645 ( .C1(n17173), .C2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n15490), .B(n15489), .ZN(n15491) );
  NAND3_X1 U18646 ( .A1(n15493), .A2(n15492), .A3(n15491), .ZN(n15494) );
  NAND2_X1 U18647 ( .A1(n15495), .A2(n15494), .ZN(n16983) );
  OAI21_X1 U18648 ( .B1(n15495), .B2(n15494), .A(n16983), .ZN(n17280) );
  OAI22_X1 U18649 ( .A1(n15497), .A2(n15496), .B1(n17251), .B2(n17280), .ZN(
        P3_U2675) );
  NAND2_X1 U18650 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18445) );
  AOI221_X1 U18651 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18445), .C1(n15499), 
        .C2(n18445), .A(n15498), .ZN(n18215) );
  NOR2_X1 U18652 ( .A1(n15500), .A2(n18699), .ZN(n15501) );
  OAI21_X1 U18653 ( .B1(n15501), .B2(n18470), .A(n18216), .ZN(n18213) );
  AOI22_X1 U18654 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18215), .B1(
        n18213), .B2(n18704), .ZN(P3_U2865) );
  NOR4_X1 U18655 ( .A1(n15502), .A2(n16346), .A3(n11014), .A4(n19851), .ZN(
        n15503) );
  NAND2_X1 U18656 ( .A1(n15506), .A2(n15503), .ZN(n15504) );
  OAI21_X1 U18657 ( .B1(n15506), .B2(n15505), .A(n15504), .ZN(P2_U3595) );
  AOI22_X1 U18658 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n15550), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15516) );
  AOI22_X1 U18659 ( .A1(n17208), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15515) );
  INV_X1 U18660 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18264) );
  AOI22_X1 U18661 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15507) );
  OAI21_X1 U18662 ( .B1(n12917), .B2(n18264), .A(n15507), .ZN(n15513) );
  AOI22_X1 U18663 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n15511) );
  AOI22_X1 U18664 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15510) );
  AOI22_X1 U18665 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15509) );
  AOI22_X1 U18666 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15508) );
  NAND4_X1 U18667 ( .A1(n15511), .A2(n15510), .A3(n15509), .A4(n15508), .ZN(
        n15512) );
  AOI211_X1 U18668 ( .C1(n17213), .C2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A(
        n15513), .B(n15512), .ZN(n15514) );
  AOI22_X1 U18669 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17205), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15520) );
  AOI22_X1 U18670 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15519) );
  AOI22_X1 U18671 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15518) );
  AOI22_X1 U18672 ( .A1(n9758), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15517) );
  NAND4_X1 U18673 ( .A1(n15520), .A2(n15519), .A3(n15518), .A4(n15517), .ZN(
        n15526) );
  AOI22_X1 U18674 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15524) );
  AOI22_X1 U18675 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15523) );
  AOI22_X1 U18676 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n15600), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15522) );
  AOI22_X1 U18677 ( .A1(n17209), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15521) );
  NAND4_X1 U18678 ( .A1(n15524), .A2(n15523), .A3(n15522), .A4(n15521), .ZN(
        n15525) );
  AOI22_X1 U18679 ( .A1(n15593), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17205), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15530) );
  AOI22_X1 U18680 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n15553), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15529) );
  AOI22_X1 U18681 ( .A1(n17209), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n15600), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15528) );
  AOI22_X1 U18682 ( .A1(n9758), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15527) );
  NAND4_X1 U18683 ( .A1(n15530), .A2(n15529), .A3(n15528), .A4(n15527), .ZN(
        n15536) );
  AOI22_X1 U18684 ( .A1(n17208), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15534) );
  AOI22_X1 U18685 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n15552), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15533) );
  AOI22_X1 U18686 ( .A1(n15435), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15532) );
  AOI22_X1 U18687 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15531) );
  NAND4_X1 U18688 ( .A1(n15534), .A2(n15533), .A3(n15532), .A4(n15531), .ZN(
        n15535) );
  AOI22_X1 U18689 ( .A1(n15552), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n15551), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15542) );
  AOI22_X1 U18690 ( .A1(n15538), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n15537), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n15541) );
  AOI22_X1 U18691 ( .A1(n15593), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n15559), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15540) );
  AOI22_X1 U18692 ( .A1(n15553), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n15595), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15539) );
  NAND4_X1 U18693 ( .A1(n15542), .A2(n15541), .A3(n15540), .A4(n15539), .ZN(
        n15543) );
  NOR2_X1 U18694 ( .A1(n15543), .A2(n10124), .ZN(n15549) );
  AOI22_X1 U18695 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15544) );
  AOI22_X1 U18696 ( .A1(n15435), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n15600), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15548) );
  AOI22_X1 U18697 ( .A1(n15554), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n15560), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15545) );
  OAI21_X1 U18698 ( .B1(n12917), .B2(n18230), .A(n15545), .ZN(n15546) );
  INV_X1 U18699 ( .A(n15546), .ZN(n15547) );
  AOI22_X1 U18700 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15550), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15569) );
  AOI22_X1 U18701 ( .A1(n15435), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15568) );
  AOI22_X1 U18702 ( .A1(n15601), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n15593), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15558) );
  AOI22_X1 U18703 ( .A1(n15552), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15551), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15557) );
  AOI22_X1 U18704 ( .A1(n15554), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n15553), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15556) );
  AOI22_X1 U18705 ( .A1(n15595), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n15600), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15555) );
  NAND4_X1 U18706 ( .A1(n15558), .A2(n15557), .A3(n15556), .A4(n15555), .ZN(
        n15566) );
  INV_X1 U18707 ( .A(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n20891) );
  AOI22_X1 U18708 ( .A1(n15560), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n15559), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15561) );
  OAI21_X1 U18709 ( .B1(n15562), .B2(n20891), .A(n15561), .ZN(n15564) );
  AND2_X1 U18710 ( .A1(n15463), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n15563) );
  NAND3_X1 U18711 ( .A1(n15569), .A2(n15568), .A3(n15567), .ZN(n15658) );
  NAND2_X1 U18712 ( .A1(n17398), .A2(n15658), .ZN(n15612) );
  AOI22_X1 U18713 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(n9758), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15579) );
  AOI22_X1 U18714 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n15600), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15578) );
  AOI22_X1 U18715 ( .A1(n17209), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n15553), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15570) );
  OAI21_X1 U18716 ( .B1(n12917), .B2(n18245), .A(n15570), .ZN(n15576) );
  AOI22_X1 U18717 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17205), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15574) );
  AOI22_X1 U18718 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15573) );
  AOI22_X1 U18719 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15572) );
  AOI22_X1 U18720 ( .A1(n15593), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15571) );
  NAND4_X1 U18721 ( .A1(n15574), .A2(n15573), .A3(n15572), .A4(n15571), .ZN(
        n15575) );
  AOI211_X1 U18722 ( .C1(n17215), .C2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n15576), .B(n15575), .ZN(n15577) );
  NAND3_X1 U18723 ( .A1(n15579), .A2(n15578), .A3(n15577), .ZN(n15649) );
  NAND2_X1 U18724 ( .A1(n15591), .A2(n15649), .ZN(n15590) );
  AOI22_X1 U18725 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n15589) );
  AOI22_X1 U18726 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n17209), .B1(
        P3_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n17122), .ZN(n15588) );
  INV_X1 U18727 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18256) );
  AOI22_X1 U18728 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n17206), .B1(
        n17205), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n15580) );
  OAI21_X1 U18729 ( .B1(n12917), .B2(n18256), .A(n15580), .ZN(n15586) );
  AOI22_X1 U18730 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n17212), .B1(
        P3_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n17117), .ZN(n15584) );
  AOI22_X1 U18731 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__6__SCAN_IN), .B2(n17217), .ZN(n15583) );
  AOI22_X1 U18732 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n9763), .B1(
        P3_INSTQUEUE_REG_14__6__SCAN_IN), .B2(n15559), .ZN(n15582) );
  AOI22_X1 U18733 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n17189), .B1(
        n9758), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n15581) );
  NAND4_X1 U18734 ( .A1(n15584), .A2(n15583), .A3(n15582), .A4(n15581), .ZN(
        n15585) );
  AOI211_X1 U18735 ( .C1(n9764), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n15586), .B(n15585), .ZN(n15587) );
  NAND3_X1 U18736 ( .A1(n15589), .A2(n15588), .A3(n15587), .ZN(n15650) );
  AOI21_X1 U18737 ( .B1(n17374), .B2(n16445), .A(n17674), .ZN(n15621) );
  INV_X1 U18738 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18145) );
  XOR2_X1 U18739 ( .A(n15590), .B(n17381), .Z(n17824) );
  INV_X1 U18740 ( .A(n15649), .ZN(n17385) );
  XNOR2_X1 U18741 ( .A(n15591), .B(n17385), .ZN(n15592) );
  NAND2_X1 U18742 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n15592), .ZN(
        n15617) );
  INV_X1 U18743 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18158) );
  XNOR2_X1 U18744 ( .A(n18158), .B(n15592), .ZN(n17841) );
  XNOR2_X1 U18745 ( .A(n17398), .B(n15658), .ZN(n15610) );
  NAND2_X1 U18746 ( .A1(n15648), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15609) );
  AOI22_X1 U18747 ( .A1(n15552), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n15550), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15599) );
  AOI22_X1 U18748 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n15554), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15598) );
  AOI22_X1 U18749 ( .A1(n15593), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15597) );
  AOI22_X1 U18750 ( .A1(n15551), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n15595), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15596) );
  NAND4_X1 U18751 ( .A1(n15599), .A2(n15598), .A3(n15597), .A4(n15596), .ZN(
        n15607) );
  AOI22_X1 U18752 ( .A1(n15559), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n15600), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15605) );
  AOI22_X1 U18753 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15604) );
  AOI22_X1 U18754 ( .A1(n15435), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15603) );
  AOI22_X1 U18755 ( .A1(n15601), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n15553), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15602) );
  NAND4_X1 U18756 ( .A1(n15605), .A2(n15604), .A3(n15603), .A4(n15602), .ZN(
        n15606) );
  INV_X1 U18757 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18851) );
  NAND2_X1 U18758 ( .A1(n17880), .A2(n17872), .ZN(n17871) );
  INV_X1 U18759 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18178) );
  OR2_X1 U18760 ( .A1(n18178), .A2(n15610), .ZN(n15611) );
  XOR2_X1 U18761 ( .A(n15612), .B(n17388), .Z(n15615) );
  INV_X1 U18762 ( .A(n15615), .ZN(n15613) );
  NAND2_X1 U18763 ( .A1(n15615), .A2(n15614), .ZN(n15616) );
  NAND2_X1 U18764 ( .A1(n17841), .A2(n17840), .ZN(n17839) );
  INV_X1 U18765 ( .A(n15650), .ZN(n17378) );
  XNOR2_X1 U18766 ( .A(n15618), .B(n17378), .ZN(n15619) );
  XOR2_X1 U18767 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n15619), .Z(
        n17812) );
  NAND2_X1 U18768 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15619), .ZN(
        n15620) );
  NAND2_X1 U18769 ( .A1(n15621), .A2(n15623), .ZN(n15624) );
  XNOR2_X1 U18770 ( .A(n15623), .B(n15622), .ZN(n17796) );
  NAND2_X2 U18771 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n15680), .ZN(
        n17993) );
  NAND2_X1 U18772 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18091) );
  NOR2_X1 U18773 ( .A1(n18091), .A2(n18058), .ZN(n18072) );
  INV_X1 U18774 ( .A(n18072), .ZN(n17732) );
  NOR3_X1 U18775 ( .A1(n17732), .A2(n17726), .A3(n18047), .ZN(n17691) );
  NAND2_X1 U18776 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17691), .ZN(
        n18039) );
  INV_X1 U18777 ( .A(n18039), .ZN(n18018) );
  NAND2_X1 U18778 ( .A1(n18018), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17672) );
  NAND2_X1 U18779 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18000) );
  INV_X1 U18780 ( .A(n18000), .ZN(n17948) );
  INV_X1 U18781 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17609) );
  INV_X1 U18782 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17951) );
  NOR2_X1 U18783 ( .A1(n17987), .A2(n17951), .ZN(n17967) );
  NAND2_X1 U18784 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17967), .ZN(
        n16440) );
  NOR2_X1 U18785 ( .A1(n17609), .A2(n17597), .ZN(n15691) );
  NAND2_X1 U18786 ( .A1(n17948), .A2(n15691), .ZN(n17937) );
  NOR2_X1 U18787 ( .A1(n17925), .A2(n17937), .ZN(n15689) );
  NAND2_X1 U18788 ( .A1(n18025), .A2(n15689), .ZN(n17581) );
  INV_X1 U18789 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17928) );
  NOR2_X1 U18790 ( .A1(n17581), .A2(n17928), .ZN(n17559) );
  NAND2_X1 U18791 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15692) );
  INV_X1 U18792 ( .A(n15692), .ZN(n17891) );
  NAND2_X1 U18793 ( .A1(n17559), .A2(n17891), .ZN(n17893) );
  NAND2_X1 U18794 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15647) );
  NOR2_X1 U18795 ( .A1(n17893), .A2(n15647), .ZN(n16455) );
  NAND2_X1 U18796 ( .A1(n18232), .A2(n16394), .ZN(n15625) );
  NOR2_X1 U18797 ( .A1(n18253), .A2(n15625), .ZN(n15630) );
  NAND2_X1 U18798 ( .A1(n15630), .A2(n15626), .ZN(n16437) );
  INV_X1 U18799 ( .A(n16437), .ZN(n18662) );
  XOR2_X1 U18800 ( .A(n18232), .B(n18227), .Z(n15628) );
  OAI21_X1 U18801 ( .B1(n15628), .B2(n15627), .A(n18875), .ZN(n16559) );
  NOR3_X1 U18802 ( .A1(n15629), .A2(n18660), .A3(n16559), .ZN(n15640) );
  INV_X1 U18803 ( .A(n15630), .ZN(n15638) );
  OAI211_X1 U18804 ( .C1(n15635), .C2(n15634), .A(n18232), .B(n18666), .ZN(
        n15636) );
  OAI211_X1 U18805 ( .C1(n15638), .C2(n18661), .A(n15637), .B(n15636), .ZN(
        n15639) );
  NOR2_X1 U18806 ( .A1(n16436), .A2(n18199), .ZN(n18050) );
  NOR2_X1 U18807 ( .A1(n18227), .A2(n15643), .ZN(n15645) );
  INV_X1 U18808 ( .A(n15647), .ZN(n15703) );
  INV_X1 U18809 ( .A(n15689), .ZN(n17907) );
  NAND2_X1 U18810 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17707) );
  INV_X1 U18811 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18080) );
  NOR2_X1 U18812 ( .A1(n18080), .A2(n17732), .ZN(n18037) );
  NOR2_X1 U18813 ( .A1(n15659), .A2(n15658), .ZN(n15656) );
  NOR2_X1 U18814 ( .A1(n17388), .A2(n15656), .ZN(n15654) );
  NAND2_X1 U18815 ( .A1(n15654), .A2(n15649), .ZN(n15652) );
  NOR2_X1 U18816 ( .A1(n17381), .A2(n15652), .ZN(n15667) );
  NAND2_X1 U18817 ( .A1(n15667), .A2(n15650), .ZN(n15651) );
  NOR2_X1 U18818 ( .A1(n17374), .A2(n15651), .ZN(n15676) );
  XNOR2_X1 U18819 ( .A(n16436), .B(n15651), .ZN(n17803) );
  XOR2_X1 U18820 ( .A(n17381), .B(n15652), .Z(n15653) );
  NOR2_X1 U18821 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n15653), .ZN(
        n15666) );
  XNOR2_X1 U18822 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n15653), .ZN(
        n17822) );
  XNOR2_X1 U18823 ( .A(n17385), .B(n15654), .ZN(n15655) );
  NAND2_X1 U18824 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n15655), .ZN(
        n15665) );
  XNOR2_X1 U18825 ( .A(n18158), .B(n15655), .ZN(n17836) );
  XOR2_X1 U18826 ( .A(n17388), .B(n15656), .Z(n15657) );
  NAND2_X1 U18827 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15657), .ZN(
        n15664) );
  XOR2_X1 U18828 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n15657), .Z(
        n17851) );
  INV_X1 U18829 ( .A(n15658), .ZN(n17393) );
  XNOR2_X1 U18830 ( .A(n17393), .B(n15659), .ZN(n15660) );
  OR2_X1 U18831 ( .A1(n18178), .A2(n15660), .ZN(n15663) );
  XNOR2_X1 U18832 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n15660), .ZN(
        n17861) );
  AOI21_X1 U18833 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n17398), .A(
        n15774), .ZN(n15662) );
  NOR2_X1 U18834 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n17398), .ZN(
        n15661) );
  AOI221_X1 U18835 ( .B1(n15774), .B2(n17398), .C1(n15662), .C2(n18851), .A(
        n15661), .ZN(n17860) );
  NAND2_X1 U18836 ( .A1(n17861), .A2(n17860), .ZN(n17859) );
  NAND2_X1 U18837 ( .A1(n15663), .A2(n17859), .ZN(n17850) );
  NAND2_X1 U18838 ( .A1(n17851), .A2(n17850), .ZN(n17849) );
  NAND2_X1 U18839 ( .A1(n15664), .A2(n17849), .ZN(n17835) );
  NAND2_X1 U18840 ( .A1(n17836), .A2(n17835), .ZN(n17834) );
  NAND2_X1 U18841 ( .A1(n15665), .A2(n17834), .ZN(n17821) );
  NOR2_X1 U18842 ( .A1(n17822), .A2(n17821), .ZN(n17820) );
  NOR2_X1 U18843 ( .A1(n15666), .A2(n17820), .ZN(n15669) );
  XNOR2_X1 U18844 ( .A(n17378), .B(n15667), .ZN(n15668) );
  NAND2_X1 U18845 ( .A1(n15669), .A2(n15668), .ZN(n15670) );
  XOR2_X1 U18846 ( .A(n15669), .B(n15668), .Z(n17809) );
  NAND2_X1 U18847 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17809), .ZN(
        n17808) );
  NAND2_X1 U18848 ( .A1(n15670), .A2(n17808), .ZN(n17802) );
  INV_X1 U18849 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15671) );
  NAND2_X1 U18850 ( .A1(n15676), .A2(n15672), .ZN(n15677) );
  INV_X1 U18851 ( .A(n15672), .ZN(n15675) );
  NAND2_X1 U18852 ( .A1(n17803), .A2(n17802), .ZN(n15674) );
  NAND2_X1 U18853 ( .A1(n15676), .A2(n15675), .ZN(n15673) );
  OAI211_X1 U18854 ( .C1(n15676), .C2(n15675), .A(n15674), .B(n15673), .ZN(
        n17788) );
  NAND2_X1 U18855 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17788), .ZN(
        n17787) );
  NAND2_X1 U18856 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17921), .ZN(
        n17565) );
  NAND2_X1 U18857 ( .A1(n15703), .A2(n17895), .ZN(n16451) );
  NAND2_X1 U18858 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17909) );
  NOR2_X1 U18859 ( .A1(n15692), .A2(n17909), .ZN(n15698) );
  NAND2_X1 U18860 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18119) );
  NOR2_X1 U18861 ( .A1(n10100), .A2(n18119), .ZN(n17992) );
  AOI21_X1 U18862 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n17989) );
  NAND3_X1 U18863 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17991) );
  NOR2_X1 U18864 ( .A1(n17989), .A2(n17991), .ZN(n18114) );
  NAND2_X1 U18865 ( .A1(n17992), .A2(n18114), .ZN(n18015) );
  NOR2_X1 U18866 ( .A1(n17672), .A2(n18015), .ZN(n17947) );
  NAND2_X1 U18867 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17990) );
  NOR2_X1 U18868 ( .A1(n17990), .A2(n17991), .ZN(n18115) );
  NAND2_X1 U18869 ( .A1(n18115), .A2(n17992), .ZN(n18097) );
  NOR2_X1 U18870 ( .A1(n17672), .A2(n18097), .ZN(n17946) );
  NOR2_X1 U18871 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18206), .ZN(
        n18192) );
  NOR2_X1 U18872 ( .A1(n18192), .A2(n18173), .ZN(n18179) );
  AOI22_X1 U18873 ( .A1(n18690), .A2(n17947), .B1(n17946), .B2(n18179), .ZN(
        n16438) );
  NOR2_X1 U18874 ( .A1(n16438), .A2(n17937), .ZN(n17911) );
  NAND4_X1 U18875 ( .A1(n15703), .A2(n18184), .A3(n15698), .A4(n17911), .ZN(
        n16425) );
  OAI21_X1 U18876 ( .B1(n18165), .B2(n16451), .A(n16425), .ZN(n15678) );
  AOI21_X1 U18877 ( .B1(n16455), .B2(n18050), .A(n15678), .ZN(n15759) );
  NAND2_X1 U18878 ( .A1(n18662), .A2(n16436), .ZN(n16446) );
  NOR2_X1 U18879 ( .A1(n17674), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17657) );
  NAND2_X1 U18880 ( .A1(n17657), .A2(n17987), .ZN(n15679) );
  NOR2_X1 U18881 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n15679), .ZN(
        n17622) );
  INV_X1 U18882 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17612) );
  NAND2_X1 U18883 ( .A1(n17622), .A2(n17612), .ZN(n17596) );
  NOR3_X1 U18884 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n17596), .ZN(n15690) );
  INV_X1 U18885 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15682) );
  NAND2_X1 U18886 ( .A1(n17745), .A2(n18058), .ZN(n17730) );
  NAND2_X1 U18887 ( .A1(n17698), .A2(n10133), .ZN(n15684) );
  NOR2_X2 U18888 ( .A1(n17754), .A2(n17780), .ZN(n17721) );
  INV_X1 U18889 ( .A(n17672), .ZN(n17995) );
  NAND2_X1 U18890 ( .A1(n15688), .A2(n15685), .ZN(n17673) );
  NAND2_X1 U18891 ( .A1(n15685), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15687) );
  INV_X1 U18892 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18023) );
  INV_X1 U18893 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18007) );
  OAI221_X1 U18894 ( .B1(n15690), .B2(n15689), .C1(n15690), .C2(n17673), .A(
        n17635), .ZN(n17574) );
  NOR2_X2 U18895 ( .A1(n17574), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17573) );
  NAND2_X1 U18896 ( .A1(n17948), .A2(n17673), .ZN(n17621) );
  NAND2_X2 U18897 ( .A1(n17635), .A2(n17621), .ZN(n17658) );
  NAND2_X1 U18898 ( .A1(n15691), .A2(n17658), .ZN(n17584) );
  INV_X1 U18899 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17568) );
  OR2_X1 U18900 ( .A1(n17674), .A2(n17573), .ZN(n17566) );
  OAI221_X1 U18901 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17781), 
        .C1(n17567), .C2(n17568), .A(n17566), .ZN(n17551) );
  NOR2_X1 U18902 ( .A1(n17567), .A2(n17781), .ZN(n15693) );
  NOR3_X1 U18903 ( .A1(n16458), .A2(n17781), .A3(n16441), .ZN(n15755) );
  NOR2_X1 U18904 ( .A1(n15754), .A2(n15755), .ZN(n15696) );
  XNOR2_X1 U18905 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B(n15696), .ZN(
        n16421) );
  INV_X1 U18906 ( .A(n17930), .ZN(n18118) );
  INV_X1 U18907 ( .A(n18098), .ZN(n18067) );
  INV_X1 U18908 ( .A(n18692), .ZN(n18680) );
  NAND2_X1 U18909 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n15698), .ZN(
        n17522) );
  NOR2_X1 U18910 ( .A1(n17609), .A2(n17522), .ZN(n16444) );
  INV_X1 U18911 ( .A(n17947), .ZN(n17906) );
  INV_X1 U18912 ( .A(n15698), .ZN(n17887) );
  OR2_X1 U18913 ( .A1(n17937), .A2(n17887), .ZN(n17543) );
  OAI21_X1 U18914 ( .B1(n17906), .B2(n17543), .A(n18690), .ZN(n17890) );
  NAND2_X1 U18915 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17946), .ZN(
        n18016) );
  NOR2_X1 U18916 ( .A1(n18000), .A2(n18001), .ZN(n17614) );
  INV_X1 U18917 ( .A(n17614), .ZN(n17963) );
  NOR2_X1 U18918 ( .A1(n16440), .A2(n17963), .ZN(n17599) );
  INV_X1 U18919 ( .A(n17599), .ZN(n17950) );
  OAI21_X1 U18920 ( .B1(n18016), .B2(n17950), .A(n18692), .ZN(n17952) );
  INV_X1 U18921 ( .A(n17946), .ZN(n17996) );
  NOR2_X1 U18922 ( .A1(n17937), .A2(n17996), .ZN(n17888) );
  INV_X1 U18923 ( .A(n17888), .ZN(n15699) );
  OAI21_X1 U18924 ( .B1(n17887), .B2(n15699), .A(n18206), .ZN(n15700) );
  AND4_X1 U18925 ( .A1(n18184), .A2(n17890), .A3(n17952), .A4(n15700), .ZN(
        n15701) );
  OAI21_X1 U18926 ( .B1(n18680), .B2(n16444), .A(n15701), .ZN(n15757) );
  INV_X1 U18927 ( .A(n15757), .ZN(n15702) );
  OAI21_X1 U18928 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18067), .A(
        n15702), .ZN(n16450) );
  AOI21_X1 U18929 ( .B1(n16458), .B2(n18118), .A(n16450), .ZN(n15705) );
  INV_X1 U18930 ( .A(n18050), .ZN(n18120) );
  NAND2_X1 U18931 ( .A1(n15703), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16399) );
  NOR2_X1 U18932 ( .A1(n17893), .A2(n16399), .ZN(n16406) );
  INV_X1 U18933 ( .A(n17895), .ZN(n17523) );
  NOR2_X1 U18934 ( .A1(n17523), .A2(n16399), .ZN(n16405) );
  OAI22_X1 U18935 ( .A1(n18120), .A2(n16406), .B1(n18165), .B2(n16405), .ZN(
        n15704) );
  INV_X1 U18936 ( .A(n15704), .ZN(n15758) );
  OAI21_X1 U18937 ( .B1(n9760), .B2(n15705), .A(n15758), .ZN(n15706) );
  AOI22_X1 U18938 ( .A1(n18083), .A2(n16421), .B1(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15706), .ZN(n15707) );
  NAND2_X1 U18939 ( .A1(n9760), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16419) );
  OAI211_X1 U18940 ( .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15759), .A(
        n15707), .B(n16419), .ZN(P3_U2833) );
  AOI22_X1 U18941 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n9882), .B1(
        P2_EBX_REG_22__SCAN_IN), .B2(n19054), .ZN(n15716) );
  INV_X1 U18942 ( .A(n15708), .ZN(n15709) );
  AOI22_X1 U18943 ( .A1(n15709), .A2(n19060), .B1(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n19003), .ZN(n15715) );
  INV_X1 U18944 ( .A(n15710), .ZN(n16190) );
  AOI22_X1 U18945 ( .A1(n16217), .A2(n19066), .B1(n18980), .B2(n16190), .ZN(
        n15714) );
  OAI211_X1 U18946 ( .C1(n15712), .C2(n16223), .A(n19050), .B(n15711), .ZN(
        n15713) );
  NAND4_X1 U18947 ( .A1(n15716), .A2(n15715), .A3(n15714), .A4(n15713), .ZN(
        P2_U2833) );
  NOR2_X1 U18948 ( .A1(n15717), .A2(n20611), .ZN(n15722) );
  AOI21_X1 U18949 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n15722), .A(
        n15718), .ZN(n15720) );
  NAND2_X1 U18950 ( .A1(n15720), .A2(n15719), .ZN(n15721) );
  OAI21_X1 U18951 ( .B1(n15722), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n15721), .ZN(n15724) );
  INV_X1 U18952 ( .A(n15724), .ZN(n15726) );
  AOI21_X1 U18953 ( .B1(n11766), .B2(n15724), .A(n15723), .ZN(n15725) );
  AOI21_X1 U18954 ( .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15726), .A(
        n15725), .ZN(n15731) );
  INV_X1 U18955 ( .A(n15731), .ZN(n15728) );
  INV_X1 U18956 ( .A(n15730), .ZN(n15727) );
  AOI21_X1 U18957 ( .B1(n15728), .B2(n15727), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n15729) );
  AOI21_X1 U18958 ( .B1(n15731), .B2(n15730), .A(n15729), .ZN(n15739) );
  OAI21_X1 U18959 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n15732), .ZN(n15734) );
  AND4_X1 U18960 ( .A1(n15736), .A2(n15735), .A3(n15734), .A4(n15733), .ZN(
        n15738) );
  OAI211_X1 U18961 ( .C1(n15739), .C2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n15738), .B(n15737), .ZN(n15746) );
  AND2_X1 U18962 ( .A1(n20838), .A2(n15740), .ZN(n15744) );
  NAND4_X1 U18963 ( .A1(n13176), .A2(n15742), .A3(n15763), .A4(n15741), .ZN(
        n15743) );
  OAI21_X1 U18964 ( .B1(n15747), .B2(n15744), .A(n15743), .ZN(n16109) );
  AOI221_X1 U18965 ( .B1(n11495), .B2(n20739), .C1(n15746), .C2(n20739), .A(
        n16109), .ZN(n16111) );
  AOI21_X1 U18966 ( .B1(n15747), .B2(n15746), .A(n15745), .ZN(n15748) );
  OAI211_X1 U18967 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n16106), .A(n15748), 
        .B(n16105), .ZN(n15749) );
  NOR2_X1 U18968 ( .A1(n16111), .A2(n15749), .ZN(n15753) );
  NAND2_X1 U18969 ( .A1(n20843), .A2(n15750), .ZN(n15751) );
  NAND2_X1 U18970 ( .A1(n11495), .A2(n15751), .ZN(n15752) );
  OAI22_X1 U18971 ( .A1(n15753), .A2(n11495), .B1(n16111), .B2(n15752), .ZN(
        P1_U3161) );
  INV_X1 U18972 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16427) );
  NAND2_X1 U18973 ( .A1(n16427), .A2(n15754), .ZN(n16381) );
  NAND2_X1 U18974 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15755), .ZN(
        n16382) );
  NAND2_X1 U18975 ( .A1(n16381), .A2(n16382), .ZN(n15756) );
  NAND2_X1 U18976 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15756), .ZN(
        n16384) );
  OAI21_X1 U18977 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15756), .A(
        n16384), .ZN(n16409) );
  OAI221_X1 U18978 ( .B1(n15757), .B2(n18118), .C1(n15757), .C2(n16399), .A(
        n15697), .ZN(n16424) );
  INV_X1 U18979 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16426) );
  AOI21_X1 U18980 ( .B1(n15758), .B2(n16424), .A(n16426), .ZN(n15761) );
  NOR3_X1 U18981 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15759), .A3(
        n16427), .ZN(n15760) );
  AOI211_X1 U18982 ( .C1(P3_REIP_REG_30__SCAN_IN), .C2(n9760), .A(n15761), .B(
        n15760), .ZN(n15762) );
  OAI21_X1 U18983 ( .B1(n18121), .B2(n16409), .A(n15762), .ZN(P3_U2832) );
  INV_X1 U18984 ( .A(HOLD), .ZN(n21002) );
  INV_X1 U18985 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n15764) );
  NAND2_X1 U18986 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n15764), .ZN(n20748) );
  INV_X1 U18987 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20746) );
  INV_X1 U18988 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20749) );
  NOR2_X1 U18989 ( .A1(n20746), .A2(n20749), .ZN(n20752) );
  AOI221_X1 U18990 ( .B1(n15764), .B2(n20752), .C1(n21002), .C2(n20752), .A(
        n15763), .ZN(n15766) );
  NAND2_X1 U18991 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20838), .ZN(n15765) );
  OAI211_X1 U18992 ( .C1(n21002), .C2(n20748), .A(n15766), .B(n15765), .ZN(
        P1_U3195) );
  AND2_X1 U18993 ( .A1(n20008), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR3_X1 U18994 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n15767) );
  NOR3_X1 U18995 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n18894), .A3(n19765), 
        .ZN(n16360) );
  NOR4_X1 U18996 ( .A1(n15767), .A2(n16367), .A3(n16377), .A4(n16360), .ZN(
        P2_U3178) );
  AOI221_X1 U18997 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16377), .C1(n15768), .C2(
        n16377), .A(n19683), .ZN(n19884) );
  INV_X1 U18998 ( .A(n19884), .ZN(n19885) );
  NOR2_X1 U18999 ( .A1(n15769), .A2(n19885), .ZN(P2_U3047) );
  NAND2_X1 U19000 ( .A1(n9796), .A2(n17260), .ZN(n17401) );
  INV_X1 U19001 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17461) );
  NAND2_X1 U19002 ( .A1(n17348), .A2(n15773), .ZN(n17397) );
  NAND2_X2 U19003 ( .A1(n18693), .A2(n17260), .ZN(n17394) );
  AOI22_X1 U19004 ( .A1(n17400), .A2(BUF2_REG_0__SCAN_IN), .B1(n17399), .B2(
        n15774), .ZN(n15775) );
  OAI221_X1 U19005 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17401), .C1(n17461), 
        .C2(n17260), .A(n15775), .ZN(P3_U2735) );
  OAI21_X1 U19006 ( .B1(n15787), .B2(n19937), .A(n15776), .ZN(n15804) );
  AOI21_X1 U19007 ( .B1(n19964), .B2(n14514), .A(n15804), .ZN(n15777) );
  NOR2_X1 U19008 ( .A1(n15777), .A2(n20788), .ZN(n15782) );
  NOR3_X1 U19009 ( .A1(n19937), .A2(P1_REIP_REG_22__SCAN_IN), .A3(n15778), 
        .ZN(n15781) );
  OAI22_X1 U19010 ( .A1(n15779), .A2(n19931), .B1(n19977), .B2(n20858), .ZN(
        n15780) );
  NOR3_X1 U19011 ( .A1(n15782), .A2(n15781), .A3(n15780), .ZN(n15786) );
  AOI22_X1 U19012 ( .A1(n15784), .A2(n19949), .B1(n15783), .B2(n15861), .ZN(
        n15785) );
  OAI211_X1 U19013 ( .C1(n19945), .C2(n15962), .A(n15786), .B(n15785), .ZN(
        P1_U2818) );
  INV_X1 U19014 ( .A(n15787), .ZN(n15788) );
  NOR3_X1 U19015 ( .A1(n19937), .A2(P1_REIP_REG_21__SCAN_IN), .A3(n15788), 
        .ZN(n15789) );
  AOI21_X1 U19016 ( .B1(P1_EBX_REG_21__SCAN_IN), .B2(n19942), .A(n15789), .ZN(
        n15790) );
  OAI21_X1 U19017 ( .B1(n12134), .B2(n19931), .A(n15790), .ZN(n15791) );
  AOI21_X1 U19018 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n15804), .A(n15791), 
        .ZN(n15796) );
  NOR2_X1 U19019 ( .A1(n15792), .A2(n19945), .ZN(n15793) );
  AOI21_X1 U19020 ( .B1(n15794), .B2(n19949), .A(n15793), .ZN(n15795) );
  OAI211_X1 U19021 ( .C1(n15797), .C2(n19983), .A(n15796), .B(n15795), .ZN(
        P1_U2819) );
  AOI22_X1 U19022 ( .A1(n19942), .A2(P1_EBX_REG_20__SCAN_IN), .B1(n15798), 
        .B2(n15861), .ZN(n15806) );
  INV_X1 U19023 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20783) );
  OR2_X1 U19024 ( .A1(n15799), .A2(n15843), .ZN(n15810) );
  INV_X1 U19025 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n20785) );
  OAI21_X1 U19026 ( .B1(n20783), .B2(n15810), .A(n20785), .ZN(n15803) );
  OAI22_X1 U19027 ( .A1(n15801), .A2(n19926), .B1(n19945), .B2(n15800), .ZN(
        n15802) );
  AOI21_X1 U19028 ( .B1(n15804), .B2(n15803), .A(n15802), .ZN(n15805) );
  OAI211_X1 U19029 ( .C1(n15807), .C2(n19931), .A(n15806), .B(n15805), .ZN(
        P1_U2820) );
  INV_X1 U19030 ( .A(n15892), .ZN(n15808) );
  AOI21_X1 U19031 ( .B1(n15861), .B2(n15808), .A(n19947), .ZN(n15809) );
  OAI21_X1 U19032 ( .B1(n12091), .B2(n19931), .A(n15809), .ZN(n15812) );
  NOR2_X1 U19033 ( .A1(n15810), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n15811) );
  AOI211_X1 U19034 ( .C1(P1_EBX_REG_19__SCAN_IN), .C2(n19942), .A(n15812), .B(
        n15811), .ZN(n15817) );
  AOI22_X1 U19035 ( .A1(n15889), .A2(n19949), .B1(n19974), .B2(n15964), .ZN(
        n15816) );
  INV_X1 U19036 ( .A(n15813), .ZN(n15814) );
  NOR3_X1 U19037 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n15814), .A3(n15843), 
        .ZN(n15823) );
  OAI21_X1 U19038 ( .B1(n15823), .B2(n15818), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n15815) );
  NAND3_X1 U19039 ( .A1(n15817), .A2(n15816), .A3(n15815), .ZN(P1_U2821) );
  NAND2_X1 U19040 ( .A1(n15818), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n15820) );
  AOI21_X1 U19041 ( .B1(n19960), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n19947), .ZN(n15819) );
  OAI211_X1 U19042 ( .C1(n15821), .C2(n19977), .A(n15820), .B(n15819), .ZN(
        n15822) );
  AOI211_X1 U19043 ( .C1(n15861), .C2(n15824), .A(n15823), .B(n15822), .ZN(
        n15827) );
  NAND2_X1 U19044 ( .A1(n15825), .A2(n19949), .ZN(n15826) );
  OAI211_X1 U19045 ( .C1(n15977), .C2(n19945), .A(n15827), .B(n15826), .ZN(
        P1_U2822) );
  AOI22_X1 U19046 ( .A1(n15837), .A2(P1_REIP_REG_16__SCAN_IN), .B1(n19942), 
        .B2(P1_EBX_REG_16__SCAN_IN), .ZN(n15828) );
  OAI211_X1 U19047 ( .C1(n19931), .C2(n15829), .A(n15828), .B(n19969), .ZN(
        n15834) );
  OAI21_X1 U19048 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(P1_REIP_REG_15__SCAN_IN), 
        .A(n15830), .ZN(n15831) );
  OAI22_X1 U19049 ( .A1(n15832), .A2(n19926), .B1(n15831), .B2(n15843), .ZN(
        n15833) );
  AOI211_X1 U19050 ( .C1(n15835), .C2(n15861), .A(n15834), .B(n15833), .ZN(
        n15836) );
  OAI21_X1 U19051 ( .B1(n19945), .B2(n15994), .A(n15836), .ZN(P1_U2824) );
  AOI22_X1 U19052 ( .A1(n15837), .A2(P1_REIP_REG_15__SCAN_IN), .B1(n19942), 
        .B2(P1_EBX_REG_15__SCAN_IN), .ZN(n15838) );
  OAI211_X1 U19053 ( .C1(n19931), .C2(n15839), .A(n15838), .B(n19969), .ZN(
        n15840) );
  AOI21_X1 U19054 ( .B1(n19974), .B2(n16003), .A(n15840), .ZN(n15842) );
  AOI22_X1 U19055 ( .A1(n15910), .A2(n19949), .B1(n15861), .B2(n15909), .ZN(
        n15841) );
  OAI211_X1 U19056 ( .C1(P1_REIP_REG_15__SCAN_IN), .C2(n15843), .A(n15842), 
        .B(n15841), .ZN(P1_U2825) );
  AOI21_X1 U19057 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n15844), .A(
        P1_REIP_REG_14__SCAN_IN), .ZN(n15853) );
  INV_X1 U19058 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n15846) );
  OAI22_X1 U19059 ( .A1(n19931), .A2(n15846), .B1(n19977), .B2(n15845), .ZN(
        n15847) );
  AOI211_X1 U19060 ( .C1(n16007), .C2(n19974), .A(n19947), .B(n15847), .ZN(
        n15852) );
  INV_X1 U19061 ( .A(n15848), .ZN(n15849) );
  AOI22_X1 U19062 ( .A1(n15850), .A2(n19949), .B1(n15849), .B2(n15861), .ZN(
        n15851) );
  OAI211_X1 U19063 ( .C1(n15854), .C2(n15853), .A(n15852), .B(n15851), .ZN(
        P1_U2826) );
  INV_X1 U19064 ( .A(n15855), .ZN(n15873) );
  AOI21_X1 U19065 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n15873), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n15864) );
  INV_X1 U19066 ( .A(n16029), .ZN(n15856) );
  NAND2_X1 U19067 ( .A1(n19974), .A2(n15856), .ZN(n15859) );
  NAND2_X1 U19068 ( .A1(n19960), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15857) );
  AND2_X1 U19069 ( .A1(n15857), .A2(n19969), .ZN(n15858) );
  OAI211_X1 U19070 ( .C1(n19977), .C2(n21094), .A(n15859), .B(n15858), .ZN(
        n15860) );
  INV_X1 U19071 ( .A(n15860), .ZN(n15863) );
  INV_X1 U19072 ( .A(n15881), .ZN(n15917) );
  AOI22_X1 U19073 ( .A1(n15918), .A2(n15861), .B1(n19949), .B2(n15917), .ZN(
        n15862) );
  OAI211_X1 U19074 ( .C1(n15865), .C2(n15864), .A(n15863), .B(n15862), .ZN(
        P1_U2828) );
  INV_X1 U19075 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n15870) );
  AOI21_X1 U19076 ( .B1(n15868), .B2(n15867), .A(n15866), .ZN(n16035) );
  AOI22_X1 U19077 ( .A1(n19942), .A2(P1_EBX_REG_11__SCAN_IN), .B1(n19974), 
        .B2(n16035), .ZN(n15869) );
  OAI211_X1 U19078 ( .C1(n19931), .C2(n15870), .A(n15869), .B(n19969), .ZN(
        n15871) );
  AOI221_X1 U19079 ( .B1(n15873), .B2(n20771), .C1(n15872), .C2(
        P1_REIP_REG_11__SCAN_IN), .A(n15871), .ZN(n15877) );
  XNOR2_X1 U19080 ( .A(n15875), .B(n15874), .ZN(n15925) );
  NAND2_X1 U19081 ( .A1(n19949), .A2(n15925), .ZN(n15876) );
  OAI211_X1 U19082 ( .C1(n19983), .C2(n15928), .A(n15877), .B(n15876), .ZN(
        P1_U2829) );
  AOI22_X1 U19083 ( .A1(n15925), .A2(n19996), .B1(n19995), .B2(n16035), .ZN(
        n15878) );
  OAI21_X1 U19084 ( .B1(n20000), .B2(n15879), .A(n15878), .ZN(P1_U2861) );
  AOI22_X1 U19085 ( .A1(P1_EAX_REG_12__SCAN_IN), .A2(n15884), .B1(n15883), 
        .B2(n20017), .ZN(n15880) );
  OAI21_X1 U19086 ( .B1(n20004), .B2(n15881), .A(n15880), .ZN(P1_U2892) );
  INV_X1 U19087 ( .A(n15925), .ZN(n15886) );
  AOI22_X1 U19088 ( .A1(P1_EAX_REG_11__SCAN_IN), .A2(n15884), .B1(n15883), 
        .B2(n15882), .ZN(n15885) );
  OAI21_X1 U19089 ( .B1(n20004), .B2(n15886), .A(n15885), .ZN(P1_U2893) );
  AOI22_X1 U19090 ( .A1(n20039), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n20099), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15891) );
  NAND2_X1 U19091 ( .A1(n14510), .A2(n15971), .ZN(n15887) );
  MUX2_X1 U19092 ( .A(n14510), .B(n15887), .S(n15893), .Z(n15888) );
  XNOR2_X1 U19093 ( .A(n15888), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15963) );
  AOI22_X1 U19094 ( .A1(n15889), .A2(n20045), .B1(n20046), .B2(n15963), .ZN(
        n15890) );
  OAI211_X1 U19095 ( .C1(n20050), .C2(n15892), .A(n15891), .B(n15890), .ZN(
        P1_U2980) );
  NAND2_X1 U19096 ( .A1(n15893), .A2(n15998), .ZN(n15899) );
  INV_X1 U19097 ( .A(n15894), .ZN(n15895) );
  AOI21_X1 U19098 ( .B1(n15897), .B2(n15896), .A(n15895), .ZN(n15898) );
  MUX2_X1 U19099 ( .A(n15899), .B(n15893), .S(n15898), .Z(n15900) );
  XNOR2_X1 U19100 ( .A(n15900), .B(n15984), .ZN(n15990) );
  AOI22_X1 U19101 ( .A1(n20039), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n20099), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n15904) );
  AOI22_X1 U19102 ( .A1(n15902), .A2(n20045), .B1(n15919), .B2(n15901), .ZN(
        n15903) );
  OAI211_X1 U19103 ( .C1(n19904), .C2(n15990), .A(n15904), .B(n15903), .ZN(
        P1_U2982) );
  INV_X1 U19104 ( .A(n15905), .ZN(n15906) );
  AOI21_X1 U19105 ( .B1(n15908), .B2(n15907), .A(n15906), .ZN(n16005) );
  AOI22_X1 U19106 ( .A1(n20039), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n20099), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n15912) );
  AOI22_X1 U19107 ( .A1(n15910), .A2(n20045), .B1(n15919), .B2(n15909), .ZN(
        n15911) );
  OAI211_X1 U19108 ( .C1(n16005), .C2(n19904), .A(n15912), .B(n15911), .ZN(
        P1_U2984) );
  OAI21_X1 U19109 ( .B1(n15915), .B2(n15914), .A(n15913), .ZN(n15916) );
  INV_X1 U19110 ( .A(n15916), .ZN(n16034) );
  AOI22_X1 U19111 ( .A1(n20039), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n20099), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15921) );
  AOI22_X1 U19112 ( .A1(n15919), .A2(n15918), .B1(n20045), .B2(n15917), .ZN(
        n15920) );
  OAI211_X1 U19113 ( .C1(n16034), .C2(n19904), .A(n15921), .B(n15920), .ZN(
        P1_U2987) );
  AOI22_X1 U19114 ( .A1(n20039), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n20099), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15927) );
  NAND3_X1 U19115 ( .A1(n11747), .A2(n14460), .A3(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15923) );
  NAND2_X1 U19116 ( .A1(n15923), .A2(n15922), .ZN(n15924) );
  XNOR2_X1 U19117 ( .A(n15924), .B(n16021), .ZN(n16036) );
  AOI22_X1 U19118 ( .A1(n20046), .A2(n16036), .B1(n20045), .B2(n15925), .ZN(
        n15926) );
  OAI211_X1 U19119 ( .C1(n20050), .C2(n15928), .A(n15927), .B(n15926), .ZN(
        P1_U2988) );
  AOI22_X1 U19120 ( .A1(n20039), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20099), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15934) );
  NAND2_X1 U19121 ( .A1(n15931), .A2(n15930), .ZN(n15932) );
  XNOR2_X1 U19122 ( .A(n15929), .B(n15932), .ZN(n16078) );
  AOI22_X1 U19123 ( .A1(n16078), .A2(n20046), .B1(n20045), .B2(n19991), .ZN(
        n15933) );
  OAI211_X1 U19124 ( .C1(n20050), .C2(n19940), .A(n15934), .B(n15933), .ZN(
        P1_U2992) );
  AOI22_X1 U19125 ( .A1(n20039), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20099), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n15940) );
  XNOR2_X1 U19126 ( .A(n15937), .B(n15936), .ZN(n15938) );
  XNOR2_X1 U19127 ( .A(n15935), .B(n15938), .ZN(n16083) );
  AOI22_X1 U19128 ( .A1(n16083), .A2(n20046), .B1(n20045), .B2(n19950), .ZN(
        n15939) );
  OAI211_X1 U19129 ( .C1(n20050), .C2(n19953), .A(n15940), .B(n15939), .ZN(
        P1_U2993) );
  AOI22_X1 U19130 ( .A1(n20039), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20099), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n15946) );
  OAI21_X1 U19131 ( .B1(n15943), .B2(n15942), .A(n15941), .ZN(n15944) );
  INV_X1 U19132 ( .A(n15944), .ZN(n16094) );
  AOI22_X1 U19133 ( .A1(n16094), .A2(n20046), .B1(n20045), .B2(n19997), .ZN(
        n15945) );
  OAI211_X1 U19134 ( .C1(n20050), .C2(n19959), .A(n15946), .B(n15945), .ZN(
        P1_U2994) );
  AOI22_X1 U19135 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n15947), .B1(
        n20099), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n15952) );
  INV_X1 U19136 ( .A(n15948), .ZN(n15950) );
  AOI22_X1 U19137 ( .A1(n15950), .A2(n20079), .B1(n15955), .B2(n15949), .ZN(
        n15951) );
  OAI211_X1 U19138 ( .C1(n20102), .C2(n15953), .A(n15952), .B(n15951), .ZN(
        P1_U3008) );
  AOI22_X1 U19139 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n20099), .B1(n15955), 
        .B2(n15954), .ZN(n15961) );
  OAI21_X1 U19140 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n15957), .A(
        n15956), .ZN(n15959) );
  AOI22_X1 U19141 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n15959), .B1(
        n20079), .B2(n15958), .ZN(n15960) );
  OAI211_X1 U19142 ( .C1(n20102), .C2(n15962), .A(n15961), .B(n15960), .ZN(
        P1_U3009) );
  AOI22_X1 U19143 ( .A1(n20076), .A2(n15964), .B1(n20079), .B2(n15963), .ZN(
        n15970) );
  NOR2_X1 U19144 ( .A1(n16045), .A2(n20783), .ZN(n15965) );
  AOI221_X1 U19145 ( .B1(n15968), .B2(n15967), .C1(n15966), .C2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n15965), .ZN(n15969) );
  NAND2_X1 U19146 ( .A1(n15970), .A2(n15969), .ZN(P1_U3012) );
  NAND2_X1 U19147 ( .A1(n15976), .A2(n15971), .ZN(n15982) );
  NOR2_X1 U19148 ( .A1(n16017), .A2(n15972), .ZN(n16009) );
  OAI21_X1 U19149 ( .B1(n16017), .B2(n15973), .A(n20054), .ZN(n15974) );
  OAI211_X1 U19150 ( .C1(n16009), .C2(n20072), .A(n20052), .B(n15974), .ZN(
        n16018) );
  AOI21_X1 U19151 ( .B1(n16008), .B2(n15975), .A(n16018), .ZN(n16000) );
  OAI21_X1 U19152 ( .B1(n20093), .B2(n15976), .A(n16000), .ZN(n15986) );
  OAI22_X1 U19153 ( .A1(n15978), .A2(n20088), .B1(n20102), .B2(n15977), .ZN(
        n15979) );
  AOI21_X1 U19154 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n15986), .A(
        n15979), .ZN(n15981) );
  NAND2_X1 U19155 ( .A1(n20099), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n15980) );
  OAI211_X1 U19156 ( .C1(n16001), .C2(n15982), .A(n15981), .B(n15980), .ZN(
        P1_U3013) );
  INV_X1 U19157 ( .A(n15983), .ZN(n15987) );
  OAI21_X1 U19158 ( .B1(n15991), .B2(n16001), .A(n15984), .ZN(n15985) );
  AOI22_X1 U19159 ( .A1(n20076), .A2(n15987), .B1(n15986), .B2(n15985), .ZN(
        n15989) );
  NAND2_X1 U19160 ( .A1(n20099), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n15988) );
  OAI211_X1 U19161 ( .C1(n15990), .C2(n20088), .A(n15989), .B(n15988), .ZN(
        P1_U3014) );
  OAI21_X1 U19162 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n15991), .ZN(n15993) );
  OAI222_X1 U19163 ( .A1(n15994), .A2(n20102), .B1(n16001), .B2(n15993), .C1(
        n20088), .C2(n15992), .ZN(n15995) );
  INV_X1 U19164 ( .A(n15995), .ZN(n15997) );
  NAND2_X1 U19165 ( .A1(n20099), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n15996) );
  OAI211_X1 U19166 ( .C1(n16000), .C2(n15998), .A(n15997), .B(n15996), .ZN(
        P1_U3015) );
  NAND2_X1 U19167 ( .A1(n20099), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n15999) );
  OAI221_X1 U19168 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16001), 
        .C1(n11740), .C2(n16000), .A(n15999), .ZN(n16002) );
  AOI21_X1 U19169 ( .B1(n20076), .B2(n16003), .A(n16002), .ZN(n16004) );
  OAI21_X1 U19170 ( .B1(n16005), .B2(n20088), .A(n16004), .ZN(P1_U3016) );
  AOI22_X1 U19171 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16018), .B1(
        n20099), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n16012) );
  AOI22_X1 U19172 ( .A1(n20076), .A2(n16007), .B1(n20079), .B2(n16006), .ZN(
        n16011) );
  INV_X1 U19173 ( .A(n20081), .ZN(n16028) );
  OAI21_X1 U19174 ( .B1(n16028), .B2(n20071), .A(n20072), .ZN(n16088) );
  NAND3_X1 U19175 ( .A1(n16009), .A2(n16008), .A3(n16088), .ZN(n16010) );
  NAND3_X1 U19176 ( .A1(n16012), .A2(n16011), .A3(n16010), .ZN(P1_U3017) );
  AOI22_X1 U19177 ( .A1(n16014), .A2(n20079), .B1(n20076), .B2(n16013), .ZN(
        n16020) );
  NOR2_X1 U19178 ( .A1(n16045), .A2(n14017), .ZN(n16015) );
  AOI221_X1 U19179 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16018), 
        .C1(n16017), .C2(n16016), .A(n16015), .ZN(n16019) );
  NAND2_X1 U19180 ( .A1(n16020), .A2(n16019), .ZN(P1_U3018) );
  NAND2_X1 U19181 ( .A1(n16022), .A2(n16088), .ZN(n16070) );
  NOR2_X1 U19182 ( .A1(n16023), .A2(n16070), .ZN(n16032) );
  NAND2_X1 U19183 ( .A1(n16026), .A2(n16021), .ZN(n16040) );
  INV_X1 U19184 ( .A(n20054), .ZN(n20053) );
  OAI21_X1 U19185 ( .B1(n16022), .B2(n20072), .A(n20052), .ZN(n16063) );
  AOI21_X1 U19186 ( .B1(n16024), .B2(n16023), .A(n16063), .ZN(n16025) );
  OAI221_X1 U19187 ( .B1(n20053), .B2(n16026), .C1(n20053), .C2(n16042), .A(
        n16025), .ZN(n16037) );
  INV_X1 U19188 ( .A(n16037), .ZN(n16027) );
  OAI21_X1 U19189 ( .B1(n16028), .B2(n16040), .A(n16027), .ZN(n16031) );
  OAI22_X1 U19190 ( .A1(n16045), .A2(n20772), .B1(n20102), .B2(n16029), .ZN(
        n16030) );
  AOI221_X1 U19191 ( .B1(n16032), .B2(n11742), .C1(n16031), .C2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n16030), .ZN(n16033) );
  OAI21_X1 U19192 ( .B1(n16034), .B2(n20088), .A(n16033), .ZN(P1_U3019) );
  AOI22_X1 U19193 ( .A1(n20099), .A2(P1_REIP_REG_11__SCAN_IN), .B1(n20076), 
        .B2(n16035), .ZN(n16039) );
  AOI22_X1 U19194 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16037), .B1(
        n20079), .B2(n16036), .ZN(n16038) );
  OAI211_X1 U19195 ( .C1(n16070), .C2(n16040), .A(n16039), .B(n16038), .ZN(
        P1_U3020) );
  INV_X1 U19196 ( .A(n16063), .ZN(n16041) );
  OAI21_X1 U19197 ( .B1(n20053), .B2(n16042), .A(n16041), .ZN(n16043) );
  OAI21_X1 U19198 ( .B1(n16048), .B2(n16043), .A(n16065), .ZN(n16058) );
  OAI22_X1 U19199 ( .A1(n16045), .A2(n20768), .B1(n20102), .B2(n16044), .ZN(
        n16046) );
  AOI21_X1 U19200 ( .B1(n20079), .B2(n16047), .A(n16046), .ZN(n16050) );
  NOR2_X1 U19201 ( .A1(n16048), .A2(n16070), .ZN(n16054) );
  OAI221_X1 U19202 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n14557), .C2(n16059), .A(
        n16054), .ZN(n16049) );
  OAI211_X1 U19203 ( .C1(n14557), .C2(n16058), .A(n16050), .B(n16049), .ZN(
        P1_U3021) );
  NAND2_X1 U19204 ( .A1(n13790), .A2(n16051), .ZN(n16052) );
  AND2_X1 U19205 ( .A1(n16053), .A2(n16052), .ZN(n19984) );
  AOI22_X1 U19206 ( .A1(n20099), .A2(P1_REIP_REG_9__SCAN_IN), .B1(n20076), 
        .B2(n19984), .ZN(n16057) );
  AOI22_X1 U19207 ( .A1(n16055), .A2(n20079), .B1(n16054), .B2(n16059), .ZN(
        n16056) );
  OAI211_X1 U19208 ( .C1(n16059), .C2(n16058), .A(n16057), .B(n16056), .ZN(
        P1_U3022) );
  NAND2_X1 U19209 ( .A1(n20055), .A2(n16060), .ZN(n16097) );
  AOI21_X1 U19210 ( .B1(n16061), .B2(n20055), .A(n20053), .ZN(n16062) );
  OR2_X1 U19211 ( .A1(n16063), .A2(n16062), .ZN(n16093) );
  INV_X1 U19212 ( .A(n16093), .ZN(n16064) );
  OAI211_X1 U19213 ( .C1(n16028), .C2(n16097), .A(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n16064), .ZN(n16084) );
  NAND2_X1 U19214 ( .A1(n16065), .A2(n16084), .ZN(n16081) );
  INV_X1 U19215 ( .A(n16066), .ZN(n16069) );
  INV_X1 U19216 ( .A(n16067), .ZN(n16068) );
  AOI222_X1 U19217 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n20099), .B1(n20076), 
        .B2(n16069), .C1(n20079), .C2(n16068), .ZN(n16072) );
  INV_X1 U19218 ( .A(n16070), .ZN(n16085) );
  AND2_X1 U19219 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16085), .ZN(
        n16077) );
  OAI221_X1 U19220 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n11729), .C2(n16082), .A(
        n16077), .ZN(n16071) );
  OAI211_X1 U19221 ( .C1(n16081), .C2(n11729), .A(n16072), .B(n16071), .ZN(
        P1_U3023) );
  NOR2_X1 U19222 ( .A1(n16074), .A2(n16073), .ZN(n16075) );
  AOI22_X1 U19223 ( .A1(n20099), .A2(P1_REIP_REG_7__SCAN_IN), .B1(n20076), 
        .B2(n9862), .ZN(n16080) );
  AOI22_X1 U19224 ( .A1(n16078), .A2(n20079), .B1(n16077), .B2(n16082), .ZN(
        n16079) );
  OAI211_X1 U19225 ( .C1(n16082), .C2(n16081), .A(n16080), .B(n16079), .ZN(
        P1_U3024) );
  AOI22_X1 U19226 ( .A1(n16083), .A2(n20079), .B1(n20099), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n16087) );
  OAI21_X1 U19227 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16085), .A(
        n16084), .ZN(n16086) );
  OAI211_X1 U19228 ( .C1(n19944), .C2(n20102), .A(n16087), .B(n16086), .ZN(
        P1_U3025) );
  NAND2_X1 U19229 ( .A1(n20051), .A2(n16088), .ZN(n20065) );
  NAND2_X1 U19230 ( .A1(n16090), .A2(n16089), .ZN(n16091) );
  AND2_X1 U19231 ( .A1(n16092), .A2(n16091), .ZN(n19994) );
  AOI22_X1 U19232 ( .A1(n20099), .A2(P1_REIP_REG_5__SCAN_IN), .B1(n20076), 
        .B2(n19994), .ZN(n16096) );
  AOI22_X1 U19233 ( .A1(n16094), .A2(n20079), .B1(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n16093), .ZN(n16095) );
  OAI211_X1 U19234 ( .C1(n16097), .C2(n20065), .A(n16096), .B(n16095), .ZN(
        P1_U3026) );
  INV_X1 U19235 ( .A(n16098), .ZN(n16099) );
  OAI22_X1 U19236 ( .A1(n16101), .A2(n20824), .B1(n16100), .B2(n16099), .ZN(
        P1_U3468) );
  NAND4_X1 U19237 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n20742), .A4(n16106), .ZN(n16102) );
  NAND2_X1 U19238 ( .A1(n16103), .A2(n16102), .ZN(n20740) );
  INV_X1 U19239 ( .A(n20843), .ZN(n16107) );
  OAI21_X1 U19240 ( .B1(n16111), .B2(n11495), .A(n20739), .ZN(n16104) );
  OAI211_X1 U19241 ( .C1(n16107), .C2(n16106), .A(n16105), .B(n16104), .ZN(
        n16108) );
  AOI221_X1 U19242 ( .B1(n16110), .B2(n16109), .C1(n20740), .C2(n16109), .A(
        n16108), .ZN(P1_U3162) );
  NOR2_X1 U19243 ( .A1(n16111), .A2(n11495), .ZN(n16113) );
  OAI22_X1 U19244 ( .A1(n21100), .A2(n16113), .B1(n16112), .B2(n11495), .ZN(
        P1_U3466) );
  OAI222_X1 U19245 ( .A1(n19028), .A2(n14141), .B1(n19042), .B2(n16114), .C1(
        n19838), .C2(n9807), .ZN(n16115) );
  AOI21_X1 U19246 ( .B1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19024), .A(
        n16115), .ZN(n16119) );
  AOI22_X1 U19247 ( .A1(n16117), .A2(n19066), .B1(n18980), .B2(n16116), .ZN(
        n16118) );
  OAI211_X1 U19248 ( .C1(n19071), .C2(n16120), .A(n16119), .B(n16118), .ZN(
        P2_U2824) );
  AOI22_X1 U19249 ( .A1(P2_REIP_REG_29__SCAN_IN), .A2(n9882), .B1(
        P2_EBX_REG_29__SCAN_IN), .B2(n19054), .ZN(n16132) );
  AOI22_X1 U19250 ( .A1(n16121), .A2(n19060), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19024), .ZN(n16131) );
  INV_X1 U19251 ( .A(n16122), .ZN(n16123) );
  OAI22_X1 U19252 ( .A1(n16124), .A2(n19036), .B1(n16123), .B2(n19063), .ZN(
        n16125) );
  INV_X1 U19253 ( .A(n16125), .ZN(n16130) );
  OAI211_X1 U19254 ( .C1(n16128), .C2(n16127), .A(n19050), .B(n16126), .ZN(
        n16129) );
  NAND4_X1 U19255 ( .A1(n16132), .A2(n16131), .A3(n16130), .A4(n16129), .ZN(
        P2_U2826) );
  INV_X1 U19256 ( .A(n16133), .ZN(n16138) );
  AOI22_X1 U19257 ( .A1(n19054), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n19024), .ZN(n16134) );
  OAI21_X1 U19258 ( .B1(n9807), .B2(n19831), .A(n16134), .ZN(n16137) );
  NOR2_X1 U19259 ( .A1(n16135), .A2(n19042), .ZN(n16136) );
  AOI211_X1 U19260 ( .C1(n19066), .C2(n16138), .A(n16137), .B(n16136), .ZN(
        n16142) );
  OAI211_X1 U19261 ( .C1(n14054), .C2(n16140), .A(n19050), .B(n16139), .ZN(
        n16141) );
  OAI211_X1 U19262 ( .C1(n19063), .C2(n16143), .A(n16142), .B(n16141), .ZN(
        P2_U2828) );
  AOI22_X1 U19263 ( .A1(P2_REIP_REG_26__SCAN_IN), .A2(n9882), .B1(
        P2_EBX_REG_26__SCAN_IN), .B2(n19054), .ZN(n16154) );
  AOI22_X1 U19264 ( .A1(n16144), .A2(n19060), .B1(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n19003), .ZN(n16153) );
  INV_X1 U19265 ( .A(n16145), .ZN(n16146) );
  AOI22_X1 U19266 ( .A1(n16147), .A2(n19066), .B1(n16146), .B2(n18980), .ZN(
        n16152) );
  OAI211_X1 U19267 ( .C1(n16150), .C2(n16149), .A(n19050), .B(n16148), .ZN(
        n16151) );
  NAND4_X1 U19268 ( .A1(n16154), .A2(n16153), .A3(n16152), .A4(n16151), .ZN(
        P2_U2829) );
  AOI22_X1 U19269 ( .A1(P2_REIP_REG_25__SCAN_IN), .A2(n9882), .B1(
        P2_EBX_REG_25__SCAN_IN), .B2(n19054), .ZN(n16167) );
  OAI22_X1 U19270 ( .A1(n16156), .A2(n19042), .B1(n16155), .B2(n19057), .ZN(
        n16157) );
  INV_X1 U19271 ( .A(n16157), .ZN(n16166) );
  INV_X1 U19272 ( .A(n16158), .ZN(n16160) );
  AOI22_X1 U19273 ( .A1(n16160), .A2(n19066), .B1(n18980), .B2(n16159), .ZN(
        n16165) );
  OAI211_X1 U19274 ( .C1(n16163), .C2(n16162), .A(n19050), .B(n16161), .ZN(
        n16164) );
  NAND4_X1 U19275 ( .A1(n16167), .A2(n16166), .A3(n16165), .A4(n16164), .ZN(
        P2_U2830) );
  AOI22_X1 U19276 ( .A1(n19054), .A2(P2_EBX_REG_24__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n19024), .ZN(n16168) );
  OAI21_X1 U19277 ( .B1(n16169), .B2(n19036), .A(n16168), .ZN(n16172) );
  NOR2_X1 U19278 ( .A1(n16170), .A2(n19042), .ZN(n16171) );
  AOI211_X1 U19279 ( .C1(n9882), .C2(P2_REIP_REG_24__SCAN_IN), .A(n16172), .B(
        n16171), .ZN(n16176) );
  OAI211_X1 U19280 ( .C1(n16213), .C2(n16174), .A(n19050), .B(n16173), .ZN(
        n16175) );
  OAI211_X1 U19281 ( .C1(n19063), .C2(n16177), .A(n16176), .B(n16175), .ZN(
        P2_U2831) );
  AOI22_X1 U19282 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n9882), .B1(
        P2_EBX_REG_23__SCAN_IN), .B2(n19054), .ZN(n16188) );
  AOI22_X1 U19283 ( .A1(n16178), .A2(n19060), .B1(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n19024), .ZN(n16187) );
  INV_X1 U19284 ( .A(n16179), .ZN(n16181) );
  AOI22_X1 U19285 ( .A1(n16181), .A2(n19066), .B1(n18980), .B2(n16180), .ZN(
        n16186) );
  OAI211_X1 U19286 ( .C1(n16184), .C2(n16183), .A(n19050), .B(n16182), .ZN(
        n16185) );
  NAND4_X1 U19287 ( .A1(n16188), .A2(n16187), .A3(n16186), .A4(n16185), .ZN(
        P2_U2832) );
  AOI22_X1 U19288 ( .A1(n19076), .A2(n16189), .B1(P2_EAX_REG_22__SCAN_IN), 
        .B2(n19126), .ZN(n16194) );
  AOI22_X1 U19289 ( .A1(n19078), .A2(BUF1_REG_22__SCAN_IN), .B1(n19077), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n16193) );
  AOI22_X1 U19290 ( .A1(n16191), .A2(n19131), .B1(n19127), .B2(n16190), .ZN(
        n16192) );
  NAND3_X1 U19291 ( .A1(n16194), .A2(n16193), .A3(n16192), .ZN(P2_U2897) );
  AOI22_X1 U19292 ( .A1(n19076), .A2(n19260), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n19126), .ZN(n16198) );
  AOI22_X1 U19293 ( .A1(n19078), .A2(BUF1_REG_20__SCAN_IN), .B1(n19077), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n16197) );
  AOI22_X1 U19294 ( .A1(n16195), .A2(n19131), .B1(n19127), .B2(n18926), .ZN(
        n16196) );
  NAND3_X1 U19295 ( .A1(n16198), .A2(n16197), .A3(n16196), .ZN(P2_U2899) );
  AOI22_X1 U19296 ( .A1(n19076), .A2(n16199), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n19126), .ZN(n16204) );
  AOI22_X1 U19297 ( .A1(n19078), .A2(BUF1_REG_18__SCAN_IN), .B1(n19077), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n16203) );
  INV_X1 U19298 ( .A(n16200), .ZN(n18951) );
  AOI22_X1 U19299 ( .A1(n16201), .A2(n19131), .B1(n19127), .B2(n18951), .ZN(
        n16202) );
  NAND3_X1 U19300 ( .A1(n16204), .A2(n16203), .A3(n16202), .ZN(P2_U2901) );
  AOI22_X1 U19301 ( .A1(n16247), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19030), .ZN(n16212) );
  NAND2_X1 U19302 ( .A1(n16205), .A2(n11305), .ZN(n16208) );
  NAND2_X1 U19303 ( .A1(n16206), .A2(n19207), .ZN(n16207) );
  OAI211_X1 U19304 ( .C1(n16209), .C2(n16265), .A(n16208), .B(n16207), .ZN(
        n16210) );
  INV_X1 U19305 ( .A(n16210), .ZN(n16211) );
  OAI211_X1 U19306 ( .C1(n16262), .C2(n16213), .A(n16212), .B(n16211), .ZN(
        P2_U2990) );
  AOI22_X1 U19307 ( .A1(n16247), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19030), .ZN(n16222) );
  NAND3_X1 U19308 ( .A1(n16215), .A2(n19204), .A3(n16214), .ZN(n16220) );
  NAND2_X1 U19309 ( .A1(n16216), .A2(n11305), .ZN(n16219) );
  NAND2_X1 U19310 ( .A1(n19207), .A2(n16217), .ZN(n16218) );
  AND3_X1 U19311 ( .A1(n16220), .A2(n16219), .A3(n16218), .ZN(n16221) );
  OAI211_X1 U19312 ( .C1(n16262), .C2(n16223), .A(n16222), .B(n16221), .ZN(
        P2_U2992) );
  AOI22_X1 U19313 ( .A1(n16247), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n19030), .ZN(n16228) );
  OAI222_X1 U19314 ( .A1(n18949), .A2(n13644), .B1(n16263), .B2(n16225), .C1(
        n16265), .C2(n16224), .ZN(n16226) );
  INV_X1 U19315 ( .A(n16226), .ZN(n16227) );
  OAI211_X1 U19316 ( .C1(n16262), .C2(n18945), .A(n16228), .B(n16227), .ZN(
        P2_U2996) );
  AOI22_X1 U19317 ( .A1(n16247), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19030), .ZN(n16236) );
  NAND2_X1 U19318 ( .A1(n16230), .A2(n16229), .ZN(n16231) );
  XNOR2_X1 U19319 ( .A(n16232), .B(n16231), .ZN(n16289) );
  AOI21_X1 U19320 ( .B1(n15088), .B2(n16233), .A(n11284), .ZN(n16288) );
  INV_X1 U19321 ( .A(n16234), .ZN(n16287) );
  AOI222_X1 U19322 ( .A1(n16289), .A2(n11305), .B1(n16288), .B2(n19204), .C1(
        n19207), .C2(n16287), .ZN(n16235) );
  OAI211_X1 U19323 ( .C1(n16262), .C2(n16237), .A(n16236), .B(n16235), .ZN(
        P2_U3000) );
  AOI22_X1 U19324 ( .A1(n16247), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19030), .ZN(n16245) );
  NOR2_X1 U19325 ( .A1(n16239), .A2(n16238), .ZN(n16241) );
  XOR2_X1 U19326 ( .A(n16241), .B(n16240), .Z(n16302) );
  OAI21_X1 U19327 ( .B1(n16242), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15089), .ZN(n16300) );
  OAI22_X1 U19328 ( .A1(n16300), .A2(n16265), .B1(n13644), .B2(n16298), .ZN(
        n16243) );
  AOI21_X1 U19329 ( .B1(n11305), .B2(n16302), .A(n16243), .ZN(n16244) );
  OAI211_X1 U19330 ( .C1(n16262), .C2(n16246), .A(n16245), .B(n16244), .ZN(
        P2_U3002) );
  AOI22_X1 U19331 ( .A1(n16247), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19030), .ZN(n16260) );
  NAND2_X1 U19332 ( .A1(n16249), .A2(n16248), .ZN(n16250) );
  NAND2_X1 U19333 ( .A1(n16251), .A2(n16250), .ZN(n16317) );
  NAND2_X1 U19334 ( .A1(n16313), .A2(n19207), .ZN(n16257) );
  NAND2_X1 U19335 ( .A1(n15303), .A2(n16252), .ZN(n16255) );
  NAND2_X1 U19336 ( .A1(n9867), .A2(n16253), .ZN(n16254) );
  XNOR2_X1 U19337 ( .A(n16255), .B(n16254), .ZN(n16314) );
  NAND2_X1 U19338 ( .A1(n16314), .A2(n11305), .ZN(n16256) );
  OAI211_X1 U19339 ( .C1(n16317), .C2(n16265), .A(n16257), .B(n16256), .ZN(
        n16258) );
  INV_X1 U19340 ( .A(n16258), .ZN(n16259) );
  OAI211_X1 U19341 ( .C1(n16262), .C2(n16261), .A(n16260), .B(n16259), .ZN(
        P2_U3004) );
  AOI22_X1 U19342 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19030), .B1(n19203), 
        .B2(n19007), .ZN(n16270) );
  OAI22_X1 U19343 ( .A1(n16266), .A2(n16265), .B1(n16264), .B2(n16263), .ZN(
        n16267) );
  AOI21_X1 U19344 ( .B1(n19207), .B2(n16268), .A(n16267), .ZN(n16269) );
  OAI211_X1 U19345 ( .C1(n19212), .C2(n16271), .A(n16270), .B(n16269), .ZN(
        P2_U3005) );
  AOI22_X1 U19346 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19030), .B1(n19203), 
        .B2(n16272), .ZN(n16281) );
  XOR2_X1 U19347 ( .A(n16273), .B(n16274), .Z(n16324) );
  INV_X1 U19348 ( .A(n16276), .ZN(n16278) );
  NOR2_X1 U19349 ( .A1(n16278), .A2(n16277), .ZN(n16279) );
  XNOR2_X1 U19350 ( .A(n16275), .B(n16279), .ZN(n16322) );
  AOI222_X1 U19351 ( .A1(n16324), .A2(n19204), .B1(n11305), .B2(n16322), .C1(
        n19207), .C2(n16321), .ZN(n16280) );
  OAI211_X1 U19352 ( .C1(n19212), .C2(n16282), .A(n16281), .B(n16280), .ZN(
        P2_U3006) );
  NOR2_X1 U19353 ( .A1(n15334), .A2(n19813), .ZN(n16286) );
  AOI21_X1 U19354 ( .B1(n16284), .B2(n16283), .A(n16233), .ZN(n16285) );
  AOI211_X1 U19355 ( .C1(n19087), .C2(n19228), .A(n16286), .B(n16285), .ZN(
        n16291) );
  AOI222_X1 U19356 ( .A1(n16289), .A2(n16323), .B1(n16288), .B2(n19233), .C1(
        n19220), .C2(n16287), .ZN(n16290) );
  OAI211_X1 U19357 ( .C1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n16292), .A(
        n16291), .B(n16290), .ZN(P2_U3032) );
  AOI21_X1 U19358 ( .B1(n16295), .B2(n16294), .A(n16293), .ZN(n16306) );
  NOR2_X1 U19359 ( .A1(n15334), .A2(n14789), .ZN(n16297) );
  AOI211_X1 U19360 ( .C1(n19093), .C2(n19228), .A(n16297), .B(n16296), .ZN(
        n16304) );
  OAI22_X1 U19361 ( .A1(n16300), .A2(n16318), .B1(n16299), .B2(n16298), .ZN(
        n16301) );
  AOI21_X1 U19362 ( .B1(n16323), .B2(n16302), .A(n16301), .ZN(n16303) );
  OAI211_X1 U19363 ( .C1(n16306), .C2(n16305), .A(n16304), .B(n16303), .ZN(
        P2_U3034) );
  NAND2_X1 U19364 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16307), .ZN(
        n16310) );
  NAND2_X1 U19365 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n19030), .ZN(n16308) );
  OAI221_X1 U19366 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16310), 
        .C1(n16248), .C2(n16309), .A(n16308), .ZN(n16311) );
  AOI21_X1 U19367 ( .B1(n16312), .B2(n19228), .A(n16311), .ZN(n16316) );
  AOI22_X1 U19368 ( .A1(n16314), .A2(n16323), .B1(n19220), .B2(n16313), .ZN(
        n16315) );
  OAI211_X1 U19369 ( .C1(n16318), .C2(n16317), .A(n16316), .B(n16315), .ZN(
        P2_U3036) );
  AOI22_X1 U19370 ( .A1(n16320), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n19228), .B2(n16319), .ZN(n16331) );
  AOI222_X1 U19371 ( .A1(n16324), .A2(n19233), .B1(n16323), .B2(n16322), .C1(
        n19220), .C2(n16321), .ZN(n16330) );
  NAND2_X1 U19372 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19030), .ZN(n16329) );
  OAI221_X1 U19373 ( .B1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16327), .C2(n16326), .A(
        n16325), .ZN(n16328) );
  NAND4_X1 U19374 ( .A1(n16331), .A2(n16330), .A3(n16329), .A4(n16328), .ZN(
        P2_U3038) );
  OAI211_X1 U19375 ( .C1(n16335), .C2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n16332), .ZN(n16333) );
  OAI21_X1 U19376 ( .B1(n16340), .B2(n19861), .A(n16333), .ZN(n16334) );
  AOI211_X1 U19377 ( .C1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n16335), .A(
        n16354), .B(n16334), .ZN(n16339) );
  MUX2_X1 U19378 ( .A(n16337), .B(n16336), .S(n16354), .Z(n16343) );
  NOR2_X1 U19379 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19347) );
  AND2_X1 U19380 ( .A1(n16343), .A2(n19347), .ZN(n16338) );
  OAI22_X1 U19381 ( .A1(n16339), .A2(n16338), .B1(n16343), .B2(n19868), .ZN(
        n16342) );
  MUX2_X1 U19382 ( .A(n16340), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n16354), .Z(n16344) );
  INV_X1 U19383 ( .A(n16344), .ZN(n16341) );
  AOI221_X1 U19384 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n16342), 
        .C1(n16341), .C2(n16342), .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n16358) );
  NAND2_X1 U19385 ( .A1(n16344), .A2(n16343), .ZN(n16356) );
  OAI21_X1 U19386 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n16345), .ZN(n16350) );
  INV_X1 U19387 ( .A(n16346), .ZN(n16347) );
  NAND3_X1 U19388 ( .A1(n16348), .A2(n9788), .A3(n16347), .ZN(n16349) );
  NAND4_X1 U19389 ( .A1(n16352), .A2(n16351), .A3(n16350), .A4(n16349), .ZN(
        n16353) );
  AOI21_X1 U19390 ( .B1(n16354), .B2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n16353), .ZN(n16355) );
  NAND2_X1 U19391 ( .A1(n16356), .A2(n16355), .ZN(n16357) );
  OR2_X1 U19392 ( .A1(n16358), .A2(n16357), .ZN(n16369) );
  INV_X1 U19393 ( .A(n16369), .ZN(n16376) );
  AOI211_X1 U19394 ( .C1(n16377), .C2(n16361), .A(n16360), .B(n16359), .ZN(
        n16374) );
  INV_X1 U19395 ( .A(n16362), .ZN(n16366) );
  NAND2_X1 U19396 ( .A1(n16363), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n16364) );
  AOI21_X1 U19397 ( .B1(n16366), .B2(n16365), .A(n16364), .ZN(n16370) );
  AOI22_X1 U19398 ( .A1(n16368), .A2(n16367), .B1(n19785), .B2(n16370), .ZN(
        n16372) );
  OAI21_X1 U19399 ( .B1(n16369), .B2(P2_STATE2_REG_1__SCAN_IN), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n16371) );
  INV_X1 U19400 ( .A(n19763), .ZN(n19766) );
  NAND2_X1 U19401 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19766), .ZN(n16378) );
  OAI21_X1 U19402 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n16372), .A(n16378), 
        .ZN(n16373) );
  OAI211_X1 U19403 ( .C1(n16376), .C2(n16375), .A(n16374), .B(n16373), .ZN(
        P2_U3176) );
  AOI21_X1 U19404 ( .B1(n16378), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n16377), 
        .ZN(n16379) );
  INV_X1 U19405 ( .A(n16379), .ZN(P2_U3593) );
  INV_X1 U19406 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18833) );
  AOI22_X1 U19407 ( .A1(n17674), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        n18833), .B2(n17781), .ZN(n16388) );
  AND2_X1 U19408 ( .A1(n17781), .A2(n16381), .ZN(n16386) );
  OAI21_X1 U19409 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n16426), .A(
        n16382), .ZN(n16383) );
  OAI22_X1 U19410 ( .A1(n16386), .A2(n16383), .B1(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18833), .ZN(n16387) );
  NAND2_X1 U19411 ( .A1(n16388), .A2(n16384), .ZN(n16385) );
  OAI22_X1 U19412 ( .A1(n16388), .A2(n16387), .B1(n16386), .B2(n16385), .ZN(
        n16435) );
  INV_X1 U19413 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18808) );
  NOR2_X1 U19414 ( .A1(n15697), .A2(n18808), .ZN(n16428) );
  INV_X1 U19415 ( .A(n17602), .ZN(n16389) );
  OR2_X1 U19416 ( .A1(n16390), .A2(n17716), .ZN(n16402) );
  INV_X1 U19417 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16599) );
  XOR2_X1 U19418 ( .A(n16599), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16392) );
  NOR2_X1 U19419 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17602), .ZN(
        n16413) );
  INV_X1 U19420 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n20928) );
  NAND2_X1 U19421 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17548), .ZN(
        n17518) );
  NOR2_X1 U19422 ( .A1(n20928), .A2(n17518), .ZN(n16581) );
  NAND3_X1 U19423 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A3(n16581), .ZN(n16577) );
  AOI22_X1 U19424 ( .A1(n17713), .A2(n16577), .B1(n18607), .B2(n16390), .ZN(
        n16391) );
  NAND2_X1 U19425 ( .A1(n16391), .A2(n17882), .ZN(n16414) );
  NOR2_X1 U19426 ( .A1(n16413), .A2(n16414), .ZN(n16401) );
  OAI22_X1 U19427 ( .A1(n16402), .A2(n16392), .B1(n16401), .B2(n16599), .ZN(
        n16393) );
  AOI211_X1 U19428 ( .C1(n17538), .C2(n16907), .A(n16428), .B(n16393), .ZN(
        n16398) );
  NAND2_X1 U19429 ( .A1(n16405), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16395) );
  XNOR2_X1 U19430 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n16395), .ZN(
        n16432) );
  NAND2_X1 U19431 ( .A1(n16406), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16396) );
  XNOR2_X1 U19432 ( .A(n16396), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16431) );
  AOI22_X1 U19433 ( .A1(n17874), .A2(n16432), .B1(n17711), .B2(n16431), .ZN(
        n16397) );
  OAI211_X1 U19434 ( .C1(n17794), .C2(n16435), .A(n16398), .B(n16397), .ZN(
        P3_U2799) );
  XOR2_X1 U19435 ( .A(n16412), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16602) );
  NOR4_X1 U19436 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16399), .A3(
        n17543), .A4(n17685), .ZN(n16404) );
  INV_X1 U19437 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16603) );
  NAND2_X1 U19438 ( .A1(n9760), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16400) );
  OAI221_X1 U19439 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16402), .C1(
        n16603), .C2(n16401), .A(n16400), .ZN(n16403) );
  AOI211_X1 U19440 ( .C1(n17538), .C2(n16602), .A(n16404), .B(n16403), .ZN(
        n16408) );
  NOR2_X1 U19441 ( .A1(n16405), .A2(n17886), .ZN(n16410) );
  NOR2_X1 U19442 ( .A1(n16406), .A2(n17789), .ZN(n16411) );
  OAI21_X1 U19443 ( .B1(n16410), .B2(n16411), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16407) );
  OAI211_X1 U19444 ( .C1(n16409), .C2(n17794), .A(n16408), .B(n16407), .ZN(
        P3_U2800) );
  INV_X1 U19445 ( .A(n16410), .ZN(n16423) );
  OAI21_X1 U19446 ( .B1(n16455), .B2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n16411), .ZN(n16418) );
  INV_X1 U19447 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16613) );
  AOI21_X1 U19448 ( .B1(n16613), .B2(n16577), .A(n16412), .ZN(n16612) );
  OAI21_X1 U19449 ( .B1(n17538), .B2(n16413), .A(n16612), .ZN(n16417) );
  OAI221_X1 U19450 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n16415), .C1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n18607), .A(n16414), .ZN(
        n16416) );
  NAND4_X1 U19451 ( .A1(n16419), .A2(n16418), .A3(n16417), .A4(n16416), .ZN(
        n16420) );
  AOI21_X1 U19452 ( .B1(n17748), .B2(n16421), .A(n16420), .ZN(n16422) );
  OAI221_X1 U19453 ( .B1(n16423), .B2(n16451), .C1(n16423), .C2(n16427), .A(
        n16422), .ZN(P3_U2801) );
  NAND2_X1 U19454 ( .A1(n18184), .A2(n18118), .ZN(n18191) );
  OAI21_X1 U19455 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18191), .A(
        n16424), .ZN(n16430) );
  NOR4_X1 U19456 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16427), .A3(
        n16426), .A4(n16425), .ZN(n16429) );
  AOI211_X1 U19457 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n16430), .A(
        n16429), .B(n16428), .ZN(n16434) );
  AOI22_X1 U19458 ( .A1(n16432), .A2(n18204), .B1(n16431), .B2(n18050), .ZN(
        n16433) );
  OAI211_X1 U19459 ( .C1(n18121), .C2(n16435), .A(n16434), .B(n16433), .ZN(
        P3_U2831) );
  NOR2_X1 U19460 ( .A1(n16437), .A2(n16436), .ZN(n18060) );
  OAI21_X1 U19461 ( .B1(n18664), .B2(n17945), .A(n16438), .ZN(n16439) );
  AOI21_X1 U19462 ( .B1(n18060), .B2(n18025), .A(n16439), .ZN(n17938) );
  NOR2_X1 U19463 ( .A1(n17938), .A2(n18205), .ZN(n17933) );
  NAND2_X1 U19464 ( .A1(n17614), .A2(n17933), .ZN(n17988) );
  NOR2_X1 U19465 ( .A1(n16440), .A2(n17988), .ZN(n17944) );
  AOI22_X1 U19466 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17781), .B1(
        n17674), .B2(n16458), .ZN(n17521) );
  AOI21_X1 U19467 ( .B1(n17944), .B2(n16444), .A(n16443), .ZN(n16465) );
  INV_X1 U19468 ( .A(n16445), .ZN(n16447) );
  INV_X1 U19469 ( .A(n16449), .ZN(n16453) );
  INV_X1 U19470 ( .A(n18664), .ZN(n18062) );
  INV_X1 U19471 ( .A(n16454), .ZN(n16457) );
  INV_X1 U19472 ( .A(n18060), .ZN(n18085) );
  OR2_X1 U19473 ( .A1(n16455), .A2(n18085), .ZN(n16456) );
  NAND2_X1 U19474 ( .A1(n16457), .A2(n16456), .ZN(n16461) );
  NOR2_X1 U19475 ( .A1(n9760), .A2(n16458), .ZN(n16460) );
  AND2_X1 U19476 ( .A1(n9760), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n16459) );
  NAND3_X1 U19477 ( .A1(n16462), .A2(n18083), .A3(n17521), .ZN(n16463) );
  OAI211_X1 U19478 ( .C1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n16465), .A(
        n16464), .B(n16463), .ZN(P3_U2834) );
  NOR3_X1 U19479 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16467) );
  NOR4_X1 U19480 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16466) );
  INV_X2 U19481 ( .A(n16544), .ZN(U215) );
  NAND4_X1 U19482 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16467), .A3(n16466), .A4(
        U215), .ZN(U213) );
  INV_X1 U19483 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n16549) );
  INV_X2 U19484 ( .A(U214), .ZN(n16510) );
  INV_X1 U19485 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16548) );
  OAI222_X1 U19486 ( .A1(U212), .A2(n16549), .B1(n16512), .B2(n20176), .C1(
        U214), .C2(n16548), .ZN(U216) );
  INV_X1 U19487 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20166) );
  AOI22_X1 U19488 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n16509), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n16510), .ZN(n16469) );
  OAI21_X1 U19489 ( .B1(n20166), .B2(n16512), .A(n16469), .ZN(U217) );
  AOI22_X1 U19490 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n16509), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n16510), .ZN(n16470) );
  OAI21_X1 U19491 ( .B1(n19264), .B2(n16512), .A(n16470), .ZN(U218) );
  INV_X1 U19492 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n19258) );
  AOI22_X1 U19493 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n16509), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n16510), .ZN(n16471) );
  OAI21_X1 U19494 ( .B1(n19258), .B2(n16512), .A(n16471), .ZN(U219) );
  AOI22_X1 U19495 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n16509), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n16510), .ZN(n16472) );
  OAI21_X1 U19496 ( .B1(n21078), .B2(n16512), .A(n16472), .ZN(U220) );
  INV_X1 U19497 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16474) );
  AOI22_X1 U19498 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n16509), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n16510), .ZN(n16473) );
  OAI21_X1 U19499 ( .B1(n16474), .B2(n16512), .A(n16473), .ZN(U221) );
  AOI22_X1 U19500 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n16509), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n16510), .ZN(n16475) );
  OAI21_X1 U19501 ( .B1(n14943), .B2(n16512), .A(n16475), .ZN(U222) );
  AOI22_X1 U19502 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n16509), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n16510), .ZN(n16476) );
  OAI21_X1 U19503 ( .B1(n20118), .B2(n16512), .A(n16476), .ZN(U223) );
  AOI22_X1 U19504 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n16509), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n16510), .ZN(n16477) );
  OAI21_X1 U19505 ( .B1(n16478), .B2(n16512), .A(n16477), .ZN(U224) );
  INV_X1 U19506 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n19270) );
  AOI22_X1 U19507 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n16509), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n16510), .ZN(n16479) );
  OAI21_X1 U19508 ( .B1(n19270), .B2(n16512), .A(n16479), .ZN(U225) );
  AOI22_X1 U19509 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n16509), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n16510), .ZN(n16480) );
  OAI21_X1 U19510 ( .B1(n14964), .B2(n16512), .A(n16480), .ZN(U226) );
  INV_X1 U19511 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n20155) );
  AOI22_X1 U19512 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n16509), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n16510), .ZN(n16481) );
  OAI21_X1 U19513 ( .B1(n20155), .B2(n16512), .A(n16481), .ZN(U227) );
  AOI22_X1 U19514 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n16509), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n16510), .ZN(n16482) );
  OAI21_X1 U19515 ( .B1(n14976), .B2(n16512), .A(n16482), .ZN(U228) );
  AOI22_X1 U19516 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n16509), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n16510), .ZN(n16483) );
  OAI21_X1 U19517 ( .B1(n20139), .B2(n16512), .A(n16483), .ZN(U229) );
  AOI22_X1 U19518 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n16509), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n16510), .ZN(n16484) );
  OAI21_X1 U19519 ( .B1(n13891), .B2(n16512), .A(n16484), .ZN(U230) );
  INV_X1 U19520 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16486) );
  AOI22_X1 U19521 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n16509), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n16510), .ZN(n16485) );
  OAI21_X1 U19522 ( .B1(n16486), .B2(n16512), .A(n16485), .ZN(U231) );
  AOI22_X1 U19523 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16510), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16509), .ZN(n16487) );
  OAI21_X1 U19524 ( .B1(n13292), .B2(n16512), .A(n16487), .ZN(U232) );
  INV_X1 U19525 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n16489) );
  AOI22_X1 U19526 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16510), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16509), .ZN(n16488) );
  OAI21_X1 U19527 ( .B1(n16489), .B2(n16512), .A(n16488), .ZN(U233) );
  AOI22_X1 U19528 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16510), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16509), .ZN(n16490) );
  OAI21_X1 U19529 ( .B1(n13094), .B2(n16512), .A(n16490), .ZN(U234) );
  INV_X1 U19530 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n21046) );
  INV_X1 U19531 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n20866) );
  OAI222_X1 U19532 ( .A1(U212), .A2(n21046), .B1(n16512), .B2(n20866), .C1(
        U214), .C2(n13535), .ZN(U235) );
  AOI22_X1 U19533 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16510), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16509), .ZN(n16491) );
  OAI21_X1 U19534 ( .B1(n13085), .B2(n16512), .A(n16491), .ZN(U236) );
  INV_X1 U19535 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16493) );
  AOI22_X1 U19536 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16510), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16509), .ZN(n16492) );
  OAI21_X1 U19537 ( .B1(n16493), .B2(n16512), .A(n16492), .ZN(U237) );
  AOI22_X1 U19538 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16510), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16509), .ZN(n16494) );
  OAI21_X1 U19539 ( .B1(n16495), .B2(n16512), .A(n16494), .ZN(U238) );
  AOI22_X1 U19540 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16510), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16509), .ZN(n16496) );
  OAI21_X1 U19541 ( .B1(n13108), .B2(n16512), .A(n16496), .ZN(U239) );
  INV_X1 U19542 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16521) );
  INV_X1 U19543 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16497) );
  OAI222_X1 U19544 ( .A1(U212), .A2(n16521), .B1(n16512), .B2(n16497), .C1(
        U214), .C2(n13542), .ZN(U240) );
  INV_X1 U19545 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n20877) );
  AOI22_X1 U19546 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16510), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16509), .ZN(n16498) );
  OAI21_X1 U19547 ( .B1(n20877), .B2(n16512), .A(n16498), .ZN(U241) );
  INV_X1 U19548 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16500) );
  AOI22_X1 U19549 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16510), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16509), .ZN(n16499) );
  OAI21_X1 U19550 ( .B1(n16500), .B2(n16512), .A(n16499), .ZN(U242) );
  AOI22_X1 U19551 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16510), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16509), .ZN(n16501) );
  OAI21_X1 U19552 ( .B1(n16502), .B2(n16512), .A(n16501), .ZN(U243) );
  INV_X1 U19553 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16504) );
  AOI22_X1 U19554 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16510), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16509), .ZN(n16503) );
  OAI21_X1 U19555 ( .B1(n16504), .B2(n16512), .A(n16503), .ZN(U244) );
  AOI22_X1 U19556 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16510), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16509), .ZN(n16505) );
  OAI21_X1 U19557 ( .B1(n16506), .B2(n16512), .A(n16505), .ZN(U245) );
  INV_X1 U19558 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16508) );
  AOI22_X1 U19559 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16510), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16509), .ZN(n16507) );
  OAI21_X1 U19560 ( .B1(n16508), .B2(n16512), .A(n16507), .ZN(U246) );
  AOI22_X1 U19561 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16510), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16509), .ZN(n16511) );
  OAI21_X1 U19562 ( .B1(n16513), .B2(n16512), .A(n16511), .ZN(U247) );
  INV_X1 U19563 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n16514) );
  AOI22_X1 U19564 ( .A1(n16544), .A2(n16514), .B1(n18218), .B2(U215), .ZN(U251) );
  OAI22_X1 U19565 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16544), .ZN(n16515) );
  INV_X1 U19566 ( .A(n16515), .ZN(U252) );
  INV_X1 U19567 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16516) );
  AOI22_X1 U19568 ( .A1(n16544), .A2(n16516), .B1(n18231), .B2(U215), .ZN(U253) );
  INV_X1 U19569 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16517) );
  INV_X1 U19570 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18237) );
  AOI22_X1 U19571 ( .A1(n16544), .A2(n16517), .B1(n18237), .B2(U215), .ZN(U254) );
  INV_X1 U19572 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16518) );
  AOI22_X1 U19573 ( .A1(n16544), .A2(n16518), .B1(n18241), .B2(U215), .ZN(U255) );
  INV_X1 U19574 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16519) );
  INV_X1 U19575 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18246) );
  AOI22_X1 U19576 ( .A1(n16544), .A2(n16519), .B1(n18246), .B2(U215), .ZN(U256) );
  INV_X1 U19577 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16520) );
  INV_X1 U19578 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18252) );
  AOI22_X1 U19579 ( .A1(n16544), .A2(n16520), .B1(n18252), .B2(U215), .ZN(U257) );
  INV_X1 U19580 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18257) );
  AOI22_X1 U19581 ( .A1(n16546), .A2(n16521), .B1(n18257), .B2(U215), .ZN(U258) );
  OAI22_X1 U19582 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16546), .ZN(n16522) );
  INV_X1 U19583 ( .A(n16522), .ZN(U259) );
  INV_X1 U19584 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16523) );
  INV_X1 U19585 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17496) );
  AOI22_X1 U19586 ( .A1(n16546), .A2(n16523), .B1(n17496), .B2(U215), .ZN(U260) );
  INV_X1 U19587 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n16524) );
  INV_X1 U19588 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17498) );
  AOI22_X1 U19589 ( .A1(n16544), .A2(n16524), .B1(n17498), .B2(U215), .ZN(U261) );
  OAI22_X1 U19590 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16544), .ZN(n16525) );
  INV_X1 U19591 ( .A(n16525), .ZN(U262) );
  INV_X1 U19592 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17503) );
  AOI22_X1 U19593 ( .A1(n16544), .A2(n21046), .B1(n17503), .B2(U215), .ZN(U263) );
  INV_X1 U19594 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16526) );
  INV_X1 U19595 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17508) );
  AOI22_X1 U19596 ( .A1(n16544), .A2(n16526), .B1(n17508), .B2(U215), .ZN(U264) );
  OAI22_X1 U19597 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16544), .ZN(n16527) );
  INV_X1 U19598 ( .A(n16527), .ZN(U265) );
  INV_X1 U19599 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n16528) );
  INV_X1 U19600 ( .A(BUF2_REG_15__SCAN_IN), .ZN(n21015) );
  AOI22_X1 U19601 ( .A1(n16544), .A2(n16528), .B1(n21015), .B2(U215), .ZN(U266) );
  OAI22_X1 U19602 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16546), .ZN(n16529) );
  INV_X1 U19603 ( .A(n16529), .ZN(U267) );
  INV_X1 U19604 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n16530) );
  AOI22_X1 U19605 ( .A1(n16546), .A2(n16530), .B1(n13890), .B2(U215), .ZN(U268) );
  INV_X1 U19606 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n16531) );
  AOI22_X1 U19607 ( .A1(n16544), .A2(n16531), .B1(n18233), .B2(U215), .ZN(U269) );
  OAI22_X1 U19608 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16546), .ZN(n16532) );
  INV_X1 U19609 ( .A(n16532), .ZN(U270) );
  OAI22_X1 U19610 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16544), .ZN(n16533) );
  INV_X1 U19611 ( .A(n16533), .ZN(U271) );
  INV_X1 U19612 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n16534) );
  AOI22_X1 U19613 ( .A1(n16546), .A2(n16534), .B1(n14963), .B2(U215), .ZN(U272) );
  INV_X1 U19614 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n16535) );
  INV_X1 U19615 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n19269) );
  AOI22_X1 U19616 ( .A1(n16544), .A2(n16535), .B1(n19269), .B2(U215), .ZN(U273) );
  OAI22_X1 U19617 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16546), .ZN(n16536) );
  INV_X1 U19618 ( .A(n16536), .ZN(U274) );
  INV_X1 U19619 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n16537) );
  AOI22_X1 U19620 ( .A1(n16546), .A2(n16537), .B1(n18223), .B2(U215), .ZN(U275) );
  OAI22_X1 U19621 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16544), .ZN(n16538) );
  INV_X1 U19622 ( .A(n16538), .ZN(U276) );
  OAI22_X1 U19623 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16544), .ZN(n16539) );
  INV_X1 U19624 ( .A(n16539), .ZN(U277) );
  INV_X1 U19625 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n16540) );
  INV_X1 U19626 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n19253) );
  AOI22_X1 U19627 ( .A1(n16544), .A2(n16540), .B1(n19253), .B2(U215), .ZN(U278) );
  INV_X1 U19628 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n16541) );
  INV_X1 U19629 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n19257) );
  AOI22_X1 U19630 ( .A1(n16544), .A2(n16541), .B1(n19257), .B2(U215), .ZN(U279) );
  INV_X1 U19631 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n16542) );
  INV_X1 U19632 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n21050) );
  AOI22_X1 U19633 ( .A1(n16544), .A2(n16542), .B1(n21050), .B2(U215), .ZN(U280) );
  INV_X1 U19634 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n16543) );
  INV_X1 U19635 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n18251) );
  AOI22_X1 U19636 ( .A1(n16544), .A2(n16543), .B1(n18251), .B2(U215), .ZN(U281) );
  INV_X1 U19637 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n21051) );
  AOI22_X1 U19638 ( .A1(n16546), .A2(n16549), .B1(n21051), .B2(U215), .ZN(U282) );
  INV_X1 U19639 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16547) );
  AOI222_X1 U19640 ( .A1(n16549), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n16548), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .C1(n16547), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16550) );
  INV_X2 U19641 ( .A(n16552), .ZN(n16551) );
  INV_X1 U19642 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18768) );
  INV_X1 U19643 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19809) );
  AOI22_X1 U19644 ( .A1(n16551), .A2(n18768), .B1(n19809), .B2(n16552), .ZN(
        U347) );
  INV_X1 U19645 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18766) );
  INV_X1 U19646 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n21079) );
  AOI22_X1 U19647 ( .A1(n16550), .A2(n18766), .B1(n21079), .B2(n16552), .ZN(
        U348) );
  INV_X1 U19648 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18763) );
  INV_X1 U19649 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19806) );
  AOI22_X1 U19650 ( .A1(n16551), .A2(n18763), .B1(n19806), .B2(n16552), .ZN(
        U349) );
  INV_X1 U19651 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18762) );
  INV_X1 U19652 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19804) );
  AOI22_X1 U19653 ( .A1(n16551), .A2(n18762), .B1(n19804), .B2(n16552), .ZN(
        U350) );
  INV_X1 U19654 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18760) );
  INV_X1 U19655 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19802) );
  AOI22_X1 U19656 ( .A1(n16551), .A2(n18760), .B1(n19802), .B2(n16552), .ZN(
        U351) );
  INV_X1 U19657 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18757) );
  INV_X1 U19658 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19800) );
  AOI22_X1 U19659 ( .A1(n16551), .A2(n18757), .B1(n19800), .B2(n16552), .ZN(
        U352) );
  INV_X1 U19660 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18756) );
  INV_X1 U19661 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20896) );
  AOI22_X1 U19662 ( .A1(n16551), .A2(n18756), .B1(n20896), .B2(n16552), .ZN(
        U353) );
  INV_X1 U19663 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18753) );
  AOI22_X1 U19664 ( .A1(n16551), .A2(n18753), .B1(n19798), .B2(n16552), .ZN(
        U354) );
  INV_X1 U19665 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18807) );
  INV_X1 U19666 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19837) );
  AOI22_X1 U19667 ( .A1(n16551), .A2(n18807), .B1(n19837), .B2(n16552), .ZN(
        U355) );
  INV_X1 U19668 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18805) );
  INV_X1 U19669 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19834) );
  AOI22_X1 U19670 ( .A1(n16551), .A2(n18805), .B1(n19834), .B2(n16552), .ZN(
        U356) );
  INV_X1 U19671 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18803) );
  INV_X1 U19672 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19832) );
  AOI22_X1 U19673 ( .A1(n16551), .A2(n18803), .B1(n19832), .B2(n16552), .ZN(
        U357) );
  INV_X1 U19674 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18799) );
  INV_X1 U19675 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19830) );
  AOI22_X1 U19676 ( .A1(n16551), .A2(n18799), .B1(n19830), .B2(n16552), .ZN(
        U358) );
  INV_X1 U19677 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18798) );
  INV_X1 U19678 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19829) );
  AOI22_X1 U19679 ( .A1(n16551), .A2(n18798), .B1(n19829), .B2(n16552), .ZN(
        U359) );
  INV_X1 U19680 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18797) );
  INV_X1 U19681 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19828) );
  AOI22_X1 U19682 ( .A1(n16551), .A2(n18797), .B1(n19828), .B2(n16552), .ZN(
        U360) );
  INV_X1 U19683 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18796) );
  INV_X1 U19684 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19827) );
  AOI22_X1 U19685 ( .A1(n16551), .A2(n18796), .B1(n19827), .B2(n16552), .ZN(
        U361) );
  INV_X1 U19686 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18793) );
  INV_X1 U19687 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19826) );
  AOI22_X1 U19688 ( .A1(n16551), .A2(n18793), .B1(n19826), .B2(n16552), .ZN(
        U362) );
  INV_X1 U19689 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18792) );
  INV_X1 U19690 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n21085) );
  AOI22_X1 U19691 ( .A1(n16551), .A2(n18792), .B1(n21085), .B2(n16552), .ZN(
        U363) );
  INV_X1 U19692 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18789) );
  INV_X1 U19693 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19824) );
  AOI22_X1 U19694 ( .A1(n16551), .A2(n18789), .B1(n19824), .B2(n16552), .ZN(
        U364) );
  INV_X1 U19695 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18752) );
  INV_X1 U19696 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19796) );
  AOI22_X1 U19697 ( .A1(n16551), .A2(n18752), .B1(n19796), .B2(n16552), .ZN(
        U365) );
  INV_X1 U19698 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18787) );
  INV_X1 U19699 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19822) );
  AOI22_X1 U19700 ( .A1(n16551), .A2(n18787), .B1(n19822), .B2(n16552), .ZN(
        U366) );
  INV_X1 U19701 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18786) );
  INV_X1 U19702 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19821) );
  AOI22_X1 U19703 ( .A1(n16551), .A2(n18786), .B1(n19821), .B2(n16552), .ZN(
        U367) );
  INV_X1 U19704 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18784) );
  INV_X1 U19705 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19820) );
  AOI22_X1 U19706 ( .A1(n16551), .A2(n18784), .B1(n19820), .B2(n16552), .ZN(
        U368) );
  INV_X1 U19707 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18782) );
  INV_X1 U19708 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19819) );
  AOI22_X1 U19709 ( .A1(n16551), .A2(n18782), .B1(n19819), .B2(n16552), .ZN(
        U369) );
  INV_X1 U19710 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18780) );
  INV_X1 U19711 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19817) );
  AOI22_X1 U19712 ( .A1(n16551), .A2(n18780), .B1(n19817), .B2(n16552), .ZN(
        U370) );
  INV_X1 U19713 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18778) );
  INV_X1 U19714 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19815) );
  AOI22_X1 U19715 ( .A1(n16550), .A2(n18778), .B1(n19815), .B2(n16552), .ZN(
        U371) );
  INV_X1 U19716 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18775) );
  INV_X1 U19717 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19814) );
  AOI22_X1 U19718 ( .A1(n16551), .A2(n18775), .B1(n19814), .B2(n16552), .ZN(
        U372) );
  INV_X1 U19719 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18774) );
  INV_X1 U19720 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19812) );
  AOI22_X1 U19721 ( .A1(n16551), .A2(n18774), .B1(n19812), .B2(n16552), .ZN(
        U373) );
  INV_X1 U19722 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18772) );
  INV_X1 U19723 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19811) );
  AOI22_X1 U19724 ( .A1(n16551), .A2(n18772), .B1(n19811), .B2(n16552), .ZN(
        U374) );
  INV_X1 U19725 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18770) );
  INV_X1 U19726 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19810) );
  AOI22_X1 U19727 ( .A1(n16550), .A2(n18770), .B1(n19810), .B2(n16552), .ZN(
        U375) );
  INV_X1 U19728 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18750) );
  INV_X1 U19729 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19794) );
  AOI22_X1 U19730 ( .A1(n16550), .A2(n18750), .B1(n19794), .B2(n16552), .ZN(
        U376) );
  INV_X1 U19731 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16554) );
  NAND2_X1 U19732 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n20848), .ZN(n18738) );
  INV_X1 U19733 ( .A(n18738), .ZN(n16553) );
  NOR2_X1 U19734 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_0__SCAN_IN), 
        .ZN(n20855) );
  AOI21_X1 U19735 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n16553), .A(n20855), 
        .ZN(n18818) );
  OAI21_X1 U19736 ( .B1(n20849), .B2(n16554), .A(n18818), .ZN(P3_U2633) );
  OAI21_X1 U19737 ( .B1(n16561), .B2(n17464), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16555) );
  OAI21_X1 U19738 ( .B1(n16556), .B2(n18729), .A(n16555), .ZN(P3_U2634) );
  AOI21_X1 U19739 ( .B1(n20849), .B2(n20848), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16557) );
  AOI22_X1 U19740 ( .A1(n18864), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16557), 
        .B2(n18882), .ZN(P3_U2635) );
  NOR2_X1 U19741 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n16558) );
  OAI21_X1 U19742 ( .B1(n16558), .B2(BS16), .A(n18821), .ZN(n18819) );
  OAI21_X1 U19743 ( .B1(n18821), .B2(n18873), .A(n18819), .ZN(P3_U2636) );
  INV_X1 U19744 ( .A(n16559), .ZN(n16560) );
  NOR3_X1 U19745 ( .A1(n16561), .A2(n16560), .A3(n18660), .ZN(n18667) );
  NOR2_X1 U19746 ( .A1(n18667), .A2(n18724), .ZN(n18865) );
  OAI21_X1 U19747 ( .B1(n18865), .B2(n18211), .A(n16562), .ZN(P3_U2637) );
  NOR4_X1 U19748 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_19__SCAN_IN), .A3(P3_DATAWIDTH_REG_20__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_21__SCAN_IN), .ZN(n16566) );
  NOR4_X1 U19749 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_15__SCAN_IN), .A3(P3_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_17__SCAN_IN), .ZN(n16565) );
  NOR4_X1 U19750 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16564) );
  NOR4_X1 U19751 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_23__SCAN_IN), .A3(P3_DATAWIDTH_REG_24__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n16563) );
  NAND4_X1 U19752 ( .A1(n16566), .A2(n16565), .A3(n16564), .A4(n16563), .ZN(
        n16572) );
  NOR4_X1 U19753 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_2__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16570) );
  AOI211_X1 U19754 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_30__SCAN_IN), .B(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16569) );
  NOR4_X1 U19755 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_12__SCAN_IN), .ZN(n16568) );
  NOR4_X1 U19756 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16567) );
  NAND4_X1 U19757 ( .A1(n16570), .A2(n16569), .A3(n16568), .A4(n16567), .ZN(
        n16571) );
  NOR2_X1 U19758 ( .A1(n16572), .A2(n16571), .ZN(n18859) );
  INV_X1 U19759 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18814) );
  NOR3_X1 U19760 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16574) );
  OAI21_X1 U19761 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16574), .A(n18859), .ZN(
        n16573) );
  OAI21_X1 U19762 ( .B1(n18859), .B2(n18814), .A(n16573), .ZN(P3_U2638) );
  INV_X1 U19763 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18820) );
  AOI21_X1 U19764 ( .B1(n18855), .B2(n18820), .A(n16574), .ZN(n16575) );
  INV_X1 U19765 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18811) );
  INV_X1 U19766 ( .A(n18859), .ZN(n18861) );
  AOI22_X1 U19767 ( .A1(n18859), .A2(n16575), .B1(n18811), .B2(n18861), .ZN(
        P3_U2639) );
  INV_X1 U19768 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18806) );
  INV_X1 U19769 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n20971) );
  INV_X1 U19770 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18794) );
  INV_X1 U19771 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18769) );
  INV_X1 U19772 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18754) );
  NAND2_X1 U19773 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n16934) );
  NOR2_X1 U19774 ( .A1(n18754), .A2(n16934), .ZN(n16882) );
  NAND3_X1 U19775 ( .A1(n16882), .A2(P3_REIP_REG_5__SCAN_IN), .A3(
        P3_REIP_REG_4__SCAN_IN), .ZN(n16847) );
  NAND2_X1 U19776 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .ZN(n16861) );
  NOR3_X1 U19777 ( .A1(n18764), .A2(n16847), .A3(n16861), .ZN(n16814) );
  INV_X1 U19778 ( .A(n16814), .ZN(n16822) );
  INV_X1 U19779 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18767) );
  INV_X1 U19780 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18765) );
  NOR4_X1 U19781 ( .A1(n18769), .A2(n16822), .A3(n18767), .A4(n18765), .ZN(
        n16803) );
  AND2_X1 U19782 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16803), .ZN(n16786) );
  NAND3_X1 U19783 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(P3_REIP_REG_13__SCAN_IN), 
        .A3(n16786), .ZN(n16741) );
  NAND3_X1 U19784 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .ZN(n16716) );
  NOR2_X1 U19785 ( .A1(n16741), .A2(n16716), .ZN(n16711) );
  NAND4_X1 U19786 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(P3_REIP_REG_19__SCAN_IN), 
        .A3(P3_REIP_REG_18__SCAN_IN), .A4(n16711), .ZN(n16685) );
  NAND2_X1 U19787 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(P3_REIP_REG_22__SCAN_IN), 
        .ZN(n16693) );
  NOR3_X1 U19788 ( .A1(n18794), .A2(n16685), .A3(n16693), .ZN(n16666) );
  NAND2_X1 U19789 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16666), .ZN(n16657) );
  NOR2_X1 U19790 ( .A1(n20971), .A2(n16657), .ZN(n16644) );
  NAND2_X1 U19791 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16644), .ZN(n16591) );
  NAND4_X1 U19792 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16622), .ZN(n16593) );
  NOR3_X1 U19793 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18806), .A3(n16593), 
        .ZN(n16576) );
  AOI21_X1 U19794 ( .B1(n16947), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16576), .ZN(
        n16598) );
  NOR3_X1 U19795 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16936) );
  INV_X1 U19796 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n16916) );
  NAND2_X1 U19797 ( .A1(n16936), .A2(n16916), .ZN(n16915) );
  NOR2_X1 U19798 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16915), .ZN(n16893) );
  NAND2_X1 U19799 ( .A1(n16893), .A2(n20968), .ZN(n16889) );
  NAND2_X1 U19800 ( .A1(n16870), .A2(n16868), .ZN(n16865) );
  NAND2_X1 U19801 ( .A1(n16843), .A2(n21019), .ZN(n16834) );
  NAND2_X1 U19802 ( .A1(n16823), .A2(n17158), .ZN(n16818) );
  NAND2_X1 U19803 ( .A1(n16805), .A2(n16796), .ZN(n16795) );
  INV_X1 U19804 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16770) );
  NAND2_X1 U19805 ( .A1(n16774), .A2(n16770), .ZN(n16769) );
  INV_X1 U19806 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17049) );
  NAND2_X1 U19807 ( .A1(n16750), .A2(n17049), .ZN(n16746) );
  NAND2_X1 U19808 ( .A1(n16729), .A2(n17062), .ZN(n16725) );
  NAND2_X1 U19809 ( .A1(n16708), .A2(n17037), .ZN(n16702) );
  NAND2_X1 U19810 ( .A1(n16686), .A2(n16681), .ZN(n16680) );
  NAND2_X1 U19811 ( .A1(n16667), .A2(n16661), .ZN(n16660) );
  NAND2_X1 U19812 ( .A1(n16645), .A2(n16639), .ZN(n16638) );
  NOR2_X1 U19813 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16638), .ZN(n16623) );
  INV_X1 U19814 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16952) );
  NAND2_X1 U19815 ( .A1(n16623), .A2(n16952), .ZN(n16600) );
  NOR2_X1 U19816 ( .A1(n16937), .A2(n16600), .ZN(n16607) );
  INV_X1 U19817 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16957) );
  INV_X1 U19818 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16579) );
  NAND2_X1 U19819 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n16581), .ZN(
        n16580) );
  INV_X1 U19820 ( .A(n16577), .ZN(n16578) );
  AOI21_X1 U19821 ( .B1(n16579), .B2(n16580), .A(n16578), .ZN(n17519) );
  OAI21_X1 U19822 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n16581), .A(
        n16580), .ZN(n17539) );
  INV_X1 U19823 ( .A(n17539), .ZN(n16634) );
  AOI21_X1 U19824 ( .B1(n20928), .B2(n17518), .A(n16581), .ZN(n17549) );
  INV_X1 U19825 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17579) );
  NAND2_X1 U19826 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17627), .ZN(
        n16751) );
  INV_X1 U19827 ( .A(n16751), .ZN(n16582) );
  NAND2_X1 U19828 ( .A1(n16583), .A2(n16582), .ZN(n16588) );
  NOR2_X1 U19829 ( .A1(n9896), .A2(n17560), .ZN(n16586) );
  INV_X1 U19830 ( .A(n16586), .ZN(n16585) );
  NOR2_X1 U19831 ( .A1(n17579), .A2(n16585), .ZN(n16584) );
  OAI21_X1 U19832 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16584), .A(
        n17518), .ZN(n17564) );
  INV_X1 U19833 ( .A(n17564), .ZN(n16655) );
  OAI22_X1 U19834 ( .A1(n17579), .A2(n16586), .B1(n16585), .B2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17575) );
  AOI21_X1 U19835 ( .B1(n9896), .B2(n17560), .A(n16586), .ZN(n17587) );
  INV_X1 U19836 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17619) );
  NOR2_X1 U19837 ( .A1(n17619), .A2(n16588), .ZN(n16587) );
  OAI21_X1 U19838 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n16587), .A(
        n17560), .ZN(n17607) );
  INV_X1 U19839 ( .A(n17607), .ZN(n16689) );
  AOI21_X1 U19840 ( .B1(n17619), .B2(n16588), .A(n16587), .ZN(n17615) );
  NOR2_X1 U19841 ( .A1(n17630), .A2(n16751), .ZN(n17600) );
  OAI21_X1 U19842 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17600), .A(
        n16588), .ZN(n16589) );
  INV_X1 U19843 ( .A(n16589), .ZN(n17633) );
  NOR2_X1 U19844 ( .A1(n17633), .A2(n16707), .ZN(n16706) );
  NOR2_X1 U19845 ( .A1(n16706), .A2(n16858), .ZN(n16699) );
  NOR2_X1 U19846 ( .A1(n16675), .A2(n16858), .ZN(n16669) );
  NOR2_X1 U19847 ( .A1(n17549), .A2(n16647), .ZN(n16646) );
  NOR2_X1 U19848 ( .A1(n16646), .A2(n16858), .ZN(n16633) );
  NOR2_X1 U19849 ( .A1(n16632), .A2(n16858), .ZN(n16625) );
  NOR3_X1 U19850 ( .A1(n16602), .A2(n16601), .A3(n16873), .ZN(n16596) );
  NAND3_X1 U19851 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16592) );
  INV_X1 U19852 ( .A(n16945), .ZN(n16923) );
  AND2_X1 U19853 ( .A1(n16935), .A2(n16591), .ZN(n16643) );
  NOR2_X1 U19854 ( .A1(n16923), .A2(n16643), .ZN(n16642) );
  INV_X1 U19855 ( .A(n16642), .ZN(n16650) );
  AOI21_X1 U19856 ( .B1(n16935), .B2(n16592), .A(n16650), .ZN(n16621) );
  NOR2_X1 U19857 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16593), .ZN(n16605) );
  INV_X1 U19858 ( .A(n16605), .ZN(n16594) );
  AOI21_X1 U19859 ( .B1(n16621), .B2(n16594), .A(n18808), .ZN(n16595) );
  AOI211_X1 U19860 ( .C1(n16607), .C2(n16957), .A(n16596), .B(n16595), .ZN(
        n16597) );
  OAI211_X1 U19861 ( .C1(n16599), .C2(n16920), .A(n16598), .B(n16597), .ZN(
        P3_U2640) );
  NAND2_X1 U19862 ( .A1(n16946), .A2(n16600), .ZN(n16617) );
  XOR2_X1 U19863 ( .A(n16602), .B(n16601), .Z(n16606) );
  OAI22_X1 U19864 ( .A1(n16621), .A2(n18806), .B1(n16603), .B2(n16920), .ZN(
        n16604) );
  AOI211_X1 U19865 ( .C1(n16606), .C2(n18733), .A(n16605), .B(n16604), .ZN(
        n16609) );
  OAI21_X1 U19866 ( .B1(n16947), .B2(n16607), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16608) );
  OAI211_X1 U19867 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16617), .A(n16609), .B(
        n16608), .ZN(P3_U2641) );
  INV_X1 U19868 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18804) );
  AOI211_X1 U19869 ( .C1(n16612), .C2(n16611), .A(n16610), .B(n16926), .ZN(
        n16616) );
  NAND3_X1 U19870 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16622), .ZN(n16614) );
  OAI22_X1 U19871 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16614), .B1(n16613), 
        .B2(n16920), .ZN(n16615) );
  AOI211_X1 U19872 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n16947), .A(n16616), .B(
        n16615), .ZN(n16620) );
  INV_X1 U19873 ( .A(n16617), .ZN(n16618) );
  OAI21_X1 U19874 ( .B1(n16623), .B2(n16952), .A(n16618), .ZN(n16619) );
  OAI211_X1 U19875 ( .C1(n16621), .C2(n18804), .A(n16620), .B(n16619), .ZN(
        P3_U2642) );
  NAND2_X1 U19876 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16622), .ZN(n16631) );
  AOI22_X1 U19877 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16930), .B1(
        n16947), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16630) );
  INV_X1 U19878 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18800) );
  NAND2_X1 U19879 ( .A1(n16622), .A2(n18800), .ZN(n16635) );
  NAND2_X1 U19880 ( .A1(n16642), .A2(n16635), .ZN(n16628) );
  AOI211_X1 U19881 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16638), .A(n16623), .B(
        n16937), .ZN(n16627) );
  AOI211_X1 U19882 ( .C1(n17519), .C2(n16625), .A(n16624), .B(n16926), .ZN(
        n16626) );
  AOI211_X1 U19883 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16628), .A(n16627), 
        .B(n16626), .ZN(n16629) );
  OAI211_X1 U19884 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16631), .A(n16630), 
        .B(n16629), .ZN(P3_U2643) );
  AOI211_X1 U19885 ( .C1(n16634), .C2(n16633), .A(n16632), .B(n16926), .ZN(
        n16637) );
  INV_X1 U19886 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n21063) );
  OAI21_X1 U19887 ( .B1(n16920), .B2(n21063), .A(n16635), .ZN(n16636) );
  AOI211_X1 U19888 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n16947), .A(n16637), .B(
        n16636), .ZN(n16641) );
  OAI211_X1 U19889 ( .C1(n16645), .C2(n16639), .A(n16946), .B(n16638), .ZN(
        n16640) );
  OAI211_X1 U19890 ( .C1(n16642), .C2(n18800), .A(n16641), .B(n16640), .ZN(
        P3_U2644) );
  AOI22_X1 U19891 ( .A1(n16947), .A2(P3_EBX_REG_26__SCAN_IN), .B1(n16644), 
        .B2(n16643), .ZN(n16652) );
  AOI211_X1 U19892 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16660), .A(n16645), .B(
        n16937), .ZN(n16649) );
  AOI211_X1 U19893 ( .C1(n17549), .C2(n16647), .A(n16646), .B(n16926), .ZN(
        n16648) );
  AOI211_X1 U19894 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n16650), .A(n16649), 
        .B(n16648), .ZN(n16651) );
  OAI211_X1 U19895 ( .C1(n20928), .C2(n16920), .A(n16652), .B(n16651), .ZN(
        P3_U2645) );
  INV_X1 U19896 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18795) );
  OAI21_X1 U19897 ( .B1(n16666), .B2(n16909), .A(n16945), .ZN(n16674) );
  AOI21_X1 U19898 ( .B1(n16935), .B2(n18795), .A(n16674), .ZN(n16664) );
  AOI211_X1 U19899 ( .C1(n16655), .C2(n16654), .A(n16653), .B(n16926), .ZN(
        n16659) );
  NAND2_X1 U19900 ( .A1(n16935), .A2(n20971), .ZN(n16656) );
  OAI22_X1 U19901 ( .A1(n16911), .A2(n16661), .B1(n16657), .B2(n16656), .ZN(
        n16658) );
  AOI211_X1 U19902 ( .C1(n16930), .C2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16659), .B(n16658), .ZN(n16663) );
  OAI211_X1 U19903 ( .C1(n16667), .C2(n16661), .A(n16946), .B(n16660), .ZN(
        n16662) );
  OAI211_X1 U19904 ( .C1(n16664), .C2(n20971), .A(n16663), .B(n16662), .ZN(
        P3_U2646) );
  NOR2_X1 U19905 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16909), .ZN(n16665) );
  AOI22_X1 U19906 ( .A1(n16947), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16666), 
        .B2(n16665), .ZN(n16673) );
  AOI211_X1 U19907 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16680), .A(n16667), .B(
        n16937), .ZN(n16671) );
  AOI211_X1 U19908 ( .C1(n17575), .C2(n16669), .A(n16668), .B(n16926), .ZN(
        n16670) );
  AOI211_X1 U19909 ( .C1(n16674), .C2(P3_REIP_REG_24__SCAN_IN), .A(n16671), 
        .B(n16670), .ZN(n16672) );
  OAI211_X1 U19910 ( .C1(n17579), .C2(n16920), .A(n16673), .B(n16672), .ZN(
        P3_U2647) );
  INV_X1 U19911 ( .A(n16674), .ZN(n16684) );
  AOI211_X1 U19912 ( .C1(n17587), .C2(n16676), .A(n16675), .B(n16926), .ZN(
        n16679) );
  NOR4_X1 U19913 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n16909), .A3(n16685), 
        .A4(n16693), .ZN(n16678) );
  OAI22_X1 U19914 ( .A1(n9896), .A2(n16920), .B1(n16911), .B2(n16681), .ZN(
        n16677) );
  NOR3_X1 U19915 ( .A1(n16679), .A2(n16678), .A3(n16677), .ZN(n16683) );
  OAI211_X1 U19916 ( .C1(n16686), .C2(n16681), .A(n16946), .B(n16680), .ZN(
        n16682) );
  OAI211_X1 U19917 ( .C1(n16684), .C2(n18794), .A(n16683), .B(n16682), .ZN(
        P3_U2648) );
  AOI22_X1 U19918 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n16930), .B1(
        n16947), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n16697) );
  INV_X1 U19919 ( .A(n16685), .ZN(n16692) );
  OAI21_X1 U19920 ( .B1(n16692), .B2(n16909), .A(n16945), .ZN(n16712) );
  AOI211_X1 U19921 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16702), .A(n16686), .B(
        n16937), .ZN(n16691) );
  AOI211_X1 U19922 ( .C1(n16689), .C2(n16688), .A(n16687), .B(n16926), .ZN(
        n16690) );
  AOI211_X1 U19923 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n16712), .A(n16691), 
        .B(n16690), .ZN(n16696) );
  NAND2_X1 U19924 ( .A1(n16935), .A2(n16692), .ZN(n16705) );
  INV_X1 U19925 ( .A(n16705), .ZN(n16694) );
  OAI211_X1 U19926 ( .C1(P3_REIP_REG_21__SCAN_IN), .C2(P3_REIP_REG_22__SCAN_IN), .A(n16694), .B(n16693), .ZN(n16695) );
  NAND3_X1 U19927 ( .A1(n16697), .A2(n16696), .A3(n16695), .ZN(P3_U2649) );
  AOI211_X1 U19928 ( .C1(n17615), .C2(n16699), .A(n16698), .B(n16926), .ZN(
        n16701) );
  OAI22_X1 U19929 ( .A1(n17619), .A2(n16920), .B1(n16911), .B2(n17037), .ZN(
        n16700) );
  AOI211_X1 U19930 ( .C1(n16712), .C2(P3_REIP_REG_21__SCAN_IN), .A(n16701), 
        .B(n16700), .ZN(n16704) );
  OAI211_X1 U19931 ( .C1(n16708), .C2(n17037), .A(n16946), .B(n16702), .ZN(
        n16703) );
  OAI211_X1 U19932 ( .C1(P3_REIP_REG_21__SCAN_IN), .C2(n16705), .A(n16704), 
        .B(n16703), .ZN(P3_U2650) );
  AOI211_X1 U19933 ( .C1(n17633), .C2(n16707), .A(n16706), .B(n16926), .ZN(
        n16710) );
  AOI211_X1 U19934 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16725), .A(n16708), .B(
        n16937), .ZN(n16709) );
  AOI211_X1 U19935 ( .C1(n16930), .C2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16710), .B(n16709), .ZN(n16714) );
  INV_X1 U19936 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18783) );
  NAND2_X1 U19937 ( .A1(n16935), .A2(n16711), .ZN(n16728) );
  NOR2_X1 U19938 ( .A1(n18783), .A2(n16728), .ZN(n16724) );
  OAI221_X1 U19939 ( .B1(P3_REIP_REG_20__SCAN_IN), .B2(P3_REIP_REG_19__SCAN_IN), .C1(P3_REIP_REG_20__SCAN_IN), .C2(n16724), .A(n16712), .ZN(n16713) );
  OAI211_X1 U19940 ( .C1(n16715), .C2(n16911), .A(n16714), .B(n16713), .ZN(
        P3_U2651) );
  INV_X1 U19941 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18785) );
  OR2_X1 U19942 ( .A1(n16741), .A2(n16923), .ZN(n16775) );
  NAND2_X1 U19943 ( .A1(n16909), .A2(n16945), .ZN(n16944) );
  OAI21_X1 U19944 ( .B1(n16716), .B2(n16775), .A(n16944), .ZN(n16740) );
  OAI21_X1 U19945 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n16728), .A(n16740), 
        .ZN(n16723) );
  INV_X1 U19946 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16721) );
  NAND2_X1 U19947 ( .A1(n17627), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17640) );
  NOR2_X1 U19948 ( .A1(n17875), .A2(n17640), .ZN(n17639) );
  NAND2_X1 U19949 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17639), .ZN(
        n16730) );
  AOI21_X1 U19950 ( .B1(n16721), .B2(n16730), .A(n17600), .ZN(n16717) );
  INV_X1 U19951 ( .A(n16717), .ZN(n17643) );
  OAI21_X1 U19952 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16730), .A(
        n16907), .ZN(n16719) );
  AOI21_X1 U19953 ( .B1(n17643), .B2(n16719), .A(n16926), .ZN(n16718) );
  OAI21_X1 U19954 ( .B1(n17643), .B2(n16719), .A(n16718), .ZN(n16720) );
  OAI211_X1 U19955 ( .C1(n16721), .C2(n16920), .A(n15697), .B(n16720), .ZN(
        n16722) );
  AOI221_X1 U19956 ( .B1(n16724), .B2(n18785), .C1(n16723), .C2(
        P3_REIP_REG_19__SCAN_IN), .A(n16722), .ZN(n16727) );
  OAI211_X1 U19957 ( .C1(n16729), .C2(n17062), .A(n16946), .B(n16725), .ZN(
        n16726) );
  OAI211_X1 U19958 ( .C1(n17062), .C2(n16911), .A(n16727), .B(n16726), .ZN(
        P3_U2652) );
  AOI22_X1 U19959 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16930), .B1(
        n16947), .B2(P3_EBX_REG_18__SCAN_IN), .ZN(n16738) );
  NOR2_X1 U19960 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n16728), .ZN(n16736) );
  AOI211_X1 U19961 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16746), .A(n16729), .B(
        n16937), .ZN(n16735) );
  OAI21_X1 U19962 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17639), .A(
        n16730), .ZN(n17652) );
  NAND2_X1 U19963 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16731), .ZN(
        n16927) );
  OAI21_X1 U19964 ( .B1(n17640), .B2(n16927), .A(n16907), .ZN(n16733) );
  OAI21_X1 U19965 ( .B1(n17652), .B2(n16733), .A(n18733), .ZN(n16732) );
  AOI21_X1 U19966 ( .B1(n17652), .B2(n16733), .A(n16732), .ZN(n16734) );
  NOR4_X1 U19967 ( .A1(n9760), .A2(n16736), .A3(n16735), .A4(n16734), .ZN(
        n16737) );
  OAI211_X1 U19968 ( .C1(n18783), .C2(n16740), .A(n16738), .B(n16737), .ZN(
        P3_U2653) );
  AOI22_X1 U19969 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n16930), .B1(
        n16947), .B2(P3_EBX_REG_17__SCAN_IN), .ZN(n16749) );
  INV_X1 U19970 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17663) );
  AOI21_X1 U19971 ( .B1(n17663), .B2(n16751), .A(n17639), .ZN(n17666) );
  OAI21_X1 U19972 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16751), .A(
        n16907), .ZN(n16739) );
  XNOR2_X1 U19973 ( .A(n17666), .B(n16739), .ZN(n16745) );
  INV_X1 U19974 ( .A(n16740), .ZN(n16744) );
  NAND2_X1 U19975 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16742) );
  OR2_X1 U19976 ( .A1(n16909), .A2(n16741), .ZN(n16757) );
  INV_X1 U19977 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18781) );
  OAI21_X1 U19978 ( .B1(n16742), .B2(n16757), .A(n18781), .ZN(n16743) );
  AOI22_X1 U19979 ( .A1(n18733), .A2(n16745), .B1(n16744), .B2(n16743), .ZN(
        n16748) );
  OAI211_X1 U19980 ( .C1(n16750), .C2(n17049), .A(n16946), .B(n16746), .ZN(
        n16747) );
  NAND4_X1 U19981 ( .A1(n16749), .A2(n16748), .A3(n15697), .A4(n16747), .ZN(
        P3_U2654) );
  AOI22_X1 U19982 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n16930), .B1(
        n16947), .B2(P3_EBX_REG_16__SCAN_IN), .ZN(n16760) );
  AOI211_X1 U19983 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16769), .A(n16750), .B(
        n16937), .ZN(n16756) );
  INV_X1 U19984 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18777) );
  NOR3_X1 U19985 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n18777), .A3(n16757), 
        .ZN(n16755) );
  NOR2_X1 U19986 ( .A1(n17875), .A2(n17677), .ZN(n17676) );
  NAND2_X1 U19987 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17676), .ZN(
        n16761) );
  INV_X1 U19988 ( .A(n16761), .ZN(n16752) );
  OAI21_X1 U19989 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16752), .A(
        n16751), .ZN(n17681) );
  OAI21_X1 U19990 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16761), .A(
        n16907), .ZN(n16763) );
  OAI21_X1 U19991 ( .B1(n17681), .B2(n16763), .A(n18733), .ZN(n16753) );
  AOI21_X1 U19992 ( .B1(n17681), .B2(n16763), .A(n16753), .ZN(n16754) );
  NOR4_X1 U19993 ( .A1(n9760), .A2(n16756), .A3(n16755), .A4(n16754), .ZN(
        n16759) );
  NAND2_X1 U19994 ( .A1(n16944), .A2(n16775), .ZN(n16781) );
  INV_X1 U19995 ( .A(n16781), .ZN(n16768) );
  NOR2_X1 U19996 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n16757), .ZN(n16767) );
  OAI21_X1 U19997 ( .B1(n16768), .B2(n16767), .A(P3_REIP_REG_16__SCAN_IN), 
        .ZN(n16758) );
  NAND3_X1 U19998 ( .A1(n16760), .A2(n16759), .A3(n16758), .ZN(P3_U2655) );
  OAI21_X1 U19999 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17676), .A(
        n16761), .ZN(n17686) );
  INV_X1 U20000 ( .A(n17676), .ZN(n16762) );
  AOI221_X1 U20001 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16907), .C1(
        n16762), .C2(n16907), .A(n16926), .ZN(n16765) );
  OAI21_X1 U20002 ( .B1(n16926), .B2(n16763), .A(n17686), .ZN(n16764) );
  OAI21_X1 U20003 ( .B1(n17686), .B2(n16765), .A(n16764), .ZN(n16773) );
  INV_X1 U20004 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17689) );
  OAI22_X1 U20005 ( .A1(n17689), .A2(n16920), .B1(n16911), .B2(n16770), .ZN(
        n16766) );
  AOI211_X1 U20006 ( .C1(n16768), .C2(P3_REIP_REG_15__SCAN_IN), .A(n16767), 
        .B(n16766), .ZN(n16772) );
  OAI211_X1 U20007 ( .C1(n16774), .C2(n16770), .A(n16946), .B(n16769), .ZN(
        n16771) );
  NAND4_X1 U20008 ( .A1(n16773), .A2(n16772), .A3(n15697), .A4(n16771), .ZN(
        P3_U2656) );
  INV_X1 U20009 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n16785) );
  AOI211_X1 U20010 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16795), .A(n16774), .B(
        n16937), .ZN(n16783) );
  INV_X1 U20011 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18776) );
  NAND4_X1 U20012 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16935), .A3(n16786), 
        .A4(n16775), .ZN(n16780) );
  INV_X1 U20013 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17702) );
  NAND2_X1 U20014 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16776), .ZN(
        n16787) );
  AOI21_X1 U20015 ( .B1(n17702), .B2(n16787), .A(n17676), .ZN(n17704) );
  OAI21_X1 U20016 ( .B1(n16787), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n16907), .ZN(n16777) );
  INV_X1 U20017 ( .A(n16777), .ZN(n16790) );
  AOI21_X1 U20018 ( .B1(n17704), .B2(n16790), .A(n16926), .ZN(n16778) );
  OAI21_X1 U20019 ( .B1(n17704), .B2(n16790), .A(n16778), .ZN(n16779) );
  OAI211_X1 U20020 ( .C1(n16781), .C2(n18776), .A(n16780), .B(n16779), .ZN(
        n16782) );
  AOI211_X1 U20021 ( .C1(n16930), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16783), .B(n16782), .ZN(n16784) );
  OAI211_X1 U20022 ( .C1(n16911), .C2(n16785), .A(n16784), .B(n15697), .ZN(
        P3_U2657) );
  INV_X1 U20023 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16799) );
  OAI21_X1 U20024 ( .B1(n16803), .B2(n16909), .A(n16945), .ZN(n16816) );
  NOR2_X1 U20025 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16909), .ZN(n16802) );
  NAND2_X1 U20026 ( .A1(n16935), .A2(n16786), .ZN(n16793) );
  OR2_X1 U20027 ( .A1(n17875), .A2(n17814), .ZN(n16883) );
  NOR2_X1 U20028 ( .A1(n17815), .A2(n16883), .ZN(n16871) );
  NAND2_X1 U20029 ( .A1(n17700), .A2(n16871), .ZN(n17712) );
  INV_X1 U20030 ( .A(n17712), .ZN(n16810) );
  NAND2_X1 U20031 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16810), .ZN(
        n16800) );
  INV_X1 U20032 ( .A(n16800), .ZN(n16788) );
  OAI21_X1 U20033 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16788), .A(
        n16787), .ZN(n17719) );
  AOI211_X1 U20034 ( .C1(n16907), .C2(n16800), .A(n16872), .B(n17719), .ZN(
        n16789) );
  AOI211_X1 U20035 ( .C1(n16947), .C2(P3_EBX_REG_13__SCAN_IN), .A(n9760), .B(
        n16789), .ZN(n16792) );
  NAND3_X1 U20036 ( .A1(n18733), .A2(n16790), .A3(n17719), .ZN(n16791) );
  OAI211_X1 U20037 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n16793), .A(n16792), 
        .B(n16791), .ZN(n16794) );
  AOI221_X1 U20038 ( .B1(n16816), .B2(P3_REIP_REG_13__SCAN_IN), .C1(n16802), 
        .C2(P3_REIP_REG_13__SCAN_IN), .A(n16794), .ZN(n16798) );
  OAI211_X1 U20039 ( .C1(n16805), .C2(n16796), .A(n16946), .B(n16795), .ZN(
        n16797) );
  OAI211_X1 U20040 ( .C1(n16920), .C2(n16799), .A(n16798), .B(n16797), .ZN(
        P3_U2658) );
  AOI22_X1 U20041 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16930), .B1(
        n16947), .B2(P3_EBX_REG_12__SCAN_IN), .ZN(n16809) );
  INV_X1 U20042 ( .A(n16844), .ZN(n17784) );
  NOR2_X1 U20043 ( .A1(n17784), .A2(n16927), .ZN(n16874) );
  AOI21_X1 U20044 ( .B1(n17700), .B2(n16874), .A(n16858), .ZN(n16801) );
  OAI21_X1 U20045 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n16810), .A(
        n16800), .ZN(n17739) );
  XNOR2_X1 U20046 ( .A(n16801), .B(n17739), .ZN(n16804) );
  AOI22_X1 U20047 ( .A1(n18733), .A2(n16804), .B1(n16803), .B2(n16802), .ZN(
        n16808) );
  AOI211_X1 U20048 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16818), .A(n16805), .B(
        n16937), .ZN(n16806) );
  AOI211_X1 U20049 ( .C1(P3_REIP_REG_12__SCAN_IN), .C2(n16816), .A(n9760), .B(
        n16806), .ZN(n16807) );
  NAND3_X1 U20050 ( .A1(n16809), .A2(n16808), .A3(n16807), .ZN(P3_U2659) );
  AOI22_X1 U20051 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n16930), .B1(
        n16947), .B2(P3_EBX_REG_11__SCAN_IN), .ZN(n16821) );
  INV_X1 U20052 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17770) );
  NAND2_X1 U20053 ( .A1(n17782), .A2(n16871), .ZN(n16845) );
  NOR2_X1 U20054 ( .A1(n17770), .A2(n16845), .ZN(n16833) );
  NAND2_X1 U20055 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n16833), .ZN(
        n16825) );
  AOI21_X1 U20056 ( .B1(n17741), .B2(n16825), .A(n16810), .ZN(n17744) );
  INV_X1 U20057 ( .A(n16874), .ZN(n16811) );
  NOR2_X1 U20058 ( .A1(n16812), .A2(n16811), .ZN(n16824) );
  AOI21_X1 U20059 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16824), .A(
        n16858), .ZN(n16813) );
  XOR2_X1 U20060 ( .A(n17744), .B(n16813), .Z(n16817) );
  NAND2_X1 U20061 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n16826) );
  NAND2_X1 U20062 ( .A1(n16935), .A2(n16814), .ZN(n16842) );
  OAI21_X1 U20063 ( .B1(n16826), .B2(n16842), .A(n18769), .ZN(n16815) );
  AOI22_X1 U20064 ( .A1(n18733), .A2(n16817), .B1(n16816), .B2(n16815), .ZN(
        n16820) );
  OAI211_X1 U20065 ( .C1(n16823), .C2(n17158), .A(n16946), .B(n16818), .ZN(
        n16819) );
  NAND4_X1 U20066 ( .A1(n16821), .A2(n16820), .A3(n15697), .A4(n16819), .ZN(
        P3_U2660) );
  AOI21_X1 U20067 ( .B1(n16935), .B2(n16822), .A(n16923), .ZN(n16854) );
  AOI21_X1 U20068 ( .B1(n16947), .B2(P3_EBX_REG_10__SCAN_IN), .A(n9760), .ZN(
        n16832) );
  AOI211_X1 U20069 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16834), .A(n16823), .B(
        n16937), .ZN(n16830) );
  NOR2_X1 U20070 ( .A1(n16824), .A2(n16858), .ZN(n16837) );
  OAI21_X1 U20071 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16833), .A(
        n16825), .ZN(n17759) );
  XOR2_X1 U20072 ( .A(n16837), .B(n17759), .Z(n16828) );
  OAI21_X1 U20073 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(P3_REIP_REG_9__SCAN_IN), 
        .A(n16826), .ZN(n16827) );
  OAI22_X1 U20074 ( .A1(n16926), .A2(n16828), .B1(n16842), .B2(n16827), .ZN(
        n16829) );
  AOI211_X1 U20075 ( .C1(n16930), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16830), .B(n16829), .ZN(n16831) );
  OAI211_X1 U20076 ( .C1(n18767), .C2(n16854), .A(n16832), .B(n16831), .ZN(
        P3_U2661) );
  AOI21_X1 U20077 ( .B1(n17770), .B2(n16845), .A(n16833), .ZN(n17774) );
  NOR2_X1 U20078 ( .A1(n16907), .A2(n16926), .ZN(n16928) );
  OAI211_X1 U20079 ( .C1(n16843), .C2(n21019), .A(n16946), .B(n16834), .ZN(
        n16835) );
  OAI21_X1 U20080 ( .B1(n21019), .B2(n16911), .A(n16835), .ZN(n16840) );
  OAI21_X1 U20081 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16845), .A(
        n17774), .ZN(n16836) );
  NAND3_X1 U20082 ( .A1(n16837), .A2(n18733), .A3(n16836), .ZN(n16838) );
  OAI211_X1 U20083 ( .C1(n17770), .C2(n16920), .A(n15697), .B(n16838), .ZN(
        n16839) );
  AOI211_X1 U20084 ( .C1(n17774), .C2(n16928), .A(n16840), .B(n16839), .ZN(
        n16841) );
  OAI221_X1 U20085 ( .B1(P3_REIP_REG_9__SCAN_IN), .B2(n16842), .C1(n18765), 
        .C2(n16854), .A(n16841), .ZN(P3_U2662) );
  AOI21_X1 U20086 ( .B1(n16947), .B2(P3_EBX_REG_8__SCAN_IN), .A(n9760), .ZN(
        n16853) );
  AOI211_X1 U20087 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16865), .A(n16843), .B(
        n16937), .ZN(n16851) );
  NAND2_X1 U20088 ( .A1(n16844), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17783) );
  NOR2_X1 U20089 ( .A1(n17875), .A2(n17783), .ZN(n16856) );
  OAI21_X1 U20090 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16856), .A(
        n16845), .ZN(n17786) );
  OAI21_X1 U20091 ( .B1(n17783), .B2(n16927), .A(n16907), .ZN(n16846) );
  XNOR2_X1 U20092 ( .A(n17786), .B(n16846), .ZN(n16849) );
  NOR2_X1 U20093 ( .A1(n16909), .A2(n16847), .ZN(n16869) );
  NAND2_X1 U20094 ( .A1(n16869), .A2(n18764), .ZN(n16848) );
  OAI22_X1 U20095 ( .A1(n16926), .A2(n16849), .B1(n16861), .B2(n16848), .ZN(
        n16850) );
  AOI211_X1 U20096 ( .C1(n16930), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16851), .B(n16850), .ZN(n16852) );
  OAI211_X1 U20097 ( .C1(n18764), .C2(n16854), .A(n16853), .B(n16852), .ZN(
        P3_U2663) );
  NAND2_X1 U20098 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(P3_REIP_REG_4__SCAN_IN), 
        .ZN(n16855) );
  NAND2_X1 U20099 ( .A1(n16882), .A2(n16945), .ZN(n16892) );
  OAI21_X1 U20100 ( .B1(n16855), .B2(n16892), .A(n16944), .ZN(n16886) );
  INV_X1 U20101 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18761) );
  INV_X1 U20102 ( .A(n16871), .ZN(n16857) );
  AOI21_X1 U20103 ( .B1(n17798), .B2(n16857), .A(n16856), .ZN(n17805) );
  NOR2_X1 U20104 ( .A1(n16874), .A2(n16858), .ZN(n16860) );
  AOI21_X1 U20105 ( .B1(n17805), .B2(n16860), .A(n16926), .ZN(n16859) );
  OAI21_X1 U20106 ( .B1(n17805), .B2(n16860), .A(n16859), .ZN(n16863) );
  OAI211_X1 U20107 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(P3_REIP_REG_6__SCAN_IN), 
        .A(n16869), .B(n16861), .ZN(n16862) );
  OAI211_X1 U20108 ( .C1(n16886), .C2(n18761), .A(n16863), .B(n16862), .ZN(
        n16864) );
  AOI211_X1 U20109 ( .C1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n16930), .A(
        n9760), .B(n16864), .ZN(n16867) );
  OAI211_X1 U20110 ( .C1(n16870), .C2(n16868), .A(n16946), .B(n16865), .ZN(
        n16866) );
  OAI211_X1 U20111 ( .C1(n16868), .C2(n16911), .A(n16867), .B(n16866), .ZN(
        P3_U2664) );
  INV_X1 U20112 ( .A(n16869), .ZN(n16881) );
  INV_X1 U20113 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18759) );
  AOI211_X1 U20114 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16889), .A(n16870), .B(
        n16937), .ZN(n16879) );
  AOI21_X1 U20115 ( .B1(n17815), .B2(n16883), .A(n16871), .ZN(n17817) );
  AOI21_X1 U20116 ( .B1(n16907), .B2(n16883), .A(n16872), .ZN(n16876) );
  NOR3_X1 U20117 ( .A1(n17817), .A2(n16874), .A3(n16873), .ZN(n16875) );
  AOI211_X1 U20118 ( .C1(n17817), .C2(n16876), .A(n9760), .B(n16875), .ZN(
        n16877) );
  OAI21_X1 U20119 ( .B1(n17815), .B2(n16920), .A(n16877), .ZN(n16878) );
  AOI211_X1 U20120 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16947), .A(n16879), .B(
        n16878), .ZN(n16880) );
  OAI221_X1 U20121 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n16881), .C1(n18759), 
        .C2(n16886), .A(n16880), .ZN(P3_U2665) );
  AND2_X1 U20122 ( .A1(n16935), .A2(n16882), .ZN(n16898) );
  AOI21_X1 U20123 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n16898), .A(
        P3_REIP_REG_5__SCAN_IN), .ZN(n16887) );
  INV_X1 U20124 ( .A(n17826), .ZN(n16884) );
  NOR2_X1 U20125 ( .A1(n17875), .A2(n16884), .ZN(n16894) );
  OAI21_X1 U20126 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n16894), .A(
        n16883), .ZN(n17829) );
  OAI21_X1 U20127 ( .B1(n16884), .B2(n16927), .A(n16907), .ZN(n16896) );
  XNOR2_X1 U20128 ( .A(n17829), .B(n16896), .ZN(n16885) );
  OAI22_X1 U20129 ( .A1(n16887), .A2(n16886), .B1(n16926), .B2(n16885), .ZN(
        n16888) );
  AOI211_X1 U20130 ( .C1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n16930), .A(
        n9760), .B(n16888), .ZN(n16891) );
  OAI211_X1 U20131 ( .C1(n16893), .C2(n20968), .A(n16946), .B(n16889), .ZN(
        n16890) );
  OAI211_X1 U20132 ( .C1(n20968), .C2(n16911), .A(n16891), .B(n16890), .ZN(
        P3_U2666) );
  INV_X1 U20133 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18755) );
  NAND2_X1 U20134 ( .A1(n16944), .A2(n16892), .ZN(n16908) );
  AOI211_X1 U20135 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16915), .A(n16893), .B(
        n16937), .ZN(n16903) );
  INV_X1 U20136 ( .A(n17842), .ZN(n16895) );
  NAND2_X1 U20137 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16895), .ZN(
        n16905) );
  AOI21_X1 U20138 ( .B1(n17844), .B2(n16905), .A(n16894), .ZN(n17846) );
  NAND2_X1 U20139 ( .A1(n17844), .A2(n16895), .ZN(n17837) );
  OAI22_X1 U20140 ( .A1(n17846), .A2(n16896), .B1(n16927), .B2(n17837), .ZN(
        n16897) );
  AOI22_X1 U20141 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n16930), .B1(
        n18733), .B2(n16897), .ZN(n16901) );
  AOI22_X1 U20142 ( .A1(n16928), .A2(n17846), .B1(n16898), .B2(n18755), .ZN(
        n16900) );
  OAI21_X1 U20143 ( .B1(n17224), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n18891), .ZN(n16899) );
  NAND4_X1 U20144 ( .A1(n16901), .A2(n16900), .A3(n15697), .A4(n16899), .ZN(
        n16902) );
  AOI211_X1 U20145 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16947), .A(n16903), .B(
        n16902), .ZN(n16904) );
  OAI21_X1 U20146 ( .B1(n18755), .B2(n16908), .A(n16904), .ZN(P3_U2667) );
  INV_X1 U20147 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16919) );
  NAND2_X1 U20148 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16924) );
  INV_X1 U20149 ( .A(n16905), .ZN(n16906) );
  AOI21_X1 U20150 ( .B1(n16919), .B2(n16924), .A(n16906), .ZN(n17857) );
  INV_X1 U20151 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17868) );
  OAI21_X1 U20152 ( .B1(n17868), .B2(n16927), .A(n16907), .ZN(n16925) );
  XNOR2_X1 U20153 ( .A(n17857), .B(n16925), .ZN(n16914) );
  AOI221_X1 U20154 ( .B1(n16909), .B2(n18754), .C1(n16934), .C2(n18754), .A(
        n16908), .ZN(n16913) );
  NAND2_X1 U20155 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18685), .ZN(
        n18676) );
  INV_X1 U20156 ( .A(n18676), .ZN(n18687) );
  OAI21_X1 U20157 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18687), .A(
        n12917), .ZN(n18827) );
  OAI22_X1 U20158 ( .A1(n16911), .A2(n16916), .B1(n16910), .B2(n18827), .ZN(
        n16912) );
  AOI211_X1 U20159 ( .C1(n16914), .C2(n18733), .A(n16913), .B(n16912), .ZN(
        n16918) );
  OAI211_X1 U20160 ( .C1(n16936), .C2(n16916), .A(n16946), .B(n16915), .ZN(
        n16917) );
  OAI211_X1 U20161 ( .C1(n16920), .C2(n16919), .A(n16918), .B(n16917), .ZN(
        P3_U2668) );
  NAND2_X1 U20162 ( .A1(n13018), .A2(n16921), .ZN(n18674) );
  NAND2_X1 U20163 ( .A1(n18676), .A2(n18674), .ZN(n18835) );
  INV_X1 U20164 ( .A(n18835), .ZN(n16922) );
  AOI22_X1 U20165 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n16923), .B1(n16922), 
        .B2(n18891), .ZN(n16943) );
  OAI21_X1 U20166 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16924), .ZN(n17865) );
  INV_X1 U20167 ( .A(n17865), .ZN(n16929) );
  AOI211_X1 U20168 ( .C1(n16929), .C2(n16927), .A(n16926), .B(n16925), .ZN(
        n16933) );
  AOI22_X1 U20169 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n16930), .B1(
        n16929), .B2(n16928), .ZN(n16931) );
  INV_X1 U20170 ( .A(n16931), .ZN(n16932) );
  AOI211_X1 U20171 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16947), .A(n16933), .B(
        n16932), .ZN(n16942) );
  OAI211_X1 U20172 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n16935), .B(n16934), .ZN(n16941) );
  AOI211_X1 U20173 ( .C1(n16938), .C2(P3_EBX_REG_2__SCAN_IN), .A(n16937), .B(
        n16936), .ZN(n16939) );
  INV_X1 U20174 ( .A(n16939), .ZN(n16940) );
  NAND4_X1 U20175 ( .A1(n16943), .A2(n16942), .A3(n16941), .A4(n16940), .ZN(
        P3_U2669) );
  AOI22_X1 U20176 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n16944), .B1(n18891), 
        .B2(n12916), .ZN(n16950) );
  NAND3_X1 U20177 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18837), .A3(
        n16945), .ZN(n16949) );
  OAI21_X1 U20178 ( .B1(n16947), .B2(n16946), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n16948) );
  NAND3_X1 U20179 ( .A1(n16950), .A2(n16949), .A3(n16948), .ZN(P3_U2671) );
  INV_X1 U20180 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n21029) );
  NAND4_X1 U20181 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(P3_EBX_REG_24__SCAN_IN), .A4(P3_EBX_REG_23__SCAN_IN), .ZN(n16951)
         );
  NOR4_X1 U20182 ( .A1(n16952), .A2(n21029), .A3(n17037), .A4(n16951), .ZN(
        n16953) );
  NAND4_X1 U20183 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(n17025), .A4(n16953), .ZN(n16956) );
  NOR2_X1 U20184 ( .A1(n16957), .A2(n16956), .ZN(n16982) );
  NAND2_X1 U20185 ( .A1(n17251), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16955) );
  NAND2_X1 U20186 ( .A1(n16982), .A2(n9796), .ZN(n16954) );
  OAI22_X1 U20187 ( .A1(n16982), .A2(n16955), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n16954), .ZN(P3_U2672) );
  NAND2_X1 U20188 ( .A1(n16957), .A2(n16956), .ZN(n16958) );
  NAND2_X1 U20189 ( .A1(n16958), .A2(n17251), .ZN(n16981) );
  AOI22_X1 U20190 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n17212), .B1(
        n17205), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16962) );
  AOI22_X1 U20191 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__6__SCAN_IN), .B2(n17213), .ZN(n16961) );
  AOI22_X1 U20192 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__6__SCAN_IN), .B2(n17117), .ZN(n16960) );
  AOI22_X1 U20193 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n17189), .ZN(n16959) );
  NAND4_X1 U20194 ( .A1(n16962), .A2(n16961), .A3(n16960), .A4(n16959), .ZN(
        n16968) );
  AOI22_X1 U20195 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n17123), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16966) );
  AOI22_X1 U20196 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n17206), .B1(
        P3_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n15559), .ZN(n16965) );
  AOI22_X1 U20197 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16964) );
  AOI22_X1 U20198 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__6__SCAN_IN), .B2(n15600), .ZN(n16963) );
  NAND4_X1 U20199 ( .A1(n16966), .A2(n16965), .A3(n16964), .A4(n16963), .ZN(
        n16967) );
  NOR2_X1 U20200 ( .A1(n16968), .A2(n16967), .ZN(n16984) );
  NOR2_X1 U20201 ( .A1(n16983), .A2(n16984), .ZN(n16980) );
  AOI22_X1 U20202 ( .A1(n17209), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16972) );
  AOI22_X1 U20203 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16971) );
  AOI22_X1 U20204 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16970) );
  AOI22_X1 U20205 ( .A1(n17207), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16969) );
  NAND4_X1 U20206 ( .A1(n16972), .A2(n16971), .A3(n16970), .A4(n16969), .ZN(
        n16978) );
  AOI22_X1 U20207 ( .A1(n15435), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16976) );
  AOI22_X1 U20208 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16975) );
  AOI22_X1 U20209 ( .A1(n9758), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16974) );
  AOI22_X1 U20210 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16973) );
  NAND4_X1 U20211 ( .A1(n16976), .A2(n16975), .A3(n16974), .A4(n16973), .ZN(
        n16977) );
  NOR2_X1 U20212 ( .A1(n16978), .A2(n16977), .ZN(n16979) );
  XOR2_X1 U20213 ( .A(n16980), .B(n16979), .Z(n17268) );
  OAI22_X1 U20214 ( .A1(n16982), .A2(n16981), .B1(n17268), .B2(n17251), .ZN(
        P3_U2673) );
  XNOR2_X1 U20215 ( .A(n16984), .B(n16983), .ZN(n17276) );
  NAND3_X1 U20216 ( .A1(n16986), .A2(P3_EBX_REG_29__SCAN_IN), .A3(n17251), 
        .ZN(n16985) );
  OAI221_X1 U20217 ( .B1(n16986), .B2(P3_EBX_REG_29__SCAN_IN), .C1(n17251), 
        .C2(n17276), .A(n16985), .ZN(P3_U2674) );
  INV_X1 U20218 ( .A(n16987), .ZN(n16995) );
  AOI21_X1 U20219 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17251), .A(n16995), .ZN(
        n16989) );
  XNOR2_X1 U20220 ( .A(n16988), .B(n16991), .ZN(n17284) );
  OAI22_X1 U20221 ( .A1(n16990), .A2(n16989), .B1(n17251), .B2(n17284), .ZN(
        P3_U2676) );
  AOI21_X1 U20222 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17251), .A(n16999), .ZN(
        n16994) );
  OAI21_X1 U20223 ( .B1(n16993), .B2(n16992), .A(n16991), .ZN(n17288) );
  OAI22_X1 U20224 ( .A1(n16995), .A2(n16994), .B1(n17251), .B2(n17288), .ZN(
        P3_U2677) );
  INV_X1 U20225 ( .A(n16996), .ZN(n17004) );
  AOI21_X1 U20226 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17251), .A(n17004), .ZN(
        n16998) );
  XNOR2_X1 U20227 ( .A(n16997), .B(n17000), .ZN(n17293) );
  OAI22_X1 U20228 ( .A1(n16999), .A2(n16998), .B1(n17251), .B2(n17293), .ZN(
        P3_U2678) );
  AOI21_X1 U20229 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17251), .A(n17009), .ZN(
        n17003) );
  OAI21_X1 U20230 ( .B1(n17002), .B2(n17001), .A(n17000), .ZN(n17299) );
  OAI22_X1 U20231 ( .A1(n17004), .A2(n17003), .B1(n17251), .B2(n17299), .ZN(
        P3_U2679) );
  INV_X1 U20232 ( .A(n17005), .ZN(n17024) );
  AOI21_X1 U20233 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17251), .A(n17024), .ZN(
        n17008) );
  XNOR2_X1 U20234 ( .A(n17007), .B(n17006), .ZN(n17305) );
  OAI22_X1 U20235 ( .A1(n17009), .A2(n17008), .B1(n17251), .B2(n17305), .ZN(
        P3_U2680) );
  AOI21_X1 U20236 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17251), .A(n17010), .ZN(
        n17023) );
  AOI22_X1 U20237 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__6__SCAN_IN), .B2(n9763), .ZN(n17021) );
  AOI22_X1 U20238 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n17117), .B1(
        P3_INSTQUEUE_REG_3__6__SCAN_IN), .B2(n17122), .ZN(n17020) );
  AOI22_X1 U20239 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n17215), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17011) );
  OAI21_X1 U20240 ( .B1(n17012), .B2(n18256), .A(n17011), .ZN(n17018) );
  AOI22_X1 U20241 ( .A1(n15435), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__6__SCAN_IN), .B2(n17205), .ZN(n17016) );
  AOI22_X1 U20242 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__6__SCAN_IN), .B2(n17212), .ZN(n17015) );
  AOI22_X1 U20243 ( .A1(n17207), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17014) );
  AOI22_X1 U20244 ( .A1(n17209), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n17189), .ZN(n17013) );
  NAND4_X1 U20245 ( .A1(n17016), .A2(n17015), .A3(n17014), .A4(n17013), .ZN(
        n17017) );
  AOI211_X1 U20246 ( .C1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .C2(n9758), .A(
        n17018), .B(n17017), .ZN(n17019) );
  NAND3_X1 U20247 ( .A1(n17021), .A2(n17020), .A3(n17019), .ZN(n17306) );
  INV_X1 U20248 ( .A(n17306), .ZN(n17022) );
  OAI22_X1 U20249 ( .A1(n17024), .A2(n17023), .B1(n17022), .B2(n17251), .ZN(
        P3_U2681) );
  OR2_X1 U20250 ( .A1(n17254), .A2(n17025), .ZN(n17050) );
  AOI22_X1 U20251 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(n9763), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17029) );
  AOI22_X1 U20252 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n15600), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17028) );
  AOI22_X1 U20253 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17027) );
  AOI22_X1 U20254 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17026) );
  NAND4_X1 U20255 ( .A1(n17029), .A2(n17028), .A3(n17027), .A4(n17026), .ZN(
        n17035) );
  AOI22_X1 U20256 ( .A1(n17207), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17033) );
  AOI22_X1 U20257 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17032) );
  AOI22_X1 U20258 ( .A1(n17209), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17031) );
  AOI22_X1 U20259 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17205), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17030) );
  NAND4_X1 U20260 ( .A1(n17033), .A2(n17032), .A3(n17031), .A4(n17030), .ZN(
        n17034) );
  NOR2_X1 U20261 ( .A1(n17035), .A2(n17034), .ZN(n17312) );
  OR2_X1 U20262 ( .A1(n17312), .A2(n17251), .ZN(n17036) );
  OAI221_X1 U20263 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n17038), .C1(n17037), 
        .C2(n17050), .A(n17036), .ZN(P3_U2682) );
  AOI22_X1 U20264 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17042) );
  AOI22_X1 U20265 ( .A1(n9763), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17041) );
  AOI22_X1 U20266 ( .A1(n17207), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9758), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17040) );
  AOI22_X1 U20267 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17039) );
  NAND4_X1 U20268 ( .A1(n17042), .A2(n17041), .A3(n17040), .A4(n17039), .ZN(
        n17048) );
  AOI22_X1 U20269 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n15600), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17046) );
  AOI22_X1 U20270 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17045) );
  AOI22_X1 U20271 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17044) );
  AOI22_X1 U20272 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17043) );
  NAND4_X1 U20273 ( .A1(n17046), .A2(n17045), .A3(n17044), .A4(n17043), .ZN(
        n17047) );
  NOR2_X1 U20274 ( .A1(n17048), .A2(n17047), .ZN(n17319) );
  INV_X1 U20275 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n20990) );
  NOR4_X1 U20276 ( .A1(n17247), .A2(n17049), .A3(n20990), .A4(n17078), .ZN(
        n17090) );
  AND2_X1 U20277 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17090), .ZN(n17063) );
  AOI21_X1 U20278 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17063), .A(
        P3_EBX_REG_20__SCAN_IN), .ZN(n17051) );
  OAI22_X1 U20279 ( .A1(n17319), .A2(n17251), .B1(n17051), .B2(n17050), .ZN(
        P3_U2683) );
  AOI22_X1 U20280 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17055) );
  AOI22_X1 U20281 ( .A1(n17207), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17054) );
  AOI22_X1 U20282 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17053) );
  AOI22_X1 U20283 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17052) );
  NAND4_X1 U20284 ( .A1(n17055), .A2(n17054), .A3(n17053), .A4(n17052), .ZN(
        n17061) );
  AOI22_X1 U20285 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17059) );
  AOI22_X1 U20286 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17058) );
  AOI22_X1 U20287 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n15600), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17057) );
  AOI22_X1 U20288 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17056) );
  NAND4_X1 U20289 ( .A1(n17059), .A2(n17058), .A3(n17057), .A4(n17056), .ZN(
        n17060) );
  NOR2_X1 U20290 ( .A1(n17061), .A2(n17060), .ZN(n17324) );
  OAI221_X1 U20291 ( .B1(n17063), .B2(P3_EBX_REG_19__SCAN_IN), .C1(n17065), 
        .C2(n17062), .A(n17251), .ZN(n17064) );
  OAI21_X1 U20292 ( .B1(n17324), .B2(n17251), .A(n17064), .ZN(P3_U2684) );
  INV_X1 U20293 ( .A(n17065), .ZN(n17077) );
  AOI21_X1 U20294 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17251), .A(n17090), .ZN(
        n17076) );
  AOI22_X1 U20295 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17069) );
  AOI22_X1 U20296 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17068) );
  AOI22_X1 U20297 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17067) );
  AOI22_X1 U20298 ( .A1(n9758), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17066) );
  NAND4_X1 U20299 ( .A1(n17069), .A2(n17068), .A3(n17067), .A4(n17066), .ZN(
        n17075) );
  AOI22_X1 U20300 ( .A1(n17207), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17224), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17073) );
  AOI22_X1 U20301 ( .A1(n17208), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n15600), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17072) );
  AOI22_X1 U20302 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17071) );
  AOI22_X1 U20303 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17070) );
  NAND4_X1 U20304 ( .A1(n17073), .A2(n17072), .A3(n17071), .A4(n17070), .ZN(
        n17074) );
  NOR2_X1 U20305 ( .A1(n17075), .A2(n17074), .ZN(n17328) );
  OAI22_X1 U20306 ( .A1(n17077), .A2(n17076), .B1(n17328), .B2(n17251), .ZN(
        P3_U2685) );
  NOR2_X1 U20307 ( .A1(n17247), .A2(n17078), .ZN(n17102) );
  AOI22_X1 U20308 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17251), .B1(
        P3_EBX_REG_16__SCAN_IN), .B2(n17102), .ZN(n17089) );
  AOI22_X1 U20309 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17082) );
  AOI22_X1 U20310 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17207), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17081) );
  AOI22_X1 U20311 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17080) );
  AOI22_X1 U20312 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n15600), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17079) );
  NAND4_X1 U20313 ( .A1(n17082), .A2(n17081), .A3(n17080), .A4(n17079), .ZN(
        n17088) );
  AOI22_X1 U20314 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17086) );
  AOI22_X1 U20315 ( .A1(n17209), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17085) );
  AOI22_X1 U20316 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17205), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17084) );
  AOI22_X1 U20317 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17083) );
  NAND4_X1 U20318 ( .A1(n17086), .A2(n17085), .A3(n17084), .A4(n17083), .ZN(
        n17087) );
  NOR2_X1 U20319 ( .A1(n17088), .A2(n17087), .ZN(n17335) );
  OAI22_X1 U20320 ( .A1(n17090), .A2(n17089), .B1(n17335), .B2(n17251), .ZN(
        P3_U2686) );
  AOI22_X1 U20321 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17094) );
  AOI22_X1 U20322 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9758), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17093) );
  AOI22_X1 U20323 ( .A1(n17207), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17092) );
  AOI22_X1 U20324 ( .A1(n17209), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17091) );
  NAND4_X1 U20325 ( .A1(n17094), .A2(n17093), .A3(n17092), .A4(n17091), .ZN(
        n17100) );
  AOI22_X1 U20326 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17098) );
  AOI22_X1 U20327 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17097) );
  AOI22_X1 U20328 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17096) );
  AOI22_X1 U20329 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17095) );
  NAND4_X1 U20330 ( .A1(n17098), .A2(n17097), .A3(n17096), .A4(n17095), .ZN(
        n17099) );
  NOR2_X1 U20331 ( .A1(n17100), .A2(n17099), .ZN(n17341) );
  NOR2_X1 U20332 ( .A1(n17254), .A2(n17101), .ZN(n17114) );
  AOI22_X1 U20333 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17114), .B1(n17102), 
        .B2(n20990), .ZN(n17103) );
  OAI21_X1 U20334 ( .B1(n17341), .B2(n17251), .A(n17103), .ZN(P3_U2687) );
  AOI22_X1 U20335 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17107) );
  AOI22_X1 U20336 ( .A1(n9758), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17106) );
  AOI22_X1 U20337 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17105) );
  AOI22_X1 U20338 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17104) );
  NAND4_X1 U20339 ( .A1(n17107), .A2(n17106), .A3(n17105), .A4(n17104), .ZN(
        n17113) );
  AOI22_X1 U20340 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17205), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17111) );
  AOI22_X1 U20341 ( .A1(n15593), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n15600), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17110) );
  AOI22_X1 U20342 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17109) );
  AOI22_X1 U20343 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17108) );
  NAND4_X1 U20344 ( .A1(n17111), .A2(n17110), .A3(n17109), .A4(n17108), .ZN(
        n17112) );
  NOR2_X1 U20345 ( .A1(n17113), .A2(n17112), .ZN(n17345) );
  OAI21_X1 U20346 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17115), .A(n17114), .ZN(
        n17116) );
  OAI21_X1 U20347 ( .B1(n17345), .B2(n17251), .A(n17116), .ZN(P3_U2688) );
  AOI22_X1 U20348 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n17213), .B1(
        P3_INSTQUEUE_REG_3__6__SCAN_IN), .B2(n17117), .ZN(n17121) );
  AOI22_X1 U20349 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__6__SCAN_IN), .B2(n17212), .ZN(n17120) );
  AOI22_X1 U20350 ( .A1(n9758), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__6__SCAN_IN), .B2(n17205), .ZN(n17119) );
  AOI22_X1 U20351 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17118) );
  NAND4_X1 U20352 ( .A1(n17121), .A2(n17120), .A3(n17119), .A4(n17118), .ZN(
        n17129) );
  AOI22_X1 U20353 ( .A1(n17207), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17127) );
  AOI22_X1 U20354 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n17217), .B1(
        P3_INSTQUEUE_REG_11__6__SCAN_IN), .B2(n9763), .ZN(n17126) );
  AOI22_X1 U20355 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n17122), .ZN(n17125) );
  AOI22_X1 U20356 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n15559), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17124) );
  NAND4_X1 U20357 ( .A1(n17127), .A2(n17126), .A3(n17125), .A4(n17124), .ZN(
        n17128) );
  NOR2_X1 U20358 ( .A1(n17129), .A2(n17128), .ZN(n17351) );
  NOR2_X1 U20359 ( .A1(n17254), .A2(n17131), .ZN(n17143) );
  NOR2_X1 U20360 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17247), .ZN(n17130) );
  AOI22_X1 U20361 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17143), .B1(n17131), 
        .B2(n17130), .ZN(n17132) );
  OAI21_X1 U20362 ( .B1(n17351), .B2(n17251), .A(n17132), .ZN(P3_U2689) );
  AOI22_X1 U20363 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17136) );
  AOI22_X1 U20364 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17135) );
  AOI22_X1 U20365 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17134) );
  AOI22_X1 U20366 ( .A1(n17209), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17133) );
  NAND4_X1 U20367 ( .A1(n17136), .A2(n17135), .A3(n17134), .A4(n17133), .ZN(
        n17142) );
  AOI22_X1 U20368 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17140) );
  AOI22_X1 U20369 ( .A1(n9758), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17205), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17139) );
  AOI22_X1 U20370 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n15600), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17138) );
  AOI22_X1 U20371 ( .A1(n9763), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17137) );
  NAND4_X1 U20372 ( .A1(n17140), .A2(n17139), .A3(n17138), .A4(n17137), .ZN(
        n17141) );
  NOR2_X1 U20373 ( .A1(n17142), .A2(n17141), .ZN(n17352) );
  INV_X1 U20374 ( .A(n17156), .ZN(n17144) );
  OAI21_X1 U20375 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n17144), .A(n17143), .ZN(
        n17145) );
  OAI21_X1 U20376 ( .B1(n17352), .B2(n17251), .A(n17145), .ZN(P3_U2690) );
  AOI22_X1 U20377 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17149) );
  AOI22_X1 U20378 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17148) );
  AOI22_X1 U20379 ( .A1(n17207), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17224), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17147) );
  AOI22_X1 U20380 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17146) );
  NAND4_X1 U20381 ( .A1(n17149), .A2(n17148), .A3(n17147), .A4(n17146), .ZN(
        n17155) );
  AOI22_X1 U20382 ( .A1(n17208), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n15600), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17153) );
  AOI22_X1 U20383 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17152) );
  AOI22_X1 U20384 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17151) );
  AOI22_X1 U20385 ( .A1(n17209), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17150) );
  NAND4_X1 U20386 ( .A1(n17153), .A2(n17152), .A3(n17151), .A4(n17150), .ZN(
        n17154) );
  NOR2_X1 U20387 ( .A1(n17155), .A2(n17154), .ZN(n17356) );
  OAI21_X1 U20388 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17172), .A(n17156), .ZN(
        n17157) );
  AOI22_X1 U20389 ( .A1(n17254), .A2(n17356), .B1(n17157), .B2(n17251), .ZN(
        P3_U2691) );
  AOI21_X1 U20390 ( .B1(n17158), .B2(n17186), .A(n17254), .ZN(n17159) );
  INV_X1 U20391 ( .A(n17159), .ZN(n17171) );
  AOI22_X1 U20392 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17169) );
  AOI22_X1 U20393 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17168) );
  INV_X1 U20394 ( .A(n17189), .ZN(n17211) );
  AOI22_X1 U20395 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17160) );
  OAI21_X1 U20396 ( .B1(n17211), .B2(n20907), .A(n17160), .ZN(n17166) );
  AOI22_X1 U20397 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17164) );
  AOI22_X1 U20398 ( .A1(n17209), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17163) );
  AOI22_X1 U20399 ( .A1(n17208), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17162) );
  AOI22_X1 U20400 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17161) );
  NAND4_X1 U20401 ( .A1(n17164), .A2(n17163), .A3(n17162), .A4(n17161), .ZN(
        n17165) );
  AOI211_X1 U20402 ( .C1(n9764), .C2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A(
        n17166), .B(n17165), .ZN(n17167) );
  NAND3_X1 U20403 ( .A1(n17169), .A2(n17168), .A3(n17167), .ZN(n17359) );
  INV_X1 U20404 ( .A(n17359), .ZN(n17170) );
  OAI22_X1 U20405 ( .A1(n17172), .A2(n17171), .B1(n17170), .B2(n17251), .ZN(
        P3_U2692) );
  AOI22_X1 U20406 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17185) );
  AOI22_X1 U20407 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17184) );
  AOI22_X1 U20408 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17174) );
  OAI21_X1 U20409 ( .B1(n17175), .B2(n20891), .A(n17174), .ZN(n17182) );
  AOI22_X1 U20410 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(n9758), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17180) );
  AOI22_X1 U20411 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17179) );
  AOI22_X1 U20412 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n15600), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17178) );
  AOI22_X1 U20413 ( .A1(n17209), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17177) );
  NAND4_X1 U20414 ( .A1(n17180), .A2(n17179), .A3(n17178), .A4(n17177), .ZN(
        n17181) );
  AOI211_X1 U20415 ( .C1(n17215), .C2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n17182), .B(n17181), .ZN(n17183) );
  NAND3_X1 U20416 ( .A1(n17185), .A2(n17184), .A3(n17183), .ZN(n17362) );
  INV_X1 U20417 ( .A(n17362), .ZN(n17188) );
  OAI21_X1 U20418 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17202), .A(n17186), .ZN(
        n17187) );
  AOI22_X1 U20419 ( .A1(n17254), .A2(n17188), .B1(n17187), .B2(n17251), .ZN(
        P3_U2693) );
  AOI22_X1 U20420 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17193) );
  AOI22_X1 U20421 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17192) );
  AOI22_X1 U20422 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17191) );
  AOI22_X1 U20423 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17190) );
  NAND4_X1 U20424 ( .A1(n17193), .A2(n17192), .A3(n17191), .A4(n17190), .ZN(
        n17200) );
  AOI22_X1 U20425 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17205), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17198) );
  AOI22_X1 U20426 ( .A1(n9763), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17197) );
  AOI22_X1 U20427 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17196) );
  AOI22_X1 U20428 ( .A1(n17207), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n15600), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17195) );
  NAND4_X1 U20429 ( .A1(n17198), .A2(n17197), .A3(n17196), .A4(n17195), .ZN(
        n17199) );
  NOR2_X1 U20430 ( .A1(n17200), .A2(n17199), .ZN(n17366) );
  NAND2_X1 U20431 ( .A1(n17251), .A2(n17201), .ZN(n17228) );
  NAND2_X1 U20432 ( .A1(n9796), .A2(n17202), .ZN(n17203) );
  OAI21_X1 U20433 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17228), .A(n17203), .ZN(
        n17204) );
  AOI21_X1 U20434 ( .B1(n17254), .B2(n17366), .A(n17204), .ZN(P3_U2694) );
  AOI22_X1 U20435 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17205), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17227) );
  AOI22_X1 U20436 ( .A1(n17207), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17226) );
  AOI22_X1 U20437 ( .A1(n17209), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17210) );
  OAI21_X1 U20438 ( .B1(n17211), .B2(n18226), .A(n17210), .ZN(n17223) );
  AOI22_X1 U20439 ( .A1(n9764), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17221) );
  AOI22_X1 U20440 ( .A1(n9758), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17220) );
  AOI22_X1 U20441 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17219) );
  AOI22_X1 U20442 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17218) );
  NAND4_X1 U20443 ( .A1(n17221), .A2(n17220), .A3(n17219), .A4(n17218), .ZN(
        n17222) );
  AOI211_X1 U20444 ( .C1(n17224), .C2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n17223), .B(n17222), .ZN(n17225) );
  NAND3_X1 U20445 ( .A1(n17227), .A2(n17226), .A3(n17225), .ZN(n17369) );
  INV_X1 U20446 ( .A(n17369), .ZN(n17230) );
  NOR2_X1 U20447 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17234), .ZN(n17229) );
  OAI22_X1 U20448 ( .A1(n17230), .A2(n17251), .B1(n17229), .B2(n17228), .ZN(
        P3_U2695) );
  INV_X1 U20449 ( .A(n17231), .ZN(n17232) );
  OAI21_X1 U20450 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n17232), .A(n17251), .ZN(
        n17233) );
  OAI22_X1 U20451 ( .A1(n17234), .A2(n17233), .B1(n18264), .B2(n17251), .ZN(
        P3_U2696) );
  NAND2_X1 U20452 ( .A1(n9796), .A2(n9756), .ZN(n17258) );
  NOR2_X1 U20453 ( .A1(n17235), .A2(n17258), .ZN(n17249) );
  NAND2_X1 U20454 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17246), .ZN(n17240) );
  NOR2_X1 U20455 ( .A1(n20968), .A2(n17240), .ZN(n17242) );
  AOI21_X1 U20456 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17251), .A(n17242), .ZN(
        n17239) );
  INV_X1 U20457 ( .A(n17236), .ZN(n17237) );
  NOR2_X1 U20458 ( .A1(n17237), .A2(n17258), .ZN(n17238) );
  OAI22_X1 U20459 ( .A1(n17239), .A2(n17238), .B1(n18256), .B2(n17251), .ZN(
        P3_U2697) );
  INV_X1 U20460 ( .A(n17240), .ZN(n17244) );
  AOI21_X1 U20461 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17251), .A(n17244), .ZN(
        n17241) );
  INV_X1 U20462 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18250) );
  OAI22_X1 U20463 ( .A1(n17242), .A2(n17241), .B1(n18250), .B2(n17251), .ZN(
        P3_U2698) );
  AOI21_X1 U20464 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17251), .A(n17246), .ZN(
        n17243) );
  OAI22_X1 U20465 ( .A1(n17244), .A2(n17243), .B1(n18245), .B2(n17251), .ZN(
        P3_U2699) );
  AOI21_X1 U20466 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17251), .A(n17249), .ZN(
        n17245) );
  OAI22_X1 U20467 ( .A1(n17246), .A2(n17245), .B1(n20907), .B2(n17251), .ZN(
        P3_U2700) );
  INV_X1 U20468 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18236) );
  NOR2_X1 U20469 ( .A1(n17257), .A2(n17252), .ZN(n17248) );
  AOI221_X1 U20470 ( .B1(n17248), .B2(n9756), .C1(n17247), .C2(n9756), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n17250) );
  AOI211_X1 U20471 ( .C1(n17254), .C2(n18236), .A(n17250), .B(n17249), .ZN(
        P3_U2701) );
  OAI222_X1 U20472 ( .A1(n17258), .A2(n17253), .B1(n17252), .B2(n9756), .C1(
        n18230), .C2(n17251), .ZN(P3_U2702) );
  NAND2_X1 U20473 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17254), .ZN(
        n17255) );
  OAI221_X1 U20474 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17258), .C1(n17257), 
        .C2(n9756), .A(n17255), .ZN(P3_U2703) );
  NAND2_X1 U20475 ( .A1(n17348), .A2(n17259), .ZN(n17311) );
  INV_X1 U20476 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17479) );
  INV_X1 U20477 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17416) );
  INV_X1 U20478 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17475) );
  INV_X1 U20479 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17419) );
  INV_X1 U20480 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17432) );
  NAND3_X1 U20481 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(P3_EAX_REG_7__SCAN_IN), 
        .A3(P3_EAX_REG_0__SCAN_IN), .ZN(n17262) );
  NAND4_X1 U20482 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(P3_EAX_REG_5__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n17261) );
  NAND2_X1 U20483 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17371), .ZN(n17370) );
  NAND3_X1 U20484 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .A3(P3_EAX_REG_11__SCAN_IN), .ZN(n17346) );
  NAND3_X1 U20485 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(P3_EAX_REG_14__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .ZN(n17263) );
  INV_X1 U20486 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n20931) );
  INV_X1 U20487 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17421) );
  INV_X1 U20488 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17428) );
  INV_X1 U20489 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17467) );
  NAND2_X1 U20490 ( .A1(n9796), .A2(n17300), .ZN(n17294) );
  NAND2_X1 U20491 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17273), .ZN(n17272) );
  NOR2_X1 U20492 ( .A1(P3_EAX_REG_31__SCAN_IN), .A2(n17272), .ZN(n17265) );
  NAND2_X1 U20493 ( .A1(n17392), .A2(n17272), .ZN(n17271) );
  OAI21_X1 U20494 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17401), .A(n17271), .ZN(
        n17264) );
  AOI22_X1 U20495 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17265), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17264), .ZN(n17266) );
  OAI21_X1 U20496 ( .B1(n21051), .B2(n17311), .A(n17266), .ZN(P3_U2704) );
  INV_X1 U20497 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17483) );
  NOR2_X2 U20498 ( .A1(n17267), .A2(n17392), .ZN(n17337) );
  OAI22_X1 U20499 ( .A1(n17268), .A2(n17394), .B1(n18251), .B2(n17311), .ZN(
        n17269) );
  AOI21_X1 U20500 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n17337), .A(n17269), .ZN(
        n17270) );
  OAI221_X1 U20501 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17272), .C1(n17483), 
        .C2(n17271), .A(n17270), .ZN(P3_U2705) );
  AOI22_X1 U20502 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17337), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17336), .ZN(n17275) );
  OAI211_X1 U20503 ( .C1(n17273), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17392), .B(
        n17272), .ZN(n17274) );
  OAI211_X1 U20504 ( .C1(n17394), .C2(n17276), .A(n17275), .B(n17274), .ZN(
        P3_U2706) );
  AOI22_X1 U20505 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17337), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17336), .ZN(n17279) );
  OAI211_X1 U20506 ( .C1(n9818), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17392), .B(
        n17277), .ZN(n17278) );
  OAI211_X1 U20507 ( .C1(n17394), .C2(n17280), .A(n17279), .B(n17278), .ZN(
        P3_U2707) );
  AOI22_X1 U20508 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17337), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17336), .ZN(n17283) );
  AOI211_X1 U20509 ( .C1(n17479), .C2(n17285), .A(n9818), .B(n17348), .ZN(
        n17281) );
  INV_X1 U20510 ( .A(n17281), .ZN(n17282) );
  OAI211_X1 U20511 ( .C1(n17394), .C2(n17284), .A(n17283), .B(n17282), .ZN(
        P3_U2708) );
  AOI22_X1 U20512 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17337), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17336), .ZN(n17287) );
  OAI211_X1 U20513 ( .C1(n17289), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17392), .B(
        n17285), .ZN(n17286) );
  OAI211_X1 U20514 ( .C1(n17288), .C2(n17394), .A(n17287), .B(n17286), .ZN(
        P3_U2709) );
  AOI22_X1 U20515 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17337), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17336), .ZN(n17292) );
  AOI211_X1 U20516 ( .C1(n17416), .C2(n17295), .A(n17289), .B(n17348), .ZN(
        n17290) );
  INV_X1 U20517 ( .A(n17290), .ZN(n17291) );
  OAI211_X1 U20518 ( .C1(n17293), .C2(n17394), .A(n17292), .B(n17291), .ZN(
        P3_U2710) );
  AOI22_X1 U20519 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17337), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17336), .ZN(n17298) );
  OAI21_X1 U20520 ( .B1(n17475), .B2(n17348), .A(n17294), .ZN(n17296) );
  NAND2_X1 U20521 ( .A1(n17296), .A2(n17295), .ZN(n17297) );
  OAI211_X1 U20522 ( .C1(n17299), .C2(n17394), .A(n17298), .B(n17297), .ZN(
        P3_U2711) );
  AOI211_X1 U20523 ( .C1(n17419), .C2(n17301), .A(n17348), .B(n17300), .ZN(
        n17302) );
  AOI21_X1 U20524 ( .B1(n17336), .B2(BUF2_REG_23__SCAN_IN), .A(n17302), .ZN(
        n17304) );
  NAND2_X1 U20525 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17337), .ZN(n17303) );
  OAI211_X1 U20526 ( .C1(n17305), .C2(n17394), .A(n17304), .B(n17303), .ZN(
        P3_U2712) );
  NAND2_X1 U20527 ( .A1(n9796), .A2(n9817), .ZN(n17329) );
  NAND2_X1 U20528 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17330), .ZN(n17325) );
  NAND3_X1 U20529 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .A3(n17320), .ZN(n17310) );
  AOI22_X1 U20530 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17336), .B1(n17399), .B2(
        n17306), .ZN(n17309) );
  NAND2_X1 U20531 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17320), .ZN(n17316) );
  NAND2_X1 U20532 ( .A1(n17392), .A2(n17316), .ZN(n17315) );
  OAI21_X1 U20533 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17401), .A(n17315), .ZN(
        n17307) );
  AOI22_X1 U20534 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17337), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17307), .ZN(n17308) );
  OAI211_X1 U20535 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n17310), .A(n17309), .B(
        n17308), .ZN(P3_U2713) );
  INV_X1 U20536 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17423) );
  OAI22_X1 U20537 ( .A1(n17312), .A2(n17394), .B1(n14963), .B2(n17311), .ZN(
        n17313) );
  AOI21_X1 U20538 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17337), .A(n17313), .ZN(
        n17314) );
  OAI221_X1 U20539 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17316), .C1(n17423), 
        .C2(n17315), .A(n17314), .ZN(P3_U2714) );
  AOI22_X1 U20540 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17337), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17336), .ZN(n17318) );
  OAI211_X1 U20541 ( .C1(n17320), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17392), .B(
        n17316), .ZN(n17317) );
  OAI211_X1 U20542 ( .C1(n17319), .C2(n17394), .A(n17318), .B(n17317), .ZN(
        P3_U2715) );
  AOI22_X1 U20543 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17337), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17336), .ZN(n17323) );
  AOI211_X1 U20544 ( .C1(n20931), .C2(n17325), .A(n17320), .B(n17348), .ZN(
        n17321) );
  INV_X1 U20545 ( .A(n17321), .ZN(n17322) );
  OAI211_X1 U20546 ( .C1(n17324), .C2(n17394), .A(n17323), .B(n17322), .ZN(
        P3_U2716) );
  AOI22_X1 U20547 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17337), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17336), .ZN(n17327) );
  OAI211_X1 U20548 ( .C1(n17330), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17392), .B(
        n17325), .ZN(n17326) );
  OAI211_X1 U20549 ( .C1(n17328), .C2(n17394), .A(n17327), .B(n17326), .ZN(
        P3_U2717) );
  AOI22_X1 U20550 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17337), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17336), .ZN(n17334) );
  OAI21_X1 U20551 ( .B1(n17467), .B2(n17348), .A(n17329), .ZN(n17332) );
  INV_X1 U20552 ( .A(n17330), .ZN(n17331) );
  NAND2_X1 U20553 ( .A1(n17332), .A2(n17331), .ZN(n17333) );
  OAI211_X1 U20554 ( .C1(n17335), .C2(n17394), .A(n17334), .B(n17333), .ZN(
        P3_U2718) );
  AOI22_X1 U20555 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17337), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17336), .ZN(n17340) );
  AOI211_X1 U20556 ( .C1(n17432), .C2(n17342), .A(n17348), .B(n9817), .ZN(
        n17338) );
  INV_X1 U20557 ( .A(n17338), .ZN(n17339) );
  OAI211_X1 U20558 ( .C1(n17341), .C2(n17394), .A(n17340), .B(n17339), .ZN(
        P3_U2719) );
  OAI211_X1 U20559 ( .C1(P3_EAX_REG_15__SCAN_IN), .C2(n17347), .A(n17392), .B(
        n17342), .ZN(n17344) );
  NAND2_X1 U20560 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17400), .ZN(n17343) );
  OAI211_X1 U20561 ( .C1(n17345), .C2(n17394), .A(n17344), .B(n17343), .ZN(
        P3_U2720) );
  NAND4_X1 U20562 ( .A1(n9796), .A2(P3_EAX_REG_9__SCAN_IN), .A3(
        P3_EAX_REG_8__SCAN_IN), .A4(n17371), .ZN(n17364) );
  INV_X1 U20563 ( .A(n17364), .ZN(n17368) );
  NAND2_X1 U20564 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17368), .ZN(n17361) );
  NOR2_X1 U20565 ( .A1(n17346), .A2(n17361), .ZN(n17353) );
  INV_X1 U20566 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17510) );
  AOI22_X1 U20567 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17400), .B1(n17353), .B2(
        n17510), .ZN(n17350) );
  OR3_X1 U20568 ( .A1(n17510), .A2(n17348), .A3(n17347), .ZN(n17349) );
  OAI211_X1 U20569 ( .C1(n17351), .C2(n17394), .A(n17350), .B(n17349), .ZN(
        P3_U2721) );
  INV_X1 U20570 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17500) );
  NOR2_X1 U20571 ( .A1(n17500), .A2(n17361), .ZN(n17355) );
  AND2_X1 U20572 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17355), .ZN(n17358) );
  AOI21_X1 U20573 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17392), .A(n17358), .ZN(
        n17354) );
  OAI222_X1 U20574 ( .A1(n17397), .A2(n17508), .B1(n17354), .B2(n17353), .C1(
        n17394), .C2(n17352), .ZN(P3_U2722) );
  AOI21_X1 U20575 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17392), .A(n17355), .ZN(
        n17357) );
  OAI222_X1 U20576 ( .A1(n17397), .A2(n17503), .B1(n17358), .B2(n17357), .C1(
        n17394), .C2(n17356), .ZN(P3_U2723) );
  NAND2_X1 U20577 ( .A1(n17392), .A2(n17361), .ZN(n17365) );
  AOI22_X1 U20578 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17400), .B1(n17399), .B2(
        n17359), .ZN(n17360) );
  OAI221_X1 U20579 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17361), .C1(n17500), 
        .C2(n17365), .A(n17360), .ZN(P3_U2724) );
  INV_X1 U20580 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17442) );
  AOI22_X1 U20581 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17400), .B1(n17399), .B2(
        n17362), .ZN(n17363) );
  OAI221_X1 U20582 ( .B1(n17365), .B2(n17442), .C1(n17365), .C2(n17364), .A(
        n17363), .ZN(P3_U2725) );
  AND2_X1 U20583 ( .A1(n9796), .A2(n17371), .ZN(n17376) );
  AOI22_X1 U20584 ( .A1(n17376), .A2(P3_EAX_REG_8__SCAN_IN), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n17392), .ZN(n17367) );
  OAI222_X1 U20585 ( .A1(n17397), .A2(n17496), .B1(n17368), .B2(n17367), .C1(
        n17394), .C2(n17366), .ZN(P3_U2726) );
  AOI22_X1 U20586 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17400), .B1(n17399), .B2(
        n17369), .ZN(n17373) );
  OAI211_X1 U20587 ( .C1(P3_EAX_REG_8__SCAN_IN), .C2(n17371), .A(n17392), .B(
        n17370), .ZN(n17372) );
  NAND2_X1 U20588 ( .A1(n17373), .A2(n17372), .ZN(P3_U2727) );
  INV_X1 U20589 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17450) );
  INV_X1 U20590 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n20861) );
  INV_X1 U20591 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17486) );
  NOR3_X1 U20592 ( .A1(n17486), .A2(n17461), .A3(n17401), .ZN(n17391) );
  NAND2_X1 U20593 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17396), .ZN(n17384) );
  NOR2_X1 U20594 ( .A1(n20861), .A2(n17384), .ZN(n17387) );
  NAND2_X1 U20595 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17387), .ZN(n17377) );
  NOR2_X1 U20596 ( .A1(n17450), .A2(n17377), .ZN(n17380) );
  AOI21_X1 U20597 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17392), .A(n17380), .ZN(
        n17375) );
  OAI222_X1 U20598 ( .A1(n17397), .A2(n18257), .B1(n17376), .B2(n17375), .C1(
        n17394), .C2(n17374), .ZN(P3_U2728) );
  INV_X1 U20599 ( .A(n17377), .ZN(n17383) );
  AOI21_X1 U20600 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17392), .A(n17383), .ZN(
        n17379) );
  OAI222_X1 U20601 ( .A1(n18252), .A2(n17397), .B1(n17380), .B2(n17379), .C1(
        n17394), .C2(n17378), .ZN(P3_U2729) );
  AOI21_X1 U20602 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17392), .A(n17387), .ZN(
        n17382) );
  OAI222_X1 U20603 ( .A1(n18246), .A2(n17397), .B1(n17383), .B2(n17382), .C1(
        n17394), .C2(n17381), .ZN(P3_U2730) );
  INV_X1 U20604 ( .A(n17384), .ZN(n17390) );
  AOI21_X1 U20605 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17392), .A(n17390), .ZN(
        n17386) );
  OAI222_X1 U20606 ( .A1(n18241), .A2(n17397), .B1(n17387), .B2(n17386), .C1(
        n17394), .C2(n17385), .ZN(P3_U2731) );
  AOI21_X1 U20607 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17392), .A(n17396), .ZN(
        n17389) );
  OAI222_X1 U20608 ( .A1(n18237), .A2(n17397), .B1(n17390), .B2(n17389), .C1(
        n17394), .C2(n17388), .ZN(P3_U2732) );
  AOI21_X1 U20609 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17392), .A(n17391), .ZN(
        n17395) );
  OAI222_X1 U20610 ( .A1(n18231), .A2(n17397), .B1(n17396), .B2(n17395), .C1(
        n17394), .C2(n17393), .ZN(P3_U2733) );
  AOI22_X1 U20611 ( .A1(n17400), .A2(BUF2_REG_1__SCAN_IN), .B1(n17399), .B2(
        n17398), .ZN(n17406) );
  NOR2_X1 U20612 ( .A1(n17461), .A2(n17401), .ZN(n17404) );
  NOR2_X1 U20613 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17401), .ZN(n17403) );
  OAI22_X1 U20614 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17404), .B1(n17403), .B2(
        n17402), .ZN(n17405) );
  NAND2_X1 U20615 ( .A1(n17406), .A2(n17405), .ZN(P3_U2734) );
  INV_X1 U20616 ( .A(n17713), .ZN(n17881) );
  INV_X2 U20617 ( .A(n18869), .ZN(n18715) );
  NOR2_X4 U20618 ( .A1(n18715), .A2(n17433), .ZN(n17448) );
  AND2_X1 U20619 ( .A1(n17448), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NAND2_X1 U20620 ( .A1(n17433), .A2(n18874), .ZN(n17431) );
  AOI22_X1 U20621 ( .A1(n18715), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17408) );
  OAI21_X1 U20622 ( .B1(n17483), .B2(n17431), .A(n17408), .ZN(P3_U2737) );
  INV_X1 U20623 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17410) );
  AOI22_X1 U20624 ( .A1(n18715), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17409) );
  OAI21_X1 U20625 ( .B1(n17410), .B2(n17431), .A(n17409), .ZN(P3_U2738) );
  INV_X1 U20626 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17412) );
  AOI22_X1 U20627 ( .A1(n18715), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17411) );
  OAI21_X1 U20628 ( .B1(n17412), .B2(n17431), .A(n17411), .ZN(P3_U2739) );
  AOI22_X1 U20629 ( .A1(n18715), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17413) );
  OAI21_X1 U20630 ( .B1(n17479), .B2(n17431), .A(n17413), .ZN(P3_U2740) );
  AOI22_X1 U20631 ( .A1(n18715), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17414) );
  OAI21_X1 U20632 ( .B1(n9985), .B2(n17431), .A(n17414), .ZN(P3_U2741) );
  AOI22_X1 U20633 ( .A1(n18715), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17415) );
  OAI21_X1 U20634 ( .B1(n17416), .B2(n17431), .A(n17415), .ZN(P3_U2742) );
  AOI22_X1 U20635 ( .A1(n18715), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17417) );
  OAI21_X1 U20636 ( .B1(n17475), .B2(n17431), .A(n17417), .ZN(P3_U2743) );
  AOI22_X1 U20637 ( .A1(n18715), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17418) );
  OAI21_X1 U20638 ( .B1(n17419), .B2(n17431), .A(n17418), .ZN(P3_U2744) );
  AOI22_X1 U20639 ( .A1(n18715), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17420) );
  OAI21_X1 U20640 ( .B1(n17421), .B2(n17431), .A(n17420), .ZN(P3_U2745) );
  AOI22_X1 U20641 ( .A1(n18715), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17422) );
  OAI21_X1 U20642 ( .B1(n17423), .B2(n17431), .A(n17422), .ZN(P3_U2746) );
  INV_X1 U20643 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17425) );
  AOI22_X1 U20644 ( .A1(n18715), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17424) );
  OAI21_X1 U20645 ( .B1(n17425), .B2(n17431), .A(n17424), .ZN(P3_U2747) );
  AOI22_X1 U20646 ( .A1(n18715), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17426) );
  OAI21_X1 U20647 ( .B1(n20931), .B2(n17431), .A(n17426), .ZN(P3_U2748) );
  AOI22_X1 U20648 ( .A1(n18715), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17427) );
  OAI21_X1 U20649 ( .B1(n17428), .B2(n17431), .A(n17427), .ZN(P3_U2749) );
  AOI22_X1 U20650 ( .A1(n18715), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17429) );
  OAI21_X1 U20651 ( .B1(n17467), .B2(n17431), .A(n17429), .ZN(P3_U2750) );
  AOI22_X1 U20652 ( .A1(n18715), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17430) );
  OAI21_X1 U20653 ( .B1(n17432), .B2(n17431), .A(n17430), .ZN(P3_U2751) );
  AOI22_X1 U20654 ( .A1(n18715), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17434) );
  OAI21_X1 U20655 ( .B1(n9982), .B2(n17460), .A(n17434), .ZN(P3_U2752) );
  AOI22_X1 U20656 ( .A1(n18715), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17435) );
  OAI21_X1 U20657 ( .B1(n17510), .B2(n17460), .A(n17435), .ZN(P3_U2753) );
  INV_X1 U20658 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17437) );
  AOI22_X1 U20659 ( .A1(n18715), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17436) );
  OAI21_X1 U20660 ( .B1(n17437), .B2(n17460), .A(n17436), .ZN(P3_U2754) );
  INV_X1 U20661 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17439) );
  AOI22_X1 U20662 ( .A1(n18715), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17438) );
  OAI21_X1 U20663 ( .B1(n17439), .B2(n17460), .A(n17438), .ZN(P3_U2755) );
  AOI22_X1 U20664 ( .A1(n18715), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17440) );
  OAI21_X1 U20665 ( .B1(n17500), .B2(n17460), .A(n17440), .ZN(P3_U2756) );
  AOI22_X1 U20666 ( .A1(n18715), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17441) );
  OAI21_X1 U20667 ( .B1(n17442), .B2(n17460), .A(n17441), .ZN(P3_U2757) );
  INV_X1 U20668 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17444) );
  AOI22_X1 U20669 ( .A1(n18715), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17443) );
  OAI21_X1 U20670 ( .B1(n17444), .B2(n17460), .A(n17443), .ZN(P3_U2758) );
  INV_X1 U20671 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17494) );
  AOI22_X1 U20672 ( .A1(n18715), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17445) );
  OAI21_X1 U20673 ( .B1(n17494), .B2(n17460), .A(n17445), .ZN(P3_U2759) );
  INV_X1 U20674 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17447) );
  AOI22_X1 U20675 ( .A1(n18715), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17446) );
  OAI21_X1 U20676 ( .B1(n17447), .B2(n17460), .A(n17446), .ZN(P3_U2760) );
  AOI22_X1 U20677 ( .A1(n18715), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17449) );
  OAI21_X1 U20678 ( .B1(n17450), .B2(n17460), .A(n17449), .ZN(P3_U2761) );
  INV_X1 U20679 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17452) );
  AOI22_X1 U20680 ( .A1(n18715), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17451) );
  OAI21_X1 U20681 ( .B1(n17452), .B2(n17460), .A(n17451), .ZN(P3_U2762) );
  AOI22_X1 U20682 ( .A1(n18715), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17453) );
  OAI21_X1 U20683 ( .B1(n20861), .B2(n17460), .A(n17453), .ZN(P3_U2763) );
  INV_X1 U20684 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17455) );
  AOI22_X1 U20685 ( .A1(n18715), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17454) );
  OAI21_X1 U20686 ( .B1(n17455), .B2(n17460), .A(n17454), .ZN(P3_U2764) );
  INV_X1 U20687 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17457) );
  AOI22_X1 U20688 ( .A1(n18715), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17456) );
  OAI21_X1 U20689 ( .B1(n17457), .B2(n17460), .A(n17456), .ZN(P3_U2765) );
  AOI22_X1 U20690 ( .A1(n18715), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17458) );
  OAI21_X1 U20691 ( .B1(n17486), .B2(n17460), .A(n17458), .ZN(P3_U2766) );
  AOI22_X1 U20692 ( .A1(n18715), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17459) );
  OAI21_X1 U20693 ( .B1(n17461), .B2(n17460), .A(n17459), .ZN(P3_U2767) );
  OAI211_X1 U20694 ( .C1(n18875), .C2(n18227), .A(n9783), .B(n17462), .ZN(
        n17504) );
  NAND2_X1 U20695 ( .A1(n18227), .A2(n9783), .ZN(n18717) );
  AOI22_X1 U20696 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17505), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17511), .ZN(n17465) );
  OAI21_X1 U20697 ( .B1(n18218), .B2(n17507), .A(n17465), .ZN(P3_U2768) );
  INV_X1 U20698 ( .A(n17505), .ZN(n17514) );
  AOI22_X1 U20699 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17512), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17511), .ZN(n17466) );
  OAI21_X1 U20700 ( .B1(n17467), .B2(n17514), .A(n17466), .ZN(P3_U2769) );
  AOI22_X1 U20701 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17501), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17511), .ZN(n17468) );
  OAI21_X1 U20702 ( .B1(n18231), .B2(n17507), .A(n17468), .ZN(P3_U2770) );
  AOI22_X1 U20703 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17501), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17511), .ZN(n17469) );
  OAI21_X1 U20704 ( .B1(n18237), .B2(n17507), .A(n17469), .ZN(P3_U2771) );
  AOI22_X1 U20705 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17505), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17511), .ZN(n17470) );
  OAI21_X1 U20706 ( .B1(n18241), .B2(n17507), .A(n17470), .ZN(P3_U2772) );
  AOI22_X1 U20707 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17505), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17511), .ZN(n17471) );
  OAI21_X1 U20708 ( .B1(n18246), .B2(n17507), .A(n17471), .ZN(P3_U2773) );
  AOI22_X1 U20709 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17505), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17511), .ZN(n17472) );
  OAI21_X1 U20710 ( .B1(n18252), .B2(n17507), .A(n17472), .ZN(P3_U2774) );
  AOI22_X1 U20711 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17501), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17511), .ZN(n17473) );
  OAI21_X1 U20712 ( .B1(n18257), .B2(n17507), .A(n17473), .ZN(P3_U2775) );
  AOI22_X1 U20713 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17512), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17511), .ZN(n17474) );
  OAI21_X1 U20714 ( .B1(n17475), .B2(n17514), .A(n17474), .ZN(P3_U2776) );
  AOI22_X1 U20715 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17505), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17511), .ZN(n17476) );
  OAI21_X1 U20716 ( .B1(n17496), .B2(n17507), .A(n17476), .ZN(P3_U2777) );
  AOI22_X1 U20717 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17505), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17511), .ZN(n17477) );
  OAI21_X1 U20718 ( .B1(n17498), .B2(n17507), .A(n17477), .ZN(P3_U2778) );
  AOI22_X1 U20719 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17512), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17511), .ZN(n17478) );
  OAI21_X1 U20720 ( .B1(n17479), .B2(n17514), .A(n17478), .ZN(P3_U2779) );
  AOI22_X1 U20721 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17501), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17511), .ZN(n17480) );
  OAI21_X1 U20722 ( .B1(n17503), .B2(n17507), .A(n17480), .ZN(P3_U2780) );
  AOI22_X1 U20723 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17501), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17511), .ZN(n17481) );
  OAI21_X1 U20724 ( .B1(n17508), .B2(n17507), .A(n17481), .ZN(P3_U2781) );
  AOI22_X1 U20725 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17512), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17511), .ZN(n17482) );
  OAI21_X1 U20726 ( .B1(n17483), .B2(n17514), .A(n17482), .ZN(P3_U2782) );
  AOI22_X1 U20727 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17501), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17511), .ZN(n17484) );
  OAI21_X1 U20728 ( .B1(n18218), .B2(n17507), .A(n17484), .ZN(P3_U2783) );
  AOI22_X1 U20729 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17512), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17511), .ZN(n17485) );
  OAI21_X1 U20730 ( .B1(n17486), .B2(n17514), .A(n17485), .ZN(P3_U2784) );
  AOI22_X1 U20731 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17505), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17511), .ZN(n17487) );
  OAI21_X1 U20732 ( .B1(n18231), .B2(n17507), .A(n17487), .ZN(P3_U2785) );
  AOI22_X1 U20733 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17501), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17504), .ZN(n17488) );
  OAI21_X1 U20734 ( .B1(n18237), .B2(n17507), .A(n17488), .ZN(P3_U2786) );
  AOI22_X1 U20735 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17501), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17504), .ZN(n17489) );
  OAI21_X1 U20736 ( .B1(n18241), .B2(n17507), .A(n17489), .ZN(P3_U2787) );
  AOI22_X1 U20737 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17501), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17504), .ZN(n17490) );
  OAI21_X1 U20738 ( .B1(n18246), .B2(n17507), .A(n17490), .ZN(P3_U2788) );
  AOI22_X1 U20739 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17505), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17504), .ZN(n17491) );
  OAI21_X1 U20740 ( .B1(n18252), .B2(n17507), .A(n17491), .ZN(P3_U2789) );
  AOI22_X1 U20741 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17505), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17504), .ZN(n17492) );
  OAI21_X1 U20742 ( .B1(n18257), .B2(n17507), .A(n17492), .ZN(P3_U2790) );
  AOI22_X1 U20743 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17512), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17504), .ZN(n17493) );
  OAI21_X1 U20744 ( .B1(n17494), .B2(n17514), .A(n17493), .ZN(P3_U2791) );
  AOI22_X1 U20745 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17501), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17504), .ZN(n17495) );
  OAI21_X1 U20746 ( .B1(n17496), .B2(n17507), .A(n17495), .ZN(P3_U2792) );
  AOI22_X1 U20747 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17501), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17504), .ZN(n17497) );
  OAI21_X1 U20748 ( .B1(n17498), .B2(n17507), .A(n17497), .ZN(P3_U2793) );
  AOI22_X1 U20749 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17512), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17511), .ZN(n17499) );
  OAI21_X1 U20750 ( .B1(n17500), .B2(n17514), .A(n17499), .ZN(P3_U2794) );
  AOI22_X1 U20751 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17501), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17504), .ZN(n17502) );
  OAI21_X1 U20752 ( .B1(n17503), .B2(n17507), .A(n17502), .ZN(P3_U2795) );
  AOI22_X1 U20753 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17505), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17504), .ZN(n17506) );
  OAI21_X1 U20754 ( .B1(n17508), .B2(n17507), .A(n17506), .ZN(P3_U2796) );
  AOI22_X1 U20755 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17512), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17511), .ZN(n17509) );
  OAI21_X1 U20756 ( .B1(n17510), .B2(n17514), .A(n17509), .ZN(P3_U2797) );
  AOI22_X1 U20757 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17512), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17511), .ZN(n17513) );
  OAI21_X1 U20758 ( .B1(n9982), .B2(n17514), .A(n17513), .ZN(P3_U2798) );
  INV_X1 U20759 ( .A(n17530), .ZN(n17516) );
  OAI21_X1 U20760 ( .B1(n17516), .B2(n17515), .A(n17882), .ZN(n17517) );
  AOI21_X1 U20761 ( .B1(n17713), .B2(n17518), .A(n17517), .ZN(n17558) );
  OAI21_X1 U20762 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17602), .A(
        n17558), .ZN(n17541) );
  AOI22_X1 U20763 ( .A1(n17538), .A2(n17519), .B1(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n17541), .ZN(n17535) );
  INV_X1 U20764 ( .A(n17520), .ZN(n17529) );
  AOI21_X1 U20765 ( .B1(n9839), .B2(n17521), .A(n17794), .ZN(n17528) );
  NOR4_X1 U20766 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17937), .A3(
        n17522), .A4(n17685), .ZN(n17526) );
  AOI22_X1 U20767 ( .A1(n17874), .A2(n17523), .B1(n17711), .B2(n17893), .ZN(
        n17553) );
  NAND2_X1 U20768 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17553), .ZN(
        n17544) );
  INV_X1 U20769 ( .A(n17544), .ZN(n17524) );
  NOR2_X1 U20770 ( .A1(n17874), .A2(n17711), .ZN(n17634) );
  NAND2_X1 U20771 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n9760), .ZN(n17533) );
  NOR2_X1 U20772 ( .A1(n17716), .A2(n17530), .ZN(n17542) );
  OAI211_X1 U20773 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17542), .B(n17531), .ZN(n17532) );
  NAND4_X1 U20774 ( .A1(n17535), .A2(n17534), .A3(n17533), .A4(n17532), .ZN(
        P3_U2802) );
  AOI21_X1 U20775 ( .B1(n17781), .B2(n17537), .A(n17536), .ZN(n17900) );
  OAI22_X1 U20776 ( .A1(n15697), .A2(n18800), .B1(n17740), .B2(n17539), .ZN(
        n17540) );
  AOI221_X1 U20777 ( .B1(n17542), .B2(n21063), .C1(n17541), .C2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(n17540), .ZN(n17547) );
  NOR2_X1 U20778 ( .A1(n17543), .A2(n17685), .ZN(n17545) );
  OAI21_X1 U20779 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17545), .A(
        n17544), .ZN(n17546) );
  OAI211_X1 U20780 ( .C1(n17900), .C2(n17794), .A(n17547), .B(n17546), .ZN(
        P3_U2803) );
  AOI21_X1 U20781 ( .B1(n17548), .B2(n18607), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17557) );
  NAND2_X1 U20782 ( .A1(n17740), .A2(n17602), .ZN(n17876) );
  AOI22_X1 U20783 ( .A1(n9760), .A2(P3_REIP_REG_26__SCAN_IN), .B1(n17549), 
        .B2(n17876), .ZN(n17556) );
  NOR4_X1 U20784 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17568), .A3(
        n17937), .A4(n17909), .ZN(n17901) );
  INV_X1 U20785 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17552) );
  AOI21_X1 U20786 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17551), .A(
        n17550), .ZN(n17905) );
  OAI22_X1 U20787 ( .A1(n17553), .A2(n17552), .B1(n17905), .B2(n17794), .ZN(
        n17554) );
  AOI21_X1 U20788 ( .B1(n17613), .B2(n17901), .A(n17554), .ZN(n17555) );
  OAI211_X1 U20789 ( .C1(n17558), .C2(n17557), .A(n17556), .B(n17555), .ZN(
        P3_U2804) );
  XNOR2_X1 U20790 ( .A(n17559), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17915) );
  INV_X1 U20791 ( .A(n17882), .ZN(n17869) );
  AND2_X1 U20792 ( .A1(n17561), .A2(n18607), .ZN(n17588) );
  AOI211_X1 U20793 ( .C1(n17713), .C2(n17560), .A(n17869), .B(n17588), .ZN(
        n17590) );
  OAI21_X1 U20794 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17602), .A(
        n17590), .ZN(n17578) );
  NOR2_X1 U20795 ( .A1(n17716), .A2(n17561), .ZN(n17580) );
  OAI211_X1 U20796 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17580), .B(n17562), .ZN(n17563) );
  NAND2_X1 U20797 ( .A1(n9760), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n17913) );
  OAI211_X1 U20798 ( .C1(n17740), .C2(n17564), .A(n17563), .B(n17913), .ZN(
        n17571) );
  XNOR2_X1 U20799 ( .A(n17568), .B(n17565), .ZN(n17920) );
  OAI21_X1 U20800 ( .B1(n17567), .B2(n17781), .A(n17566), .ZN(n17569) );
  XNOR2_X1 U20801 ( .A(n17569), .B(n17568), .ZN(n17916) );
  OAI22_X1 U20802 ( .A1(n17886), .A2(n17920), .B1(n17794), .B2(n17916), .ZN(
        n17570) );
  AOI211_X1 U20803 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17578), .A(
        n17571), .B(n17570), .ZN(n17572) );
  OAI21_X1 U20804 ( .B1(n17789), .B2(n17915), .A(n17572), .ZN(P3_U2805) );
  AOI21_X1 U20805 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17574), .A(
        n17573), .ZN(n17936) );
  INV_X1 U20806 ( .A(n17575), .ZN(n17576) );
  OAI22_X1 U20807 ( .A1(n15697), .A2(n18795), .B1(n17740), .B2(n17576), .ZN(
        n17577) );
  AOI221_X1 U20808 ( .B1(n17580), .B2(n17579), .C1(n17578), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17577), .ZN(n17583) );
  INV_X1 U20809 ( .A(n17581), .ZN(n17922) );
  OAI22_X1 U20810 ( .A1(n17921), .A2(n17886), .B1(n17922), .B2(n17789), .ZN(
        n17592) );
  NOR2_X1 U20811 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17907), .ZN(
        n17932) );
  AOI22_X1 U20812 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17592), .B1(
        n17613), .B2(n17932), .ZN(n17582) );
  OAI211_X1 U20813 ( .C1(n17936), .C2(n17794), .A(n17583), .B(n17582), .ZN(
        P3_U2806) );
  AOI22_X1 U20814 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17781), .B1(
        n17584), .B2(n17596), .ZN(n17585) );
  NAND2_X1 U20815 ( .A1(n17635), .A2(n17585), .ZN(n17586) );
  XNOR2_X1 U20816 ( .A(n17586), .B(n17925), .ZN(n17943) );
  NOR2_X1 U20817 ( .A1(n17937), .A2(n17685), .ZN(n17593) );
  AOI22_X1 U20818 ( .A1(n9879), .A2(n17588), .B1(n17587), .B2(n17876), .ZN(
        n17589) );
  NAND2_X1 U20819 ( .A1(n9760), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17942) );
  OAI211_X1 U20820 ( .C1(n17590), .C2(n9896), .A(n17589), .B(n17942), .ZN(
        n17591) );
  AOI221_X1 U20821 ( .B1(n17593), .B2(n17925), .C1(n17592), .C2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n17591), .ZN(n17594) );
  OAI21_X1 U20822 ( .B1(n17794), .B2(n17943), .A(n17594), .ZN(P3_U2807) );
  INV_X1 U20823 ( .A(n17635), .ZN(n17595) );
  AOI221_X1 U20824 ( .B1(n17597), .B2(n17596), .C1(n17621), .C2(n17596), .A(
        n17595), .ZN(n17598) );
  XNOR2_X1 U20825 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n17598), .ZN(
        n17955) );
  NOR2_X1 U20826 ( .A1(n17950), .A2(n17685), .ZN(n17610) );
  NOR2_X1 U20827 ( .A1(n18025), .A2(n17789), .ZN(n17694) );
  AOI21_X1 U20828 ( .B1(n17874), .B2(n17945), .A(n17694), .ZN(n17684) );
  OAI21_X1 U20829 ( .B1(n17599), .B2(n17634), .A(n17684), .ZN(n17624) );
  OAI21_X1 U20830 ( .B1(n17600), .B2(n17881), .A(n17882), .ZN(n17601) );
  AOI21_X1 U20831 ( .B1(n17843), .B2(n17603), .A(n17601), .ZN(n17628) );
  OAI21_X1 U20832 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17602), .A(
        n17628), .ZN(n17618) );
  AOI22_X1 U20833 ( .A1(n9760), .A2(P3_REIP_REG_22__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n17618), .ZN(n17606) );
  NOR2_X1 U20834 ( .A1(n17716), .A2(n17603), .ZN(n17620) );
  OAI211_X1 U20835 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17620), .B(n17604), .ZN(n17605) );
  OAI211_X1 U20836 ( .C1(n17740), .C2(n17607), .A(n17606), .B(n17605), .ZN(
        n17608) );
  AOI221_X1 U20837 ( .B1(n17610), .B2(n17609), .C1(n17624), .C2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n17608), .ZN(n17611) );
  OAI21_X1 U20838 ( .B1(n17794), .B2(n17955), .A(n17611), .ZN(P3_U2808) );
  NAND2_X1 U20839 ( .A1(n17967), .A2(n17612), .ZN(n17971) );
  NAND2_X1 U20840 ( .A1(n17614), .A2(n17613), .ZN(n17651) );
  INV_X1 U20841 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18790) );
  INV_X1 U20842 ( .A(n17615), .ZN(n17616) );
  OAI22_X1 U20843 ( .A1(n15697), .A2(n18790), .B1(n17740), .B2(n17616), .ZN(
        n17617) );
  AOI221_X1 U20844 ( .B1(n17620), .B2(n17619), .C1(n17618), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17617), .ZN(n17626) );
  NOR3_X1 U20845 ( .A1(n17781), .A2(n18001), .A3(n17621), .ZN(n17645) );
  INV_X1 U20846 ( .A(n17658), .ZN(n17646) );
  AOI22_X1 U20847 ( .A1(n17967), .A2(n17645), .B1(n17646), .B2(n17622), .ZN(
        n17623) );
  XNOR2_X1 U20848 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17623), .ZN(
        n17961) );
  AOI22_X1 U20849 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17624), .B1(
        n17748), .B2(n17961), .ZN(n17625) );
  OAI211_X1 U20850 ( .C1(n17971), .C2(n17651), .A(n17626), .B(n17625), .ZN(
        P3_U2809) );
  NAND2_X1 U20851 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17951), .ZN(
        n17981) );
  NAND2_X1 U20852 ( .A1(n9760), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n17979) );
  INV_X1 U20853 ( .A(n17979), .ZN(n17632) );
  NAND2_X1 U20854 ( .A1(n17627), .A2(n18607), .ZN(n17662) );
  AOI221_X1 U20855 ( .B1(n17630), .B2(n17629), .C1(n17662), .C2(n17629), .A(
        n17628), .ZN(n17631) );
  AOI211_X1 U20856 ( .C1(n17633), .C2(n17876), .A(n17632), .B(n17631), .ZN(
        n17638) );
  NOR2_X1 U20857 ( .A1(n17987), .A2(n17963), .ZN(n17972) );
  OAI21_X1 U20858 ( .B1(n17634), .B2(n17972), .A(n17684), .ZN(n17648) );
  OAI221_X1 U20859 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17657), 
        .C1(n17987), .C2(n17645), .A(n17635), .ZN(n17636) );
  XNOR2_X1 U20860 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17636), .ZN(
        n17977) );
  AOI22_X1 U20861 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17648), .B1(
        n17748), .B2(n17977), .ZN(n17637) );
  OAI211_X1 U20862 ( .C1(n17981), .C2(n17651), .A(n17638), .B(n17637), .ZN(
        P3_U2810) );
  AOI21_X1 U20863 ( .B1(n17843), .B2(n17640), .A(n17869), .ZN(n17664) );
  OAI21_X1 U20864 ( .B1(n17639), .B2(n17881), .A(n17664), .ZN(n17654) );
  NOR2_X1 U20865 ( .A1(n17716), .A2(n17640), .ZN(n17656) );
  NAND2_X1 U20866 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17641) );
  OAI211_X1 U20867 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17656), .B(n17641), .ZN(n17642) );
  NAND2_X1 U20868 ( .A1(n9760), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n17982) );
  OAI211_X1 U20869 ( .C1(n17740), .C2(n17643), .A(n17642), .B(n17982), .ZN(
        n17644) );
  AOI21_X1 U20870 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17654), .A(
        n17644), .ZN(n17650) );
  AOI21_X1 U20871 ( .B1(n17657), .B2(n17646), .A(n17645), .ZN(n17647) );
  XNOR2_X1 U20872 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n17647), .ZN(
        n17984) );
  AOI22_X1 U20873 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17648), .B1(
        n17748), .B2(n17984), .ZN(n17649) );
  OAI211_X1 U20874 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17651), .A(
        n17650), .B(n17649), .ZN(P3_U2811) );
  NAND2_X1 U20875 ( .A1(n17948), .A2(n18001), .ZN(n18006) );
  INV_X1 U20876 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17655) );
  OAI22_X1 U20877 ( .A1(n15697), .A2(n18783), .B1(n17740), .B2(n17652), .ZN(
        n17653) );
  AOI221_X1 U20878 ( .B1(n17656), .B2(n17655), .C1(n17654), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17653), .ZN(n17661) );
  OAI21_X1 U20879 ( .B1(n17948), .B2(n17685), .A(n17684), .ZN(n17669) );
  AOI21_X1 U20880 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n17674), .A(
        n17657), .ZN(n17659) );
  XNOR2_X1 U20881 ( .A(n17659), .B(n17658), .ZN(n18003) );
  AOI22_X1 U20882 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17669), .B1(
        n17748), .B2(n18003), .ZN(n17660) );
  OAI211_X1 U20883 ( .C1(n17685), .C2(n18006), .A(n17661), .B(n17660), .ZN(
        P3_U2812) );
  NAND2_X1 U20884 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18007), .ZN(
        n18013) );
  NAND2_X1 U20885 ( .A1(n9760), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n18011) );
  OAI221_X1 U20886 ( .B1(n17664), .B2(n17663), .C1(n17664), .C2(n17662), .A(
        n18011), .ZN(n17665) );
  AOI21_X1 U20887 ( .B1(n17666), .B2(n17876), .A(n17665), .ZN(n17671) );
  OAI21_X1 U20888 ( .B1(n17668), .B2(n18007), .A(n17667), .ZN(n18010) );
  AOI22_X1 U20889 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17669), .B1(
        n17748), .B2(n18010), .ZN(n17670) );
  OAI211_X1 U20890 ( .C1(n17685), .C2(n18013), .A(n17671), .B(n17670), .ZN(
        P3_U2813) );
  NAND2_X1 U20891 ( .A1(n17674), .A2(n18086), .ZN(n17766) );
  OAI22_X1 U20892 ( .A1(n17674), .A2(n17673), .B1(n17766), .B2(n17672), .ZN(
        n17675) );
  XNOR2_X1 U20893 ( .A(n18023), .B(n17675), .ZN(n18020) );
  AOI21_X1 U20894 ( .B1(n17843), .B2(n17677), .A(n17869), .ZN(n17701) );
  OAI21_X1 U20895 ( .B1(n17676), .B2(n17881), .A(n17701), .ZN(n17688) );
  AOI22_X1 U20896 ( .A1(n9760), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17688), .ZN(n17680) );
  NOR2_X1 U20897 ( .A1(n17716), .A2(n17677), .ZN(n17690) );
  OAI211_X1 U20898 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17690), .B(n17678), .ZN(n17679) );
  OAI211_X1 U20899 ( .C1(n17740), .C2(n17681), .A(n17680), .B(n17679), .ZN(
        n17682) );
  AOI21_X1 U20900 ( .B1(n17748), .B2(n18020), .A(n17682), .ZN(n17683) );
  OAI221_X1 U20901 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17685), 
        .C1(n18023), .C2(n17684), .A(n17683), .ZN(P3_U2814) );
  NOR2_X1 U20902 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17706), .ZN(
        n18030) );
  NAND2_X1 U20903 ( .A1(n17874), .A2(n17945), .ZN(n17697) );
  OAI22_X1 U20904 ( .A1(n15697), .A2(n18777), .B1(n17740), .B2(n17686), .ZN(
        n17687) );
  AOI221_X1 U20905 ( .B1(n17690), .B2(n17689), .C1(n17688), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17687), .ZN(n17696) );
  AOI21_X1 U20906 ( .B1(n17691), .B2(n17721), .A(n17698), .ZN(n17692) );
  AOI221_X1 U20907 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18080), 
        .C1(n17781), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n17692), .ZN(
        n17693) );
  XNOR2_X1 U20908 ( .A(n17693), .B(n15683), .ZN(n18034) );
  NAND2_X1 U20909 ( .A1(n18086), .A2(n18037), .ZN(n18061) );
  OAI21_X1 U20910 ( .B1(n17707), .B2(n18061), .A(n15683), .ZN(n18028) );
  AOI22_X1 U20911 ( .A1(n17748), .A2(n18034), .B1(n17694), .B2(n18028), .ZN(
        n17695) );
  OAI211_X1 U20912 ( .C1(n18030), .C2(n17697), .A(n17696), .B(n17695), .ZN(
        P3_U2815) );
  INV_X1 U20913 ( .A(n18037), .ZN(n18038) );
  NOR2_X1 U20914 ( .A1(n17726), .A2(n18038), .ZN(n17705) );
  INV_X1 U20915 ( .A(n17766), .ZN(n17746) );
  AOI22_X1 U20916 ( .A1(n17705), .A2(n17746), .B1(n17698), .B2(n18080), .ZN(
        n17699) );
  XNOR2_X1 U20917 ( .A(n17699), .B(n18047), .ZN(n18055) );
  NOR3_X1 U20918 ( .A1(n17814), .A2(n17815), .A3(n18260), .ZN(n17799) );
  NAND2_X1 U20919 ( .A1(n17700), .A2(n17799), .ZN(n17743) );
  AOI221_X1 U20920 ( .B1(n17717), .B2(n17702), .C1(n17743), .C2(n17702), .A(
        n17701), .ZN(n17703) );
  NOR2_X1 U20921 ( .A1(n15697), .A2(n18776), .ZN(n18049) );
  AOI211_X1 U20922 ( .C1(n17704), .C2(n17876), .A(n17703), .B(n18049), .ZN(
        n17710) );
  INV_X1 U20923 ( .A(n17705), .ZN(n18043) );
  AOI221_X1 U20924 ( .B1(n17994), .B2(n18047), .C1(n18043), .C2(n18047), .A(
        n17706), .ZN(n18052) );
  NOR2_X1 U20925 ( .A1(n17707), .A2(n18061), .ZN(n17708) );
  AOI221_X1 U20926 ( .B1(n17726), .B2(n18047), .C1(n18061), .C2(n18047), .A(
        n17708), .ZN(n18051) );
  AOI22_X1 U20927 ( .A1(n17874), .A2(n18052), .B1(n17711), .B2(n18051), .ZN(
        n17709) );
  OAI211_X1 U20928 ( .C1(n18055), .C2(n17794), .A(n17710), .B(n17709), .ZN(
        P3_U2816) );
  AOI22_X1 U20929 ( .A1(n17711), .A2(n18061), .B1(n17874), .B2(n18063), .ZN(
        n17733) );
  AOI22_X1 U20930 ( .A1(n17843), .A2(n17715), .B1(n17713), .B2(n17712), .ZN(
        n17714) );
  NAND2_X1 U20931 ( .A1(n17714), .A2(n17882), .ZN(n17727) );
  NOR2_X1 U20932 ( .A1(n17716), .A2(n17715), .ZN(n17729) );
  OAI211_X1 U20933 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17729), .B(n17717), .ZN(n17718) );
  NAND2_X1 U20934 ( .A1(n9760), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n18070) );
  OAI211_X1 U20935 ( .C1(n17740), .C2(n17719), .A(n17718), .B(n18070), .ZN(
        n17720) );
  AOI21_X1 U20936 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17727), .A(
        n17720), .ZN(n17725) );
  AOI22_X1 U20937 ( .A1(n17721), .A2(n18037), .B1(n17781), .B2(n18080), .ZN(
        n17722) );
  AOI21_X1 U20938 ( .B1(n17730), .B2(n17781), .A(n17722), .ZN(n17723) );
  XNOR2_X1 U20939 ( .A(n17723), .B(n17726), .ZN(n18057) );
  NOR2_X1 U20940 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18038), .ZN(
        n18056) );
  AOI22_X1 U20941 ( .A1(n17748), .A2(n18057), .B1(n18056), .B2(n9754), .ZN(
        n17724) );
  OAI211_X1 U20942 ( .C1(n17733), .C2(n17726), .A(n17725), .B(n17724), .ZN(
        P3_U2817) );
  INV_X1 U20943 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17728) );
  INV_X1 U20944 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18771) );
  NOR2_X1 U20945 ( .A1(n15697), .A2(n18771), .ZN(n18077) );
  AOI221_X1 U20946 ( .B1(n17729), .B2(n17728), .C1(n17727), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n18077), .ZN(n17738) );
  OAI21_X1 U20947 ( .B1(n17732), .B2(n17766), .A(n17730), .ZN(n17731) );
  XNOR2_X1 U20948 ( .A(n17731), .B(n18080), .ZN(n18078) );
  INV_X1 U20949 ( .A(n9754), .ZN(n17749) );
  NOR2_X1 U20950 ( .A1(n17749), .A2(n17732), .ZN(n17735) );
  INV_X1 U20951 ( .A(n17733), .ZN(n17734) );
  MUX2_X1 U20952 ( .A(n17735), .B(n17734), .S(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n17736) );
  AOI21_X1 U20953 ( .B1(n17748), .B2(n18078), .A(n17736), .ZN(n17737) );
  OAI211_X1 U20954 ( .C1(n17740), .C2(n17739), .A(n17738), .B(n17737), .ZN(
        P3_U2818) );
  INV_X1 U20955 ( .A(n17877), .ZN(n17769) );
  NAND2_X1 U20956 ( .A1(n17782), .A2(n17799), .ZN(n17771) );
  NOR2_X1 U20957 ( .A1(n17770), .A2(n17771), .ZN(n17768) );
  NAND2_X1 U20958 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17768), .ZN(
        n17757) );
  OAI21_X1 U20959 ( .B1(n17769), .B2(n17741), .A(n17757), .ZN(n17742) );
  AOI22_X1 U20960 ( .A1(n17744), .A2(n17876), .B1(n17743), .B2(n17742), .ZN(
        n17753) );
  INV_X1 U20961 ( .A(n18091), .ZN(n17750) );
  AOI21_X1 U20962 ( .B1(n17750), .B2(n17746), .A(n17745), .ZN(n17747) );
  XNOR2_X1 U20963 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n17747), .ZN(
        n18082) );
  NOR2_X1 U20964 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18091), .ZN(
        n18081) );
  AOI22_X1 U20965 ( .A1(n17748), .A2(n18082), .B1(n18081), .B2(n9754), .ZN(
        n17752) );
  NOR2_X1 U20966 ( .A1(n17750), .A2(n17749), .ZN(n17762) );
  OAI22_X1 U20967 ( .A1(n18086), .A2(n17789), .B1(n17886), .B2(n18084), .ZN(
        n17776) );
  OAI21_X1 U20968 ( .B1(n17762), .B2(n17776), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17751) );
  NAND2_X1 U20969 ( .A1(n9760), .A2(P3_REIP_REG_11__SCAN_IN), .ZN(n18095) );
  NAND4_X1 U20970 ( .A1(n17753), .A2(n17752), .A3(n17751), .A4(n18095), .ZN(
        P3_U2819) );
  OAI221_X1 U20971 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17765), .C1(
        n15682), .C2(n17766), .A(n15681), .ZN(n17756) );
  NAND4_X1 U20972 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17754), .A3(
        n17781), .A4(n15682), .ZN(n17755) );
  OAI211_X1 U20973 ( .C1(n17766), .C2(n18091), .A(n17756), .B(n17755), .ZN(
        n18105) );
  INV_X1 U20974 ( .A(n17876), .ZN(n17866) );
  OAI211_X1 U20975 ( .C1(n17768), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n17877), .B(n17757), .ZN(n17758) );
  OAI21_X1 U20976 ( .B1(n17866), .B2(n17759), .A(n17758), .ZN(n17760) );
  AOI21_X1 U20977 ( .B1(n9760), .B2(P3_REIP_REG_10__SCAN_IN), .A(n17760), .ZN(
        n17764) );
  AOI22_X1 U20978 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17776), .B1(
        n17762), .B2(n17761), .ZN(n17763) );
  OAI211_X1 U20979 ( .C1(n17794), .C2(n18105), .A(n17764), .B(n17763), .ZN(
        P3_U2820) );
  NAND2_X1 U20980 ( .A1(n17766), .A2(n17765), .ZN(n17767) );
  XNOR2_X1 U20981 ( .A(n17767), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n18113) );
  AOI211_X1 U20982 ( .C1(n17771), .C2(n17770), .A(n17769), .B(n17768), .ZN(
        n17773) );
  NOR2_X1 U20983 ( .A1(n15697), .A2(n18765), .ZN(n17772) );
  AOI211_X1 U20984 ( .C1(n17774), .C2(n17876), .A(n17773), .B(n17772), .ZN(
        n17778) );
  AOI22_X1 U20985 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17776), .B1(
        n9754), .B2(n15682), .ZN(n17777) );
  OAI211_X1 U20986 ( .C1(n18113), .C2(n17794), .A(n17778), .B(n17777), .ZN(
        P3_U2821) );
  AOI21_X1 U20987 ( .B1(n17781), .B2(n17779), .A(n17780), .ZN(n18122) );
  NOR2_X1 U20988 ( .A1(n15697), .A2(n18764), .ZN(n18126) );
  AOI211_X1 U20989 ( .C1(n17785), .C2(n17783), .A(n17782), .B(n18260), .ZN(
        n17792) );
  AOI21_X1 U20990 ( .B1(n17843), .B2(n17784), .A(n17869), .ZN(n17797) );
  OAI22_X1 U20991 ( .A1(n17866), .A2(n17786), .B1(n17785), .B2(n17797), .ZN(
        n17791) );
  OAI21_X1 U20992 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17788), .A(
        n17787), .ZN(n18128) );
  OAI22_X1 U20993 ( .A1(n17779), .A2(n17789), .B1(n17886), .B2(n18128), .ZN(
        n17790) );
  NOR4_X1 U20994 ( .A1(n18126), .A2(n17792), .A3(n17791), .A4(n17790), .ZN(
        n17793) );
  OAI21_X1 U20995 ( .B1(n18122), .B2(n17794), .A(n17793), .ZN(P3_U2822) );
  OAI21_X1 U20996 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17796), .A(
        n17795), .ZN(n18137) );
  INV_X1 U20997 ( .A(n17797), .ZN(n17800) );
  NOR2_X1 U20998 ( .A1(n15697), .A2(n18761), .ZN(n18129) );
  AOI221_X1 U20999 ( .B1(n17800), .B2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C1(
        n17799), .C2(n17798), .A(n18129), .ZN(n17807) );
  AOI21_X1 U21000 ( .B1(n17803), .B2(n17802), .A(n17801), .ZN(n17804) );
  XOR2_X1 U21001 ( .A(n17804), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n18133) );
  AOI22_X1 U21002 ( .A1(n17874), .A2(n18133), .B1(n17805), .B2(n17876), .ZN(
        n17806) );
  OAI211_X1 U21003 ( .C1(n17885), .C2(n18137), .A(n17807), .B(n17806), .ZN(
        P3_U2823) );
  OAI21_X1 U21004 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17809), .A(
        n17808), .ZN(n18139) );
  NOR2_X1 U21005 ( .A1(n17814), .A2(n18260), .ZN(n17810) );
  AOI22_X1 U21006 ( .A1(n9760), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n17810), .B2(
        n17815), .ZN(n17819) );
  OAI21_X1 U21007 ( .B1(n17813), .B2(n17812), .A(n17811), .ZN(n18140) );
  OAI21_X1 U21008 ( .B1(n17814), .B2(n18260), .A(n17877), .ZN(n17827) );
  OAI22_X1 U21009 ( .A1(n17885), .A2(n18140), .B1(n17815), .B2(n17827), .ZN(
        n17816) );
  AOI21_X1 U21010 ( .B1(n17817), .B2(n17876), .A(n17816), .ZN(n17818) );
  OAI211_X1 U21011 ( .C1(n17886), .C2(n18139), .A(n17819), .B(n17818), .ZN(
        P3_U2824) );
  AOI21_X1 U21012 ( .B1(n17822), .B2(n17821), .A(n17820), .ZN(n18148) );
  AOI21_X1 U21013 ( .B1(n17824), .B2(n17823), .A(n9869), .ZN(n17825) );
  XOR2_X1 U21014 ( .A(n17825), .B(n18145), .Z(n18152) );
  INV_X1 U21015 ( .A(n18152), .ZN(n17831) );
  AOI21_X1 U21016 ( .B1(n17826), .B2(n17882), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17828) );
  OAI22_X1 U21017 ( .A1(n17866), .A2(n17829), .B1(n17828), .B2(n17827), .ZN(
        n17830) );
  AOI21_X1 U21018 ( .B1(n17832), .B2(n17831), .A(n17830), .ZN(n17833) );
  NAND2_X1 U21019 ( .A1(n9760), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n18147) );
  OAI211_X1 U21020 ( .C1(n18148), .C2(n17886), .A(n17833), .B(n18147), .ZN(
        P3_U2825) );
  OAI21_X1 U21021 ( .B1(n17836), .B2(n17835), .A(n17834), .ZN(n18161) );
  INV_X1 U21022 ( .A(n17837), .ZN(n17838) );
  AOI22_X1 U21023 ( .A1(n9760), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18607), .B2(
        n17838), .ZN(n17848) );
  OAI21_X1 U21024 ( .B1(n17841), .B2(n17840), .A(n17839), .ZN(n18155) );
  AOI21_X1 U21025 ( .B1(n17843), .B2(n17842), .A(n17869), .ZN(n17854) );
  OAI22_X1 U21026 ( .A1(n17885), .A2(n18155), .B1(n17844), .B2(n17854), .ZN(
        n17845) );
  AOI21_X1 U21027 ( .B1(n17846), .B2(n17876), .A(n17845), .ZN(n17847) );
  OAI211_X1 U21028 ( .C1(n17886), .C2(n18161), .A(n17848), .B(n17847), .ZN(
        P3_U2826) );
  OAI21_X1 U21029 ( .B1(n17851), .B2(n17850), .A(n17849), .ZN(n18164) );
  AOI21_X1 U21030 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17882), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17855) );
  OAI21_X1 U21031 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n17853), .A(
        n17852), .ZN(n18166) );
  OAI22_X1 U21032 ( .A1(n17855), .A2(n17854), .B1(n17885), .B2(n18166), .ZN(
        n17856) );
  AOI21_X1 U21033 ( .B1(n17857), .B2(n17876), .A(n17856), .ZN(n17858) );
  NAND2_X1 U21034 ( .A1(n9760), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n18169) );
  OAI211_X1 U21035 ( .C1(n17886), .C2(n18164), .A(n17858), .B(n18169), .ZN(
        P3_U2827) );
  OAI21_X1 U21036 ( .B1(n17861), .B2(n17860), .A(n17859), .ZN(n18182) );
  OAI21_X1 U21037 ( .B1(n17864), .B2(n17863), .A(n17862), .ZN(n18188) );
  OAI22_X1 U21038 ( .A1(n17866), .A2(n17865), .B1(n17885), .B2(n18188), .ZN(
        n17867) );
  AOI221_X1 U21039 ( .B1(n17869), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C1(
        n18607), .C2(n17868), .A(n17867), .ZN(n17870) );
  NAND2_X1 U21040 ( .A1(n9760), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18186) );
  OAI211_X1 U21041 ( .C1(n17886), .C2(n18182), .A(n17870), .B(n18186), .ZN(
        P3_U2828) );
  OAI21_X1 U21042 ( .B1(n17880), .B2(n17872), .A(n17871), .ZN(n18198) );
  XNOR2_X1 U21043 ( .A(n17873), .B(n17872), .ZN(n18195) );
  AOI22_X1 U21044 ( .A1(n9760), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n17874), .B2(
        n18195), .ZN(n17879) );
  AOI22_X1 U21045 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17877), .B1(
        n17876), .B2(n17875), .ZN(n17878) );
  OAI211_X1 U21046 ( .C1(n17885), .C2(n18198), .A(n17879), .B(n17878), .ZN(
        P3_U2829) );
  INV_X1 U21047 ( .A(n18201), .ZN(n18203) );
  NAND3_X1 U21048 ( .A1(n18834), .A2(n17882), .A3(n17881), .ZN(n17883) );
  AOI22_X1 U21049 ( .A1(n9760), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17883), .ZN(n17884) );
  OAI221_X1 U21050 ( .B1(n18201), .B2(n17886), .C1(n18203), .C2(n17885), .A(
        n17884), .ZN(P3_U2830) );
  AOI22_X1 U21051 ( .A1(n9760), .A2(P3_REIP_REG_27__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18185), .ZN(n17899) );
  NOR3_X1 U21052 ( .A1(n17938), .A2(n17887), .A3(n17937), .ZN(n17897) );
  INV_X1 U21053 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17896) );
  INV_X1 U21054 ( .A(n18173), .ZN(n17889) );
  OAI21_X1 U21055 ( .B1(n17888), .B2(n18173), .A(n17952), .ZN(n17924) );
  AOI21_X1 U21056 ( .B1(n17909), .B2(n17889), .A(n17924), .ZN(n17908) );
  OAI211_X1 U21057 ( .C1(n17891), .C2(n18173), .A(n17908), .B(n17890), .ZN(
        n17892) );
  AOI21_X1 U21058 ( .B1(n18060), .B2(n17893), .A(n17892), .ZN(n17894) );
  OAI21_X1 U21059 ( .B1(n17895), .B2(n18664), .A(n17894), .ZN(n17902) );
  OAI221_X1 U21060 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17897), 
        .C1(n17896), .C2(n17902), .A(n18184), .ZN(n17898) );
  OAI211_X1 U21061 ( .C1(n17900), .C2(n18121), .A(n17899), .B(n17898), .ZN(
        P3_U2835) );
  AOI22_X1 U21062 ( .A1(n9760), .A2(P3_REIP_REG_26__SCAN_IN), .B1(n17933), 
        .B2(n17901), .ZN(n17904) );
  OAI211_X1 U21063 ( .C1(n18205), .C2(n17902), .A(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n15697), .ZN(n17903) );
  OAI211_X1 U21064 ( .C1(n17905), .C2(n18121), .A(n17904), .B(n17903), .ZN(
        P3_U2836) );
  NOR2_X1 U21065 ( .A1(n17907), .A2(n17906), .ZN(n17927) );
  OAI221_X1 U21066 ( .B1(n18665), .B2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), 
        .C1(n18665), .C2(n17927), .A(n17908), .ZN(n17912) );
  NOR2_X1 U21067 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17909), .ZN(
        n17910) );
  AOI22_X1 U21068 ( .A1(n17912), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n17911), .B2(n17910), .ZN(n17914) );
  OAI21_X1 U21069 ( .B1(n18205), .B2(n17914), .A(n17913), .ZN(n17918) );
  OAI22_X1 U21070 ( .A1(n18121), .A2(n17916), .B1(n18120), .B2(n17915), .ZN(
        n17917) );
  AOI211_X1 U21071 ( .C1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n18185), .A(
        n17918), .B(n17917), .ZN(n17919) );
  OAI21_X1 U21072 ( .B1(n18165), .B2(n17920), .A(n17919), .ZN(P3_U2837) );
  OAI22_X1 U21073 ( .A1(n17922), .A2(n18085), .B1(n17921), .B2(n18664), .ZN(
        n17923) );
  NOR3_X1 U21074 ( .A1(n18185), .A2(n17924), .A3(n17923), .ZN(n17929) );
  NOR2_X1 U21075 ( .A1(n18690), .A2(n17925), .ZN(n17926) );
  AOI221_X1 U21076 ( .B1(n17927), .B2(n17929), .C1(n17926), .C2(n17929), .A(
        n9760), .ZN(n17939) );
  AOI21_X1 U21077 ( .B1(n17930), .B2(n17929), .A(n17928), .ZN(n17931) );
  AOI22_X1 U21078 ( .A1(n17933), .A2(n17932), .B1(n17939), .B2(n17931), .ZN(
        n17935) );
  NAND2_X1 U21079 ( .A1(n9760), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n17934) );
  OAI211_X1 U21080 ( .C1(n17936), .C2(n18121), .A(n17935), .B(n17934), .ZN(
        P3_U2838) );
  NOR2_X1 U21081 ( .A1(n17938), .A2(n17937), .ZN(n17940) );
  OAI221_X1 U21082 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17940), 
        .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n18190), .A(n17939), .ZN(
        n17941) );
  OAI211_X1 U21083 ( .C1(n17943), .C2(n18121), .A(n17942), .B(n17941), .ZN(
        P3_U2839) );
  AOI21_X1 U21084 ( .B1(n18184), .B2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n17944), .ZN(n17960) );
  INV_X1 U21085 ( .A(n17945), .ZN(n18031) );
  OAI22_X1 U21086 ( .A1(n18025), .A2(n18085), .B1(n18031), .B2(n18664), .ZN(
        n17962) );
  AOI21_X1 U21087 ( .B1(n17946), .B2(n17972), .A(n18694), .ZN(n17949) );
  AOI21_X1 U21088 ( .B1(n17948), .B2(n17947), .A(n18665), .ZN(n17999) );
  AOI211_X1 U21089 ( .C1(n18690), .C2(n18001), .A(n17949), .B(n17999), .ZN(
        n17965) );
  OAI211_X1 U21090 ( .C1(n17967), .C2(n18665), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n17965), .ZN(n17954) );
  NAND2_X1 U21091 ( .A1(n18085), .A2(n18664), .ZN(n18090) );
  AOI22_X1 U21092 ( .A1(n17951), .A2(n18206), .B1(n17950), .B2(n18090), .ZN(
        n17966) );
  OAI211_X1 U21093 ( .C1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n18067), .A(
        n17966), .B(n17952), .ZN(n17953) );
  NOR3_X1 U21094 ( .A1(n17962), .A2(n17954), .A3(n17953), .ZN(n17959) );
  INV_X1 U21095 ( .A(n17955), .ZN(n17956) );
  AOI22_X1 U21096 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18185), .B1(
        n18083), .B2(n17956), .ZN(n17958) );
  NAND2_X1 U21097 ( .A1(n9760), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17957) );
  OAI211_X1 U21098 ( .C1(n17960), .C2(n17959), .A(n17958), .B(n17957), .ZN(
        P3_U2840) );
  AOI22_X1 U21099 ( .A1(n9760), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n18083), 
        .B2(n17961), .ZN(n17970) );
  NOR2_X1 U21100 ( .A1(n18205), .A2(n17962), .ZN(n18014) );
  OAI21_X1 U21101 ( .B1(n18016), .B2(n17963), .A(n18692), .ZN(n17964) );
  NAND3_X1 U21102 ( .A1(n18014), .A2(n17965), .A3(n17964), .ZN(n17974) );
  NOR2_X1 U21103 ( .A1(n18690), .A2(n18692), .ZN(n18189) );
  OAI21_X1 U21104 ( .B1(n17967), .B2(n18189), .A(n17966), .ZN(n17968) );
  OAI211_X1 U21105 ( .C1(n17974), .C2(n17968), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n15697), .ZN(n17969) );
  OAI211_X1 U21106 ( .C1(n17971), .C2(n17988), .A(n17970), .B(n17969), .ZN(
        P3_U2841) );
  INV_X1 U21107 ( .A(n17972), .ZN(n17973) );
  OAI221_X1 U21108 ( .B1(n17974), .B2(n18090), .C1(n17974), .C2(n17973), .A(
        n15697), .ZN(n17986) );
  INV_X1 U21109 ( .A(n18189), .ZN(n17975) );
  NAND3_X1 U21110 ( .A1(n17975), .A2(n17987), .A3(P3_STATE2_REG_2__SCAN_IN), 
        .ZN(n17976) );
  NAND2_X1 U21111 ( .A1(n17986), .A2(n17976), .ZN(n17978) );
  AOI22_X1 U21112 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17978), .B1(
        n18083), .B2(n17977), .ZN(n17980) );
  OAI211_X1 U21113 ( .C1(n17988), .C2(n17981), .A(n17980), .B(n17979), .ZN(
        P3_U2842) );
  INV_X1 U21114 ( .A(n17982), .ZN(n17983) );
  AOI21_X1 U21115 ( .B1(n18083), .B2(n17984), .A(n17983), .ZN(n17985) );
  OAI221_X1 U21116 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17988), 
        .C1(n17987), .C2(n17986), .A(n17985), .ZN(P3_U2843) );
  INV_X1 U21117 ( .A(n17989), .ZN(n18174) );
  INV_X1 U21118 ( .A(n17990), .ZN(n18153) );
  AOI22_X1 U21119 ( .A1(n18690), .A2(n18174), .B1(n18153), .B2(n18179), .ZN(
        n18163) );
  NOR2_X1 U21120 ( .A1(n18163), .A2(n17991), .ZN(n18130) );
  NAND2_X1 U21121 ( .A1(n17992), .A2(n18130), .ZN(n18044) );
  OAI222_X1 U21122 ( .A1(n18044), .A2(n18205), .B1(n18165), .B2(n17994), .C1(
        n17993), .C2(n18120), .ZN(n18106) );
  NAND2_X1 U21123 ( .A1(n17995), .A2(n18106), .ZN(n18024) );
  NOR2_X1 U21124 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18680), .ZN(
        n18177) );
  NOR3_X1 U21125 ( .A1(n18177), .A2(n17996), .A3(n18023), .ZN(n17997) );
  OAI21_X1 U21126 ( .B1(n18173), .B2(n17997), .A(n18014), .ZN(n17998) );
  AOI211_X1 U21127 ( .C1(n18000), .C2(n18090), .A(n17999), .B(n17998), .ZN(
        n18008) );
  AOI221_X1 U21128 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18008), 
        .C1(n18173), .C2(n18008), .A(n18001), .ZN(n18002) );
  AOI22_X1 U21129 ( .A1(n18003), .A2(n18083), .B1(n18002), .B2(n15697), .ZN(
        n18005) );
  NAND2_X1 U21130 ( .A1(n9760), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18004) );
  OAI211_X1 U21131 ( .C1(n18006), .C2(n18024), .A(n18005), .B(n18004), .ZN(
        P3_U2844) );
  NOR3_X1 U21132 ( .A1(n9760), .A2(n18008), .A3(n18007), .ZN(n18009) );
  AOI21_X1 U21133 ( .B1(n18083), .B2(n18010), .A(n18009), .ZN(n18012) );
  OAI211_X1 U21134 ( .C1(n18024), .C2(n18013), .A(n18012), .B(n18011), .ZN(
        P3_U2845) );
  INV_X1 U21135 ( .A(n18014), .ZN(n18019) );
  AND2_X1 U21136 ( .A1(n18690), .A2(n18015), .ZN(n18089) );
  AOI21_X1 U21137 ( .B1(n18206), .B2(n18097), .A(n18089), .ZN(n18108) );
  OAI21_X1 U21138 ( .B1(n18692), .B2(n15683), .A(n18016), .ZN(n18017) );
  OAI211_X1 U21139 ( .C1(n18018), .C2(n18067), .A(n18108), .B(n18017), .ZN(
        n18027) );
  OAI221_X1 U21140 ( .B1(n18019), .B2(n18118), .C1(n18019), .C2(n18027), .A(
        n15697), .ZN(n18022) );
  AOI22_X1 U21141 ( .A1(n9760), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n18083), 
        .B2(n18020), .ZN(n18021) );
  OAI221_X1 U21142 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18024), 
        .C1(n18023), .C2(n18022), .A(n18021), .ZN(P3_U2846) );
  NOR2_X1 U21143 ( .A1(n18025), .A2(n18085), .ZN(n18029) );
  OAI21_X1 U21144 ( .B1(n18039), .B2(n18044), .A(n15683), .ZN(n18026) );
  AOI22_X1 U21145 ( .A1(n18029), .A2(n18028), .B1(n18027), .B2(n18026), .ZN(
        n18036) );
  NOR3_X1 U21146 ( .A1(n18031), .A2(n18030), .A3(n18165), .ZN(n18033) );
  OAI22_X1 U21147 ( .A1(n15697), .A2(n18777), .B1(n15683), .B2(n18190), .ZN(
        n18032) );
  AOI211_X1 U21148 ( .C1(n18034), .C2(n18083), .A(n18033), .B(n18032), .ZN(
        n18035) );
  OAI21_X1 U21149 ( .B1(n18036), .B2(n18205), .A(n18035), .ZN(P3_U2847) );
  NOR2_X1 U21150 ( .A1(n18851), .A2(n18097), .ZN(n18109) );
  AOI21_X1 U21151 ( .B1(n18037), .B2(n18109), .A(n18680), .ZN(n18066) );
  AOI211_X1 U21152 ( .C1(n18690), .C2(n18038), .A(n18089), .B(n18066), .ZN(
        n18041) );
  OAI22_X1 U21153 ( .A1(n18047), .A2(n18206), .B1(n18039), .B2(n18097), .ZN(
        n18040) );
  OAI211_X1 U21154 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n18189), .A(
        n18041), .B(n18040), .ZN(n18042) );
  NAND2_X1 U21155 ( .A1(n18184), .A2(n18042), .ZN(n18046) );
  OR2_X1 U21156 ( .A1(n18044), .A2(n18043), .ZN(n18045) );
  AOI222_X1 U21157 ( .A1(n18047), .A2(n18046), .B1(n18047), .B2(n18045), .C1(
        n18046), .C2(n18190), .ZN(n18048) );
  AOI211_X1 U21158 ( .C1(n18051), .C2(n18050), .A(n18049), .B(n18048), .ZN(
        n18054) );
  NAND2_X1 U21159 ( .A1(n18204), .A2(n18052), .ZN(n18053) );
  OAI211_X1 U21160 ( .C1(n18055), .C2(n18121), .A(n18054), .B(n18053), .ZN(
        P3_U2848) );
  AOI22_X1 U21161 ( .A1(n18083), .A2(n18057), .B1(n18056), .B2(n18106), .ZN(
        n18071) );
  AOI21_X1 U21162 ( .B1(n18058), .B2(n18206), .A(n18080), .ZN(n18075) );
  OAI21_X1 U21163 ( .B1(n18091), .B2(n18097), .A(n18206), .ZN(n18059) );
  OAI21_X1 U21164 ( .B1(n18072), .B2(n18665), .A(n18059), .ZN(n18093) );
  AOI22_X1 U21165 ( .A1(n18063), .A2(n18062), .B1(n18061), .B2(n18060), .ZN(
        n18064) );
  INV_X1 U21166 ( .A(n18064), .ZN(n18065) );
  NOR4_X1 U21167 ( .A1(n18089), .A2(n18066), .A3(n18093), .A4(n18065), .ZN(
        n18074) );
  OAI211_X1 U21168 ( .C1(n18067), .C2(n18075), .A(n18184), .B(n18074), .ZN(
        n18068) );
  NAND3_X1 U21169 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15697), .A3(
        n18068), .ZN(n18069) );
  NAND3_X1 U21170 ( .A1(n18071), .A2(n18070), .A3(n18069), .ZN(P3_U2849) );
  AOI22_X1 U21171 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18184), .B1(
        n18072), .B2(n18106), .ZN(n18073) );
  AOI21_X1 U21172 ( .B1(n18075), .B2(n18074), .A(n18073), .ZN(n18076) );
  AOI211_X1 U21173 ( .C1(n18083), .C2(n18078), .A(n18077), .B(n18076), .ZN(
        n18079) );
  OAI21_X1 U21174 ( .B1(n18080), .B2(n18190), .A(n18079), .ZN(P3_U2850) );
  AOI22_X1 U21175 ( .A1(n18083), .A2(n18082), .B1(n18081), .B2(n18106), .ZN(
        n18096) );
  OAI22_X1 U21176 ( .A1(n18086), .A2(n18085), .B1(n18664), .B2(n18084), .ZN(
        n18087) );
  NOR2_X1 U21177 ( .A1(n18205), .A2(n18087), .ZN(n18107) );
  OAI221_X1 U21178 ( .B1(n18680), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(
        n18680), .C2(n18109), .A(n18107), .ZN(n18088) );
  AOI211_X1 U21179 ( .C1(n18091), .C2(n18090), .A(n18089), .B(n18088), .ZN(
        n18100) );
  OAI21_X1 U21180 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n18680), .A(
        n18100), .ZN(n18092) );
  OAI211_X1 U21181 ( .C1(n18093), .C2(n18092), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n15697), .ZN(n18094) );
  NAND3_X1 U21182 ( .A1(n18096), .A2(n18095), .A3(n18094), .ZN(P3_U2851) );
  NOR2_X1 U21183 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n15682), .ZN(
        n18102) );
  AOI22_X1 U21184 ( .A1(n15682), .A2(n18098), .B1(n18206), .B2(n18097), .ZN(
        n18099) );
  AOI211_X1 U21185 ( .C1(n18100), .C2(n18099), .A(n9760), .B(n15681), .ZN(
        n18101) );
  AOI21_X1 U21186 ( .B1(n18102), .B2(n18106), .A(n18101), .ZN(n18104) );
  NAND2_X1 U21187 ( .A1(n9760), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n18103) );
  OAI211_X1 U21188 ( .C1(n18105), .C2(n18121), .A(n18104), .B(n18103), .ZN(
        P3_U2852) );
  AOI22_X1 U21189 ( .A1(n9760), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n15682), .B2(
        n18106), .ZN(n18112) );
  OAI211_X1 U21190 ( .C1(n18109), .C2(n18680), .A(n18108), .B(n18107), .ZN(
        n18110) );
  NAND3_X1 U21191 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15697), .A3(
        n18110), .ZN(n18111) );
  OAI211_X1 U21192 ( .C1(n18113), .C2(n18121), .A(n18112), .B(n18111), .ZN(
        P3_U2853) );
  OAI22_X1 U21193 ( .A1(n18115), .A2(n18173), .B1(n18114), .B2(n18665), .ZN(
        n18116) );
  NOR2_X1 U21194 ( .A1(n18177), .A2(n18116), .ZN(n18138) );
  INV_X1 U21195 ( .A(n18138), .ZN(n18117) );
  AOI21_X1 U21196 ( .B1(n18119), .B2(n18118), .A(n18117), .ZN(n18132) );
  AOI221_X1 U21197 ( .B1(n18132), .B2(n18190), .C1(n18191), .C2(n18190), .A(
        n10100), .ZN(n18125) );
  INV_X1 U21198 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18171) );
  NOR3_X1 U21199 ( .A1(n18163), .A2(n18205), .A3(n18171), .ZN(n18159) );
  NAND3_X1 U21200 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n18159), .ZN(n18144) );
  NOR3_X1 U21201 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18119), .A3(
        n18144), .ZN(n18124) );
  OAI22_X1 U21202 ( .A1(n18122), .A2(n18121), .B1(n17779), .B2(n18120), .ZN(
        n18123) );
  NOR4_X1 U21203 ( .A1(n18126), .A2(n18125), .A3(n18124), .A4(n18123), .ZN(
        n18127) );
  OAI21_X1 U21204 ( .B1(n18165), .B2(n18128), .A(n18127), .ZN(P3_U2854) );
  AOI21_X1 U21205 ( .B1(n18185), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18129), .ZN(n18136) );
  AOI21_X1 U21206 ( .B1(n18130), .B2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18131) );
  NOR2_X1 U21207 ( .A1(n18132), .A2(n18131), .ZN(n18134) );
  AOI22_X1 U21208 ( .A1(n18184), .A2(n18134), .B1(n18204), .B2(n18133), .ZN(
        n18135) );
  OAI211_X1 U21209 ( .C1(n18199), .C2(n18137), .A(n18136), .B(n18135), .ZN(
        P3_U2855) );
  OAI21_X1 U21210 ( .B1(n18138), .B2(n18205), .A(n18190), .ZN(n18150) );
  NOR2_X1 U21211 ( .A1(n15697), .A2(n18759), .ZN(n18142) );
  OAI22_X1 U21212 ( .A1(n18199), .A2(n18140), .B1(n18165), .B2(n18139), .ZN(
        n18141) );
  AOI211_X1 U21213 ( .C1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n18150), .A(
        n18142), .B(n18141), .ZN(n18143) );
  OAI21_X1 U21214 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18144), .A(
        n18143), .ZN(P3_U2856) );
  NAND3_X1 U21215 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18159), .A3(
        n18145), .ZN(n18146) );
  OAI211_X1 U21216 ( .C1(n18148), .C2(n18165), .A(n18147), .B(n18146), .ZN(
        n18149) );
  AOI21_X1 U21217 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n18150), .A(
        n18149), .ZN(n18151) );
  OAI21_X1 U21218 ( .B1(n18199), .B2(n18152), .A(n18151), .ZN(P3_U2857) );
  OAI22_X1 U21219 ( .A1(n18153), .A2(n18173), .B1(n18665), .B2(n18174), .ZN(
        n18154) );
  NOR3_X1 U21220 ( .A1(n18177), .A2(n18171), .A3(n18154), .ZN(n18162) );
  OAI21_X1 U21221 ( .B1(n18162), .B2(n18191), .A(n18190), .ZN(n18157) );
  OAI22_X1 U21222 ( .A1(n15697), .A2(n18755), .B1(n18199), .B2(n18155), .ZN(
        n18156) );
  AOI221_X1 U21223 ( .B1(n18159), .B2(n18158), .C1(n18157), .C2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n18156), .ZN(n18160) );
  OAI21_X1 U21224 ( .B1(n18165), .B2(n18161), .A(n18160), .ZN(P3_U2858) );
  AOI211_X1 U21225 ( .C1(n18163), .C2(n18171), .A(n18162), .B(n18205), .ZN(
        n18168) );
  OAI22_X1 U21226 ( .A1(n18199), .A2(n18166), .B1(n18165), .B2(n18164), .ZN(
        n18167) );
  NOR2_X1 U21227 ( .A1(n18168), .A2(n18167), .ZN(n18170) );
  OAI211_X1 U21228 ( .C1(n18190), .C2(n18171), .A(n18170), .B(n18169), .ZN(
        P3_U2859) );
  NAND2_X1 U21229 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18172) );
  OAI22_X1 U21230 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18173), .B1(
        n18172), .B2(n18665), .ZN(n18176) );
  NOR2_X1 U21231 ( .A1(n18665), .A2(n18174), .ZN(n18175) );
  AOI221_X1 U21232 ( .B1(n18177), .B2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .C1(
        n18176), .C2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(n18175), .ZN(
        n18181) );
  NAND3_X1 U21233 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18179), .A3(
        n18178), .ZN(n18180) );
  OAI211_X1 U21234 ( .C1(n18182), .C2(n18664), .A(n18181), .B(n18180), .ZN(
        n18183) );
  AOI22_X1 U21235 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18185), .B1(
        n18184), .B2(n18183), .ZN(n18187) );
  OAI211_X1 U21236 ( .C1(n18188), .C2(n18199), .A(n18187), .B(n18186), .ZN(
        P3_U2860) );
  OR3_X1 U21237 ( .A1(n18205), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n18189), .ZN(n18208) );
  AOI21_X1 U21238 ( .B1(n18190), .B2(n18208), .A(n15608), .ZN(n18194) );
  NOR3_X1 U21239 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18192), .A3(
        n18191), .ZN(n18193) );
  AOI211_X1 U21240 ( .C1(n18204), .C2(n18195), .A(n18194), .B(n18193), .ZN(
        n18197) );
  NAND2_X1 U21241 ( .A1(n9760), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18196) );
  OAI211_X1 U21242 ( .C1(n18198), .C2(n18199), .A(n18197), .B(n18196), .ZN(
        P3_U2861) );
  INV_X1 U21243 ( .A(n18199), .ZN(n18202) );
  INV_X1 U21244 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n20867) );
  NOR2_X1 U21245 ( .A1(n15697), .A2(n20867), .ZN(n18200) );
  AOI221_X1 U21246 ( .B1(n18204), .B2(n18203), .C1(n18202), .C2(n18201), .A(
        n18200), .ZN(n18209) );
  OAI211_X1 U21247 ( .C1(n18206), .C2(n18205), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n15697), .ZN(n18207) );
  NAND3_X1 U21248 ( .A1(n18209), .A2(n18208), .A3(n18207), .ZN(P3_U2862) );
  AOI211_X1 U21249 ( .C1(n18211), .C2(n18210), .A(n18888), .B(n18834), .ZN(
        n18719) );
  OAI21_X1 U21250 ( .B1(n18719), .B2(n18265), .A(n18216), .ZN(n18212) );
  OAI221_X1 U21251 ( .B1(n18217), .B2(n18867), .C1(n18217), .C2(n18216), .A(
        n18212), .ZN(P3_U2863) );
  INV_X1 U21252 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18707) );
  NOR2_X1 U21253 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18704), .ZN(
        n18400) );
  INV_X1 U21254 ( .A(n18470), .ZN(n18564) );
  NOR2_X1 U21255 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18707), .ZN(
        n18493) );
  INV_X1 U21256 ( .A(n18493), .ZN(n18491) );
  NOR2_X1 U21257 ( .A1(n18564), .A2(n18491), .ZN(n18518) );
  NOR2_X1 U21258 ( .A1(n18400), .A2(n18518), .ZN(n18214) );
  OAI22_X1 U21259 ( .A1(n18215), .A2(n18707), .B1(n18214), .B2(n18213), .ZN(
        P3_U2866) );
  NOR2_X1 U21260 ( .A1(n18708), .A2(n18216), .ZN(P3_U2867) );
  NOR2_X1 U21261 ( .A1(n18699), .A2(n18217), .ZN(n18308) );
  NOR2_X1 U21262 ( .A1(n18704), .A2(n18707), .ZN(n18222) );
  NAND2_X1 U21263 ( .A1(n18308), .A2(n18222), .ZN(n18658) );
  NAND2_X1 U21264 ( .A1(n18699), .A2(n18217), .ZN(n18700) );
  NAND2_X1 U21265 ( .A1(n18704), .A2(n18707), .ZN(n18352) );
  NOR2_X1 U21266 ( .A1(n18700), .A2(n18352), .ZN(n18326) );
  CLKBUF_X1 U21267 ( .A(n18326), .Z(n18302) );
  NOR2_X1 U21268 ( .A1(n18303), .A2(n18302), .ZN(n18285) );
  OAI21_X1 U21269 ( .B1(n18824), .B2(n18217), .A(n18331), .ZN(n18563) );
  NOR2_X1 U21270 ( .A1(n18699), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18467) );
  NOR2_X1 U21271 ( .A1(n18217), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18444) );
  OR2_X1 U21272 ( .A1(n18467), .A2(n18444), .ZN(n18517) );
  NAND2_X1 U21273 ( .A1(n18222), .A2(n18517), .ZN(n18566) );
  OAI22_X1 U21274 ( .A1(n18285), .A2(n18563), .B1(n18260), .B2(n18566), .ZN(
        n18263) );
  NOR2_X2 U21275 ( .A1(n18515), .A2(n18218), .ZN(n18602) );
  NOR2_X1 U21276 ( .A1(n9746), .A2(n18285), .ZN(n18258) );
  AOI22_X1 U21277 ( .A1(n18608), .A2(n18597), .B1(n18602), .B2(n18258), .ZN(
        n18225) );
  NAND2_X1 U21278 ( .A1(n18220), .A2(n18219), .ZN(n18259) );
  NOR2_X1 U21279 ( .A1(n18221), .A2(n18259), .ZN(n18567) );
  NAND2_X1 U21280 ( .A1(n18222), .A2(n18699), .ZN(n18541) );
  INV_X1 U21281 ( .A(n18541), .ZN(n18606) );
  NAND2_X1 U21282 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18606), .ZN(
        n18562) );
  INV_X1 U21283 ( .A(n18562), .ZN(n18653) );
  NOR2_X2 U21284 ( .A1(n18223), .A2(n18260), .ZN(n18603) );
  AOI22_X1 U21285 ( .A1(n18302), .A2(n18567), .B1(n18653), .B2(n18603), .ZN(
        n18224) );
  OAI211_X1 U21286 ( .C1(n18226), .C2(n18263), .A(n18225), .B(n18224), .ZN(
        P3_U2868) );
  NOR2_X2 U21287 ( .A1(n18260), .A2(n13890), .ZN(n18614) );
  AND2_X1 U21288 ( .A1(n18331), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18612) );
  AOI22_X1 U21289 ( .A1(n18597), .A2(n18614), .B1(n18258), .B2(n18612), .ZN(
        n18229) );
  NOR2_X1 U21290 ( .A1(n18227), .A2(n18259), .ZN(n18570) );
  AND2_X1 U21291 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18607), .ZN(n18613) );
  AOI22_X1 U21292 ( .A1(n18302), .A2(n18570), .B1(n18653), .B2(n18613), .ZN(
        n18228) );
  OAI211_X1 U21293 ( .C1(n18230), .C2(n18263), .A(n18229), .B(n18228), .ZN(
        P3_U2869) );
  AND2_X1 U21294 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18607), .ZN(n18620) );
  NOR2_X2 U21295 ( .A1(n18515), .A2(n18231), .ZN(n18618) );
  AOI22_X1 U21296 ( .A1(n18653), .A2(n18620), .B1(n18258), .B2(n18618), .ZN(
        n18235) );
  NOR2_X1 U21297 ( .A1(n18232), .A2(n18259), .ZN(n18574) );
  NOR2_X2 U21298 ( .A1(n18260), .A2(n18233), .ZN(n18619) );
  AOI22_X1 U21299 ( .A1(n18302), .A2(n18574), .B1(n18597), .B2(n18619), .ZN(
        n18234) );
  OAI211_X1 U21300 ( .C1(n18236), .C2(n18263), .A(n18235), .B(n18234), .ZN(
        P3_U2870) );
  NOR2_X2 U21301 ( .A1(n19253), .A2(n18260), .ZN(n18625) );
  NOR2_X2 U21302 ( .A1(n18515), .A2(n18237), .ZN(n18624) );
  AOI22_X1 U21303 ( .A1(n18653), .A2(n18625), .B1(n18258), .B2(n18624), .ZN(
        n18240) );
  NOR2_X1 U21304 ( .A1(n18238), .A2(n18259), .ZN(n18578) );
  AOI22_X1 U21305 ( .A1(n18302), .A2(n18578), .B1(n18597), .B2(n18626), .ZN(
        n18239) );
  OAI211_X1 U21306 ( .C1(n20907), .C2(n18263), .A(n18240), .B(n18239), .ZN(
        P3_U2871) );
  NOR2_X2 U21307 ( .A1(n19257), .A2(n18260), .ZN(n18632) );
  NOR2_X2 U21308 ( .A1(n18515), .A2(n18241), .ZN(n18630) );
  AOI22_X1 U21309 ( .A1(n18653), .A2(n18632), .B1(n18258), .B2(n18630), .ZN(
        n18244) );
  NOR2_X1 U21310 ( .A1(n18242), .A2(n18259), .ZN(n18582) );
  AND2_X1 U21311 ( .A1(n18607), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18631) );
  AOI22_X1 U21312 ( .A1(n18302), .A2(n18582), .B1(n18597), .B2(n18631), .ZN(
        n18243) );
  OAI211_X1 U21313 ( .C1(n18245), .C2(n18263), .A(n18244), .B(n18243), .ZN(
        P3_U2872) );
  NOR2_X2 U21314 ( .A1(n21050), .A2(n18260), .ZN(n18638) );
  NOR2_X2 U21315 ( .A1(n18515), .A2(n18246), .ZN(n18636) );
  AOI22_X1 U21316 ( .A1(n18653), .A2(n18638), .B1(n18258), .B2(n18636), .ZN(
        n18249) );
  NOR2_X1 U21317 ( .A1(n18247), .A2(n18259), .ZN(n18586) );
  NOR2_X2 U21318 ( .A1(n18260), .A2(n14963), .ZN(n18637) );
  AOI22_X1 U21319 ( .A1(n18302), .A2(n18586), .B1(n18597), .B2(n18637), .ZN(
        n18248) );
  OAI211_X1 U21320 ( .C1(n18250), .C2(n18263), .A(n18249), .B(n18248), .ZN(
        P3_U2873) );
  NOR2_X2 U21321 ( .A1(n18251), .A2(n18260), .ZN(n18644) );
  NOR2_X2 U21322 ( .A1(n18515), .A2(n18252), .ZN(n18642) );
  AOI22_X1 U21323 ( .A1(n18653), .A2(n18644), .B1(n18258), .B2(n18642), .ZN(
        n18255) );
  NOR2_X1 U21324 ( .A1(n18253), .A2(n18259), .ZN(n18590) );
  NOR2_X2 U21325 ( .A1(n18260), .A2(n19269), .ZN(n18643) );
  AOI22_X1 U21326 ( .A1(n18302), .A2(n18590), .B1(n18597), .B2(n18643), .ZN(
        n18254) );
  OAI211_X1 U21327 ( .C1(n18256), .C2(n18263), .A(n18255), .B(n18254), .ZN(
        P3_U2874) );
  AND2_X1 U21328 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18607), .ZN(n18652) );
  NOR2_X2 U21329 ( .A1(n18257), .A2(n18515), .ZN(n18649) );
  AOI22_X1 U21330 ( .A1(n18597), .A2(n18652), .B1(n18258), .B2(n18649), .ZN(
        n18262) );
  NOR2_X1 U21331 ( .A1(n9796), .A2(n18259), .ZN(n18596) );
  NOR2_X2 U21332 ( .A1(n18260), .A2(n21051), .ZN(n18651) );
  AOI22_X1 U21333 ( .A1(n18302), .A2(n18596), .B1(n18653), .B2(n18651), .ZN(
        n18261) );
  OAI211_X1 U21334 ( .C1(n18264), .C2(n18263), .A(n18262), .B(n18261), .ZN(
        P3_U2875) );
  INV_X1 U21335 ( .A(n18352), .ZN(n18310) );
  NAND2_X1 U21336 ( .A1(n18310), .A2(n18444), .ZN(n18284) );
  AOI22_X1 U21337 ( .A1(n18303), .A2(n18608), .B1(n18602), .B2(n18280), .ZN(
        n18267) );
  NOR2_X1 U21338 ( .A1(n18707), .A2(n18445), .ZN(n18604) );
  NOR2_X1 U21339 ( .A1(n18515), .A2(n18265), .ZN(n18605) );
  INV_X1 U21340 ( .A(n18605), .ZN(n18309) );
  NOR2_X1 U21341 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18309), .ZN(
        n18353) );
  AOI22_X1 U21342 ( .A1(n18607), .A2(n18604), .B1(n18310), .B2(n18353), .ZN(
        n18281) );
  AOI22_X1 U21343 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18281), .B1(
        n18603), .B2(n18597), .ZN(n18266) );
  OAI211_X1 U21344 ( .C1(n18611), .C2(n18284), .A(n18267), .B(n18266), .ZN(
        P3_U2876) );
  INV_X1 U21345 ( .A(n18570), .ZN(n18617) );
  AOI22_X1 U21346 ( .A1(n18597), .A2(n18613), .B1(n18612), .B2(n18280), .ZN(
        n18269) );
  AOI22_X1 U21347 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18281), .B1(
        n18303), .B2(n18614), .ZN(n18268) );
  OAI211_X1 U21348 ( .C1(n18617), .C2(n18284), .A(n18269), .B(n18268), .ZN(
        P3_U2877) );
  INV_X1 U21349 ( .A(n18574), .ZN(n18623) );
  AOI22_X1 U21350 ( .A1(n18597), .A2(n18620), .B1(n18618), .B2(n18280), .ZN(
        n18271) );
  AOI22_X1 U21351 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18281), .B1(
        n18303), .B2(n18619), .ZN(n18270) );
  OAI211_X1 U21352 ( .C1(n18623), .C2(n18284), .A(n18271), .B(n18270), .ZN(
        P3_U2878) );
  INV_X1 U21353 ( .A(n18578), .ZN(n18629) );
  AOI22_X1 U21354 ( .A1(n18303), .A2(n18626), .B1(n18624), .B2(n18280), .ZN(
        n18273) );
  AOI22_X1 U21355 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18281), .B1(
        n18597), .B2(n18625), .ZN(n18272) );
  OAI211_X1 U21356 ( .C1(n18629), .C2(n18284), .A(n18273), .B(n18272), .ZN(
        P3_U2879) );
  AOI22_X1 U21357 ( .A1(n18597), .A2(n18632), .B1(n18630), .B2(n18280), .ZN(
        n18275) );
  AOI22_X1 U21358 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18281), .B1(
        n18303), .B2(n18631), .ZN(n18274) );
  OAI211_X1 U21359 ( .C1(n18635), .C2(n18284), .A(n18275), .B(n18274), .ZN(
        P3_U2880) );
  INV_X1 U21360 ( .A(n18586), .ZN(n18641) );
  AOI22_X1 U21361 ( .A1(n18303), .A2(n18637), .B1(n18636), .B2(n18280), .ZN(
        n18277) );
  AOI22_X1 U21362 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18281), .B1(
        n18597), .B2(n18638), .ZN(n18276) );
  OAI211_X1 U21363 ( .C1(n18641), .C2(n18284), .A(n18277), .B(n18276), .ZN(
        P3_U2881) );
  INV_X1 U21364 ( .A(n18590), .ZN(n18647) );
  AOI22_X1 U21365 ( .A1(n18597), .A2(n18644), .B1(n18642), .B2(n18280), .ZN(
        n18279) );
  AOI22_X1 U21366 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18281), .B1(
        n18303), .B2(n18643), .ZN(n18278) );
  OAI211_X1 U21367 ( .C1(n18647), .C2(n18284), .A(n18279), .B(n18278), .ZN(
        P3_U2882) );
  INV_X1 U21368 ( .A(n18596), .ZN(n18657) );
  AOI22_X1 U21369 ( .A1(n18303), .A2(n18652), .B1(n18649), .B2(n18280), .ZN(
        n18283) );
  AOI22_X1 U21370 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18281), .B1(
        n18597), .B2(n18651), .ZN(n18282) );
  OAI211_X1 U21371 ( .C1(n18657), .C2(n18284), .A(n18283), .B(n18282), .ZN(
        P3_U2883) );
  NAND2_X1 U21372 ( .A1(n18310), .A2(n18467), .ZN(n18307) );
  NOR2_X1 U21373 ( .A1(n18348), .A2(n18370), .ZN(n18330) );
  NOR2_X1 U21374 ( .A1(n9746), .A2(n18330), .ZN(n18301) );
  AOI22_X1 U21375 ( .A1(n18303), .A2(n18603), .B1(n18602), .B2(n18301), .ZN(
        n18288) );
  AOI221_X1 U21376 ( .B1(n18330), .B2(n18564), .C1(n18330), .C2(n18285), .A(
        n18563), .ZN(n18286) );
  INV_X1 U21377 ( .A(n18286), .ZN(n18304) );
  AOI22_X1 U21378 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18304), .B1(
        n18326), .B2(n18608), .ZN(n18287) );
  OAI211_X1 U21379 ( .C1(n18611), .C2(n18307), .A(n18288), .B(n18287), .ZN(
        P3_U2884) );
  AOI22_X1 U21380 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18304), .B1(
        n18612), .B2(n18301), .ZN(n18290) );
  AOI22_X1 U21381 ( .A1(n18303), .A2(n18613), .B1(n18302), .B2(n18614), .ZN(
        n18289) );
  OAI211_X1 U21382 ( .C1(n18617), .C2(n18307), .A(n18290), .B(n18289), .ZN(
        P3_U2885) );
  AOI22_X1 U21383 ( .A1(n18302), .A2(n18619), .B1(n18618), .B2(n18301), .ZN(
        n18292) );
  AOI22_X1 U21384 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18304), .B1(
        n18303), .B2(n18620), .ZN(n18291) );
  OAI211_X1 U21385 ( .C1(n18623), .C2(n18307), .A(n18292), .B(n18291), .ZN(
        P3_U2886) );
  AOI22_X1 U21386 ( .A1(n18303), .A2(n18625), .B1(n18624), .B2(n18301), .ZN(
        n18294) );
  AOI22_X1 U21387 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18304), .B1(
        n18302), .B2(n18626), .ZN(n18293) );
  OAI211_X1 U21388 ( .C1(n18629), .C2(n18307), .A(n18294), .B(n18293), .ZN(
        P3_U2887) );
  AOI22_X1 U21389 ( .A1(n18302), .A2(n18631), .B1(n18630), .B2(n18301), .ZN(
        n18296) );
  AOI22_X1 U21390 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18304), .B1(
        n18303), .B2(n18632), .ZN(n18295) );
  OAI211_X1 U21391 ( .C1(n18635), .C2(n18307), .A(n18296), .B(n18295), .ZN(
        P3_U2888) );
  AOI22_X1 U21392 ( .A1(n18303), .A2(n18638), .B1(n18636), .B2(n18301), .ZN(
        n18298) );
  AOI22_X1 U21393 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18304), .B1(
        n18302), .B2(n18637), .ZN(n18297) );
  OAI211_X1 U21394 ( .C1(n18641), .C2(n18307), .A(n18298), .B(n18297), .ZN(
        P3_U2889) );
  AOI22_X1 U21395 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18304), .B1(
        n18642), .B2(n18301), .ZN(n18300) );
  AOI22_X1 U21396 ( .A1(n18303), .A2(n18644), .B1(n18302), .B2(n18643), .ZN(
        n18299) );
  OAI211_X1 U21397 ( .C1(n18647), .C2(n18307), .A(n18300), .B(n18299), .ZN(
        P3_U2890) );
  AOI22_X1 U21398 ( .A1(n18302), .A2(n18652), .B1(n18649), .B2(n18301), .ZN(
        n18306) );
  AOI22_X1 U21399 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18304), .B1(
        n18303), .B2(n18651), .ZN(n18305) );
  OAI211_X1 U21400 ( .C1(n18657), .C2(n18307), .A(n18306), .B(n18305), .ZN(
        P3_U2891) );
  INV_X1 U21401 ( .A(n18308), .ZN(n18698) );
  NOR2_X2 U21402 ( .A1(n18698), .A2(n18352), .ZN(n18394) );
  AOI22_X1 U21403 ( .A1(n18326), .A2(n18603), .B1(n18602), .B2(n18325), .ZN(
        n18312) );
  AOI21_X1 U21404 ( .B1(n18699), .B2(n18564), .A(n18309), .ZN(n18401) );
  NAND2_X1 U21405 ( .A1(n18310), .A2(n18401), .ZN(n18327) );
  AOI22_X1 U21406 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18327), .B1(
        n18608), .B2(n18348), .ZN(n18311) );
  OAI211_X1 U21407 ( .C1(n18611), .C2(n18377), .A(n18312), .B(n18311), .ZN(
        P3_U2892) );
  AOI22_X1 U21408 ( .A1(n18326), .A2(n18613), .B1(n18612), .B2(n18325), .ZN(
        n18314) );
  AOI22_X1 U21409 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18327), .B1(
        n18614), .B2(n18348), .ZN(n18313) );
  OAI211_X1 U21410 ( .C1(n18617), .C2(n18377), .A(n18314), .B(n18313), .ZN(
        P3_U2893) );
  AOI22_X1 U21411 ( .A1(n18326), .A2(n18620), .B1(n18618), .B2(n18325), .ZN(
        n18316) );
  AOI22_X1 U21412 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18327), .B1(
        n18619), .B2(n18348), .ZN(n18315) );
  OAI211_X1 U21413 ( .C1(n18623), .C2(n18377), .A(n18316), .B(n18315), .ZN(
        P3_U2894) );
  AOI22_X1 U21414 ( .A1(n18326), .A2(n18625), .B1(n18624), .B2(n18325), .ZN(
        n18318) );
  AOI22_X1 U21415 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18327), .B1(
        n18626), .B2(n18348), .ZN(n18317) );
  OAI211_X1 U21416 ( .C1(n18629), .C2(n18377), .A(n18318), .B(n18317), .ZN(
        P3_U2895) );
  AOI22_X1 U21417 ( .A1(n18631), .A2(n18348), .B1(n18630), .B2(n18325), .ZN(
        n18320) );
  AOI22_X1 U21418 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18327), .B1(
        n18326), .B2(n18632), .ZN(n18319) );
  OAI211_X1 U21419 ( .C1(n18635), .C2(n18377), .A(n18320), .B(n18319), .ZN(
        P3_U2896) );
  AOI22_X1 U21420 ( .A1(n18637), .A2(n18348), .B1(n18636), .B2(n18325), .ZN(
        n18322) );
  AOI22_X1 U21421 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18327), .B1(
        n18326), .B2(n18638), .ZN(n18321) );
  OAI211_X1 U21422 ( .C1(n18641), .C2(n18377), .A(n18322), .B(n18321), .ZN(
        P3_U2897) );
  AOI22_X1 U21423 ( .A1(n18643), .A2(n18348), .B1(n18642), .B2(n18325), .ZN(
        n18324) );
  AOI22_X1 U21424 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18327), .B1(
        n18326), .B2(n18644), .ZN(n18323) );
  OAI211_X1 U21425 ( .C1(n18647), .C2(n18377), .A(n18324), .B(n18323), .ZN(
        P3_U2898) );
  AOI22_X1 U21426 ( .A1(n18649), .A2(n18325), .B1(n18652), .B2(n18348), .ZN(
        n18329) );
  AOI22_X1 U21427 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18327), .B1(
        n18326), .B2(n18651), .ZN(n18328) );
  OAI211_X1 U21428 ( .C1(n18657), .C2(n18377), .A(n18329), .B(n18328), .ZN(
        P3_U2899) );
  INV_X1 U21429 ( .A(n18400), .ZN(n18399) );
  NOR2_X2 U21430 ( .A1(n18700), .A2(n18399), .ZN(n18417) );
  AOI21_X1 U21431 ( .B1(n18377), .B2(n18376), .A(n9746), .ZN(n18347) );
  AOI22_X1 U21432 ( .A1(n18608), .A2(n18370), .B1(n18602), .B2(n18347), .ZN(
        n18334) );
  AOI221_X1 U21433 ( .B1(n18330), .B2(n18377), .C1(n18564), .C2(n18377), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18332) );
  OAI21_X1 U21434 ( .B1(n18417), .B2(n18332), .A(n18331), .ZN(n18349) );
  AOI22_X1 U21435 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18349), .B1(
        n18603), .B2(n18348), .ZN(n18333) );
  OAI211_X1 U21436 ( .C1(n18611), .C2(n18376), .A(n18334), .B(n18333), .ZN(
        P3_U2900) );
  AOI22_X1 U21437 ( .A1(n18614), .A2(n18370), .B1(n18612), .B2(n18347), .ZN(
        n18336) );
  AOI22_X1 U21438 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18349), .B1(
        n18613), .B2(n18348), .ZN(n18335) );
  OAI211_X1 U21439 ( .C1(n18617), .C2(n18376), .A(n18336), .B(n18335), .ZN(
        P3_U2901) );
  AOI22_X1 U21440 ( .A1(n18620), .A2(n18348), .B1(n18618), .B2(n18347), .ZN(
        n18338) );
  AOI22_X1 U21441 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18349), .B1(
        n18619), .B2(n18370), .ZN(n18337) );
  OAI211_X1 U21442 ( .C1(n18623), .C2(n18376), .A(n18338), .B(n18337), .ZN(
        P3_U2902) );
  AOI22_X1 U21443 ( .A1(n18626), .A2(n18370), .B1(n18624), .B2(n18347), .ZN(
        n18340) );
  AOI22_X1 U21444 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18349), .B1(
        n18625), .B2(n18348), .ZN(n18339) );
  OAI211_X1 U21445 ( .C1(n18629), .C2(n18376), .A(n18340), .B(n18339), .ZN(
        P3_U2903) );
  AOI22_X1 U21446 ( .A1(n18632), .A2(n18348), .B1(n18630), .B2(n18347), .ZN(
        n18342) );
  AOI22_X1 U21447 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18349), .B1(
        n18631), .B2(n18370), .ZN(n18341) );
  OAI211_X1 U21448 ( .C1(n18635), .C2(n18376), .A(n18342), .B(n18341), .ZN(
        P3_U2904) );
  AOI22_X1 U21449 ( .A1(n18636), .A2(n18347), .B1(n18638), .B2(n18348), .ZN(
        n18344) );
  AOI22_X1 U21450 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18349), .B1(
        n18637), .B2(n18370), .ZN(n18343) );
  OAI211_X1 U21451 ( .C1(n18641), .C2(n18376), .A(n18344), .B(n18343), .ZN(
        P3_U2905) );
  AOI22_X1 U21452 ( .A1(n18643), .A2(n18370), .B1(n18642), .B2(n18347), .ZN(
        n18346) );
  AOI22_X1 U21453 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18349), .B1(
        n18644), .B2(n18348), .ZN(n18345) );
  OAI211_X1 U21454 ( .C1(n18647), .C2(n18376), .A(n18346), .B(n18345), .ZN(
        P3_U2906) );
  AOI22_X1 U21455 ( .A1(n18649), .A2(n18347), .B1(n18652), .B2(n18370), .ZN(
        n18351) );
  AOI22_X1 U21456 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18349), .B1(
        n18651), .B2(n18348), .ZN(n18350) );
  OAI211_X1 U21457 ( .C1(n18657), .C2(n18376), .A(n18351), .B(n18350), .ZN(
        P3_U2907) );
  NAND2_X1 U21458 ( .A1(n18444), .A2(n18400), .ZN(n18374) );
  AOI22_X1 U21459 ( .A1(n18603), .A2(n18370), .B1(n18602), .B2(n18369), .ZN(
        n18356) );
  NOR2_X1 U21460 ( .A1(n18699), .A2(n18352), .ZN(n18354) );
  AOI22_X1 U21461 ( .A1(n18607), .A2(n18354), .B1(n18353), .B2(n18400), .ZN(
        n18371) );
  AOI22_X1 U21462 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18371), .B1(
        n18608), .B2(n18394), .ZN(n18355) );
  OAI211_X1 U21463 ( .C1(n18611), .C2(n18374), .A(n18356), .B(n18355), .ZN(
        P3_U2908) );
  AOI22_X1 U21464 ( .A1(n18613), .A2(n18370), .B1(n18612), .B2(n18369), .ZN(
        n18358) );
  AOI22_X1 U21465 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18371), .B1(
        n18614), .B2(n18394), .ZN(n18357) );
  OAI211_X1 U21466 ( .C1(n18617), .C2(n18374), .A(n18358), .B(n18357), .ZN(
        P3_U2909) );
  AOI22_X1 U21467 ( .A1(n18619), .A2(n18394), .B1(n18618), .B2(n18369), .ZN(
        n18360) );
  AOI22_X1 U21468 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18371), .B1(
        n18620), .B2(n18370), .ZN(n18359) );
  OAI211_X1 U21469 ( .C1(n18623), .C2(n18374), .A(n18360), .B(n18359), .ZN(
        P3_U2910) );
  AOI22_X1 U21470 ( .A1(n18625), .A2(n18370), .B1(n18624), .B2(n18369), .ZN(
        n18362) );
  AOI22_X1 U21471 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18371), .B1(
        n18626), .B2(n18394), .ZN(n18361) );
  OAI211_X1 U21472 ( .C1(n18629), .C2(n18374), .A(n18362), .B(n18361), .ZN(
        P3_U2911) );
  AOI22_X1 U21473 ( .A1(n18632), .A2(n18370), .B1(n18630), .B2(n18369), .ZN(
        n18364) );
  AOI22_X1 U21474 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18371), .B1(
        n18631), .B2(n18394), .ZN(n18363) );
  OAI211_X1 U21475 ( .C1(n18635), .C2(n18374), .A(n18364), .B(n18363), .ZN(
        P3_U2912) );
  AOI22_X1 U21476 ( .A1(n18637), .A2(n18394), .B1(n18636), .B2(n18369), .ZN(
        n18366) );
  AOI22_X1 U21477 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18371), .B1(
        n18638), .B2(n18370), .ZN(n18365) );
  OAI211_X1 U21478 ( .C1(n18641), .C2(n18374), .A(n18366), .B(n18365), .ZN(
        P3_U2913) );
  AOI22_X1 U21479 ( .A1(n18644), .A2(n18370), .B1(n18642), .B2(n18369), .ZN(
        n18368) );
  AOI22_X1 U21480 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18371), .B1(
        n18643), .B2(n18394), .ZN(n18367) );
  OAI211_X1 U21481 ( .C1(n18647), .C2(n18374), .A(n18368), .B(n18367), .ZN(
        P3_U2914) );
  AOI22_X1 U21482 ( .A1(n18649), .A2(n18369), .B1(n18652), .B2(n18394), .ZN(
        n18373) );
  AOI22_X1 U21483 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18371), .B1(
        n18651), .B2(n18370), .ZN(n18372) );
  OAI211_X1 U21484 ( .C1(n18657), .C2(n18374), .A(n18373), .B(n18372), .ZN(
        P3_U2915) );
  NAND2_X1 U21485 ( .A1(n18467), .A2(n18400), .ZN(n18398) );
  INV_X1 U21486 ( .A(n18374), .ZN(n18440) );
  NOR2_X1 U21487 ( .A1(n18440), .A2(n18463), .ZN(n18375) );
  NOR2_X1 U21488 ( .A1(n9746), .A2(n18375), .ZN(n18393) );
  AOI22_X1 U21489 ( .A1(n18603), .A2(n18394), .B1(n18602), .B2(n18393), .ZN(
        n18380) );
  INV_X1 U21490 ( .A(n18375), .ZN(n18423) );
  NAND2_X1 U21491 ( .A1(n18377), .A2(n18376), .ZN(n18378) );
  INV_X1 U21492 ( .A(n18563), .ZN(n18468) );
  OAI221_X1 U21493 ( .B1(n18423), .B2(n18470), .C1(n18423), .C2(n18378), .A(
        n18468), .ZN(n18395) );
  AOI22_X1 U21494 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18395), .B1(
        n18608), .B2(n18417), .ZN(n18379) );
  OAI211_X1 U21495 ( .C1(n18611), .C2(n18398), .A(n18380), .B(n18379), .ZN(
        P3_U2916) );
  AOI22_X1 U21496 ( .A1(n18614), .A2(n18417), .B1(n18612), .B2(n18393), .ZN(
        n18382) );
  AOI22_X1 U21497 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18395), .B1(
        n18613), .B2(n18394), .ZN(n18381) );
  OAI211_X1 U21498 ( .C1(n18617), .C2(n18398), .A(n18382), .B(n18381), .ZN(
        P3_U2917) );
  AOI22_X1 U21499 ( .A1(n18619), .A2(n18417), .B1(n18618), .B2(n18393), .ZN(
        n18384) );
  AOI22_X1 U21500 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18395), .B1(
        n18620), .B2(n18394), .ZN(n18383) );
  OAI211_X1 U21501 ( .C1(n18623), .C2(n18398), .A(n18384), .B(n18383), .ZN(
        P3_U2918) );
  AOI22_X1 U21502 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18395), .B1(
        n18624), .B2(n18393), .ZN(n18386) );
  AOI22_X1 U21503 ( .A1(n18626), .A2(n18417), .B1(n18625), .B2(n18394), .ZN(
        n18385) );
  OAI211_X1 U21504 ( .C1(n18629), .C2(n18398), .A(n18386), .B(n18385), .ZN(
        P3_U2919) );
  AOI22_X1 U21505 ( .A1(n18632), .A2(n18394), .B1(n18630), .B2(n18393), .ZN(
        n18388) );
  AOI22_X1 U21506 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18395), .B1(
        n18631), .B2(n18417), .ZN(n18387) );
  OAI211_X1 U21507 ( .C1(n18635), .C2(n18398), .A(n18388), .B(n18387), .ZN(
        P3_U2920) );
  AOI22_X1 U21508 ( .A1(n18637), .A2(n18417), .B1(n18636), .B2(n18393), .ZN(
        n18390) );
  AOI22_X1 U21509 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18395), .B1(
        n18638), .B2(n18394), .ZN(n18389) );
  OAI211_X1 U21510 ( .C1(n18641), .C2(n18398), .A(n18390), .B(n18389), .ZN(
        P3_U2921) );
  AOI22_X1 U21511 ( .A1(n18644), .A2(n18394), .B1(n18642), .B2(n18393), .ZN(
        n18392) );
  AOI22_X1 U21512 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18395), .B1(
        n18643), .B2(n18417), .ZN(n18391) );
  OAI211_X1 U21513 ( .C1(n18647), .C2(n18398), .A(n18392), .B(n18391), .ZN(
        P3_U2922) );
  AOI22_X1 U21514 ( .A1(n18649), .A2(n18393), .B1(n18652), .B2(n18417), .ZN(
        n18397) );
  AOI22_X1 U21515 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18395), .B1(
        n18651), .B2(n18394), .ZN(n18396) );
  OAI211_X1 U21516 ( .C1(n18657), .C2(n18398), .A(n18397), .B(n18396), .ZN(
        P3_U2923) );
  NOR2_X2 U21517 ( .A1(n18698), .A2(n18399), .ZN(n18488) );
  INV_X1 U21518 ( .A(n18488), .ZN(n18421) );
  AOI22_X1 U21519 ( .A1(n18608), .A2(n18440), .B1(n18602), .B2(n18416), .ZN(
        n18403) );
  NAND2_X1 U21520 ( .A1(n18401), .A2(n18400), .ZN(n18418) );
  AOI22_X1 U21521 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18418), .B1(
        n18603), .B2(n18417), .ZN(n18402) );
  OAI211_X1 U21522 ( .C1(n18611), .C2(n18421), .A(n18403), .B(n18402), .ZN(
        P3_U2924) );
  AOI22_X1 U21523 ( .A1(n18613), .A2(n18417), .B1(n18612), .B2(n18416), .ZN(
        n18405) );
  AOI22_X1 U21524 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18418), .B1(
        n18614), .B2(n18440), .ZN(n18404) );
  OAI211_X1 U21525 ( .C1(n18617), .C2(n18421), .A(n18405), .B(n18404), .ZN(
        P3_U2925) );
  AOI22_X1 U21526 ( .A1(n18619), .A2(n18440), .B1(n18618), .B2(n18416), .ZN(
        n18407) );
  AOI22_X1 U21527 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18418), .B1(
        n18620), .B2(n18417), .ZN(n18406) );
  OAI211_X1 U21528 ( .C1(n18623), .C2(n18421), .A(n18407), .B(n18406), .ZN(
        P3_U2926) );
  AOI22_X1 U21529 ( .A1(n18626), .A2(n18440), .B1(n18624), .B2(n18416), .ZN(
        n18409) );
  AOI22_X1 U21530 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18418), .B1(
        n18625), .B2(n18417), .ZN(n18408) );
  OAI211_X1 U21531 ( .C1(n18629), .C2(n18421), .A(n18409), .B(n18408), .ZN(
        P3_U2927) );
  AOI22_X1 U21532 ( .A1(n18632), .A2(n18417), .B1(n18630), .B2(n18416), .ZN(
        n18411) );
  AOI22_X1 U21533 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18418), .B1(
        n18631), .B2(n18440), .ZN(n18410) );
  OAI211_X1 U21534 ( .C1(n18635), .C2(n18421), .A(n18411), .B(n18410), .ZN(
        P3_U2928) );
  AOI22_X1 U21535 ( .A1(n18636), .A2(n18416), .B1(n18638), .B2(n18417), .ZN(
        n18413) );
  AOI22_X1 U21536 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18418), .B1(
        n18637), .B2(n18440), .ZN(n18412) );
  OAI211_X1 U21537 ( .C1(n18641), .C2(n18421), .A(n18413), .B(n18412), .ZN(
        P3_U2929) );
  AOI22_X1 U21538 ( .A1(n18644), .A2(n18417), .B1(n18642), .B2(n18416), .ZN(
        n18415) );
  AOI22_X1 U21539 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18418), .B1(
        n18643), .B2(n18440), .ZN(n18414) );
  OAI211_X1 U21540 ( .C1(n18647), .C2(n18421), .A(n18415), .B(n18414), .ZN(
        P3_U2930) );
  AOI22_X1 U21541 ( .A1(n18651), .A2(n18417), .B1(n18649), .B2(n18416), .ZN(
        n18420) );
  AOI22_X1 U21542 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18418), .B1(
        n18652), .B2(n18440), .ZN(n18419) );
  OAI211_X1 U21543 ( .C1(n18657), .C2(n18421), .A(n18420), .B(n18419), .ZN(
        P3_U2931) );
  NOR2_X2 U21544 ( .A1(n18700), .A2(n18491), .ZN(n18510) );
  INV_X1 U21545 ( .A(n18510), .ZN(n18443) );
  NOR2_X1 U21546 ( .A1(n18488), .A2(n18510), .ZN(n18422) );
  NOR2_X1 U21547 ( .A1(n9746), .A2(n18422), .ZN(n18438) );
  AOI22_X1 U21548 ( .A1(n18603), .A2(n18440), .B1(n18602), .B2(n18438), .ZN(
        n18425) );
  INV_X1 U21549 ( .A(n18422), .ZN(n18469) );
  OAI221_X1 U21550 ( .B1(n18469), .B2(n18470), .C1(n18469), .C2(n18423), .A(
        n18468), .ZN(n18439) );
  AOI22_X1 U21551 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18439), .B1(
        n18608), .B2(n18463), .ZN(n18424) );
  OAI211_X1 U21552 ( .C1(n18611), .C2(n18443), .A(n18425), .B(n18424), .ZN(
        P3_U2932) );
  AOI22_X1 U21553 ( .A1(n18613), .A2(n18440), .B1(n18612), .B2(n18438), .ZN(
        n18427) );
  AOI22_X1 U21554 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18439), .B1(
        n18614), .B2(n18463), .ZN(n18426) );
  OAI211_X1 U21555 ( .C1(n18617), .C2(n18443), .A(n18427), .B(n18426), .ZN(
        P3_U2933) );
  AOI22_X1 U21556 ( .A1(n18619), .A2(n18463), .B1(n18618), .B2(n18438), .ZN(
        n18429) );
  AOI22_X1 U21557 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18439), .B1(
        n18620), .B2(n18440), .ZN(n18428) );
  OAI211_X1 U21558 ( .C1(n18623), .C2(n18443), .A(n18429), .B(n18428), .ZN(
        P3_U2934) );
  AOI22_X1 U21559 ( .A1(n18626), .A2(n18463), .B1(n18624), .B2(n18438), .ZN(
        n18431) );
  AOI22_X1 U21560 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18439), .B1(
        n18625), .B2(n18440), .ZN(n18430) );
  OAI211_X1 U21561 ( .C1(n18629), .C2(n18443), .A(n18431), .B(n18430), .ZN(
        P3_U2935) );
  AOI22_X1 U21562 ( .A1(n18631), .A2(n18463), .B1(n18630), .B2(n18438), .ZN(
        n18433) );
  AOI22_X1 U21563 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18439), .B1(
        n18632), .B2(n18440), .ZN(n18432) );
  OAI211_X1 U21564 ( .C1(n18635), .C2(n18443), .A(n18433), .B(n18432), .ZN(
        P3_U2936) );
  AOI22_X1 U21565 ( .A1(n18636), .A2(n18438), .B1(n18638), .B2(n18440), .ZN(
        n18435) );
  AOI22_X1 U21566 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18439), .B1(
        n18637), .B2(n18463), .ZN(n18434) );
  OAI211_X1 U21567 ( .C1(n18641), .C2(n18443), .A(n18435), .B(n18434), .ZN(
        P3_U2937) );
  AOI22_X1 U21568 ( .A1(n18643), .A2(n18463), .B1(n18642), .B2(n18438), .ZN(
        n18437) );
  AOI22_X1 U21569 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18439), .B1(
        n18644), .B2(n18440), .ZN(n18436) );
  OAI211_X1 U21570 ( .C1(n18647), .C2(n18443), .A(n18437), .B(n18436), .ZN(
        P3_U2938) );
  AOI22_X1 U21571 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18439), .B1(
        n18649), .B2(n18438), .ZN(n18442) );
  AOI22_X1 U21572 ( .A1(n18651), .A2(n18440), .B1(n18652), .B2(n18463), .ZN(
        n18441) );
  OAI211_X1 U21573 ( .C1(n18657), .C2(n18443), .A(n18442), .B(n18441), .ZN(
        P3_U2939) );
  NAND2_X1 U21574 ( .A1(n18444), .A2(n18493), .ZN(n18494) );
  AOI22_X1 U21575 ( .A1(n18608), .A2(n18488), .B1(n18602), .B2(n18462), .ZN(
        n18449) );
  NOR2_X1 U21576 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18445), .ZN(
        n18447) );
  NOR2_X1 U21577 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18491), .ZN(
        n18446) );
  AOI22_X1 U21578 ( .A1(n18607), .A2(n18447), .B1(n18605), .B2(n18446), .ZN(
        n18464) );
  AOI22_X1 U21579 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18464), .B1(
        n18603), .B2(n18463), .ZN(n18448) );
  OAI211_X1 U21580 ( .C1(n18611), .C2(n18494), .A(n18449), .B(n18448), .ZN(
        P3_U2940) );
  AOI22_X1 U21581 ( .A1(n18614), .A2(n18488), .B1(n18612), .B2(n18462), .ZN(
        n18451) );
  AOI22_X1 U21582 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18464), .B1(
        n18613), .B2(n18463), .ZN(n18450) );
  OAI211_X1 U21583 ( .C1(n18617), .C2(n18494), .A(n18451), .B(n18450), .ZN(
        P3_U2941) );
  AOI22_X1 U21584 ( .A1(n18620), .A2(n18463), .B1(n18618), .B2(n18462), .ZN(
        n18453) );
  AOI22_X1 U21585 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18464), .B1(
        n18619), .B2(n18488), .ZN(n18452) );
  OAI211_X1 U21586 ( .C1(n18623), .C2(n18494), .A(n18453), .B(n18452), .ZN(
        P3_U2942) );
  AOI22_X1 U21587 ( .A1(n18625), .A2(n18463), .B1(n18624), .B2(n18462), .ZN(
        n18455) );
  AOI22_X1 U21588 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18464), .B1(
        n18626), .B2(n18488), .ZN(n18454) );
  OAI211_X1 U21589 ( .C1(n18629), .C2(n18494), .A(n18455), .B(n18454), .ZN(
        P3_U2943) );
  AOI22_X1 U21590 ( .A1(n18631), .A2(n18488), .B1(n18630), .B2(n18462), .ZN(
        n18457) );
  AOI22_X1 U21591 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18464), .B1(
        n18632), .B2(n18463), .ZN(n18456) );
  OAI211_X1 U21592 ( .C1(n18635), .C2(n18494), .A(n18457), .B(n18456), .ZN(
        P3_U2944) );
  AOI22_X1 U21593 ( .A1(n18636), .A2(n18462), .B1(n18638), .B2(n18463), .ZN(
        n18459) );
  AOI22_X1 U21594 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18464), .B1(
        n18637), .B2(n18488), .ZN(n18458) );
  OAI211_X1 U21595 ( .C1(n18641), .C2(n18494), .A(n18459), .B(n18458), .ZN(
        P3_U2945) );
  AOI22_X1 U21596 ( .A1(n18644), .A2(n18463), .B1(n18642), .B2(n18462), .ZN(
        n18461) );
  AOI22_X1 U21597 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18464), .B1(
        n18643), .B2(n18488), .ZN(n18460) );
  OAI211_X1 U21598 ( .C1(n18647), .C2(n18494), .A(n18461), .B(n18460), .ZN(
        P3_U2946) );
  AOI22_X1 U21599 ( .A1(n18651), .A2(n18463), .B1(n18649), .B2(n18462), .ZN(
        n18466) );
  AOI22_X1 U21600 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18464), .B1(
        n18652), .B2(n18488), .ZN(n18465) );
  OAI211_X1 U21601 ( .C1(n18657), .C2(n18494), .A(n18466), .B(n18465), .ZN(
        P3_U2947) );
  NAND2_X1 U21602 ( .A1(n18467), .A2(n18493), .ZN(n18520) );
  NAND2_X1 U21603 ( .A1(n18494), .A2(n18520), .ZN(n18471) );
  OAI221_X1 U21604 ( .B1(n18471), .B2(n18470), .C1(n18471), .C2(n18469), .A(
        n18468), .ZN(n18487) );
  AOI21_X1 U21605 ( .B1(n18494), .B2(n18520), .A(n9746), .ZN(n18486) );
  AOI22_X1 U21606 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18487), .B1(
        n18602), .B2(n18486), .ZN(n18473) );
  AOI22_X1 U21607 ( .A1(n18603), .A2(n18488), .B1(n18608), .B2(n18510), .ZN(
        n18472) );
  OAI211_X1 U21608 ( .C1(n18611), .C2(n18520), .A(n18473), .B(n18472), .ZN(
        P3_U2948) );
  AOI22_X1 U21609 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18487), .B1(
        n18612), .B2(n18486), .ZN(n18475) );
  AOI22_X1 U21610 ( .A1(n18613), .A2(n18488), .B1(n18614), .B2(n18510), .ZN(
        n18474) );
  OAI211_X1 U21611 ( .C1(n18617), .C2(n18520), .A(n18475), .B(n18474), .ZN(
        P3_U2949) );
  AOI22_X1 U21612 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18487), .B1(
        n18618), .B2(n18486), .ZN(n18477) );
  AOI22_X1 U21613 ( .A1(n18619), .A2(n18510), .B1(n18620), .B2(n18488), .ZN(
        n18476) );
  OAI211_X1 U21614 ( .C1(n18623), .C2(n18520), .A(n18477), .B(n18476), .ZN(
        P3_U2950) );
  AOI22_X1 U21615 ( .A1(n18626), .A2(n18510), .B1(n18624), .B2(n18486), .ZN(
        n18479) );
  AOI22_X1 U21616 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18487), .B1(
        n18625), .B2(n18488), .ZN(n18478) );
  OAI211_X1 U21617 ( .C1(n18629), .C2(n18520), .A(n18479), .B(n18478), .ZN(
        P3_U2951) );
  AOI22_X1 U21618 ( .A1(n18631), .A2(n18510), .B1(n18630), .B2(n18486), .ZN(
        n18481) );
  AOI22_X1 U21619 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18487), .B1(
        n18632), .B2(n18488), .ZN(n18480) );
  OAI211_X1 U21620 ( .C1(n18635), .C2(n18520), .A(n18481), .B(n18480), .ZN(
        P3_U2952) );
  AOI22_X1 U21621 ( .A1(n18636), .A2(n18486), .B1(n18638), .B2(n18488), .ZN(
        n18483) );
  AOI22_X1 U21622 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18487), .B1(
        n18637), .B2(n18510), .ZN(n18482) );
  OAI211_X1 U21623 ( .C1(n18641), .C2(n18520), .A(n18483), .B(n18482), .ZN(
        P3_U2953) );
  AOI22_X1 U21624 ( .A1(n18643), .A2(n18510), .B1(n18642), .B2(n18486), .ZN(
        n18485) );
  AOI22_X1 U21625 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18487), .B1(
        n18644), .B2(n18488), .ZN(n18484) );
  OAI211_X1 U21626 ( .C1(n18647), .C2(n18520), .A(n18485), .B(n18484), .ZN(
        P3_U2954) );
  AOI22_X1 U21627 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18487), .B1(
        n18649), .B2(n18486), .ZN(n18490) );
  AOI22_X1 U21628 ( .A1(n18651), .A2(n18488), .B1(n18652), .B2(n18510), .ZN(
        n18489) );
  OAI211_X1 U21629 ( .C1(n18657), .C2(n18520), .A(n18490), .B(n18489), .ZN(
        P3_U2955) );
  NOR2_X2 U21630 ( .A1(n18698), .A2(n18491), .ZN(n18595) );
  INV_X1 U21631 ( .A(n18595), .ZN(n18514) );
  NOR2_X1 U21632 ( .A1(n18699), .A2(n18491), .ZN(n18542) );
  INV_X1 U21633 ( .A(n18542), .ZN(n18492) );
  NOR2_X1 U21634 ( .A1(n9746), .A2(n18492), .ZN(n18509) );
  AOI22_X1 U21635 ( .A1(n18603), .A2(n18510), .B1(n18602), .B2(n18509), .ZN(
        n18496) );
  OAI211_X1 U21636 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n18607), .A(
        n18605), .B(n18493), .ZN(n18511) );
  AOI22_X1 U21637 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18511), .B1(
        n18608), .B2(n18536), .ZN(n18495) );
  OAI211_X1 U21638 ( .C1(n18611), .C2(n18514), .A(n18496), .B(n18495), .ZN(
        P3_U2956) );
  AOI22_X1 U21639 ( .A1(n18614), .A2(n18536), .B1(n18612), .B2(n18509), .ZN(
        n18498) );
  AOI22_X1 U21640 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18511), .B1(
        n18613), .B2(n18510), .ZN(n18497) );
  OAI211_X1 U21641 ( .C1(n18617), .C2(n18514), .A(n18498), .B(n18497), .ZN(
        P3_U2957) );
  AOI22_X1 U21642 ( .A1(n18620), .A2(n18510), .B1(n18618), .B2(n18509), .ZN(
        n18500) );
  AOI22_X1 U21643 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18511), .B1(
        n18619), .B2(n18536), .ZN(n18499) );
  OAI211_X1 U21644 ( .C1(n18623), .C2(n18514), .A(n18500), .B(n18499), .ZN(
        P3_U2958) );
  AOI22_X1 U21645 ( .A1(n18625), .A2(n18510), .B1(n18624), .B2(n18509), .ZN(
        n18502) );
  AOI22_X1 U21646 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18511), .B1(
        n18626), .B2(n18536), .ZN(n18501) );
  OAI211_X1 U21647 ( .C1(n18629), .C2(n18514), .A(n18502), .B(n18501), .ZN(
        P3_U2959) );
  AOI22_X1 U21648 ( .A1(n18631), .A2(n18536), .B1(n18630), .B2(n18509), .ZN(
        n18504) );
  AOI22_X1 U21649 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18511), .B1(
        n18632), .B2(n18510), .ZN(n18503) );
  OAI211_X1 U21650 ( .C1(n18635), .C2(n18514), .A(n18504), .B(n18503), .ZN(
        P3_U2960) );
  AOI22_X1 U21651 ( .A1(n18636), .A2(n18509), .B1(n18638), .B2(n18510), .ZN(
        n18506) );
  AOI22_X1 U21652 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18511), .B1(
        n18637), .B2(n18536), .ZN(n18505) );
  OAI211_X1 U21653 ( .C1(n18641), .C2(n18514), .A(n18506), .B(n18505), .ZN(
        P3_U2961) );
  AOI22_X1 U21654 ( .A1(n18643), .A2(n18536), .B1(n18642), .B2(n18509), .ZN(
        n18508) );
  AOI22_X1 U21655 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18511), .B1(
        n18644), .B2(n18510), .ZN(n18507) );
  OAI211_X1 U21656 ( .C1(n18647), .C2(n18514), .A(n18508), .B(n18507), .ZN(
        P3_U2962) );
  AOI22_X1 U21657 ( .A1(n18651), .A2(n18510), .B1(n18649), .B2(n18509), .ZN(
        n18513) );
  AOI22_X1 U21658 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18511), .B1(
        n18652), .B2(n18536), .ZN(n18512) );
  OAI211_X1 U21659 ( .C1(n18657), .C2(n18514), .A(n18513), .B(n18512), .ZN(
        P3_U2963) );
  NOR2_X2 U21660 ( .A1(n18541), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18650) );
  INV_X1 U21661 ( .A(n18650), .ZN(n18540) );
  NOR2_X1 U21662 ( .A1(n18595), .A2(n18650), .ZN(n18565) );
  NOR2_X1 U21663 ( .A1(n9746), .A2(n18565), .ZN(n18535) );
  AOI22_X1 U21664 ( .A1(n18603), .A2(n18536), .B1(n18602), .B2(n18535), .ZN(
        n18522) );
  INV_X1 U21665 ( .A(n18565), .ZN(n18519) );
  AOI21_X1 U21666 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18540), .A(n18515), 
        .ZN(n18516) );
  OAI221_X1 U21667 ( .B1(n18519), .B2(n18518), .C1(n18519), .C2(n18517), .A(
        n18516), .ZN(n18537) );
  INV_X1 U21668 ( .A(n18520), .ZN(n18558) );
  AOI22_X1 U21669 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18537), .B1(
        n18608), .B2(n18558), .ZN(n18521) );
  OAI211_X1 U21670 ( .C1(n18611), .C2(n18540), .A(n18522), .B(n18521), .ZN(
        P3_U2964) );
  AOI22_X1 U21671 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18537), .B1(
        n18612), .B2(n18535), .ZN(n18524) );
  AOI22_X1 U21672 ( .A1(n18613), .A2(n18536), .B1(n18614), .B2(n18558), .ZN(
        n18523) );
  OAI211_X1 U21673 ( .C1(n18617), .C2(n18540), .A(n18524), .B(n18523), .ZN(
        P3_U2965) );
  AOI22_X1 U21674 ( .A1(n18619), .A2(n18558), .B1(n18618), .B2(n18535), .ZN(
        n18526) );
  AOI22_X1 U21675 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18537), .B1(
        n18620), .B2(n18536), .ZN(n18525) );
  OAI211_X1 U21676 ( .C1(n18623), .C2(n18540), .A(n18526), .B(n18525), .ZN(
        P3_U2966) );
  AOI22_X1 U21677 ( .A1(n18625), .A2(n18536), .B1(n18624), .B2(n18535), .ZN(
        n18528) );
  AOI22_X1 U21678 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18537), .B1(
        n18626), .B2(n18558), .ZN(n18527) );
  OAI211_X1 U21679 ( .C1(n18629), .C2(n18540), .A(n18528), .B(n18527), .ZN(
        P3_U2967) );
  AOI22_X1 U21680 ( .A1(n18631), .A2(n18558), .B1(n18630), .B2(n18535), .ZN(
        n18530) );
  AOI22_X1 U21681 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18537), .B1(
        n18632), .B2(n18536), .ZN(n18529) );
  OAI211_X1 U21682 ( .C1(n18635), .C2(n18540), .A(n18530), .B(n18529), .ZN(
        P3_U2968) );
  AOI22_X1 U21683 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18537), .B1(
        n18636), .B2(n18535), .ZN(n18532) );
  AOI22_X1 U21684 ( .A1(n18637), .A2(n18558), .B1(n18638), .B2(n18536), .ZN(
        n18531) );
  OAI211_X1 U21685 ( .C1(n18641), .C2(n18540), .A(n18532), .B(n18531), .ZN(
        P3_U2969) );
  AOI22_X1 U21686 ( .A1(n18644), .A2(n18536), .B1(n18642), .B2(n18535), .ZN(
        n18534) );
  AOI22_X1 U21687 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18537), .B1(
        n18643), .B2(n18558), .ZN(n18533) );
  OAI211_X1 U21688 ( .C1(n18647), .C2(n18540), .A(n18534), .B(n18533), .ZN(
        P3_U2970) );
  AOI22_X1 U21689 ( .A1(n18651), .A2(n18536), .B1(n18649), .B2(n18535), .ZN(
        n18539) );
  AOI22_X1 U21690 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18537), .B1(
        n18652), .B2(n18558), .ZN(n18538) );
  OAI211_X1 U21691 ( .C1(n18657), .C2(n18540), .A(n18539), .B(n18538), .ZN(
        P3_U2971) );
  NOR2_X1 U21692 ( .A1(n9746), .A2(n18541), .ZN(n18557) );
  AOI22_X1 U21693 ( .A1(n18603), .A2(n18558), .B1(n18602), .B2(n18557), .ZN(
        n18544) );
  AOI22_X1 U21694 ( .A1(n18607), .A2(n18542), .B1(n18606), .B2(n18605), .ZN(
        n18559) );
  AOI22_X1 U21695 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18559), .B1(
        n18608), .B2(n18595), .ZN(n18543) );
  OAI211_X1 U21696 ( .C1(n18562), .C2(n18611), .A(n18544), .B(n18543), .ZN(
        P3_U2972) );
  AOI22_X1 U21697 ( .A1(n18613), .A2(n18558), .B1(n18612), .B2(n18557), .ZN(
        n18546) );
  AOI22_X1 U21698 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18559), .B1(
        n18614), .B2(n18595), .ZN(n18545) );
  OAI211_X1 U21699 ( .C1(n18562), .C2(n18617), .A(n18546), .B(n18545), .ZN(
        P3_U2973) );
  AOI22_X1 U21700 ( .A1(n18620), .A2(n18558), .B1(n18618), .B2(n18557), .ZN(
        n18548) );
  AOI22_X1 U21701 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18559), .B1(
        n18619), .B2(n18595), .ZN(n18547) );
  OAI211_X1 U21702 ( .C1(n18562), .C2(n18623), .A(n18548), .B(n18547), .ZN(
        P3_U2974) );
  AOI22_X1 U21703 ( .A1(n18625), .A2(n18558), .B1(n18624), .B2(n18557), .ZN(
        n18550) );
  AOI22_X1 U21704 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18559), .B1(
        n18626), .B2(n18595), .ZN(n18549) );
  OAI211_X1 U21705 ( .C1(n18562), .C2(n18629), .A(n18550), .B(n18549), .ZN(
        P3_U2975) );
  AOI22_X1 U21706 ( .A1(n18632), .A2(n18558), .B1(n18630), .B2(n18557), .ZN(
        n18552) );
  AOI22_X1 U21707 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18559), .B1(
        n18631), .B2(n18595), .ZN(n18551) );
  OAI211_X1 U21708 ( .C1(n18562), .C2(n18635), .A(n18552), .B(n18551), .ZN(
        P3_U2976) );
  AOI22_X1 U21709 ( .A1(n18637), .A2(n18595), .B1(n18636), .B2(n18557), .ZN(
        n18554) );
  AOI22_X1 U21710 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18559), .B1(
        n18638), .B2(n18558), .ZN(n18553) );
  OAI211_X1 U21711 ( .C1(n18562), .C2(n18641), .A(n18554), .B(n18553), .ZN(
        P3_U2977) );
  AOI22_X1 U21712 ( .A1(n18644), .A2(n18558), .B1(n18642), .B2(n18557), .ZN(
        n18556) );
  AOI22_X1 U21713 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18559), .B1(
        n18643), .B2(n18595), .ZN(n18555) );
  OAI211_X1 U21714 ( .C1(n18562), .C2(n18647), .A(n18556), .B(n18555), .ZN(
        P3_U2978) );
  AOI22_X1 U21715 ( .A1(n18649), .A2(n18557), .B1(n18652), .B2(n18595), .ZN(
        n18561) );
  AOI22_X1 U21716 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18559), .B1(
        n18651), .B2(n18558), .ZN(n18560) );
  OAI211_X1 U21717 ( .C1(n18562), .C2(n18657), .A(n18561), .B(n18560), .ZN(
        P3_U2979) );
  INV_X1 U21718 ( .A(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n20989) );
  NOR2_X1 U21719 ( .A1(n9746), .A2(n18566), .ZN(n18594) );
  AOI22_X1 U21720 ( .A1(n18603), .A2(n18595), .B1(n18602), .B2(n18594), .ZN(
        n18569) );
  AOI22_X1 U21721 ( .A1(n18567), .A2(n18597), .B1(n18608), .B2(n18650), .ZN(
        n18568) );
  OAI211_X1 U21722 ( .C1(n18600), .C2(n20989), .A(n18569), .B(n18568), .ZN(
        P3_U2980) );
  INV_X1 U21723 ( .A(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n18573) );
  AOI22_X1 U21724 ( .A1(n18614), .A2(n18650), .B1(n18612), .B2(n18594), .ZN(
        n18572) );
  AOI22_X1 U21725 ( .A1(n18597), .A2(n18570), .B1(n18613), .B2(n18595), .ZN(
        n18571) );
  OAI211_X1 U21726 ( .C1(n18600), .C2(n18573), .A(n18572), .B(n18571), .ZN(
        P3_U2981) );
  INV_X1 U21727 ( .A(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n18577) );
  AOI22_X1 U21728 ( .A1(n18620), .A2(n18595), .B1(n18618), .B2(n18594), .ZN(
        n18576) );
  AOI22_X1 U21729 ( .A1(n18597), .A2(n18574), .B1(n18619), .B2(n18650), .ZN(
        n18575) );
  OAI211_X1 U21730 ( .C1(n18600), .C2(n18577), .A(n18576), .B(n18575), .ZN(
        P3_U2982) );
  INV_X1 U21731 ( .A(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18581) );
  AOI22_X1 U21732 ( .A1(n18626), .A2(n18650), .B1(n18624), .B2(n18594), .ZN(
        n18580) );
  AOI22_X1 U21733 ( .A1(n18597), .A2(n18578), .B1(n18625), .B2(n18595), .ZN(
        n18579) );
  OAI211_X1 U21734 ( .C1(n18600), .C2(n18581), .A(n18580), .B(n18579), .ZN(
        P3_U2983) );
  INV_X1 U21735 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n18585) );
  AOI22_X1 U21736 ( .A1(n18632), .A2(n18595), .B1(n18630), .B2(n18594), .ZN(
        n18584) );
  AOI22_X1 U21737 ( .A1(n18597), .A2(n18582), .B1(n18631), .B2(n18650), .ZN(
        n18583) );
  OAI211_X1 U21738 ( .C1(n18600), .C2(n18585), .A(n18584), .B(n18583), .ZN(
        P3_U2984) );
  INV_X1 U21739 ( .A(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n18589) );
  AOI22_X1 U21740 ( .A1(n18636), .A2(n18594), .B1(n18638), .B2(n18595), .ZN(
        n18588) );
  AOI22_X1 U21741 ( .A1(n18597), .A2(n18586), .B1(n18637), .B2(n18650), .ZN(
        n18587) );
  OAI211_X1 U21742 ( .C1(n18600), .C2(n18589), .A(n18588), .B(n18587), .ZN(
        P3_U2985) );
  INV_X1 U21743 ( .A(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18593) );
  AOI22_X1 U21744 ( .A1(n18643), .A2(n18650), .B1(n18642), .B2(n18594), .ZN(
        n18592) );
  AOI22_X1 U21745 ( .A1(n18597), .A2(n18590), .B1(n18644), .B2(n18595), .ZN(
        n18591) );
  OAI211_X1 U21746 ( .C1(n18600), .C2(n18593), .A(n18592), .B(n18591), .ZN(
        P3_U2986) );
  INV_X1 U21747 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n20889) );
  AOI22_X1 U21748 ( .A1(n18651), .A2(n18595), .B1(n18649), .B2(n18594), .ZN(
        n18599) );
  AOI22_X1 U21749 ( .A1(n18597), .A2(n18596), .B1(n18652), .B2(n18650), .ZN(
        n18598) );
  OAI211_X1 U21750 ( .C1(n18600), .C2(n20889), .A(n18599), .B(n18598), .ZN(
        P3_U2987) );
  INV_X1 U21751 ( .A(n18604), .ZN(n18601) );
  NOR2_X1 U21752 ( .A1(n9746), .A2(n18601), .ZN(n18648) );
  AOI22_X1 U21753 ( .A1(n18603), .A2(n18650), .B1(n18602), .B2(n18648), .ZN(
        n18610) );
  AOI22_X1 U21754 ( .A1(n18607), .A2(n18606), .B1(n18605), .B2(n18604), .ZN(
        n18654) );
  AOI22_X1 U21755 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18654), .B1(
        n18653), .B2(n18608), .ZN(n18609) );
  OAI211_X1 U21756 ( .C1(n18658), .C2(n18611), .A(n18610), .B(n18609), .ZN(
        P3_U2988) );
  AOI22_X1 U21757 ( .A1(n18613), .A2(n18650), .B1(n18612), .B2(n18648), .ZN(
        n18616) );
  AOI22_X1 U21758 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18654), .B1(
        n18653), .B2(n18614), .ZN(n18615) );
  OAI211_X1 U21759 ( .C1(n18658), .C2(n18617), .A(n18616), .B(n18615), .ZN(
        P3_U2989) );
  AOI22_X1 U21760 ( .A1(n18653), .A2(n18619), .B1(n18618), .B2(n18648), .ZN(
        n18622) );
  AOI22_X1 U21761 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18654), .B1(
        n18620), .B2(n18650), .ZN(n18621) );
  OAI211_X1 U21762 ( .C1(n18658), .C2(n18623), .A(n18622), .B(n18621), .ZN(
        P3_U2990) );
  AOI22_X1 U21763 ( .A1(n18625), .A2(n18650), .B1(n18624), .B2(n18648), .ZN(
        n18628) );
  AOI22_X1 U21764 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18654), .B1(
        n18653), .B2(n18626), .ZN(n18627) );
  OAI211_X1 U21765 ( .C1(n18658), .C2(n18629), .A(n18628), .B(n18627), .ZN(
        P3_U2991) );
  AOI22_X1 U21766 ( .A1(n18653), .A2(n18631), .B1(n18630), .B2(n18648), .ZN(
        n18634) );
  AOI22_X1 U21767 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18654), .B1(
        n18632), .B2(n18650), .ZN(n18633) );
  OAI211_X1 U21768 ( .C1(n18658), .C2(n18635), .A(n18634), .B(n18633), .ZN(
        P3_U2992) );
  AOI22_X1 U21769 ( .A1(n18653), .A2(n18637), .B1(n18636), .B2(n18648), .ZN(
        n18640) );
  AOI22_X1 U21770 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18654), .B1(
        n18638), .B2(n18650), .ZN(n18639) );
  OAI211_X1 U21771 ( .C1(n18658), .C2(n18641), .A(n18640), .B(n18639), .ZN(
        P3_U2993) );
  AOI22_X1 U21772 ( .A1(n18653), .A2(n18643), .B1(n18642), .B2(n18648), .ZN(
        n18646) );
  AOI22_X1 U21773 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18654), .B1(
        n18644), .B2(n18650), .ZN(n18645) );
  OAI211_X1 U21774 ( .C1(n18658), .C2(n18647), .A(n18646), .B(n18645), .ZN(
        P3_U2994) );
  AOI22_X1 U21775 ( .A1(n18651), .A2(n18650), .B1(n18649), .B2(n18648), .ZN(
        n18656) );
  AOI22_X1 U21776 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18654), .B1(
        n18653), .B2(n18652), .ZN(n18655) );
  OAI211_X1 U21777 ( .C1(n18658), .C2(n18657), .A(n18656), .B(n18655), .ZN(
        P3_U2995) );
  NAND2_X1 U21778 ( .A1(n9819), .A2(n18684), .ZN(n18659) );
  AOI22_X1 U21779 ( .A1(n18662), .A2(n18661), .B1(n18660), .B2(n18659), .ZN(
        n18663) );
  OAI221_X1 U21780 ( .B1(n18666), .B2(n18665), .C1(n18666), .C2(n18664), .A(
        n18663), .ZN(n18866) );
  INV_X1 U21781 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18670) );
  OAI21_X1 U21782 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18667), .ZN(n18668) );
  OAI211_X1 U21783 ( .C1(n18691), .C2(n18670), .A(n18669), .B(n18668), .ZN(
        n18713) );
  NAND2_X1 U21784 ( .A1(n18694), .A2(n12916), .ZN(n18695) );
  AOI22_X1 U21785 ( .A1(n18685), .A2(n18695), .B1(n18690), .B2(n18674), .ZN(
        n18829) );
  NOR2_X1 U21786 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18829), .ZN(
        n18678) );
  OAI21_X1 U21787 ( .B1(n18673), .B2(n18672), .A(n18671), .ZN(n18682) );
  OAI21_X1 U21788 ( .B1(n18685), .B2(n18694), .A(n18674), .ZN(n18675) );
  AOI21_X1 U21789 ( .B1(n18676), .B2(n18682), .A(n18675), .ZN(n18825) );
  NAND2_X1 U21790 ( .A1(n18691), .A2(n18825), .ZN(n18677) );
  AOI22_X1 U21791 ( .A1(n18691), .A2(n18678), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18677), .ZN(n18711) );
  INV_X1 U21792 ( .A(n18691), .ZN(n18702) );
  NAND2_X1 U21793 ( .A1(n13018), .A2(n18848), .ZN(n18689) );
  OAI21_X1 U21794 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18679), .A(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18683) );
  OAI211_X1 U21795 ( .C1(n18680), .C2(n12916), .A(n18679), .B(n13018), .ZN(
        n18681) );
  OAI21_X1 U21796 ( .B1(n18683), .B2(n18682), .A(n18681), .ZN(n18686) );
  OAI22_X1 U21797 ( .A1(n18687), .A2(n18686), .B1(n18685), .B2(n18684), .ZN(
        n18688) );
  AOI22_X1 U21798 ( .A1(n18690), .A2(n18835), .B1(n18689), .B2(n18688), .ZN(
        n18838) );
  AOI22_X1 U21799 ( .A1(n18702), .A2(n13018), .B1(n18838), .B2(n18691), .ZN(
        n18706) );
  NOR2_X1 U21800 ( .A1(n18693), .A2(n18692), .ZN(n18697) );
  AOI22_X1 U21801 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18694), .B1(
        n18697), .B2(n12916), .ZN(n18850) );
  INV_X1 U21802 ( .A(n18695), .ZN(n18696) );
  OAI22_X1 U21803 ( .A1(n18697), .A2(n18841), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18696), .ZN(n18846) );
  AOI222_X1 U21804 ( .A1(n18850), .A2(n18846), .B1(n18850), .B2(n18699), .C1(
        n18846), .C2(n18698), .ZN(n18701) );
  OAI21_X1 U21805 ( .B1(n18702), .B2(n18701), .A(n18700), .ZN(n18705) );
  AND2_X1 U21806 ( .A1(n18706), .A2(n18705), .ZN(n18703) );
  OAI221_X1 U21807 ( .B1(n18706), .B2(n18705), .C1(n18704), .C2(n18703), .A(
        n18708), .ZN(n18710) );
  AOI21_X1 U21808 ( .B1(n18708), .B2(n18707), .A(n18706), .ZN(n18709) );
  AOI222_X1 U21809 ( .A1(n18711), .A2(n18710), .B1(n18711), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18710), .C2(n18709), .ZN(
        n18712) );
  NOR4_X1 U21810 ( .A1(n18714), .A2(n18866), .A3(n18713), .A4(n18712), .ZN(
        n18725) );
  NOR2_X1 U21811 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18877) );
  AOI22_X1 U21812 ( .A1(n18870), .A2(n18715), .B1(n18849), .B2(n18877), .ZN(
        n18716) );
  INV_X1 U21813 ( .A(n18716), .ZN(n18721) );
  OAI211_X1 U21814 ( .C1(n18718), .C2(n18717), .A(n18868), .B(n18725), .ZN(
        n18823) );
  NAND2_X1 U21815 ( .A1(n18870), .A2(n18888), .ZN(n18726) );
  NAND2_X1 U21816 ( .A1(n18823), .A2(n18726), .ZN(n18728) );
  NOR2_X1 U21817 ( .A1(n18719), .A2(n18728), .ZN(n18720) );
  MUX2_X1 U21818 ( .A(n18721), .B(n18720), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18723) );
  OAI211_X1 U21819 ( .C1(n18725), .C2(n18724), .A(n18723), .B(n18722), .ZN(
        P3_U2996) );
  NOR2_X1 U21820 ( .A1(n18875), .A2(n18869), .ZN(n18732) );
  NOR3_X1 U21821 ( .A1(n18834), .A2(n18727), .A3(n18726), .ZN(n18735) );
  NOR3_X1 U21822 ( .A1(n9746), .A2(n18729), .A3(n18728), .ZN(n18731) );
  OR4_X1 U21823 ( .A1(n18733), .A2(n18732), .A3(n18735), .A4(n18731), .ZN(
        P3_U2997) );
  NOR3_X1 U21824 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .ZN(n18736) );
  INV_X1 U21825 ( .A(n18822), .ZN(n18734) );
  NOR4_X1 U21826 ( .A1(n18877), .A2(n18736), .A3(n18735), .A4(n18734), .ZN(
        P3_U2998) );
  AND2_X1 U21827 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18818), .ZN(
        P3_U2999) );
  AND2_X1 U21828 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18737), .ZN(
        P3_U3000) );
  AND2_X1 U21829 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18737), .ZN(
        P3_U3001) );
  AND2_X1 U21830 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18737), .ZN(
        P3_U3002) );
  AND2_X1 U21831 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18737), .ZN(
        P3_U3003) );
  AND2_X1 U21832 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18737), .ZN(
        P3_U3004) );
  INV_X1 U21833 ( .A(P3_DATAWIDTH_REG_25__SCAN_IN), .ZN(n21082) );
  NOR2_X1 U21834 ( .A1(n21082), .A2(n18821), .ZN(P3_U3005) );
  AND2_X1 U21835 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18737), .ZN(
        P3_U3006) );
  AND2_X1 U21836 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18737), .ZN(
        P3_U3007) );
  AND2_X1 U21837 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18737), .ZN(
        P3_U3008) );
  AND2_X1 U21838 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18737), .ZN(
        P3_U3009) );
  AND2_X1 U21839 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18737), .ZN(
        P3_U3010) );
  AND2_X1 U21840 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18737), .ZN(
        P3_U3011) );
  AND2_X1 U21841 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18737), .ZN(
        P3_U3012) );
  AND2_X1 U21842 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18737), .ZN(
        P3_U3013) );
  AND2_X1 U21843 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18737), .ZN(
        P3_U3014) );
  AND2_X1 U21844 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18737), .ZN(
        P3_U3015) );
  AND2_X1 U21845 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18737), .ZN(
        P3_U3016) );
  AND2_X1 U21846 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18737), .ZN(
        P3_U3017) );
  AND2_X1 U21847 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18818), .ZN(
        P3_U3018) );
  AND2_X1 U21848 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18737), .ZN(
        P3_U3019) );
  AND2_X1 U21849 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18737), .ZN(
        P3_U3020) );
  AND2_X1 U21850 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18737), .ZN(P3_U3021) );
  AND2_X1 U21851 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18818), .ZN(P3_U3022) );
  AND2_X1 U21852 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18737), .ZN(P3_U3023) );
  AND2_X1 U21853 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18818), .ZN(P3_U3024) );
  AND2_X1 U21854 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18818), .ZN(P3_U3025) );
  AND2_X1 U21855 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18818), .ZN(P3_U3026) );
  AND2_X1 U21856 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18818), .ZN(P3_U3027) );
  AND2_X1 U21857 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18818), .ZN(P3_U3028) );
  AOI21_X1 U21858 ( .B1(HOLD), .B2(n18738), .A(n20855), .ZN(n18741) );
  NAND2_X1 U21859 ( .A1(n18870), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18744) );
  INV_X1 U21860 ( .A(n18744), .ZN(n20850) );
  NAND2_X1 U21861 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n20852) );
  OAI21_X1 U21862 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(n20852), .A(n18739), 
        .ZN(n18740) );
  AOI211_X1 U21863 ( .C1(P3_REQUESTPENDING_REG_SCAN_IN), .C2(n18741), .A(
        n20850), .B(n18740), .ZN(n18742) );
  OAI22_X1 U21864 ( .A1(n18749), .A2(n18742), .B1(n18875), .B2(n18882), .ZN(
        P3_U3030) );
  NAND2_X1 U21865 ( .A1(n20855), .A2(NA), .ZN(n18743) );
  AOI21_X1 U21866 ( .B1(n20849), .B2(n18743), .A(n20850), .ZN(n18748) );
  NAND2_X1 U21867 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n20851) );
  INV_X1 U21868 ( .A(n20851), .ZN(n18746) );
  OAI22_X1 U21869 ( .A1(NA), .A2(n18744), .B1(P3_STATE_REG_1__SCAN_IN), .B2(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18745) );
  OAI22_X1 U21870 ( .A1(n18746), .A2(n18745), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18747) );
  OAI22_X1 U21871 ( .A1(n18748), .A2(n20848), .B1(n20849), .B2(n18747), .ZN(
        P3_U3031) );
  INV_X1 U21872 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18751) );
  NAND2_X2 U21873 ( .A1(n18864), .A2(n20848), .ZN(n18809) );
  OAI222_X1 U21874 ( .A1(n18855), .A2(n18801), .B1(n18750), .B2(n18864), .C1(
        n18751), .C2(n18809), .ZN(P3_U3032) );
  OAI222_X1 U21875 ( .A1(n18809), .A2(n18754), .B1(n18752), .B2(n18864), .C1(
        n18751), .C2(n18801), .ZN(P3_U3033) );
  OAI222_X1 U21876 ( .A1(n18754), .A2(n18801), .B1(n18753), .B2(n18864), .C1(
        n18755), .C2(n18809), .ZN(P3_U3034) );
  INV_X1 U21877 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18758) );
  OAI222_X1 U21878 ( .A1(n18809), .A2(n18758), .B1(n18756), .B2(n18864), .C1(
        n18755), .C2(n18801), .ZN(P3_U3035) );
  OAI222_X1 U21879 ( .A1(n18758), .A2(n18801), .B1(n18757), .B2(n18864), .C1(
        n18759), .C2(n18809), .ZN(P3_U3036) );
  OAI222_X1 U21880 ( .A1(n18809), .A2(n18761), .B1(n18760), .B2(n18864), .C1(
        n18759), .C2(n18801), .ZN(P3_U3037) );
  OAI222_X1 U21881 ( .A1(n18809), .A2(n18764), .B1(n18762), .B2(n18864), .C1(
        n18761), .C2(n18801), .ZN(P3_U3038) );
  OAI222_X1 U21882 ( .A1(n18764), .A2(n18801), .B1(n18763), .B2(n18864), .C1(
        n18765), .C2(n18809), .ZN(P3_U3039) );
  OAI222_X1 U21883 ( .A1(n18809), .A2(n18767), .B1(n18766), .B2(n18864), .C1(
        n18765), .C2(n18801), .ZN(P3_U3040) );
  OAI222_X1 U21884 ( .A1(n18809), .A2(n18769), .B1(n18768), .B2(n18864), .C1(
        n18767), .C2(n18801), .ZN(P3_U3041) );
  OAI222_X1 U21885 ( .A1(n18809), .A2(n18771), .B1(n18770), .B2(n18864), .C1(
        n18769), .C2(n18801), .ZN(P3_U3042) );
  INV_X1 U21886 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18773) );
  OAI222_X1 U21887 ( .A1(n18809), .A2(n18773), .B1(n18772), .B2(n18864), .C1(
        n18771), .C2(n18801), .ZN(P3_U3043) );
  OAI222_X1 U21888 ( .A1(n18809), .A2(n18776), .B1(n18774), .B2(n18864), .C1(
        n18773), .C2(n18801), .ZN(P3_U3044) );
  OAI222_X1 U21889 ( .A1(n18776), .A2(n18801), .B1(n18775), .B2(n18864), .C1(
        n18777), .C2(n18809), .ZN(P3_U3045) );
  INV_X1 U21890 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18779) );
  OAI222_X1 U21891 ( .A1(n18809), .A2(n18779), .B1(n18778), .B2(n18864), .C1(
        n18777), .C2(n18801), .ZN(P3_U3046) );
  OAI222_X1 U21892 ( .A1(n18809), .A2(n18781), .B1(n18780), .B2(n18864), .C1(
        n18779), .C2(n18801), .ZN(P3_U3047) );
  OAI222_X1 U21893 ( .A1(n18809), .A2(n18783), .B1(n18782), .B2(n18864), .C1(
        n18781), .C2(n18801), .ZN(P3_U3048) );
  OAI222_X1 U21894 ( .A1(n18809), .A2(n18785), .B1(n18784), .B2(n18864), .C1(
        n18783), .C2(n18801), .ZN(P3_U3049) );
  INV_X1 U21895 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18788) );
  OAI222_X1 U21896 ( .A1(n18809), .A2(n18788), .B1(n18786), .B2(n18864), .C1(
        n18785), .C2(n18801), .ZN(P3_U3050) );
  OAI222_X1 U21897 ( .A1(n18788), .A2(n18801), .B1(n18787), .B2(n18864), .C1(
        n18790), .C2(n18809), .ZN(P3_U3051) );
  INV_X1 U21898 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18791) );
  OAI222_X1 U21899 ( .A1(n18790), .A2(n18801), .B1(n18789), .B2(n18864), .C1(
        n18791), .C2(n18809), .ZN(P3_U3052) );
  OAI222_X1 U21900 ( .A1(n18809), .A2(n18794), .B1(n18792), .B2(n18864), .C1(
        n18791), .C2(n18801), .ZN(P3_U3053) );
  OAI222_X1 U21901 ( .A1(n18794), .A2(n18801), .B1(n18793), .B2(n18864), .C1(
        n18795), .C2(n18809), .ZN(P3_U3054) );
  OAI222_X1 U21902 ( .A1(n18809), .A2(n20971), .B1(n18796), .B2(n18864), .C1(
        n18795), .C2(n18801), .ZN(P3_U3055) );
  INV_X1 U21903 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n20942) );
  OAI222_X1 U21904 ( .A1(n18809), .A2(n20942), .B1(n18797), .B2(n18864), .C1(
        n20971), .C2(n18801), .ZN(P3_U3056) );
  OAI222_X1 U21905 ( .A1(n18809), .A2(n18800), .B1(n18798), .B2(n18864), .C1(
        n20942), .C2(n18801), .ZN(P3_U3057) );
  INV_X1 U21906 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18802) );
  OAI222_X1 U21907 ( .A1(n18801), .A2(n18800), .B1(n18799), .B2(n18864), .C1(
        n18802), .C2(n18809), .ZN(P3_U3058) );
  OAI222_X1 U21908 ( .A1(n18809), .A2(n18804), .B1(n18803), .B2(n18864), .C1(
        n18802), .C2(n18801), .ZN(P3_U3059) );
  OAI222_X1 U21909 ( .A1(n18809), .A2(n18806), .B1(n18805), .B2(n18864), .C1(
        n18804), .C2(n18801), .ZN(P3_U3060) );
  OAI222_X1 U21910 ( .A1(n18809), .A2(n18808), .B1(n18807), .B2(n18864), .C1(
        n18806), .C2(n18801), .ZN(P3_U3061) );
  INV_X1 U21911 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n18810) );
  AOI22_X1 U21912 ( .A1(n18864), .A2(n18811), .B1(n18810), .B2(n18882), .ZN(
        P3_U3274) );
  INV_X1 U21913 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18857) );
  INV_X1 U21914 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n18812) );
  AOI22_X1 U21915 ( .A1(n18864), .A2(n18857), .B1(n18812), .B2(n18882), .ZN(
        P3_U3275) );
  INV_X1 U21916 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n18813) );
  AOI22_X1 U21917 ( .A1(n18864), .A2(n18814), .B1(n18813), .B2(n18882), .ZN(
        P3_U3276) );
  INV_X1 U21918 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18862) );
  INV_X1 U21919 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n18815) );
  AOI22_X1 U21920 ( .A1(n18864), .A2(n18862), .B1(n18815), .B2(n18882), .ZN(
        P3_U3277) );
  INV_X1 U21921 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18817) );
  INV_X1 U21922 ( .A(n18819), .ZN(n18816) );
  AOI21_X1 U21923 ( .B1(n18818), .B2(n18817), .A(n18816), .ZN(P3_U3280) );
  OAI21_X1 U21924 ( .B1(n18821), .B2(n18820), .A(n18819), .ZN(P3_U3281) );
  OAI221_X1 U21925 ( .B1(n18824), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18824), 
        .C2(n18823), .A(n18822), .ZN(P3_U3282) );
  INV_X1 U21926 ( .A(n18854), .ZN(n18852) );
  OAI21_X1 U21927 ( .B1(n18825), .B2(n18837), .A(n18852), .ZN(n18831) );
  INV_X1 U21928 ( .A(n18837), .ZN(n18889) );
  NAND2_X1 U21929 ( .A1(n18889), .A2(n18826), .ZN(n18828) );
  OAI22_X1 U21930 ( .A1(n18829), .A2(n18828), .B1(n18836), .B2(n18827), .ZN(
        n18830) );
  AOI22_X1 U21931 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18831), .B1(
        n18852), .B2(n18830), .ZN(n18832) );
  INV_X1 U21932 ( .A(n18832), .ZN(P3_U3285) );
  AOI22_X1 U21933 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n18833), .B2(n15608), .ZN(
        n18842) );
  NOR2_X1 U21934 ( .A1(n18834), .A2(n18851), .ZN(n18843) );
  OAI22_X1 U21935 ( .A1(n18838), .A2(n18837), .B1(n18836), .B2(n18835), .ZN(
        n18839) );
  AOI21_X1 U21936 ( .B1(n18842), .B2(n18843), .A(n18839), .ZN(n18840) );
  AOI22_X1 U21937 ( .A1(n18854), .A2(n13018), .B1(n18840), .B2(n18852), .ZN(
        P3_U3288) );
  INV_X1 U21938 ( .A(n18841), .ZN(n18845) );
  INV_X1 U21939 ( .A(n18842), .ZN(n18844) );
  AOI222_X1 U21940 ( .A1(n18846), .A2(n18889), .B1(n18849), .B2(n18845), .C1(
        n18844), .C2(n18843), .ZN(n18847) );
  AOI22_X1 U21941 ( .A1(n18854), .A2(n18848), .B1(n18847), .B2(n18852), .ZN(
        P3_U3289) );
  AOI222_X1 U21942 ( .A1(n18851), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18889), 
        .B2(n18850), .C1(n12916), .C2(n18849), .ZN(n18853) );
  AOI22_X1 U21943 ( .A1(n18854), .A2(n12916), .B1(n18853), .B2(n18852), .ZN(
        P3_U3290) );
  AOI21_X1 U21944 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18856) );
  AOI22_X1 U21945 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18856), .B2(n18855), .ZN(n18858) );
  AOI22_X1 U21946 ( .A1(n18859), .A2(n18858), .B1(n18857), .B2(n18861), .ZN(
        P3_U3292) );
  NOR2_X1 U21947 ( .A1(n18861), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18860) );
  AOI22_X1 U21948 ( .A1(n18862), .A2(n18861), .B1(n20867), .B2(n18860), .ZN(
        P3_U3293) );
  INV_X1 U21949 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18863) );
  AOI22_X1 U21950 ( .A1(n18864), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18863), 
        .B2(n18882), .ZN(P3_U3294) );
  MUX2_X1 U21951 ( .A(P3_MORE_REG_SCAN_IN), .B(n18866), .S(n18865), .Z(
        P3_U3295) );
  OAI22_X1 U21952 ( .A1(n18870), .A2(n18869), .B1(n18868), .B2(n18867), .ZN(
        n18871) );
  NOR2_X1 U21953 ( .A1(n18887), .A2(n18871), .ZN(n18881) );
  AOI21_X1 U21954 ( .B1(n18874), .B2(n18873), .A(n18872), .ZN(n18876) );
  OAI211_X1 U21955 ( .C1(n18876), .C2(n18884), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n18875), .ZN(n18878) );
  AOI21_X1 U21956 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18878), .A(n18877), 
        .ZN(n18880) );
  NAND2_X1 U21957 ( .A1(n18881), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n18879) );
  OAI21_X1 U21958 ( .B1(n18881), .B2(n18880), .A(n18879), .ZN(P3_U3296) );
  INV_X1 U21959 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n20986) );
  INV_X1 U21960 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n18883) );
  AOI22_X1 U21961 ( .A1(n18864), .A2(n20986), .B1(n18883), .B2(n18882), .ZN(
        P3_U3297) );
  AOI21_X1 U21962 ( .B1(n18889), .B2(n18888), .A(P3_READREQUEST_REG_SCAN_IN), 
        .ZN(n18886) );
  AOI22_X1 U21963 ( .A1(n18887), .A2(n9977), .B1(n18886), .B2(n18885), .ZN(
        P3_U3298) );
  AOI211_X1 U21964 ( .C1(n18889), .C2(n18888), .A(n18887), .B(
        P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18890) );
  NOR2_X1 U21965 ( .A1(n18891), .A2(n18890), .ZN(P3_U3299) );
  INV_X1 U21966 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n18897) );
  INV_X1 U21967 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n18892) );
  NAND2_X1 U21968 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19792), .ZN(n19782) );
  NAND2_X1 U21969 ( .A1(n18897), .A2(n18896), .ZN(n19779) );
  OAI21_X1 U21970 ( .B1(n18897), .B2(n19782), .A(n19779), .ZN(n19849) );
  OAI21_X1 U21971 ( .B1(n18897), .B2(n18892), .A(n19772), .ZN(P2_U2815) );
  INV_X1 U21972 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n20897) );
  OAI22_X1 U21973 ( .A1(n18895), .A2(n20897), .B1(n18894), .B2(n18893), .ZN(
        P2_U2816) );
  OR2_X1 U21974 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n18896), .ZN(n19888) );
  INV_X2 U21975 ( .A(n19888), .ZN(n19891) );
  AOI21_X1 U21976 ( .B1(n18897), .B2(n19792), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n18898) );
  AOI22_X1 U21977 ( .A1(n19891), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n18898), 
        .B2(n19888), .ZN(P2_U2817) );
  OAI21_X1 U21978 ( .B1(n19773), .B2(BS16), .A(n19849), .ZN(n19847) );
  OAI21_X1 U21979 ( .B1(n19849), .B2(n19420), .A(n19847), .ZN(P2_U2818) );
  OAI21_X1 U21980 ( .B1(n18900), .B2(n10762), .A(n18899), .ZN(P2_U2819) );
  NOR4_X1 U21981 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18904) );
  NOR4_X1 U21982 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18903) );
  NOR4_X1 U21983 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_30__SCAN_IN), .ZN(n18902) );
  NOR4_X1 U21984 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n18901) );
  NAND4_X1 U21985 ( .A1(n18904), .A2(n18903), .A3(n18902), .A4(n18901), .ZN(
        n18910) );
  NOR4_X1 U21986 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18908) );
  AOI211_X1 U21987 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_31__SCAN_IN), .B(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18907) );
  NOR4_X1 U21988 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18906) );
  NOR4_X1 U21989 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18905) );
  NAND4_X1 U21990 ( .A1(n18908), .A2(n18907), .A3(n18906), .A4(n18905), .ZN(
        n18909) );
  NOR2_X1 U21991 ( .A1(n18910), .A2(n18909), .ZN(n18918) );
  INV_X1 U21992 ( .A(n18918), .ZN(n18917) );
  NOR2_X1 U21993 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18917), .ZN(n18911) );
  INV_X1 U21994 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19845) );
  AOI22_X1 U21995 ( .A1(n18911), .A2(n18912), .B1(n18917), .B2(n19845), .ZN(
        P2_U2820) );
  OR3_X1 U21996 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18916) );
  INV_X1 U21997 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19843) );
  AOI22_X1 U21998 ( .A1(n18911), .A2(n18916), .B1(n18917), .B2(n19843), .ZN(
        P2_U2821) );
  INV_X1 U21999 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19848) );
  NAND2_X1 U22000 ( .A1(n18911), .A2(n19848), .ZN(n18915) );
  OAI21_X1 U22001 ( .B1(n19793), .B2(n18912), .A(n18918), .ZN(n18913) );
  OAI21_X1 U22002 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18918), .A(n18913), 
        .ZN(n18914) );
  OAI221_X1 U22003 ( .B1(n18915), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18915), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18914), .ZN(P2_U2822) );
  INV_X1 U22004 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19841) );
  OAI221_X1 U22005 ( .B1(n18918), .B2(n19841), .C1(n18917), .C2(n18916), .A(
        n18915), .ZN(P2_U2823) );
  AOI21_X1 U22006 ( .B1(n18923), .B2(n18920), .A(n18919), .ZN(n18921) );
  AOI21_X1 U22007 ( .B1(n19060), .B2(n18922), .A(n18921), .ZN(n18930) );
  AOI22_X1 U22008 ( .A1(P2_REIP_REG_20__SCAN_IN), .A2(n9882), .B1(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n19024), .ZN(n18929) );
  AOI22_X1 U22009 ( .A1(P2_EBX_REG_20__SCAN_IN), .A2(n19054), .B1(n18923), 
        .B2(n19055), .ZN(n18928) );
  INV_X1 U22010 ( .A(n18924), .ZN(n18925) );
  AOI22_X1 U22011 ( .A1(n18980), .A2(n18926), .B1(n18925), .B2(n19066), .ZN(
        n18927) );
  NAND4_X1 U22012 ( .A1(n18930), .A2(n18929), .A3(n18928), .A4(n18927), .ZN(
        P2_U2835) );
  OAI21_X1 U22013 ( .B1(n10873), .B2(n9807), .A(n18957), .ZN(n18934) );
  INV_X1 U22014 ( .A(n18931), .ZN(n18932) );
  OAI22_X1 U22015 ( .A1(n18932), .A2(n19042), .B1(n21034), .B2(n19057), .ZN(
        n18933) );
  AOI211_X1 U22016 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n19054), .A(n18934), .B(
        n18933), .ZN(n18942) );
  NOR2_X1 U22017 ( .A1(n14704), .A2(n18935), .ZN(n18937) );
  XNOR2_X1 U22018 ( .A(n18937), .B(n18936), .ZN(n18940) );
  AOI22_X1 U22019 ( .A1(n18940), .A2(n18939), .B1(n18938), .B2(n19066), .ZN(
        n18941) );
  OAI211_X1 U22020 ( .C1(n18943), .C2(n19063), .A(n18942), .B(n18941), .ZN(
        P2_U2836) );
  NAND2_X1 U22021 ( .A1(n19032), .A2(n18944), .ZN(n18965) );
  XNOR2_X1 U22022 ( .A(n18945), .B(n18965), .ZN(n18954) );
  AOI222_X1 U22023 ( .A1(n18946), .A2(n19060), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n19054), .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n19024), .ZN(
        n18947) );
  INV_X1 U22024 ( .A(n18947), .ZN(n18948) );
  AOI211_X1 U22025 ( .C1(P2_REIP_REG_18__SCAN_IN), .C2(n9882), .A(n19030), .B(
        n18948), .ZN(n18953) );
  INV_X1 U22026 ( .A(n18949), .ZN(n18950) );
  AOI22_X1 U22027 ( .A1(n18980), .A2(n18951), .B1(n18950), .B2(n19066), .ZN(
        n18952) );
  OAI211_X1 U22028 ( .C1(n19771), .C2(n18954), .A(n18953), .B(n18952), .ZN(
        P2_U2837) );
  INV_X1 U22029 ( .A(n18955), .ZN(n18964) );
  INV_X1 U22030 ( .A(n18967), .ZN(n18961) );
  INV_X1 U22031 ( .A(n18956), .ZN(n18959) );
  AOI22_X1 U22032 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19024), .B1(
        P2_EBX_REG_17__SCAN_IN), .B2(n19054), .ZN(n18958) );
  OAI211_X1 U22033 ( .C1(n18959), .C2(n19036), .A(n18958), .B(n18957), .ZN(
        n18960) );
  AOI21_X1 U22034 ( .B1(n19055), .B2(n18961), .A(n18960), .ZN(n18962) );
  OAI21_X1 U22035 ( .B1(n9807), .B2(n19818), .A(n18962), .ZN(n18963) );
  AOI21_X1 U22036 ( .B1(n18964), .B2(n19060), .A(n18963), .ZN(n18970) );
  INV_X1 U22037 ( .A(n18965), .ZN(n18966) );
  OAI211_X1 U22038 ( .C1(n18968), .C2(n18967), .A(n19050), .B(n18966), .ZN(
        n18969) );
  OAI211_X1 U22039 ( .C1(n19063), .C2(n18971), .A(n18970), .B(n18969), .ZN(
        P2_U2838) );
  NAND2_X1 U22040 ( .A1(n19032), .A2(n18972), .ZN(n18973) );
  XOR2_X1 U22041 ( .A(n18974), .B(n18973), .Z(n18983) );
  OAI21_X1 U22042 ( .B1(n19816), .B2(n9807), .A(n15334), .ZN(n18978) );
  OAI22_X1 U22043 ( .A1(n18976), .A2(n19042), .B1(n18975), .B2(n19057), .ZN(
        n18977) );
  AOI211_X1 U22044 ( .C1(P2_EBX_REG_16__SCAN_IN), .C2(n19054), .A(n18978), .B(
        n18977), .ZN(n18982) );
  AOI22_X1 U22045 ( .A1(n19079), .A2(n18980), .B1(n18979), .B2(n19066), .ZN(
        n18981) );
  OAI211_X1 U22046 ( .C1(n19771), .C2(n18983), .A(n18982), .B(n18981), .ZN(
        P2_U2839) );
  OAI22_X1 U22047 ( .A1(n18984), .A2(n19042), .B1(n10861), .B2(n19028), .ZN(
        n18985) );
  AOI211_X1 U22048 ( .C1(P2_REIP_REG_15__SCAN_IN), .C2(n9882), .A(n19030), .B(
        n18985), .ZN(n18993) );
  NOR2_X1 U22049 ( .A1(n14704), .A2(n18986), .ZN(n18987) );
  XNOR2_X1 U22050 ( .A(n18988), .B(n18987), .ZN(n18991) );
  OAI22_X1 U22051 ( .A1(n19086), .A2(n19063), .B1(n18989), .B2(n19036), .ZN(
        n18990) );
  AOI21_X1 U22052 ( .B1(n18991), .B2(n19050), .A(n18990), .ZN(n18992) );
  OAI211_X1 U22053 ( .C1(n18994), .C2(n19057), .A(n18993), .B(n18992), .ZN(
        P2_U2840) );
  NOR2_X1 U22054 ( .A1(n14704), .A2(n18995), .ZN(n18996) );
  XNOR2_X1 U22055 ( .A(n18997), .B(n18996), .ZN(n19005) );
  AOI22_X1 U22056 ( .A1(n18998), .A2(n19060), .B1(P2_EBX_REG_11__SCAN_IN), 
        .B2(n19054), .ZN(n18999) );
  OAI211_X1 U22057 ( .C1(n15101), .C2(n9807), .A(n18999), .B(n18957), .ZN(
        n19002) );
  OAI22_X1 U22058 ( .A1(n19000), .A2(n19036), .B1(n19063), .B2(n19098), .ZN(
        n19001) );
  AOI211_X1 U22059 ( .C1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n19003), .A(
        n19002), .B(n19001), .ZN(n19004) );
  OAI21_X1 U22060 ( .B1(n19771), .B2(n19005), .A(n19004), .ZN(P2_U2844) );
  NOR2_X1 U22061 ( .A1(n14704), .A2(n19006), .ZN(n19008) );
  XNOR2_X1 U22062 ( .A(n19008), .B(n19007), .ZN(n19015) );
  AOI22_X1 U22063 ( .A1(n19009), .A2(n19060), .B1(P2_EBX_REG_9__SCAN_IN), .B2(
        n19054), .ZN(n19010) );
  OAI211_X1 U22064 ( .C1(n19807), .C2(n9807), .A(n19010), .B(n15334), .ZN(
        n19013) );
  OAI22_X1 U22065 ( .A1(n19105), .A2(n19063), .B1(n19036), .B2(n19011), .ZN(
        n19012) );
  AOI211_X1 U22066 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n19024), .A(
        n19013), .B(n19012), .ZN(n19014) );
  OAI21_X1 U22067 ( .B1(n19771), .B2(n19015), .A(n19014), .ZN(P2_U2846) );
  NOR2_X1 U22068 ( .A1(n14704), .A2(n19016), .ZN(n19017) );
  XOR2_X1 U22069 ( .A(n19018), .B(n19017), .Z(n19026) );
  AOI22_X1 U22070 ( .A1(n19019), .A2(n19060), .B1(P2_EBX_REG_7__SCAN_IN), .B2(
        n19054), .ZN(n19020) );
  OAI211_X1 U22071 ( .C1(n19803), .C2(n9807), .A(n19020), .B(n18957), .ZN(
        n19023) );
  OAI22_X1 U22072 ( .A1(n19108), .A2(n19063), .B1(n19036), .B2(n19021), .ZN(
        n19022) );
  AOI211_X1 U22073 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19024), .A(
        n19023), .B(n19022), .ZN(n19025) );
  OAI21_X1 U22074 ( .B1(n19771), .B2(n19026), .A(n19025), .ZN(P2_U2848) );
  OAI22_X1 U22075 ( .A1(n20987), .A2(n19028), .B1(n19027), .B2(n19042), .ZN(
        n19029) );
  AOI211_X1 U22076 ( .C1(P2_REIP_REG_6__SCAN_IN), .C2(n9882), .A(n19030), .B(
        n19029), .ZN(n19040) );
  NAND2_X1 U22077 ( .A1(n19032), .A2(n19031), .ZN(n19033) );
  XNOR2_X1 U22078 ( .A(n19034), .B(n19033), .ZN(n19038) );
  OAI22_X1 U22079 ( .A1(n19109), .A2(n19063), .B1(n19036), .B2(n19035), .ZN(
        n19037) );
  AOI21_X1 U22080 ( .B1(n19050), .B2(n19038), .A(n19037), .ZN(n19039) );
  OAI211_X1 U22081 ( .C1(n19041), .C2(n19057), .A(n19040), .B(n19039), .ZN(
        P2_U2849) );
  OAI21_X1 U22082 ( .B1(n13857), .B2(n9807), .A(n18957), .ZN(n19045) );
  OAI22_X1 U22083 ( .A1(n19043), .A2(n19042), .B1(n10071), .B2(n19057), .ZN(
        n19044) );
  AOI211_X1 U22084 ( .C1(P2_EBX_REG_5__SCAN_IN), .C2(n19054), .A(n19045), .B(
        n19044), .ZN(n19053) );
  NOR2_X1 U22085 ( .A1(n14704), .A2(n19046), .ZN(n19048) );
  XNOR2_X1 U22086 ( .A(n19048), .B(n19047), .ZN(n19051) );
  AOI22_X1 U22087 ( .A1(n19051), .A2(n19050), .B1(n19066), .B2(n19049), .ZN(
        n19052) );
  OAI211_X1 U22088 ( .C1(n19063), .C2(n19117), .A(n19053), .B(n19052), .ZN(
        P2_U2850) );
  NAND2_X1 U22089 ( .A1(n19054), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n19062) );
  INV_X1 U22090 ( .A(n19055), .ZN(n19056) );
  INV_X1 U22091 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n20970) );
  AOI21_X1 U22092 ( .B1(n19057), .B2(n19056), .A(n20970), .ZN(n19058) );
  AOI21_X1 U22093 ( .B1(n19060), .B2(n19059), .A(n19058), .ZN(n19061) );
  OAI211_X1 U22094 ( .C1(n19064), .C2(n19063), .A(n19062), .B(n19061), .ZN(
        n19065) );
  AOI21_X1 U22095 ( .B1(n13216), .B2(n19066), .A(n19065), .ZN(n19067) );
  OAI21_X1 U22096 ( .B1(n19068), .B2(n19881), .A(n19067), .ZN(n19069) );
  AOI21_X1 U22097 ( .B1(n9882), .B2(P2_REIP_REG_0__SCAN_IN), .A(n19069), .ZN(
        n19070) );
  OAI21_X1 U22098 ( .B1(n19072), .B2(n19071), .A(n19070), .ZN(P2_U2855) );
  AOI22_X1 U22099 ( .A1(n19127), .A2(n16116), .B1(n19077), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n19074) );
  AOI22_X1 U22100 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19126), .B1(n19078), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n19073) );
  NAND2_X1 U22101 ( .A1(n19074), .A2(n19073), .ZN(P2_U2888) );
  AOI22_X1 U22102 ( .A1(n19076), .A2(n19075), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n19126), .ZN(n19083) );
  AOI22_X1 U22103 ( .A1(n19078), .A2(BUF1_REG_16__SCAN_IN), .B1(n19077), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n19082) );
  AOI22_X1 U22104 ( .A1(n19080), .A2(n19131), .B1(n19127), .B2(n19079), .ZN(
        n19081) );
  NAND3_X1 U22105 ( .A1(n19083), .A2(n19082), .A3(n19081), .ZN(P2_U2903) );
  OAI222_X1 U22106 ( .A1(n19086), .A2(n19118), .B1(n13053), .B2(n19110), .C1(
        n19085), .C2(n19135), .ZN(P2_U2904) );
  INV_X1 U22107 ( .A(n19087), .ZN(n19090) );
  AOI22_X1 U22108 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19126), .B1(n19088), 
        .B2(n19102), .ZN(n19089) );
  OAI21_X1 U22109 ( .B1(n19118), .B2(n19090), .A(n19089), .ZN(P2_U2905) );
  INV_X1 U22110 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19173) );
  OAI222_X1 U22111 ( .A1(n19092), .A2(n19118), .B1(n19173), .B2(n19110), .C1(
        n19135), .C2(n19091), .ZN(P2_U2906) );
  INV_X1 U22112 ( .A(n19093), .ZN(n19096) );
  AOI22_X1 U22113 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n19126), .B1(n19094), 
        .B2(n19102), .ZN(n19095) );
  OAI21_X1 U22114 ( .B1(n19118), .B2(n19096), .A(n19095), .ZN(P2_U2907) );
  INV_X1 U22115 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19177) );
  OAI222_X1 U22116 ( .A1(n19098), .A2(n19118), .B1(n19177), .B2(n19110), .C1(
        n19135), .C2(n19097), .ZN(P2_U2908) );
  AOI22_X1 U22117 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19126), .B1(n19099), 
        .B2(n19102), .ZN(n19100) );
  OAI21_X1 U22118 ( .B1(n19118), .B2(n19101), .A(n19100), .ZN(P2_U2909) );
  AOI22_X1 U22119 ( .A1(P2_EAX_REG_9__SCAN_IN), .A2(n19126), .B1(n19103), .B2(
        n19102), .ZN(n19104) );
  OAI21_X1 U22120 ( .B1(n19118), .B2(n19105), .A(n19104), .ZN(P2_U2910) );
  INV_X1 U22121 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19183) );
  OAI222_X1 U22122 ( .A1(n19107), .A2(n19118), .B1(n19183), .B2(n19110), .C1(
        n19135), .C2(n19106), .ZN(P2_U2911) );
  OAI222_X1 U22123 ( .A1(n19108), .A2(n19118), .B1(n19185), .B2(n19110), .C1(
        n19135), .C2(n19281), .ZN(P2_U2912) );
  INV_X1 U22124 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19188) );
  OAI222_X1 U22125 ( .A1(n19109), .A2(n19118), .B1(n19188), .B2(n19110), .C1(
        n19135), .C2(n19271), .ZN(P2_U2913) );
  INV_X1 U22126 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19190) );
  OAI22_X1 U22127 ( .A1(n19190), .A2(n19110), .B1(n19266), .B2(n19135), .ZN(
        n19111) );
  INV_X1 U22128 ( .A(n19111), .ZN(n19116) );
  OR3_X1 U22129 ( .A1(n19114), .A2(n19113), .A3(n19112), .ZN(n19115) );
  OAI211_X1 U22130 ( .C1(n19118), .C2(n19117), .A(n19116), .B(n19115), .ZN(
        P2_U2914) );
  INV_X1 U22131 ( .A(n19119), .ZN(n19857) );
  AOI22_X1 U22132 ( .A1(n19857), .A2(n19127), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19126), .ZN(n19125) );
  OAI21_X1 U22133 ( .B1(n19122), .B2(n19121), .A(n19120), .ZN(n19123) );
  NAND2_X1 U22134 ( .A1(n19123), .A2(n19131), .ZN(n19124) );
  OAI211_X1 U22135 ( .C1(n19254), .C2(n19135), .A(n19125), .B(n19124), .ZN(
        P2_U2916) );
  AOI22_X1 U22136 ( .A1(n19127), .A2(n19875), .B1(n19126), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19134) );
  OAI21_X1 U22137 ( .B1(n19130), .B2(n19129), .A(n19128), .ZN(n19132) );
  NAND2_X1 U22138 ( .A1(n19132), .A2(n19131), .ZN(n19133) );
  OAI211_X1 U22139 ( .C1(n19248), .C2(n19135), .A(n19134), .B(n19133), .ZN(
        P2_U2918) );
  OAI21_X1 U22140 ( .B1(n19138), .B2(n19137), .A(n19136), .ZN(n19139) );
  NOR2_X4 U22141 ( .A1(n19169), .A2(n19178), .ZN(n19186) );
  AND2_X1 U22142 ( .A1(n19186), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  AOI22_X1 U22143 ( .A1(n19178), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19186), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n19141) );
  OAI21_X1 U22144 ( .B1(n12894), .B2(n19167), .A(n19141), .ZN(P2_U2921) );
  AOI22_X1 U22145 ( .A1(n19178), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19186), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n19142) );
  OAI21_X1 U22146 ( .B1(n19143), .B2(n19167), .A(n19142), .ZN(P2_U2922) );
  AOI22_X1 U22147 ( .A1(n19178), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19186), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n19144) );
  OAI21_X1 U22148 ( .B1(n20973), .B2(n19167), .A(n19144), .ZN(P2_U2923) );
  AOI22_X1 U22149 ( .A1(n19178), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19186), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n19145) );
  OAI21_X1 U22150 ( .B1(n19146), .B2(n19167), .A(n19145), .ZN(P2_U2924) );
  AOI22_X1 U22151 ( .A1(n19178), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19186), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n19147) );
  OAI21_X1 U22152 ( .B1(n20984), .B2(n19167), .A(n19147), .ZN(P2_U2925) );
  AOI22_X1 U22153 ( .A1(n19178), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19186), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n19148) );
  OAI21_X1 U22154 ( .B1(n19149), .B2(n19167), .A(n19148), .ZN(P2_U2926) );
  AOI22_X1 U22155 ( .A1(n19178), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19186), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n19150) );
  OAI21_X1 U22156 ( .B1(n19151), .B2(n19167), .A(n19150), .ZN(P2_U2927) );
  AOI22_X1 U22157 ( .A1(n19178), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19186), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n19152) );
  OAI21_X1 U22158 ( .B1(n19153), .B2(n19167), .A(n19152), .ZN(P2_U2928) );
  INV_X1 U22159 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n19155) );
  AOI22_X1 U22160 ( .A1(n19178), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19186), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n19154) );
  OAI21_X1 U22161 ( .B1(n19155), .B2(n19167), .A(n19154), .ZN(P2_U2929) );
  AOI22_X1 U22162 ( .A1(n19178), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19186), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n19156) );
  OAI21_X1 U22163 ( .B1(n19157), .B2(n19167), .A(n19156), .ZN(P2_U2930) );
  INV_X1 U22164 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n19159) );
  AOI22_X1 U22165 ( .A1(n19178), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19186), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n19158) );
  OAI21_X1 U22166 ( .B1(n19159), .B2(n19167), .A(n19158), .ZN(P2_U2931) );
  AOI22_X1 U22167 ( .A1(n19178), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19186), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n19160) );
  OAI21_X1 U22168 ( .B1(n19161), .B2(n19167), .A(n19160), .ZN(P2_U2932) );
  INV_X1 U22169 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n19163) );
  AOI22_X1 U22170 ( .A1(n19178), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19186), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n19162) );
  OAI21_X1 U22171 ( .B1(n19163), .B2(n19167), .A(n19162), .ZN(P2_U2933) );
  AOI22_X1 U22172 ( .A1(n19178), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19186), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n19164) );
  OAI21_X1 U22173 ( .B1(n19165), .B2(n19167), .A(n19164), .ZN(P2_U2934) );
  AOI22_X1 U22174 ( .A1(n19178), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19186), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n19166) );
  OAI21_X1 U22175 ( .B1(n19168), .B2(n19167), .A(n19166), .ZN(P2_U2935) );
  AOI22_X1 U22176 ( .A1(n19178), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19186), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19170) );
  OAI21_X1 U22177 ( .B1(n13053), .B2(n19201), .A(n19170), .ZN(P2_U2936) );
  AOI22_X1 U22178 ( .A1(n19178), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19186), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19171) );
  OAI21_X1 U22179 ( .B1(n11197), .B2(n19201), .A(n19171), .ZN(P2_U2937) );
  AOI22_X1 U22180 ( .A1(n19178), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19186), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19172) );
  OAI21_X1 U22181 ( .B1(n19173), .B2(n19201), .A(n19172), .ZN(P2_U2938) );
  AOI22_X1 U22182 ( .A1(n19178), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19186), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19174) );
  OAI21_X1 U22183 ( .B1(n19175), .B2(n19201), .A(n19174), .ZN(P2_U2939) );
  AOI22_X1 U22184 ( .A1(n19178), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19186), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19176) );
  OAI21_X1 U22185 ( .B1(n19177), .B2(n19201), .A(n19176), .ZN(P2_U2940) );
  AOI22_X1 U22186 ( .A1(n19178), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19186), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19179) );
  OAI21_X1 U22187 ( .B1(n19180), .B2(n19201), .A(n19179), .ZN(P2_U2941) );
  AOI22_X1 U22188 ( .A1(n19199), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19186), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19181) );
  OAI21_X1 U22189 ( .B1(n21066), .B2(n19201), .A(n19181), .ZN(P2_U2942) );
  AOI22_X1 U22190 ( .A1(n19199), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19186), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19182) );
  OAI21_X1 U22191 ( .B1(n19183), .B2(n19201), .A(n19182), .ZN(P2_U2943) );
  AOI22_X1 U22192 ( .A1(n19199), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19186), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19184) );
  OAI21_X1 U22193 ( .B1(n19185), .B2(n19201), .A(n19184), .ZN(P2_U2944) );
  AOI22_X1 U22194 ( .A1(n19199), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19186), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19187) );
  OAI21_X1 U22195 ( .B1(n19188), .B2(n19201), .A(n19187), .ZN(P2_U2945) );
  AOI22_X1 U22196 ( .A1(n19199), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19186), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19189) );
  OAI21_X1 U22197 ( .B1(n19190), .B2(n19201), .A(n19189), .ZN(P2_U2946) );
  INV_X1 U22198 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19192) );
  AOI22_X1 U22199 ( .A1(n19199), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19186), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19191) );
  OAI21_X1 U22200 ( .B1(n19192), .B2(n19201), .A(n19191), .ZN(P2_U2947) );
  INV_X1 U22201 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19194) );
  AOI22_X1 U22202 ( .A1(n19199), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19186), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19193) );
  OAI21_X1 U22203 ( .B1(n19194), .B2(n19201), .A(n19193), .ZN(P2_U2948) );
  INV_X1 U22204 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19196) );
  AOI22_X1 U22205 ( .A1(n19199), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19186), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19195) );
  OAI21_X1 U22206 ( .B1(n19196), .B2(n19201), .A(n19195), .ZN(P2_U2949) );
  INV_X1 U22207 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19198) );
  AOI22_X1 U22208 ( .A1(n19199), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19186), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19197) );
  OAI21_X1 U22209 ( .B1(n19198), .B2(n19201), .A(n19197), .ZN(P2_U2950) );
  AOI22_X1 U22210 ( .A1(n19199), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19186), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19200) );
  OAI21_X1 U22211 ( .B1(n13050), .B2(n19201), .A(n19200), .ZN(P2_U2951) );
  AOI22_X1 U22212 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19030), .B1(n19203), 
        .B2(n19202), .ZN(n19210) );
  AOI222_X1 U22213 ( .A1(n19208), .A2(n11305), .B1(n19207), .B2(n19206), .C1(
        n19205), .C2(n19204), .ZN(n19209) );
  OAI211_X1 U22214 ( .C1(n19212), .C2(n19211), .A(n19210), .B(n19209), .ZN(
        P2_U3010) );
  INV_X1 U22215 ( .A(n19213), .ZN(n19222) );
  NOR2_X1 U22216 ( .A1(n19214), .A2(n19217), .ZN(n19215) );
  AOI211_X1 U22217 ( .C1(n19217), .C2(n19222), .A(n19216), .B(n19215), .ZN(
        n19236) );
  INV_X1 U22218 ( .A(n19218), .ZN(n19231) );
  NOR2_X1 U22219 ( .A1(n18957), .A2(n19795), .ZN(n19219) );
  AOI21_X1 U22220 ( .B1(n19220), .B2(n13265), .A(n19219), .ZN(n19224) );
  NAND3_X1 U22221 ( .A1(n19222), .A2(n19221), .A3(n19235), .ZN(n19223) );
  OAI211_X1 U22222 ( .C1(n19226), .C2(n19225), .A(n19224), .B(n19223), .ZN(
        n19227) );
  AOI21_X1 U22223 ( .B1(n19866), .B2(n19228), .A(n19227), .ZN(n19229) );
  INV_X1 U22224 ( .A(n19229), .ZN(n19230) );
  AOI211_X1 U22225 ( .C1(n19233), .C2(n19232), .A(n19231), .B(n19230), .ZN(
        n19234) );
  OAI21_X1 U22226 ( .B1(n19236), .B2(n19235), .A(n19234), .ZN(P2_U3044) );
  NAND2_X1 U22227 ( .A1(n19347), .A2(n19877), .ZN(n19292) );
  NOR2_X1 U22228 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19292), .ZN(
        n19280) );
  AOI22_X1 U22229 ( .A1(n19677), .A2(n19740), .B1(n19676), .B2(n19280), .ZN(
        n19246) );
  NAND2_X1 U22230 ( .A1(n19856), .A2(n19311), .ZN(n19237) );
  NAND2_X1 U22231 ( .A1(n19856), .A2(n19420), .ZN(n19678) );
  OAI21_X1 U22232 ( .B1(n19740), .B2(n19237), .A(n19678), .ZN(n19241) );
  AOI21_X1 U22233 ( .B1(n19242), .B2(n19680), .A(n19856), .ZN(n19238) );
  AOI21_X1 U22234 ( .B1(n19241), .B2(n19239), .A(n19238), .ZN(n19240) );
  OAI21_X1 U22235 ( .B1(n19752), .B2(n19280), .A(n19241), .ZN(n19244) );
  OAI21_X1 U22236 ( .B1(n19242), .B2(n19280), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19243) );
  NAND2_X1 U22237 ( .A1(n19244), .A2(n19243), .ZN(n19282) );
  AOI22_X1 U22238 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19283), .B1(
        n19690), .B2(n19282), .ZN(n19245) );
  OAI211_X1 U22239 ( .C1(n19693), .C2(n19311), .A(n19246), .B(n19245), .ZN(
        P2_U3048) );
  OAI22_X2 U22240 ( .A1(n13891), .A2(n19277), .B1(n13890), .B2(n19276), .ZN(
        n19720) );
  AOI22_X1 U22241 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19275), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19274), .ZN(n19696) );
  INV_X1 U22242 ( .A(n19696), .ZN(n19719) );
  AOI22_X1 U22243 ( .A1(n19719), .A2(n19740), .B1(n19280), .B2(n19247), .ZN(
        n19250) );
  NOR2_X2 U22244 ( .A1(n19248), .A2(n19424), .ZN(n19718) );
  AOI22_X1 U22245 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19283), .B1(
        n19718), .B2(n19282), .ZN(n19249) );
  OAI211_X1 U22246 ( .C1(n19658), .C2(n19311), .A(n19250), .B(n19249), .ZN(
        P2_U3049) );
  AOI22_X1 U22247 ( .A1(n19620), .A2(n19740), .B1(n19697), .B2(n19280), .ZN(
        n19252) );
  AOI22_X1 U22248 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19283), .B1(
        n19699), .B2(n19282), .ZN(n19251) );
  OAI211_X1 U22249 ( .C1(n19623), .C2(n19311), .A(n19252), .B(n19251), .ZN(
        P2_U3050) );
  AOI22_X1 U22250 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19275), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19274), .ZN(n19730) );
  OAI22_X2 U22251 ( .A1(n19253), .A2(n19276), .B1(n21078), .B2(n19277), .ZN(
        n19727) );
  NOR2_X2 U22252 ( .A1(n10282), .A2(n19278), .ZN(n19725) );
  AOI22_X1 U22253 ( .A1(n19727), .A2(n19740), .B1(n19280), .B2(n19725), .ZN(
        n19256) );
  NOR2_X2 U22254 ( .A1(n19254), .A2(n19424), .ZN(n19726) );
  AOI22_X1 U22255 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19283), .B1(
        n19726), .B2(n19282), .ZN(n19255) );
  OAI211_X1 U22256 ( .C1(n19730), .C2(n19311), .A(n19256), .B(n19255), .ZN(
        P2_U3051) );
  AOI22_X1 U22257 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19275), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19274), .ZN(n19736) );
  OAI22_X2 U22258 ( .A1(n19258), .A2(n19277), .B1(n19257), .B2(n19276), .ZN(
        n19733) );
  NOR2_X2 U22259 ( .A1(n19259), .A2(n19278), .ZN(n19731) );
  AOI22_X1 U22260 ( .A1(n19733), .A2(n19740), .B1(n19280), .B2(n19731), .ZN(
        n19263) );
  INV_X1 U22261 ( .A(n19260), .ZN(n19261) );
  NOR2_X2 U22262 ( .A1(n19261), .A2(n19424), .ZN(n19732) );
  AOI22_X1 U22263 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19283), .B1(
        n19732), .B2(n19282), .ZN(n19262) );
  OAI211_X1 U22264 ( .C1(n19736), .C2(n19311), .A(n19263), .B(n19262), .ZN(
        P2_U3052) );
  AOI22_X1 U22265 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19275), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19274), .ZN(n19631) );
  NOR2_X2 U22266 ( .A1(n19265), .A2(n19278), .ZN(n19737) );
  AOI22_X1 U22267 ( .A1(n19628), .A2(n19740), .B1(n19737), .B2(n19280), .ZN(
        n19268) );
  NOR2_X2 U22268 ( .A1(n19266), .A2(n19424), .ZN(n19738) );
  AOI22_X1 U22269 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19283), .B1(
        n19738), .B2(n19282), .ZN(n19267) );
  OAI211_X1 U22270 ( .C1(n19631), .C2(n19311), .A(n19268), .B(n19267), .ZN(
        P2_U3053) );
  AOI22_X1 U22271 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19275), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19274), .ZN(n19599) );
  INV_X1 U22272 ( .A(n19599), .ZN(n19747) );
  NOR2_X2 U22273 ( .A1(n10251), .A2(n19278), .ZN(n19745) );
  AOI22_X1 U22274 ( .A1(n19747), .A2(n19740), .B1(n19280), .B2(n19745), .ZN(
        n19273) );
  NOR2_X2 U22275 ( .A1(n19271), .A2(n19424), .ZN(n19746) );
  AOI22_X1 U22276 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19283), .B1(
        n19746), .B2(n19282), .ZN(n19272) );
  OAI211_X1 U22277 ( .C1(n19750), .C2(n19311), .A(n19273), .B(n19272), .ZN(
        P2_U3054) );
  AOI22_X2 U22278 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19275), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19274), .ZN(n19761) );
  OAI22_X2 U22279 ( .A1(n20176), .A2(n19277), .B1(n21051), .B2(n19276), .ZN(
        n19755) );
  NOR2_X2 U22280 ( .A1(n19279), .A2(n19278), .ZN(n19751) );
  AOI22_X1 U22281 ( .A1(n19755), .A2(n19740), .B1(n19280), .B2(n19751), .ZN(
        n19285) );
  NOR2_X2 U22282 ( .A1(n19281), .A2(n19424), .ZN(n19753) );
  AOI22_X1 U22283 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19283), .B1(
        n19753), .B2(n19282), .ZN(n19284) );
  OAI211_X1 U22284 ( .C1(n19761), .C2(n19311), .A(n19285), .B(n19284), .ZN(
        P2_U3055) );
  NAND2_X1 U22285 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19877), .ZN(
        n19510) );
  INV_X1 U22286 ( .A(n19347), .ZN(n19345) );
  NOR2_X1 U22287 ( .A1(n19510), .A2(n19345), .ZN(n19309) );
  OR2_X1 U22288 ( .A1(n19309), .A2(n19544), .ZN(n19286) );
  NOR2_X1 U22289 ( .A1(n19287), .A2(n19286), .ZN(n19291) );
  INV_X1 U22290 ( .A(n19292), .ZN(n19288) );
  AOI21_X1 U22291 ( .B1(n19680), .B2(n19288), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19289) );
  AOI22_X1 U22292 ( .A1(n19310), .A2(n19690), .B1(n19676), .B2(n19309), .ZN(
        n19296) );
  INV_X1 U22293 ( .A(n19452), .ZN(n19290) );
  NAND2_X1 U22294 ( .A1(n19290), .A2(n19509), .ZN(n19293) );
  AOI21_X1 U22295 ( .B1(n19293), .B2(n19292), .A(n19291), .ZN(n19294) );
  OAI211_X1 U22296 ( .C1(n19309), .C2(n19680), .A(n19294), .B(n19683), .ZN(
        n19313) );
  NAND2_X1 U22297 ( .A1(n19509), .A2(n19448), .ZN(n19319) );
  AOI22_X1 U22298 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19313), .B1(
        n19341), .B2(n19652), .ZN(n19295) );
  OAI211_X1 U22299 ( .C1(n19655), .C2(n19311), .A(n19296), .B(n19295), .ZN(
        P2_U3056) );
  AOI22_X1 U22300 ( .A1(n19310), .A2(n19718), .B1(n19247), .B2(n19309), .ZN(
        n19298) );
  AOI22_X1 U22301 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19313), .B1(
        n19341), .B2(n19720), .ZN(n19297) );
  OAI211_X1 U22302 ( .C1(n19696), .C2(n19311), .A(n19298), .B(n19297), .ZN(
        P2_U3057) );
  AOI22_X1 U22303 ( .A1(n19310), .A2(n19699), .B1(n19697), .B2(n19309), .ZN(
        n19300) );
  AOI22_X1 U22304 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19313), .B1(
        n19341), .B2(n19698), .ZN(n19299) );
  OAI211_X1 U22305 ( .C1(n19702), .C2(n19311), .A(n19300), .B(n19299), .ZN(
        P2_U3058) );
  AOI22_X1 U22306 ( .A1(n19310), .A2(n19726), .B1(n19725), .B2(n19309), .ZN(
        n19302) );
  INV_X1 U22307 ( .A(n19730), .ZN(n19585) );
  AOI22_X1 U22308 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19313), .B1(
        n19341), .B2(n19585), .ZN(n19301) );
  OAI211_X1 U22309 ( .C1(n19588), .C2(n19311), .A(n19302), .B(n19301), .ZN(
        P2_U3059) );
  AOI22_X1 U22310 ( .A1(n19310), .A2(n19732), .B1(n19731), .B2(n19309), .ZN(
        n19304) );
  INV_X1 U22311 ( .A(n19736), .ZN(n19589) );
  AOI22_X1 U22312 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19313), .B1(
        n19341), .B2(n19589), .ZN(n19303) );
  OAI211_X1 U22313 ( .C1(n19592), .C2(n19311), .A(n19304), .B(n19303), .ZN(
        P2_U3060) );
  AOI22_X1 U22314 ( .A1(n19310), .A2(n19738), .B1(n19737), .B2(n19309), .ZN(
        n19306) );
  AOI22_X1 U22315 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19313), .B1(
        n19341), .B2(n19739), .ZN(n19305) );
  OAI211_X1 U22316 ( .C1(n19744), .C2(n19311), .A(n19306), .B(n19305), .ZN(
        P2_U3061) );
  AOI22_X1 U22317 ( .A1(n19310), .A2(n19746), .B1(n19745), .B2(n19309), .ZN(
        n19308) );
  AOI22_X1 U22318 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19313), .B1(
        n19341), .B2(n19595), .ZN(n19307) );
  OAI211_X1 U22319 ( .C1(n19599), .C2(n19311), .A(n19308), .B(n19307), .ZN(
        P2_U3062) );
  AOI22_X1 U22320 ( .A1(n19310), .A2(n19753), .B1(n19751), .B2(n19309), .ZN(
        n19315) );
  INV_X1 U22321 ( .A(n19311), .ZN(n19312) );
  AOI22_X1 U22322 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19313), .B1(
        n19312), .B2(n19755), .ZN(n19314) );
  OAI211_X1 U22323 ( .C1(n19761), .C2(n19319), .A(n19315), .B(n19314), .ZN(
        P2_U3063) );
  NOR2_X1 U22324 ( .A1(n19877), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19541) );
  AND2_X1 U22325 ( .A1(n19541), .A2(n19347), .ZN(n19339) );
  OAI21_X1 U22326 ( .B1(n10490), .B2(n19339), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19318) );
  NOR2_X1 U22327 ( .A1(n19543), .A2(n19345), .ZN(n19320) );
  INV_X1 U22328 ( .A(n19320), .ZN(n19317) );
  NAND2_X1 U22329 ( .A1(n19318), .A2(n19317), .ZN(n19340) );
  AOI22_X1 U22330 ( .A1(n19340), .A2(n19690), .B1(n19676), .B2(n19339), .ZN(
        n19326) );
  AOI21_X1 U22331 ( .B1(n10490), .B2(n19680), .A(n19339), .ZN(n19323) );
  AOI21_X1 U22332 ( .B1(n19368), .B2(n19319), .A(n19420), .ZN(n19321) );
  NOR2_X1 U22333 ( .A1(n19321), .A2(n19320), .ZN(n19322) );
  MUX2_X1 U22334 ( .A(n19323), .B(n19322), .S(n19856), .Z(n19324) );
  OR2_X1 U22335 ( .A1(n19324), .A2(n19424), .ZN(n19342) );
  AOI22_X1 U22336 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19342), .B1(
        n19341), .B2(n19677), .ZN(n19325) );
  OAI211_X1 U22337 ( .C1(n19693), .C2(n19368), .A(n19326), .B(n19325), .ZN(
        P2_U3064) );
  AOI22_X1 U22338 ( .A1(n19340), .A2(n19718), .B1(n19247), .B2(n19339), .ZN(
        n19328) );
  AOI22_X1 U22339 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19342), .B1(
        n19341), .B2(n19719), .ZN(n19327) );
  OAI211_X1 U22340 ( .C1(n19658), .C2(n19368), .A(n19328), .B(n19327), .ZN(
        P2_U3065) );
  AOI22_X1 U22341 ( .A1(n19340), .A2(n19699), .B1(n19697), .B2(n19339), .ZN(
        n19330) );
  AOI22_X1 U22342 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19342), .B1(
        n19341), .B2(n19620), .ZN(n19329) );
  OAI211_X1 U22343 ( .C1(n19623), .C2(n19368), .A(n19330), .B(n19329), .ZN(
        P2_U3066) );
  AOI22_X1 U22344 ( .A1(n19340), .A2(n19726), .B1(n19725), .B2(n19339), .ZN(
        n19332) );
  AOI22_X1 U22345 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19342), .B1(
        n19341), .B2(n19727), .ZN(n19331) );
  OAI211_X1 U22346 ( .C1(n19730), .C2(n19368), .A(n19332), .B(n19331), .ZN(
        P2_U3067) );
  AOI22_X1 U22347 ( .A1(n19340), .A2(n19732), .B1(n19731), .B2(n19339), .ZN(
        n19334) );
  AOI22_X1 U22348 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19342), .B1(
        n19341), .B2(n19733), .ZN(n19333) );
  OAI211_X1 U22349 ( .C1(n19736), .C2(n19368), .A(n19334), .B(n19333), .ZN(
        P2_U3068) );
  AOI22_X1 U22350 ( .A1(n19340), .A2(n19738), .B1(n19737), .B2(n19339), .ZN(
        n19336) );
  AOI22_X1 U22351 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19342), .B1(
        n19341), .B2(n19628), .ZN(n19335) );
  OAI211_X1 U22352 ( .C1(n19631), .C2(n19368), .A(n19336), .B(n19335), .ZN(
        P2_U3069) );
  AOI22_X1 U22353 ( .A1(n19340), .A2(n19746), .B1(n19745), .B2(n19339), .ZN(
        n19338) );
  AOI22_X1 U22354 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19342), .B1(
        n19341), .B2(n19747), .ZN(n19337) );
  OAI211_X1 U22355 ( .C1(n19750), .C2(n19368), .A(n19338), .B(n19337), .ZN(
        P2_U3070) );
  AOI22_X1 U22356 ( .A1(n19340), .A2(n19753), .B1(n19751), .B2(n19339), .ZN(
        n19344) );
  AOI22_X1 U22357 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19342), .B1(
        n19341), .B2(n19755), .ZN(n19343) );
  OAI211_X1 U22358 ( .C1(n19761), .C2(n19368), .A(n19344), .B(n19343), .ZN(
        P2_U3071) );
  NOR2_X1 U22359 ( .A1(n19570), .A2(n19345), .ZN(n19369) );
  AOI22_X1 U22360 ( .A1(n19652), .A2(n19390), .B1(n19676), .B2(n19369), .ZN(
        n19355) );
  OR2_X1 U22361 ( .A1(n19452), .A2(n19578), .ZN(n19346) );
  NAND2_X1 U22362 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19347), .ZN(
        n19352) );
  NOR2_X1 U22363 ( .A1(n19348), .A2(n19369), .ZN(n19351) );
  AOI22_X1 U22364 ( .A1(n19350), .A2(n19352), .B1(P2_STATE2_REG_2__SCAN_IN), 
        .B2(n19351), .ZN(n19349) );
  OAI211_X1 U22365 ( .C1(n19369), .C2(n19680), .A(n19349), .B(n19683), .ZN(
        n19372) );
  INV_X1 U22366 ( .A(n19350), .ZN(n19353) );
  OAI22_X1 U22367 ( .A1(n19353), .A2(n19352), .B1(n19544), .B2(n19351), .ZN(
        n19371) );
  AOI22_X1 U22368 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19372), .B1(
        n19690), .B2(n19371), .ZN(n19354) );
  OAI211_X1 U22369 ( .C1(n19655), .C2(n19368), .A(n19355), .B(n19354), .ZN(
        P2_U3072) );
  AOI22_X1 U22370 ( .A1(n19720), .A2(n19390), .B1(n19369), .B2(n19247), .ZN(
        n19357) );
  AOI22_X1 U22371 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19372), .B1(
        n19718), .B2(n19371), .ZN(n19356) );
  OAI211_X1 U22372 ( .C1(n19696), .C2(n19368), .A(n19357), .B(n19356), .ZN(
        P2_U3073) );
  INV_X1 U22373 ( .A(n19368), .ZN(n19370) );
  AOI22_X1 U22374 ( .A1(n19620), .A2(n19370), .B1(n19697), .B2(n19369), .ZN(
        n19359) );
  AOI22_X1 U22375 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19372), .B1(
        n19699), .B2(n19371), .ZN(n19358) );
  OAI211_X1 U22376 ( .C1(n19623), .C2(n19387), .A(n19359), .B(n19358), .ZN(
        P2_U3074) );
  AOI22_X1 U22377 ( .A1(n19585), .A2(n19390), .B1(n19369), .B2(n19725), .ZN(
        n19361) );
  AOI22_X1 U22378 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19372), .B1(
        n19726), .B2(n19371), .ZN(n19360) );
  OAI211_X1 U22379 ( .C1(n19588), .C2(n19368), .A(n19361), .B(n19360), .ZN(
        P2_U3075) );
  AOI22_X1 U22380 ( .A1(n19589), .A2(n19390), .B1(n19369), .B2(n19731), .ZN(
        n19363) );
  AOI22_X1 U22381 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19372), .B1(
        n19732), .B2(n19371), .ZN(n19362) );
  OAI211_X1 U22382 ( .C1(n19592), .C2(n19368), .A(n19363), .B(n19362), .ZN(
        P2_U3076) );
  AOI22_X1 U22383 ( .A1(n19739), .A2(n19390), .B1(n19737), .B2(n19369), .ZN(
        n19365) );
  AOI22_X1 U22384 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19372), .B1(
        n19738), .B2(n19371), .ZN(n19364) );
  OAI211_X1 U22385 ( .C1(n19744), .C2(n19368), .A(n19365), .B(n19364), .ZN(
        P2_U3077) );
  AOI22_X1 U22386 ( .A1(n19595), .A2(n19390), .B1(n19369), .B2(n19745), .ZN(
        n19367) );
  AOI22_X1 U22387 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19372), .B1(
        n19746), .B2(n19371), .ZN(n19366) );
  OAI211_X1 U22388 ( .C1(n19599), .C2(n19368), .A(n19367), .B(n19366), .ZN(
        P2_U3078) );
  AOI22_X1 U22389 ( .A1(n19755), .A2(n19370), .B1(n19369), .B2(n19751), .ZN(
        n19374) );
  AOI22_X1 U22390 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19372), .B1(
        n19753), .B2(n19371), .ZN(n19373) );
  OAI211_X1 U22391 ( .C1(n19761), .C2(n19387), .A(n19374), .B(n19373), .ZN(
        P2_U3079) );
  AOI22_X1 U22392 ( .A1(n19389), .A2(n19718), .B1(n19247), .B2(n19388), .ZN(
        n19376) );
  AOI22_X1 U22393 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19391), .B1(
        n19409), .B2(n19720), .ZN(n19375) );
  OAI211_X1 U22394 ( .C1(n19696), .C2(n19387), .A(n19376), .B(n19375), .ZN(
        P2_U3081) );
  AOI22_X1 U22395 ( .A1(n19389), .A2(n19699), .B1(n19697), .B2(n19388), .ZN(
        n19378) );
  AOI22_X1 U22396 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19391), .B1(
        n19409), .B2(n19698), .ZN(n19377) );
  OAI211_X1 U22397 ( .C1(n19702), .C2(n19387), .A(n19378), .B(n19377), .ZN(
        P2_U3082) );
  AOI22_X1 U22398 ( .A1(n19389), .A2(n19726), .B1(n19725), .B2(n19388), .ZN(
        n19380) );
  AOI22_X1 U22399 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19391), .B1(
        n19409), .B2(n19585), .ZN(n19379) );
  OAI211_X1 U22400 ( .C1(n19588), .C2(n19387), .A(n19380), .B(n19379), .ZN(
        P2_U3083) );
  AOI22_X1 U22401 ( .A1(n19389), .A2(n19732), .B1(n19731), .B2(n19388), .ZN(
        n19382) );
  AOI22_X1 U22402 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19391), .B1(
        n19409), .B2(n19589), .ZN(n19381) );
  OAI211_X1 U22403 ( .C1(n19592), .C2(n19387), .A(n19382), .B(n19381), .ZN(
        P2_U3084) );
  AOI22_X1 U22404 ( .A1(n19389), .A2(n19738), .B1(n19737), .B2(n19388), .ZN(
        n19384) );
  AOI22_X1 U22405 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19391), .B1(
        n19409), .B2(n19739), .ZN(n19383) );
  OAI211_X1 U22406 ( .C1(n19744), .C2(n19387), .A(n19384), .B(n19383), .ZN(
        P2_U3085) );
  AOI22_X1 U22407 ( .A1(n19389), .A2(n19746), .B1(n19745), .B2(n19388), .ZN(
        n19386) );
  AOI22_X1 U22408 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19391), .B1(
        n19409), .B2(n19595), .ZN(n19385) );
  OAI211_X1 U22409 ( .C1(n19599), .C2(n19387), .A(n19386), .B(n19385), .ZN(
        P2_U3086) );
  AOI22_X1 U22410 ( .A1(n19389), .A2(n19753), .B1(n19751), .B2(n19388), .ZN(
        n19393) );
  AOI22_X1 U22411 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19391), .B1(
        n19390), .B2(n19755), .ZN(n19392) );
  OAI211_X1 U22412 ( .C1(n19761), .C2(n19396), .A(n19393), .B(n19392), .ZN(
        P2_U3087) );
  AOI22_X1 U22413 ( .A1(n19720), .A2(n19443), .B1(n19422), .B2(n19247), .ZN(
        n19395) );
  AOI22_X1 U22414 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19407), .B1(
        n19718), .B2(n19410), .ZN(n19394) );
  OAI211_X1 U22415 ( .C1(n19696), .C2(n19396), .A(n19395), .B(n19394), .ZN(
        P2_U3089) );
  AOI22_X1 U22416 ( .A1(n19620), .A2(n19409), .B1(n19422), .B2(n19697), .ZN(
        n19398) );
  AOI22_X1 U22417 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19407), .B1(
        n19699), .B2(n19410), .ZN(n19397) );
  OAI211_X1 U22418 ( .C1(n19623), .C2(n19440), .A(n19398), .B(n19397), .ZN(
        P2_U3090) );
  AOI22_X1 U22419 ( .A1(n19727), .A2(n19409), .B1(n19422), .B2(n19725), .ZN(
        n19400) );
  AOI22_X1 U22420 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19407), .B1(
        n19726), .B2(n19410), .ZN(n19399) );
  OAI211_X1 U22421 ( .C1(n19730), .C2(n19440), .A(n19400), .B(n19399), .ZN(
        P2_U3091) );
  AOI22_X1 U22422 ( .A1(n19733), .A2(n19409), .B1(n19422), .B2(n19731), .ZN(
        n19402) );
  AOI22_X1 U22423 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19407), .B1(
        n19732), .B2(n19410), .ZN(n19401) );
  OAI211_X1 U22424 ( .C1(n19736), .C2(n19440), .A(n19402), .B(n19401), .ZN(
        P2_U3092) );
  AOI22_X1 U22425 ( .A1(n19628), .A2(n19409), .B1(n19422), .B2(n19737), .ZN(
        n19404) );
  AOI22_X1 U22426 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19407), .B1(
        n19738), .B2(n19410), .ZN(n19403) );
  OAI211_X1 U22427 ( .C1(n19631), .C2(n19440), .A(n19404), .B(n19403), .ZN(
        P2_U3093) );
  AOI22_X1 U22428 ( .A1(n19747), .A2(n19409), .B1(n19422), .B2(n19745), .ZN(
        n19406) );
  AOI22_X1 U22429 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19407), .B1(
        n19746), .B2(n19410), .ZN(n19405) );
  OAI211_X1 U22430 ( .C1(n19750), .C2(n19440), .A(n19406), .B(n19405), .ZN(
        P2_U3094) );
  INV_X1 U22431 ( .A(n19407), .ZN(n19414) );
  INV_X1 U22432 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n19413) );
  INV_X1 U22433 ( .A(n19761), .ZN(n19408) );
  AOI22_X1 U22434 ( .A1(n19408), .A2(n19443), .B1(n19422), .B2(n19751), .ZN(
        n19412) );
  AOI22_X1 U22435 ( .A1(n19753), .A2(n19410), .B1(n19409), .B2(n19755), .ZN(
        n19411) );
  OAI211_X1 U22436 ( .C1(n19414), .C2(n19413), .A(n19412), .B(n19411), .ZN(
        P2_U3095) );
  NOR2_X1 U22437 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19415), .ZN(
        n19455) );
  INV_X1 U22438 ( .A(n19455), .ZN(n19450) );
  NOR2_X1 U22439 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19450), .ZN(
        n19441) );
  NOR2_X1 U22440 ( .A1(n19422), .A2(n19441), .ZN(n19416) );
  OR2_X1 U22441 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19416), .ZN(n19418) );
  NOR3_X1 U22442 ( .A1(n19417), .A2(n19544), .A3(n19441), .ZN(n19423) );
  AOI21_X1 U22443 ( .B1(n19544), .B2(n19418), .A(n19423), .ZN(n19442) );
  AOI22_X1 U22444 ( .A1(n19442), .A2(n19690), .B1(n19676), .B2(n19441), .ZN(
        n19427) );
  AOI21_X1 U22445 ( .B1(n19440), .B2(n19470), .A(n19420), .ZN(n19421) );
  AOI221_X1 U22446 ( .B1(n19680), .B2(n19422), .C1(n19680), .C2(n19421), .A(
        n19441), .ZN(n19425) );
  OR3_X1 U22447 ( .A1(n19425), .A2(n19424), .A3(n19423), .ZN(n19444) );
  AOI22_X1 U22448 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19444), .B1(
        n19473), .B2(n19652), .ZN(n19426) );
  OAI211_X1 U22449 ( .C1(n19655), .C2(n19440), .A(n19427), .B(n19426), .ZN(
        P2_U3096) );
  AOI22_X1 U22450 ( .A1(n19442), .A2(n19718), .B1(n19247), .B2(n19441), .ZN(
        n19429) );
  AOI22_X1 U22451 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19444), .B1(
        n19473), .B2(n19720), .ZN(n19428) );
  OAI211_X1 U22452 ( .C1(n19696), .C2(n19440), .A(n19429), .B(n19428), .ZN(
        P2_U3097) );
  AOI22_X1 U22453 ( .A1(n19442), .A2(n19699), .B1(n19697), .B2(n19441), .ZN(
        n19431) );
  AOI22_X1 U22454 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19444), .B1(
        n19473), .B2(n19698), .ZN(n19430) );
  OAI211_X1 U22455 ( .C1(n19702), .C2(n19440), .A(n19431), .B(n19430), .ZN(
        P2_U3098) );
  AOI22_X1 U22456 ( .A1(n19442), .A2(n19726), .B1(n19725), .B2(n19441), .ZN(
        n19433) );
  AOI22_X1 U22457 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19444), .B1(
        n19473), .B2(n19585), .ZN(n19432) );
  OAI211_X1 U22458 ( .C1(n19588), .C2(n19440), .A(n19433), .B(n19432), .ZN(
        P2_U3099) );
  AOI22_X1 U22459 ( .A1(n19442), .A2(n19732), .B1(n19731), .B2(n19441), .ZN(
        n19435) );
  AOI22_X1 U22460 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19444), .B1(
        n19473), .B2(n19589), .ZN(n19434) );
  OAI211_X1 U22461 ( .C1(n19592), .C2(n19440), .A(n19435), .B(n19434), .ZN(
        P2_U3100) );
  AOI22_X1 U22462 ( .A1(n19442), .A2(n19738), .B1(n19737), .B2(n19441), .ZN(
        n19437) );
  AOI22_X1 U22463 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19444), .B1(
        n19473), .B2(n19739), .ZN(n19436) );
  OAI211_X1 U22464 ( .C1(n19744), .C2(n19440), .A(n19437), .B(n19436), .ZN(
        P2_U3101) );
  AOI22_X1 U22465 ( .A1(n19442), .A2(n19746), .B1(n19745), .B2(n19441), .ZN(
        n19439) );
  AOI22_X1 U22466 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19444), .B1(
        n19473), .B2(n19595), .ZN(n19438) );
  OAI211_X1 U22467 ( .C1(n19599), .C2(n19440), .A(n19439), .B(n19438), .ZN(
        P2_U3102) );
  AOI22_X1 U22468 ( .A1(n19442), .A2(n19753), .B1(n19751), .B2(n19441), .ZN(
        n19446) );
  AOI22_X1 U22469 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19444), .B1(
        n19443), .B2(n19755), .ZN(n19445) );
  OAI211_X1 U22470 ( .C1(n19761), .C2(n19470), .A(n19446), .B(n19445), .ZN(
        P2_U3103) );
  INV_X1 U22471 ( .A(n19451), .ZN(n19447) );
  NAND2_X1 U22472 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19455), .ZN(
        n19486) );
  INV_X1 U22473 ( .A(n19486), .ZN(n19471) );
  OAI21_X1 U22474 ( .B1(n10478), .B2(n19471), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19449) );
  OAI21_X1 U22475 ( .B1(n19450), .B2(n19513), .A(n19449), .ZN(n19472) );
  AOI22_X1 U22476 ( .A1(n19472), .A2(n19690), .B1(n19676), .B2(n19471), .ZN(
        n19457) );
  NOR2_X1 U22477 ( .A1(n19452), .A2(n19451), .ZN(n19855) );
  NAND2_X1 U22478 ( .A1(n10478), .A2(n19680), .ZN(n19453) );
  NAND3_X1 U22479 ( .A1(n19453), .A2(n19486), .A3(n19513), .ZN(n19454) );
  OAI211_X1 U22480 ( .C1(n19855), .C2(n19455), .A(n19683), .B(n19454), .ZN(
        n19474) );
  AOI22_X1 U22481 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19474), .B1(
        n19473), .B2(n19677), .ZN(n19456) );
  OAI211_X1 U22482 ( .C1(n19693), .C2(n19502), .A(n19457), .B(n19456), .ZN(
        P2_U3104) );
  AOI22_X1 U22483 ( .A1(n19472), .A2(n19718), .B1(n19247), .B2(n19471), .ZN(
        n19459) );
  AOI22_X1 U22484 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19474), .B1(
        n19504), .B2(n19720), .ZN(n19458) );
  OAI211_X1 U22485 ( .C1(n19696), .C2(n19470), .A(n19459), .B(n19458), .ZN(
        P2_U3105) );
  AOI22_X1 U22486 ( .A1(n19472), .A2(n19699), .B1(n19697), .B2(n19471), .ZN(
        n19461) );
  AOI22_X1 U22487 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19474), .B1(
        n19473), .B2(n19620), .ZN(n19460) );
  OAI211_X1 U22488 ( .C1(n19623), .C2(n19502), .A(n19461), .B(n19460), .ZN(
        P2_U3106) );
  AOI22_X1 U22489 ( .A1(n19472), .A2(n19726), .B1(n19725), .B2(n19471), .ZN(
        n19463) );
  AOI22_X1 U22490 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19474), .B1(
        n19504), .B2(n19585), .ZN(n19462) );
  OAI211_X1 U22491 ( .C1(n19588), .C2(n19470), .A(n19463), .B(n19462), .ZN(
        P2_U3107) );
  AOI22_X1 U22492 ( .A1(n19472), .A2(n19732), .B1(n19731), .B2(n19471), .ZN(
        n19465) );
  AOI22_X1 U22493 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19474), .B1(
        n19504), .B2(n19589), .ZN(n19464) );
  OAI211_X1 U22494 ( .C1(n19592), .C2(n19470), .A(n19465), .B(n19464), .ZN(
        P2_U3108) );
  AOI22_X1 U22495 ( .A1(n19472), .A2(n19738), .B1(n19737), .B2(n19471), .ZN(
        n19467) );
  AOI22_X1 U22496 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19474), .B1(
        n19504), .B2(n19739), .ZN(n19466) );
  OAI211_X1 U22497 ( .C1(n19744), .C2(n19470), .A(n19467), .B(n19466), .ZN(
        P2_U3109) );
  AOI22_X1 U22498 ( .A1(n19472), .A2(n19746), .B1(n19745), .B2(n19471), .ZN(
        n19469) );
  AOI22_X1 U22499 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19474), .B1(
        n19504), .B2(n19595), .ZN(n19468) );
  OAI211_X1 U22500 ( .C1(n19599), .C2(n19470), .A(n19469), .B(n19468), .ZN(
        P2_U3110) );
  AOI22_X1 U22501 ( .A1(n19472), .A2(n19753), .B1(n19751), .B2(n19471), .ZN(
        n19476) );
  AOI22_X1 U22502 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19474), .B1(
        n19473), .B2(n19755), .ZN(n19475) );
  OAI211_X1 U22503 ( .C1(n19761), .C2(n19502), .A(n19476), .B(n19475), .ZN(
        P2_U3111) );
  NOR2_X1 U22504 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19861), .ZN(
        n19569) );
  NAND2_X1 U22505 ( .A1(n19569), .A2(n19877), .ZN(n19518) );
  NOR2_X1 U22506 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19518), .ZN(
        n19503) );
  AOI22_X1 U22507 ( .A1(n19677), .A2(n19504), .B1(n19676), .B2(n19503), .ZN(
        n19489) );
  NOR3_X1 U22508 ( .A1(n19535), .A2(n19504), .A3(n19513), .ZN(n19479) );
  INV_X1 U22509 ( .A(n19678), .ZN(n19478) );
  NOR2_X1 U22510 ( .A1(n19479), .A2(n19478), .ZN(n19487) );
  INV_X1 U22511 ( .A(n19487), .ZN(n19482) );
  OAI21_X1 U22512 ( .B1(n19483), .B2(n19544), .A(n19680), .ZN(n19480) );
  AOI21_X1 U22513 ( .B1(n19482), .B2(n19486), .A(n19480), .ZN(n19481) );
  NOR2_X1 U22514 ( .A1(n19482), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19485) );
  AOI21_X1 U22515 ( .B1(n19483), .B2(P2_STATE2_REG_2__SCAN_IN), .A(n19503), 
        .ZN(n19484) );
  AOI22_X1 U22516 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19506), .B1(
        n19690), .B2(n19505), .ZN(n19488) );
  OAI211_X1 U22517 ( .C1(n19693), .C2(n19532), .A(n19489), .B(n19488), .ZN(
        P2_U3112) );
  AOI22_X1 U22518 ( .A1(n19720), .A2(n19535), .B1(n19503), .B2(n19247), .ZN(
        n19491) );
  AOI22_X1 U22519 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19506), .B1(
        n19505), .B2(n19718), .ZN(n19490) );
  OAI211_X1 U22520 ( .C1(n19696), .C2(n19502), .A(n19491), .B(n19490), .ZN(
        P2_U3113) );
  AOI22_X1 U22521 ( .A1(n19698), .A2(n19535), .B1(n19697), .B2(n19503), .ZN(
        n19493) );
  AOI22_X1 U22522 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19506), .B1(
        n19505), .B2(n19699), .ZN(n19492) );
  OAI211_X1 U22523 ( .C1(n19702), .C2(n19502), .A(n19493), .B(n19492), .ZN(
        P2_U3114) );
  AOI22_X1 U22524 ( .A1(n19727), .A2(n19504), .B1(n19503), .B2(n19725), .ZN(
        n19495) );
  AOI22_X1 U22525 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19506), .B1(
        n19505), .B2(n19726), .ZN(n19494) );
  OAI211_X1 U22526 ( .C1(n19730), .C2(n19532), .A(n19495), .B(n19494), .ZN(
        P2_U3115) );
  AOI22_X1 U22527 ( .A1(n19733), .A2(n19504), .B1(n19503), .B2(n19731), .ZN(
        n19497) );
  AOI22_X1 U22528 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19506), .B1(
        n19505), .B2(n19732), .ZN(n19496) );
  OAI211_X1 U22529 ( .C1(n19736), .C2(n19532), .A(n19497), .B(n19496), .ZN(
        P2_U3116) );
  AOI22_X1 U22530 ( .A1(n19628), .A2(n19504), .B1(n19737), .B2(n19503), .ZN(
        n19499) );
  AOI22_X1 U22531 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19506), .B1(
        n19505), .B2(n19738), .ZN(n19498) );
  OAI211_X1 U22532 ( .C1(n19631), .C2(n19532), .A(n19499), .B(n19498), .ZN(
        P2_U3117) );
  AOI22_X1 U22533 ( .A1(n19595), .A2(n19535), .B1(n19503), .B2(n19745), .ZN(
        n19501) );
  AOI22_X1 U22534 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19506), .B1(
        n19505), .B2(n19746), .ZN(n19500) );
  OAI211_X1 U22535 ( .C1(n19599), .C2(n19502), .A(n19501), .B(n19500), .ZN(
        P2_U3118) );
  AOI22_X1 U22536 ( .A1(n19755), .A2(n19504), .B1(n19503), .B2(n19751), .ZN(
        n19508) );
  AOI22_X1 U22537 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19506), .B1(
        n19505), .B2(n19753), .ZN(n19507) );
  OAI211_X1 U22538 ( .C1(n19761), .C2(n19532), .A(n19508), .B(n19507), .ZN(
        P2_U3119) );
  INV_X1 U22539 ( .A(n19569), .ZN(n19575) );
  NOR2_X1 U22540 ( .A1(n19510), .A2(n19575), .ZN(n19545) );
  AOI22_X1 U22541 ( .A1(n19652), .A2(n19565), .B1(n19676), .B2(n19545), .ZN(
        n19521) );
  OAI21_X1 U22542 ( .B1(n19643), .B2(n19511), .A(n19856), .ZN(n19519) );
  INV_X1 U22543 ( .A(n19518), .ZN(n19516) );
  INV_X1 U22544 ( .A(n19545), .ZN(n19512) );
  OAI211_X1 U22545 ( .C1(n19514), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19513), 
        .B(n19512), .ZN(n19515) );
  OAI211_X1 U22546 ( .C1(n19519), .C2(n19516), .A(n19683), .B(n19515), .ZN(
        n19537) );
  OAI21_X1 U22547 ( .B1(n10477), .B2(n19545), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19517) );
  AOI22_X1 U22548 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19537), .B1(
        n19690), .B2(n19536), .ZN(n19520) );
  OAI211_X1 U22549 ( .C1(n19655), .C2(n19532), .A(n19521), .B(n19520), .ZN(
        P2_U3120) );
  INV_X1 U22550 ( .A(n19565), .ZN(n19540) );
  AOI22_X1 U22551 ( .A1(n19719), .A2(n19535), .B1(n19545), .B2(n19247), .ZN(
        n19523) );
  AOI22_X1 U22552 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19537), .B1(
        n19718), .B2(n19536), .ZN(n19522) );
  OAI211_X1 U22553 ( .C1(n19658), .C2(n19540), .A(n19523), .B(n19522), .ZN(
        P2_U3121) );
  AOI22_X1 U22554 ( .A1(n19698), .A2(n19565), .B1(n19697), .B2(n19545), .ZN(
        n19525) );
  AOI22_X1 U22555 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19537), .B1(
        n19699), .B2(n19536), .ZN(n19524) );
  OAI211_X1 U22556 ( .C1(n19702), .C2(n19532), .A(n19525), .B(n19524), .ZN(
        P2_U3122) );
  AOI22_X1 U22557 ( .A1(n19727), .A2(n19535), .B1(n19545), .B2(n19725), .ZN(
        n19527) );
  AOI22_X1 U22558 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19537), .B1(
        n19726), .B2(n19536), .ZN(n19526) );
  OAI211_X1 U22559 ( .C1(n19730), .C2(n19540), .A(n19527), .B(n19526), .ZN(
        P2_U3123) );
  AOI22_X1 U22560 ( .A1(n19733), .A2(n19535), .B1(n19545), .B2(n19731), .ZN(
        n19529) );
  AOI22_X1 U22561 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19537), .B1(
        n19732), .B2(n19536), .ZN(n19528) );
  OAI211_X1 U22562 ( .C1(n19736), .C2(n19540), .A(n19529), .B(n19528), .ZN(
        P2_U3124) );
  AOI22_X1 U22563 ( .A1(n19739), .A2(n19565), .B1(n19737), .B2(n19545), .ZN(
        n19531) );
  AOI22_X1 U22564 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19537), .B1(
        n19738), .B2(n19536), .ZN(n19530) );
  OAI211_X1 U22565 ( .C1(n19744), .C2(n19532), .A(n19531), .B(n19530), .ZN(
        P2_U3125) );
  AOI22_X1 U22566 ( .A1(n19747), .A2(n19535), .B1(n19745), .B2(n19545), .ZN(
        n19534) );
  AOI22_X1 U22567 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19537), .B1(
        n19746), .B2(n19536), .ZN(n19533) );
  OAI211_X1 U22568 ( .C1(n19750), .C2(n19540), .A(n19534), .B(n19533), .ZN(
        P2_U3126) );
  AOI22_X1 U22569 ( .A1(n19755), .A2(n19535), .B1(n19545), .B2(n19751), .ZN(
        n19539) );
  AOI22_X1 U22570 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19537), .B1(
        n19753), .B2(n19536), .ZN(n19538) );
  OAI211_X1 U22571 ( .C1(n19761), .C2(n19540), .A(n19539), .B(n19538), .ZN(
        P2_U3127) );
  AND2_X1 U22572 ( .A1(n19541), .A2(n19569), .ZN(n19563) );
  OAI21_X1 U22573 ( .B1(n10491), .B2(n19563), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19542) );
  AOI22_X1 U22574 ( .A1(n19564), .A2(n19690), .B1(n19676), .B2(n19563), .ZN(
        n19550) );
  INV_X1 U22575 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19544) );
  NOR2_X1 U22576 ( .A1(n10491), .A2(n19544), .ZN(n19547) );
  INV_X1 U22577 ( .A(n19598), .ZN(n19602) );
  AOI221_X1 U22578 ( .B1(n19602), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19565), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19545), .ZN(n19546) );
  NOR3_X1 U22579 ( .A1(n19547), .A2(n19546), .A3(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n19548) );
  AOI22_X1 U22580 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19566), .B1(
        n19565), .B2(n19677), .ZN(n19549) );
  OAI211_X1 U22581 ( .C1(n19693), .C2(n19598), .A(n19550), .B(n19549), .ZN(
        P2_U3128) );
  AOI22_X1 U22582 ( .A1(n19564), .A2(n19718), .B1(n19247), .B2(n19563), .ZN(
        n19552) );
  AOI22_X1 U22583 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19566), .B1(
        n19565), .B2(n19719), .ZN(n19551) );
  OAI211_X1 U22584 ( .C1(n19658), .C2(n19598), .A(n19552), .B(n19551), .ZN(
        P2_U3129) );
  AOI22_X1 U22585 ( .A1(n19564), .A2(n19699), .B1(n19697), .B2(n19563), .ZN(
        n19554) );
  AOI22_X1 U22586 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19566), .B1(
        n19565), .B2(n19620), .ZN(n19553) );
  OAI211_X1 U22587 ( .C1(n19623), .C2(n19598), .A(n19554), .B(n19553), .ZN(
        P2_U3130) );
  AOI22_X1 U22588 ( .A1(n19564), .A2(n19726), .B1(n19725), .B2(n19563), .ZN(
        n19556) );
  AOI22_X1 U22589 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19566), .B1(
        n19565), .B2(n19727), .ZN(n19555) );
  OAI211_X1 U22590 ( .C1(n19730), .C2(n19598), .A(n19556), .B(n19555), .ZN(
        P2_U3131) );
  AOI22_X1 U22591 ( .A1(n19564), .A2(n19732), .B1(n19731), .B2(n19563), .ZN(
        n19558) );
  AOI22_X1 U22592 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19566), .B1(
        n19565), .B2(n19733), .ZN(n19557) );
  OAI211_X1 U22593 ( .C1(n19736), .C2(n19598), .A(n19558), .B(n19557), .ZN(
        P2_U3132) );
  AOI22_X1 U22594 ( .A1(n19564), .A2(n19738), .B1(n19737), .B2(n19563), .ZN(
        n19560) );
  AOI22_X1 U22595 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19566), .B1(
        n19565), .B2(n19628), .ZN(n19559) );
  OAI211_X1 U22596 ( .C1(n19631), .C2(n19598), .A(n19560), .B(n19559), .ZN(
        P2_U3133) );
  AOI22_X1 U22597 ( .A1(n19564), .A2(n19746), .B1(n19745), .B2(n19563), .ZN(
        n19562) );
  AOI22_X1 U22598 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19566), .B1(
        n19565), .B2(n19747), .ZN(n19561) );
  OAI211_X1 U22599 ( .C1(n19750), .C2(n19598), .A(n19562), .B(n19561), .ZN(
        P2_U3134) );
  AOI22_X1 U22600 ( .A1(n19564), .A2(n19753), .B1(n19751), .B2(n19563), .ZN(
        n19568) );
  AOI22_X1 U22601 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19566), .B1(
        n19565), .B2(n19755), .ZN(n19567) );
  OAI211_X1 U22602 ( .C1(n19761), .C2(n19598), .A(n19568), .B(n19567), .ZN(
        P2_U3135) );
  NAND3_X1 U22603 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19569), .A3(
        n19680), .ZN(n19572) );
  NOR2_X1 U22604 ( .A1(n19575), .A2(n19570), .ZN(n19600) );
  NOR3_X1 U22605 ( .A1(n19573), .A2(n19544), .A3(n19600), .ZN(n19571) );
  AOI21_X1 U22606 ( .B1(n19544), .B2(n19572), .A(n19571), .ZN(n19601) );
  AOI22_X1 U22607 ( .A1(n19601), .A2(n19690), .B1(n19676), .B2(n19600), .ZN(
        n19580) );
  INV_X1 U22608 ( .A(n19573), .ZN(n19574) );
  AOI21_X1 U22609 ( .B1(n19574), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19577) );
  OAI22_X1 U22610 ( .A1(n19643), .A2(n19578), .B1(n19575), .B2(n19877), .ZN(
        n19576) );
  OAI211_X1 U22611 ( .C1(n19600), .C2(n19577), .A(n19576), .B(n19683), .ZN(
        n19603) );
  AOI22_X1 U22612 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19603), .B1(
        n19636), .B2(n19652), .ZN(n19579) );
  OAI211_X1 U22613 ( .C1(n19655), .C2(n19598), .A(n19580), .B(n19579), .ZN(
        P2_U3136) );
  AOI22_X1 U22614 ( .A1(n19601), .A2(n19718), .B1(n19247), .B2(n19600), .ZN(
        n19582) );
  AOI22_X1 U22615 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19603), .B1(
        n19636), .B2(n19720), .ZN(n19581) );
  OAI211_X1 U22616 ( .C1(n19696), .C2(n19598), .A(n19582), .B(n19581), .ZN(
        P2_U3137) );
  AOI22_X1 U22617 ( .A1(n19601), .A2(n19699), .B1(n19697), .B2(n19600), .ZN(
        n19584) );
  AOI22_X1 U22618 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19603), .B1(
        n19636), .B2(n19698), .ZN(n19583) );
  OAI211_X1 U22619 ( .C1(n19702), .C2(n19598), .A(n19584), .B(n19583), .ZN(
        P2_U3138) );
  AOI22_X1 U22620 ( .A1(n19601), .A2(n19726), .B1(n19725), .B2(n19600), .ZN(
        n19587) );
  AOI22_X1 U22621 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19603), .B1(
        n19636), .B2(n19585), .ZN(n19586) );
  OAI211_X1 U22622 ( .C1(n19588), .C2(n19598), .A(n19587), .B(n19586), .ZN(
        P2_U3139) );
  AOI22_X1 U22623 ( .A1(n19601), .A2(n19732), .B1(n19731), .B2(n19600), .ZN(
        n19591) );
  AOI22_X1 U22624 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19603), .B1(
        n19636), .B2(n19589), .ZN(n19590) );
  OAI211_X1 U22625 ( .C1(n19592), .C2(n19598), .A(n19591), .B(n19590), .ZN(
        P2_U3140) );
  AOI22_X1 U22626 ( .A1(n19601), .A2(n19738), .B1(n19737), .B2(n19600), .ZN(
        n19594) );
  AOI22_X1 U22627 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19603), .B1(
        n19636), .B2(n19739), .ZN(n19593) );
  OAI211_X1 U22628 ( .C1(n19744), .C2(n19598), .A(n19594), .B(n19593), .ZN(
        P2_U3141) );
  AOI22_X1 U22629 ( .A1(n19601), .A2(n19746), .B1(n19745), .B2(n19600), .ZN(
        n19597) );
  AOI22_X1 U22630 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19603), .B1(
        n19636), .B2(n19595), .ZN(n19596) );
  OAI211_X1 U22631 ( .C1(n19599), .C2(n19598), .A(n19597), .B(n19596), .ZN(
        P2_U3142) );
  INV_X1 U22632 ( .A(n19636), .ZN(n19606) );
  AOI22_X1 U22633 ( .A1(n19601), .A2(n19753), .B1(n19751), .B2(n19600), .ZN(
        n19605) );
  AOI22_X1 U22634 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19603), .B1(
        n19602), .B2(n19755), .ZN(n19604) );
  OAI211_X1 U22635 ( .C1(n19761), .C2(n19606), .A(n19605), .B(n19604), .ZN(
        P2_U3143) );
  NAND3_X1 U22636 ( .A1(n19877), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19647) );
  NOR2_X1 U22637 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19647), .ZN(
        n19634) );
  INV_X1 U22638 ( .A(n19634), .ZN(n19613) );
  NAND3_X1 U22639 ( .A1(n19608), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19613), 
        .ZN(n19614) );
  NAND2_X1 U22640 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19609), .ZN(
        n19612) );
  OAI21_X1 U22641 ( .B1(n19612), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19544), 
        .ZN(n19610) );
  AND2_X1 U22642 ( .A1(n19614), .A2(n19610), .ZN(n19635) );
  AOI22_X1 U22643 ( .A1(n19635), .A2(n19690), .B1(n19676), .B2(n19634), .ZN(
        n19617) );
  OAI21_X1 U22644 ( .B1(n19671), .B2(n19636), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19611) );
  AOI22_X1 U22645 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19613), .B1(n19612), 
        .B2(n19611), .ZN(n19615) );
  NAND3_X1 U22646 ( .A1(n19615), .A2(n19683), .A3(n19614), .ZN(n19637) );
  AOI22_X1 U22647 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19637), .B1(
        n19636), .B2(n19677), .ZN(n19616) );
  OAI211_X1 U22648 ( .C1(n19693), .C2(n19667), .A(n19617), .B(n19616), .ZN(
        P2_U3144) );
  AOI22_X1 U22649 ( .A1(n19635), .A2(n19718), .B1(n19247), .B2(n19634), .ZN(
        n19619) );
  AOI22_X1 U22650 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19637), .B1(
        n19636), .B2(n19719), .ZN(n19618) );
  OAI211_X1 U22651 ( .C1(n19658), .C2(n19667), .A(n19619), .B(n19618), .ZN(
        P2_U3145) );
  AOI22_X1 U22652 ( .A1(n19635), .A2(n19699), .B1(n19697), .B2(n19634), .ZN(
        n19622) );
  AOI22_X1 U22653 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19637), .B1(
        n19636), .B2(n19620), .ZN(n19621) );
  OAI211_X1 U22654 ( .C1(n19623), .C2(n19667), .A(n19622), .B(n19621), .ZN(
        P2_U3146) );
  AOI22_X1 U22655 ( .A1(n19635), .A2(n19726), .B1(n19725), .B2(n19634), .ZN(
        n19625) );
  AOI22_X1 U22656 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19637), .B1(
        n19636), .B2(n19727), .ZN(n19624) );
  OAI211_X1 U22657 ( .C1(n19730), .C2(n19667), .A(n19625), .B(n19624), .ZN(
        P2_U3147) );
  AOI22_X1 U22658 ( .A1(n19635), .A2(n19732), .B1(n19731), .B2(n19634), .ZN(
        n19627) );
  AOI22_X1 U22659 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19637), .B1(
        n19636), .B2(n19733), .ZN(n19626) );
  OAI211_X1 U22660 ( .C1(n19736), .C2(n19667), .A(n19627), .B(n19626), .ZN(
        P2_U3148) );
  AOI22_X1 U22661 ( .A1(n19635), .A2(n19738), .B1(n19737), .B2(n19634), .ZN(
        n19630) );
  AOI22_X1 U22662 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19637), .B1(
        n19636), .B2(n19628), .ZN(n19629) );
  OAI211_X1 U22663 ( .C1(n19631), .C2(n19667), .A(n19630), .B(n19629), .ZN(
        P2_U3149) );
  AOI22_X1 U22664 ( .A1(n19635), .A2(n19746), .B1(n19745), .B2(n19634), .ZN(
        n19633) );
  AOI22_X1 U22665 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19637), .B1(
        n19636), .B2(n19747), .ZN(n19632) );
  OAI211_X1 U22666 ( .C1(n19750), .C2(n19667), .A(n19633), .B(n19632), .ZN(
        P2_U3150) );
  AOI22_X1 U22667 ( .A1(n19635), .A2(n19753), .B1(n19751), .B2(n19634), .ZN(
        n19639) );
  AOI22_X1 U22668 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19637), .B1(
        n19636), .B2(n19755), .ZN(n19638) );
  OAI211_X1 U22669 ( .C1(n19761), .C2(n19667), .A(n19639), .B(n19638), .ZN(
        P2_U3151) );
  NOR2_X1 U22670 ( .A1(n19886), .A2(n19647), .ZN(n19686) );
  NOR3_X1 U22671 ( .A1(n19640), .A2(n19544), .A3(n19686), .ZN(n19646) );
  INV_X1 U22672 ( .A(n19647), .ZN(n19641) );
  AOI21_X1 U22673 ( .B1(n19680), .B2(n19641), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19642) );
  AOI22_X1 U22674 ( .A1(n19670), .A2(n19690), .B1(n19676), .B2(n19686), .ZN(
        n19654) );
  INV_X1 U22675 ( .A(n19643), .ZN(n19645) );
  NAND2_X1 U22676 ( .A1(n19645), .A2(n19644), .ZN(n19648) );
  AOI21_X1 U22677 ( .B1(n19648), .B2(n19647), .A(n19646), .ZN(n19649) );
  OAI211_X1 U22678 ( .C1(n19686), .C2(n19680), .A(n19649), .B(n19683), .ZN(
        n19672) );
  AOI22_X1 U22679 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19672), .B1(
        n19713), .B2(n19652), .ZN(n19653) );
  OAI211_X1 U22680 ( .C1(n19655), .C2(n19667), .A(n19654), .B(n19653), .ZN(
        P2_U3152) );
  AOI22_X1 U22681 ( .A1(n19670), .A2(n19718), .B1(n19247), .B2(n19686), .ZN(
        n19657) );
  AOI22_X1 U22682 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19672), .B1(
        n19671), .B2(n19719), .ZN(n19656) );
  OAI211_X1 U22683 ( .C1(n19658), .C2(n19709), .A(n19657), .B(n19656), .ZN(
        P2_U3153) );
  AOI22_X1 U22684 ( .A1(n19670), .A2(n19699), .B1(n19697), .B2(n19686), .ZN(
        n19660) );
  AOI22_X1 U22685 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19672), .B1(
        n19713), .B2(n19698), .ZN(n19659) );
  OAI211_X1 U22686 ( .C1(n19702), .C2(n19667), .A(n19660), .B(n19659), .ZN(
        P2_U3154) );
  AOI22_X1 U22687 ( .A1(n19670), .A2(n19726), .B1(n19725), .B2(n19686), .ZN(
        n19662) );
  AOI22_X1 U22688 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19672), .B1(
        n19671), .B2(n19727), .ZN(n19661) );
  OAI211_X1 U22689 ( .C1(n19730), .C2(n19709), .A(n19662), .B(n19661), .ZN(
        P2_U3155) );
  AOI22_X1 U22690 ( .A1(n19670), .A2(n19732), .B1(n19731), .B2(n19686), .ZN(
        n19664) );
  AOI22_X1 U22691 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19672), .B1(
        n19671), .B2(n19733), .ZN(n19663) );
  OAI211_X1 U22692 ( .C1(n19736), .C2(n19709), .A(n19664), .B(n19663), .ZN(
        P2_U3156) );
  AOI22_X1 U22693 ( .A1(n19670), .A2(n19738), .B1(n19737), .B2(n19686), .ZN(
        n19666) );
  AOI22_X1 U22694 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19672), .B1(
        n19713), .B2(n19739), .ZN(n19665) );
  OAI211_X1 U22695 ( .C1(n19744), .C2(n19667), .A(n19666), .B(n19665), .ZN(
        P2_U3157) );
  AOI22_X1 U22696 ( .A1(n19670), .A2(n19746), .B1(n19745), .B2(n19686), .ZN(
        n19669) );
  AOI22_X1 U22697 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19672), .B1(
        n19671), .B2(n19747), .ZN(n19668) );
  OAI211_X1 U22698 ( .C1(n19750), .C2(n19709), .A(n19669), .B(n19668), .ZN(
        P2_U3158) );
  AOI22_X1 U22699 ( .A1(n19670), .A2(n19753), .B1(n19751), .B2(n19686), .ZN(
        n19674) );
  AOI22_X1 U22700 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19672), .B1(
        n19671), .B2(n19755), .ZN(n19673) );
  OAI211_X1 U22701 ( .C1(n19761), .C2(n19709), .A(n19674), .B(n19673), .ZN(
        P2_U3159) );
  NOR2_X1 U22702 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19675), .ZN(
        n19712) );
  AOI22_X1 U22703 ( .A1(n19677), .A2(n19713), .B1(n19676), .B2(n19712), .ZN(
        n19692) );
  NAND3_X1 U22704 ( .A1(n19743), .A2(n19709), .A3(n19856), .ZN(n19679) );
  NAND2_X1 U22705 ( .A1(n19679), .A2(n19678), .ZN(n19685) );
  INV_X1 U22706 ( .A(n19686), .ZN(n19682) );
  OAI21_X1 U22707 ( .B1(n19687), .B2(n19544), .A(n19680), .ZN(n19681) );
  AOI21_X1 U22708 ( .B1(n19685), .B2(n19682), .A(n19681), .ZN(n19684) );
  OAI21_X1 U22709 ( .B1(n19712), .B2(n19686), .A(n19685), .ZN(n19689) );
  OAI21_X1 U22710 ( .B1(n19687), .B2(n19712), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19688) );
  AOI22_X1 U22711 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19715), .B1(
        n19690), .B2(n19714), .ZN(n19691) );
  OAI211_X1 U22712 ( .C1(n19693), .C2(n19743), .A(n19692), .B(n19691), .ZN(
        P2_U3160) );
  AOI22_X1 U22713 ( .A1(n19720), .A2(n19756), .B1(n19712), .B2(n19247), .ZN(
        n19695) );
  AOI22_X1 U22714 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19715), .B1(
        n19718), .B2(n19714), .ZN(n19694) );
  OAI211_X1 U22715 ( .C1(n19696), .C2(n19709), .A(n19695), .B(n19694), .ZN(
        P2_U3161) );
  AOI22_X1 U22716 ( .A1(n19698), .A2(n19756), .B1(n19697), .B2(n19712), .ZN(
        n19701) );
  AOI22_X1 U22717 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19715), .B1(
        n19699), .B2(n19714), .ZN(n19700) );
  OAI211_X1 U22718 ( .C1(n19702), .C2(n19709), .A(n19701), .B(n19700), .ZN(
        P2_U3162) );
  AOI22_X1 U22719 ( .A1(n19727), .A2(n19713), .B1(n19712), .B2(n19725), .ZN(
        n19704) );
  AOI22_X1 U22720 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19715), .B1(
        n19726), .B2(n19714), .ZN(n19703) );
  OAI211_X1 U22721 ( .C1(n19730), .C2(n19743), .A(n19704), .B(n19703), .ZN(
        P2_U3163) );
  AOI22_X1 U22722 ( .A1(n19733), .A2(n19713), .B1(n19712), .B2(n19731), .ZN(
        n19706) );
  AOI22_X1 U22723 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19715), .B1(
        n19732), .B2(n19714), .ZN(n19705) );
  OAI211_X1 U22724 ( .C1(n19736), .C2(n19743), .A(n19706), .B(n19705), .ZN(
        P2_U3164) );
  AOI22_X1 U22725 ( .A1(n19739), .A2(n19756), .B1(n19737), .B2(n19712), .ZN(
        n19708) );
  AOI22_X1 U22726 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19715), .B1(
        n19738), .B2(n19714), .ZN(n19707) );
  OAI211_X1 U22727 ( .C1(n19744), .C2(n19709), .A(n19708), .B(n19707), .ZN(
        P2_U3165) );
  AOI22_X1 U22728 ( .A1(n19747), .A2(n19713), .B1(n19745), .B2(n19712), .ZN(
        n19711) );
  AOI22_X1 U22729 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19715), .B1(
        n19746), .B2(n19714), .ZN(n19710) );
  OAI211_X1 U22730 ( .C1(n19750), .C2(n19743), .A(n19711), .B(n19710), .ZN(
        P2_U3166) );
  AOI22_X1 U22731 ( .A1(n19755), .A2(n19713), .B1(n19712), .B2(n19751), .ZN(
        n19717) );
  AOI22_X1 U22732 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19715), .B1(
        n19753), .B2(n19714), .ZN(n19716) );
  OAI211_X1 U22733 ( .C1(n19761), .C2(n19743), .A(n19717), .B(n19716), .ZN(
        P2_U3167) );
  AOI22_X1 U22734 ( .A1(n19754), .A2(n19718), .B1(n19752), .B2(n19247), .ZN(
        n19722) );
  AOI22_X1 U22735 ( .A1(n19740), .A2(n19720), .B1(n19756), .B2(n19719), .ZN(
        n19721) );
  OAI211_X1 U22736 ( .C1(n19724), .C2(n19723), .A(n19722), .B(n19721), .ZN(
        P2_U3169) );
  INV_X1 U22737 ( .A(n19740), .ZN(n19760) );
  AOI22_X1 U22738 ( .A1(n19754), .A2(n19726), .B1(n19752), .B2(n19725), .ZN(
        n19729) );
  AOI22_X1 U22739 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19757), .B1(
        n19756), .B2(n19727), .ZN(n19728) );
  OAI211_X1 U22740 ( .C1(n19730), .C2(n19760), .A(n19729), .B(n19728), .ZN(
        P2_U3171) );
  AOI22_X1 U22741 ( .A1(n19754), .A2(n19732), .B1(n19752), .B2(n19731), .ZN(
        n19735) );
  AOI22_X1 U22742 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19757), .B1(
        n19756), .B2(n19733), .ZN(n19734) );
  OAI211_X1 U22743 ( .C1(n19736), .C2(n19760), .A(n19735), .B(n19734), .ZN(
        P2_U3172) );
  AOI22_X1 U22744 ( .A1(n19754), .A2(n19738), .B1(n19752), .B2(n19737), .ZN(
        n19742) );
  AOI22_X1 U22745 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19757), .B1(
        n19740), .B2(n19739), .ZN(n19741) );
  OAI211_X1 U22746 ( .C1(n19744), .C2(n19743), .A(n19742), .B(n19741), .ZN(
        P2_U3173) );
  AOI22_X1 U22747 ( .A1(n19754), .A2(n19746), .B1(n19752), .B2(n19745), .ZN(
        n19749) );
  AOI22_X1 U22748 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19757), .B1(
        n19756), .B2(n19747), .ZN(n19748) );
  OAI211_X1 U22749 ( .C1(n19750), .C2(n19760), .A(n19749), .B(n19748), .ZN(
        P2_U3174) );
  AOI22_X1 U22750 ( .A1(n19754), .A2(n19753), .B1(n19752), .B2(n19751), .ZN(
        n19759) );
  AOI22_X1 U22751 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19757), .B1(
        n19756), .B2(n19755), .ZN(n19758) );
  OAI211_X1 U22752 ( .C1(n19761), .C2(n19760), .A(n19759), .B(n19758), .ZN(
        P2_U3175) );
  NOR2_X1 U22753 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n18894), .ZN(n19762) );
  OAI211_X1 U22754 ( .C1(n19763), .C2(n19762), .A(n19785), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19770) );
  AND3_X1 U22755 ( .A1(n19765), .A2(n19764), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n19767) );
  OAI21_X1 U22756 ( .B1(n19768), .B2(n19767), .A(n19766), .ZN(n19769) );
  NAND3_X1 U22757 ( .A1(n19771), .A2(n19770), .A3(n19769), .ZN(P2_U3177) );
  AND2_X1 U22758 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19772), .ZN(
        P2_U3179) );
  AND2_X1 U22759 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19772), .ZN(
        P2_U3180) );
  AND2_X1 U22760 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19772), .ZN(
        P2_U3181) );
  AND2_X1 U22761 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19772), .ZN(
        P2_U3182) );
  AND2_X1 U22762 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19772), .ZN(
        P2_U3183) );
  AND2_X1 U22763 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19772), .ZN(
        P2_U3184) );
  AND2_X1 U22764 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19772), .ZN(
        P2_U3185) );
  AND2_X1 U22765 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19772), .ZN(
        P2_U3186) );
  AND2_X1 U22766 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19772), .ZN(
        P2_U3187) );
  AND2_X1 U22767 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19772), .ZN(
        P2_U3188) );
  AND2_X1 U22768 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19772), .ZN(
        P2_U3189) );
  AND2_X1 U22769 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19772), .ZN(
        P2_U3190) );
  AND2_X1 U22770 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19772), .ZN(
        P2_U3191) );
  AND2_X1 U22771 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19772), .ZN(
        P2_U3192) );
  AND2_X1 U22772 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19772), .ZN(
        P2_U3193) );
  AND2_X1 U22773 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19772), .ZN(
        P2_U3194) );
  AND2_X1 U22774 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19772), .ZN(
        P2_U3195) );
  AND2_X1 U22775 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19772), .ZN(
        P2_U3196) );
  AND2_X1 U22776 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19772), .ZN(
        P2_U3197) );
  AND2_X1 U22777 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19772), .ZN(
        P2_U3198) );
  AND2_X1 U22778 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19772), .ZN(
        P2_U3199) );
  AND2_X1 U22779 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19772), .ZN(
        P2_U3200) );
  AND2_X1 U22780 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19772), .ZN(P2_U3201) );
  AND2_X1 U22781 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19772), .ZN(P2_U3202) );
  AND2_X1 U22782 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19772), .ZN(P2_U3203) );
  AND2_X1 U22783 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19772), .ZN(P2_U3204) );
  AND2_X1 U22784 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19772), .ZN(P2_U3205) );
  AND2_X1 U22785 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19772), .ZN(P2_U3206) );
  AND2_X1 U22786 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19772), .ZN(P2_U3207) );
  AND2_X1 U22787 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19772), .ZN(P2_U3208) );
  NAND2_X1 U22788 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19785), .ZN(n19786) );
  NAND3_X1 U22789 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n19786), .ZN(n19775) );
  AOI211_X1 U22790 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n21002), .A(
        n19773), .B(n19891), .ZN(n19774) );
  INV_X1 U22791 ( .A(NA), .ZN(n20753) );
  NOR2_X1 U22792 ( .A1(n20753), .A2(n19779), .ZN(n19791) );
  AOI211_X1 U22793 ( .C1(n19792), .C2(n19775), .A(n19774), .B(n19791), .ZN(
        n19776) );
  INV_X1 U22794 ( .A(n19776), .ZN(P2_U3209) );
  INV_X1 U22795 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19777) );
  AOI21_X1 U22796 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21002), .A(n19792), 
        .ZN(n19783) );
  NOR2_X1 U22797 ( .A1(n19777), .A2(n19783), .ZN(n19780) );
  AOI21_X1 U22798 ( .B1(n19780), .B2(n19779), .A(n19778), .ZN(n19781) );
  OAI211_X1 U22799 ( .C1(n21002), .C2(n19782), .A(n19781), .B(n19786), .ZN(
        P2_U3210) );
  AOI21_X1 U22800 ( .B1(n19785), .B2(n19784), .A(n19783), .ZN(n19790) );
  OAI22_X1 U22801 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19787), .B1(NA), 
        .B2(n19786), .ZN(n19788) );
  OAI211_X1 U22802 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19788), .ZN(n19789) );
  OAI21_X1 U22803 ( .B1(n19791), .B2(n19790), .A(n19789), .ZN(P2_U3211) );
  OAI222_X1 U22804 ( .A1(n19839), .A2(n19795), .B1(n19794), .B2(n19891), .C1(
        n19793), .C2(n19835), .ZN(P2_U3212) );
  OAI222_X1 U22805 ( .A1(n19839), .A2(n19797), .B1(n19796), .B2(n19891), .C1(
        n19795), .C2(n19835), .ZN(P2_U3213) );
  OAI222_X1 U22806 ( .A1(n19839), .A2(n19799), .B1(n19798), .B2(n19891), .C1(
        n19797), .C2(n19835), .ZN(P2_U3214) );
  OAI222_X1 U22807 ( .A1(n19839), .A2(n13857), .B1(n20896), .B2(n19891), .C1(
        n19799), .C2(n19835), .ZN(P2_U3215) );
  OAI222_X1 U22808 ( .A1(n19839), .A2(n19801), .B1(n19800), .B2(n19891), .C1(
        n13857), .C2(n19835), .ZN(P2_U3216) );
  OAI222_X1 U22809 ( .A1(n19839), .A2(n19803), .B1(n19802), .B2(n19891), .C1(
        n19801), .C2(n19835), .ZN(P2_U3217) );
  INV_X1 U22810 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n19805) );
  OAI222_X1 U22811 ( .A1(n19839), .A2(n19805), .B1(n19804), .B2(n19891), .C1(
        n19803), .C2(n19835), .ZN(P2_U3218) );
  OAI222_X1 U22812 ( .A1(n19839), .A2(n19807), .B1(n19806), .B2(n19891), .C1(
        n19805), .C2(n19835), .ZN(P2_U3219) );
  INV_X1 U22813 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n19808) );
  OAI222_X1 U22814 ( .A1(n19839), .A2(n19808), .B1(n21079), .B2(n19891), .C1(
        n19807), .C2(n19835), .ZN(P2_U3220) );
  OAI222_X1 U22815 ( .A1(n19839), .A2(n15101), .B1(n19809), .B2(n19891), .C1(
        n19808), .C2(n19835), .ZN(P2_U3221) );
  OAI222_X1 U22816 ( .A1(n19839), .A2(n14789), .B1(n19810), .B2(n19891), .C1(
        n15101), .C2(n19835), .ZN(P2_U3222) );
  OAI222_X1 U22817 ( .A1(n19839), .A2(n10855), .B1(n19811), .B2(n19891), .C1(
        n14789), .C2(n19835), .ZN(P2_U3223) );
  OAI222_X1 U22818 ( .A1(n19839), .A2(n19813), .B1(n19812), .B2(n19891), .C1(
        n10855), .C2(n19835), .ZN(P2_U3224) );
  OAI222_X1 U22819 ( .A1(n19839), .A2(n15073), .B1(n19814), .B2(n19891), .C1(
        n19813), .C2(n19835), .ZN(P2_U3225) );
  OAI222_X1 U22820 ( .A1(n19839), .A2(n19816), .B1(n19815), .B2(n19891), .C1(
        n15073), .C2(n19835), .ZN(P2_U3226) );
  OAI222_X1 U22821 ( .A1(n19839), .A2(n19818), .B1(n19817), .B2(n19891), .C1(
        n19816), .C2(n19835), .ZN(P2_U3227) );
  INV_X1 U22822 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n21091) );
  OAI222_X1 U22823 ( .A1(n19839), .A2(n21091), .B1(n19819), .B2(n19891), .C1(
        n19818), .C2(n19835), .ZN(P2_U3228) );
  OAI222_X1 U22824 ( .A1(n19839), .A2(n10873), .B1(n19820), .B2(n19891), .C1(
        n21091), .C2(n19835), .ZN(P2_U3229) );
  OAI222_X1 U22825 ( .A1(n19839), .A2(n11289), .B1(n19821), .B2(n19891), .C1(
        n10873), .C2(n19835), .ZN(P2_U3230) );
  OAI222_X1 U22826 ( .A1(n19839), .A2(n19823), .B1(n19822), .B2(n19891), .C1(
        n11289), .C2(n19835), .ZN(P2_U3231) );
  OAI222_X1 U22827 ( .A1(n19839), .A2(n11236), .B1(n19824), .B2(n19891), .C1(
        n19823), .C2(n19835), .ZN(P2_U3232) );
  OAI222_X1 U22828 ( .A1(n19839), .A2(n19825), .B1(n21085), .B2(n19891), .C1(
        n11236), .C2(n19835), .ZN(P2_U3233) );
  OAI222_X1 U22829 ( .A1(n19839), .A2(n11240), .B1(n19826), .B2(n19891), .C1(
        n19825), .C2(n19835), .ZN(P2_U3234) );
  OAI222_X1 U22830 ( .A1(n19839), .A2(n21016), .B1(n19827), .B2(n19891), .C1(
        n11240), .C2(n19835), .ZN(P2_U3235) );
  OAI222_X1 U22831 ( .A1(n19839), .A2(n15000), .B1(n19828), .B2(n19891), .C1(
        n21016), .C2(n19835), .ZN(P2_U3236) );
  OAI222_X1 U22832 ( .A1(n19839), .A2(n19831), .B1(n19829), .B2(n19891), .C1(
        n15000), .C2(n19835), .ZN(P2_U3237) );
  OAI222_X1 U22833 ( .A1(n19835), .A2(n19831), .B1(n19830), .B2(n19891), .C1(
        n12478), .C2(n19839), .ZN(P2_U3238) );
  OAI222_X1 U22834 ( .A1(n19839), .A2(n19833), .B1(n19832), .B2(n19891), .C1(
        n12478), .C2(n19835), .ZN(P2_U3239) );
  OAI222_X1 U22835 ( .A1(n19839), .A2(n19836), .B1(n19834), .B2(n19891), .C1(
        n19833), .C2(n19835), .ZN(P2_U3240) );
  OAI222_X1 U22836 ( .A1(n19839), .A2(n19838), .B1(n19837), .B2(n19891), .C1(
        n19836), .C2(n19835), .ZN(P2_U3241) );
  INV_X1 U22837 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n19840) );
  AOI22_X1 U22838 ( .A1(n19891), .A2(n19841), .B1(n19840), .B2(n19888), .ZN(
        P2_U3585) );
  MUX2_X1 U22839 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n19891), .Z(P2_U3586) );
  INV_X1 U22840 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n19842) );
  AOI22_X1 U22841 ( .A1(n19891), .A2(n19843), .B1(n19842), .B2(n19888), .ZN(
        P2_U3587) );
  INV_X1 U22842 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n19844) );
  AOI22_X1 U22843 ( .A1(n19891), .A2(n19845), .B1(n19844), .B2(n19888), .ZN(
        P2_U3588) );
  OAI21_X1 U22844 ( .B1(n19849), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19847), 
        .ZN(n19846) );
  INV_X1 U22845 ( .A(n19846), .ZN(P2_U3591) );
  OAI21_X1 U22846 ( .B1(n19849), .B2(n19848), .A(n19847), .ZN(P2_U3592) );
  AND2_X1 U22847 ( .A1(n19856), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19872) );
  NAND2_X1 U22848 ( .A1(n19850), .A2(n19872), .ZN(n19862) );
  NAND3_X1 U22849 ( .A1(n19852), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19851), 
        .ZN(n19853) );
  NAND2_X1 U22850 ( .A1(n19853), .A2(n19869), .ZN(n19863) );
  NAND2_X1 U22851 ( .A1(n19862), .A2(n19863), .ZN(n19859) );
  INV_X1 U22852 ( .A(n19854), .ZN(n19858) );
  AOI222_X1 U22853 ( .A1(n19859), .A2(n19858), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n19857), .C1(n19856), .C2(n19855), .ZN(n19860) );
  AOI22_X1 U22854 ( .A1(n19884), .A2(n19861), .B1(n19860), .B2(n19885), .ZN(
        P2_U3602) );
  OAI21_X1 U22855 ( .B1(n19864), .B2(n19863), .A(n19862), .ZN(n19865) );
  AOI21_X1 U22856 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19866), .A(n19865), 
        .ZN(n19867) );
  AOI22_X1 U22857 ( .A1(n19884), .A2(n19868), .B1(n19867), .B2(n19885), .ZN(
        P2_U3603) );
  INV_X1 U22858 ( .A(n19869), .ZN(n19880) );
  AND2_X1 U22859 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19870) );
  NOR2_X1 U22860 ( .A1(n19880), .A2(n19870), .ZN(n19873) );
  MUX2_X1 U22861 ( .A(n19873), .B(n19872), .S(n19871), .Z(n19874) );
  AOI21_X1 U22862 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19875), .A(n19874), 
        .ZN(n19876) );
  AOI22_X1 U22863 ( .A1(n19884), .A2(n19877), .B1(n19876), .B2(n19885), .ZN(
        P2_U3604) );
  NAND3_X1 U22864 ( .A1(n19878), .A2(P2_STATE2_REG_1__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n19879) );
  OAI21_X1 U22865 ( .B1(n19881), .B2(n19880), .A(n19879), .ZN(n19882) );
  AOI21_X1 U22866 ( .B1(n19886), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19882), 
        .ZN(n19883) );
  OAI22_X1 U22867 ( .A1(n19886), .A2(n19885), .B1(n19884), .B2(n19883), .ZN(
        P2_U3605) );
  INV_X1 U22868 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19887) );
  AOI22_X1 U22869 ( .A1(n19891), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19887), 
        .B2(n19888), .ZN(P2_U3608) );
  INV_X1 U22870 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n19889) );
  AOI22_X1 U22871 ( .A1(n19891), .A2(n19890), .B1(n19889), .B2(n19888), .ZN(
        P2_U3611) );
  INV_X1 U22872 ( .A(n19892), .ZN(n19901) );
  INV_X1 U22873 ( .A(n19893), .ZN(n19894) );
  AOI21_X1 U22874 ( .B1(P1_MEMORYFETCH_REG_SCAN_IN), .B2(n19895), .A(n19894), 
        .ZN(n19896) );
  NAND2_X1 U22875 ( .A1(n19901), .A2(n19896), .ZN(P1_U2801) );
  AND2_X1 U22876 ( .A1(n20748), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n19898) );
  INV_X1 U22877 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19897) );
  INV_X2 U22878 ( .A(n20833), .ZN(n20800) );
  AOI21_X1 U22879 ( .B1(n19898), .B2(n19897), .A(n20800), .ZN(P1_U2802) );
  OAI21_X1 U22880 ( .B1(n10129), .B2(n19899), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19900) );
  OAI21_X1 U22881 ( .B1(n19901), .B2(n11495), .A(n19900), .ZN(P1_U2803) );
  NOR2_X1 U22882 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19903) );
  OAI21_X1 U22883 ( .B1(n19903), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20833), .ZN(
        n19902) );
  OAI21_X1 U22884 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20833), .A(n19902), 
        .ZN(P1_U2804) );
  AOI21_X1 U22885 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20748), .A(n20800), 
        .ZN(n20818) );
  OAI21_X1 U22886 ( .B1(BS16), .B2(n19903), .A(n20818), .ZN(n20816) );
  OAI21_X1 U22887 ( .B1(n20818), .B2(n20643), .A(n20816), .ZN(P1_U2805) );
  INV_X1 U22888 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19905) );
  OAI21_X1 U22889 ( .B1(n19906), .B2(n19905), .A(n19904), .ZN(P1_U2806) );
  NOR4_X1 U22890 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_19__SCAN_IN), .A3(P1_DATAWIDTH_REG_20__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_21__SCAN_IN), .ZN(n19910) );
  NOR4_X1 U22891 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_14__SCAN_IN), .A3(P1_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_17__SCAN_IN), .ZN(n19909) );
  NOR4_X1 U22892 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19908) );
  NOR4_X1 U22893 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_23__SCAN_IN), .A3(P1_DATAWIDTH_REG_24__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_25__SCAN_IN), .ZN(n19907) );
  NAND4_X1 U22894 ( .A1(n19910), .A2(n19909), .A3(n19908), .A4(n19907), .ZN(
        n19916) );
  NOR4_X1 U22895 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_27__SCAN_IN), .A3(P1_DATAWIDTH_REG_2__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n19914) );
  AOI211_X1 U22896 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_26__SCAN_IN), .B(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n19913) );
  NOR4_X1 U22897 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_12__SCAN_IN), .ZN(n19912) );
  NOR4_X1 U22898 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19911) );
  NAND4_X1 U22899 ( .A1(n19914), .A2(n19913), .A3(n19912), .A4(n19911), .ZN(
        n19915) );
  NOR2_X1 U22900 ( .A1(n19916), .A2(n19915), .ZN(n20832) );
  INV_X1 U22901 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20811) );
  NOR3_X1 U22902 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19918) );
  OAI21_X1 U22903 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19918), .A(n20832), .ZN(
        n19917) );
  OAI21_X1 U22904 ( .B1(n20832), .B2(n20811), .A(n19917), .ZN(P1_U2807) );
  INV_X1 U22905 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20817) );
  AOI21_X1 U22906 ( .B1(n13735), .B2(n20817), .A(n19918), .ZN(n19919) );
  INV_X1 U22907 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21081) );
  INV_X1 U22908 ( .A(n20832), .ZN(n20827) );
  AOI22_X1 U22909 ( .A1(n20832), .A2(n19919), .B1(n21081), .B2(n20827), .ZN(
        P1_U2808) );
  AOI22_X1 U22910 ( .A1(n19942), .A2(P1_EBX_REG_9__SCAN_IN), .B1(n19974), .B2(
        n19984), .ZN(n19920) );
  OAI211_X1 U22911 ( .C1(n19931), .C2(n19921), .A(n19920), .B(n19969), .ZN(
        n19922) );
  AOI221_X1 U22912 ( .B1(n19924), .B2(P1_REIP_REG_9__SCAN_IN), .C1(n19923), 
        .C2(n13899), .A(n19922), .ZN(n19929) );
  OAI22_X1 U22913 ( .A1(n19987), .A2(n19926), .B1(n19983), .B2(n19925), .ZN(
        n19927) );
  INV_X1 U22914 ( .A(n19927), .ZN(n19928) );
  NAND2_X1 U22915 ( .A1(n19929), .A2(n19928), .ZN(P1_U2831) );
  NAND2_X1 U22916 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n19934) );
  NOR3_X1 U22917 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19954), .A3(n19934), .ZN(
        n19933) );
  AOI22_X1 U22918 ( .A1(n19942), .A2(P1_EBX_REG_7__SCAN_IN), .B1(n19974), .B2(
        n9862), .ZN(n19930) );
  OAI211_X1 U22919 ( .C1(n19931), .C2(n21005), .A(n19930), .B(n19969), .ZN(
        n19932) );
  NOR2_X1 U22920 ( .A1(n19933), .A2(n19932), .ZN(n19939) );
  INV_X1 U22921 ( .A(n19934), .ZN(n19936) );
  AOI21_X1 U22922 ( .B1(n19964), .B2(n19963), .A(n19935), .ZN(n19967) );
  OAI21_X1 U22923 ( .B1(n19937), .B2(n19936), .A(n19967), .ZN(n19948) );
  AOI22_X1 U22924 ( .A1(n19991), .A2(n19949), .B1(P1_REIP_REG_7__SCAN_IN), 
        .B2(n19948), .ZN(n19938) );
  OAI211_X1 U22925 ( .C1(n19940), .C2(n19983), .A(n19939), .B(n19938), .ZN(
        P1_U2833) );
  NOR2_X1 U22926 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n19954), .ZN(n19941) );
  AOI22_X1 U22927 ( .A1(n19942), .A2(P1_EBX_REG_6__SCAN_IN), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n19941), .ZN(n19943) );
  OAI21_X1 U22928 ( .B1(n19945), .B2(n19944), .A(n19943), .ZN(n19946) );
  AOI211_X1 U22929 ( .C1(n19960), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n19947), .B(n19946), .ZN(n19952) );
  AOI22_X1 U22930 ( .A1(n19950), .A2(n19949), .B1(P1_REIP_REG_6__SCAN_IN), 
        .B2(n19948), .ZN(n19951) );
  OAI211_X1 U22931 ( .C1(n19953), .C2(n19983), .A(n19952), .B(n19951), .ZN(
        P1_U2834) );
  OAI22_X1 U22932 ( .A1(n19954), .A2(P1_REIP_REG_5__SCAN_IN), .B1(n19999), 
        .B2(n19977), .ZN(n19957) );
  INV_X1 U22933 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20763) );
  AOI22_X1 U22934 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n19960), .B1(
        n19974), .B2(n19994), .ZN(n19955) );
  OAI211_X1 U22935 ( .C1(n19967), .C2(n20763), .A(n19955), .B(n19969), .ZN(
        n19956) );
  AOI211_X1 U22936 ( .C1(n19997), .C2(n19980), .A(n19957), .B(n19956), .ZN(
        n19958) );
  OAI21_X1 U22937 ( .B1(n19959), .B2(n19983), .A(n19958), .ZN(P1_U2835) );
  NAND2_X1 U22938 ( .A1(n19960), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19972) );
  NAND2_X1 U22939 ( .A1(n19962), .A2(n19961), .ZN(n19971) );
  INV_X1 U22940 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20761) );
  NAND2_X1 U22941 ( .A1(n19964), .A2(n19963), .ZN(n19966) );
  NAND3_X1 U22942 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n19965) );
  OAI22_X1 U22943 ( .A1(n20761), .A2(n19967), .B1(n19966), .B2(n19965), .ZN(
        n19968) );
  INV_X1 U22944 ( .A(n19968), .ZN(n19970) );
  AND4_X1 U22945 ( .A1(n19972), .A2(n19971), .A3(n19970), .A4(n19969), .ZN(
        n19976) );
  INV_X1 U22946 ( .A(n20058), .ZN(n19973) );
  NAND2_X1 U22947 ( .A1(n19974), .A2(n19973), .ZN(n19975) );
  OAI211_X1 U22948 ( .C1(n19978), .C2(n19977), .A(n19976), .B(n19975), .ZN(
        n19979) );
  INV_X1 U22949 ( .A(n19979), .ZN(n19982) );
  NAND2_X1 U22950 ( .A1(n20044), .A2(n19980), .ZN(n19981) );
  OAI211_X1 U22951 ( .C1(n19983), .C2(n20049), .A(n19982), .B(n19981), .ZN(
        P1_U2836) );
  INV_X1 U22952 ( .A(n19984), .ZN(n19985) );
  OAI22_X1 U22953 ( .A1(n19987), .A2(n14389), .B1(n19986), .B2(n19985), .ZN(
        n19988) );
  INV_X1 U22954 ( .A(n19988), .ZN(n19989) );
  OAI21_X1 U22955 ( .B1(n20000), .B2(n19990), .A(n19989), .ZN(P1_U2863) );
  AOI22_X1 U22956 ( .A1(n19991), .A2(n19996), .B1(n19995), .B2(n9862), .ZN(
        n19992) );
  OAI21_X1 U22957 ( .B1(n20000), .B2(n19993), .A(n19992), .ZN(P1_U2865) );
  AOI22_X1 U22958 ( .A1(n19997), .A2(n19996), .B1(n19995), .B2(n19994), .ZN(
        n19998) );
  OAI21_X1 U22959 ( .B1(n20000), .B2(n19999), .A(n19998), .ZN(P1_U2867) );
  OAI222_X1 U22960 ( .A1(n20005), .A2(n20004), .B1(n20003), .B2(n20122), .C1(
        n20002), .C2(n20001), .ZN(P1_U2904) );
  AOI22_X1 U22961 ( .A1(n20008), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(
        P1_EAX_REG_15__SCAN_IN), .B2(n20007), .ZN(n20009) );
  OAI21_X1 U22962 ( .B1(n20010), .B2(n20837), .A(n20009), .ZN(P1_U2921) );
  AOI22_X1 U22963 ( .A1(n20036), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n9761), .ZN(n20012) );
  NAND2_X1 U22964 ( .A1(n20022), .A2(n20011), .ZN(n20024) );
  NAND2_X1 U22965 ( .A1(n20012), .A2(n20024), .ZN(P1_U2945) );
  AOI22_X1 U22966 ( .A1(n20036), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n9761), .ZN(n20014) );
  NAND2_X1 U22967 ( .A1(n20022), .A2(n20013), .ZN(n20026) );
  NAND2_X1 U22968 ( .A1(n20014), .A2(n20026), .ZN(P1_U2946) );
  AOI22_X1 U22969 ( .A1(n20036), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n9761), .ZN(n20016) );
  NAND2_X1 U22970 ( .A1(n20022), .A2(n20015), .ZN(n20028) );
  NAND2_X1 U22971 ( .A1(n20016), .A2(n20028), .ZN(P1_U2947) );
  AOI22_X1 U22972 ( .A1(n20036), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n9761), .ZN(n20018) );
  NAND2_X1 U22973 ( .A1(n20022), .A2(n20017), .ZN(n20032) );
  NAND2_X1 U22974 ( .A1(n20018), .A2(n20032), .ZN(P1_U2949) );
  AOI22_X1 U22975 ( .A1(n20036), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n9761), .ZN(n20020) );
  NAND2_X1 U22976 ( .A1(n20022), .A2(n20019), .ZN(n20034) );
  NAND2_X1 U22977 ( .A1(n20020), .A2(n20034), .ZN(P1_U2950) );
  AOI22_X1 U22978 ( .A1(n20036), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n9761), .ZN(n20023) );
  NAND2_X1 U22979 ( .A1(n20022), .A2(n20021), .ZN(n20037) );
  NAND2_X1 U22980 ( .A1(n20023), .A2(n20037), .ZN(P1_U2951) );
  AOI22_X1 U22981 ( .A1(n20036), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n9761), .ZN(n20025) );
  NAND2_X1 U22982 ( .A1(n20025), .A2(n20024), .ZN(P1_U2960) );
  AOI22_X1 U22983 ( .A1(n20036), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n9761), .ZN(n20027) );
  NAND2_X1 U22984 ( .A1(n20027), .A2(n20026), .ZN(P1_U2961) );
  AOI22_X1 U22985 ( .A1(n20036), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n9761), .ZN(n20029) );
  NAND2_X1 U22986 ( .A1(n20029), .A2(n20028), .ZN(P1_U2962) );
  AOI22_X1 U22987 ( .A1(n20036), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n9761), .ZN(n20031) );
  NAND2_X1 U22988 ( .A1(n20031), .A2(n20030), .ZN(P1_U2963) );
  AOI22_X1 U22989 ( .A1(n20036), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n9761), .ZN(n20033) );
  NAND2_X1 U22990 ( .A1(n20033), .A2(n20032), .ZN(P1_U2964) );
  AOI22_X1 U22991 ( .A1(n20036), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n9761), .ZN(n20035) );
  NAND2_X1 U22992 ( .A1(n20035), .A2(n20034), .ZN(P1_U2965) );
  AOI22_X1 U22993 ( .A1(n20036), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n9761), .ZN(n20038) );
  NAND2_X1 U22994 ( .A1(n20038), .A2(n20037), .ZN(P1_U2966) );
  AOI22_X1 U22995 ( .A1(n20039), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20099), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20048) );
  OAI21_X1 U22996 ( .B1(n20042), .B2(n20041), .A(n20040), .ZN(n20043) );
  INV_X1 U22997 ( .A(n20043), .ZN(n20060) );
  AOI22_X1 U22998 ( .A1(n20060), .A2(n20046), .B1(n20045), .B2(n20044), .ZN(
        n20047) );
  OAI211_X1 U22999 ( .C1(n20050), .C2(n20049), .A(n20048), .B(n20047), .ZN(
        P1_U2995) );
  NOR2_X1 U23000 ( .A1(n20072), .A2(n20051), .ZN(n20074) );
  OAI21_X1 U23001 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n20053), .A(
        n20052), .ZN(n20080) );
  AOI211_X1 U23002 ( .C1(n20082), .C2(n20054), .A(n20074), .B(n20080), .ZN(
        n20070) );
  AOI211_X1 U23003 ( .C1(n20062), .C2(n20069), .A(n20055), .B(n20065), .ZN(
        n20056) );
  AOI21_X1 U23004 ( .B1(n20099), .B2(P1_REIP_REG_4__SCAN_IN), .A(n20056), .ZN(
        n20057) );
  OAI21_X1 U23005 ( .B1(n20102), .B2(n20058), .A(n20057), .ZN(n20059) );
  AOI21_X1 U23006 ( .B1(n20060), .B2(n20079), .A(n20059), .ZN(n20061) );
  OAI21_X1 U23007 ( .B1(n20070), .B2(n20062), .A(n20061), .ZN(P1_U3027) );
  AOI22_X1 U23008 ( .A1(n20099), .A2(P1_REIP_REG_3__SCAN_IN), .B1(n20076), 
        .B2(n20063), .ZN(n20068) );
  OAI22_X1 U23009 ( .A1(n20065), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        n20064), .B2(n20088), .ZN(n20066) );
  INV_X1 U23010 ( .A(n20066), .ZN(n20067) );
  OAI211_X1 U23011 ( .C1(n20070), .C2(n20069), .A(n20068), .B(n20067), .ZN(
        P1_U3028) );
  NOR3_X1 U23012 ( .A1(n20095), .A2(n20072), .A3(n20071), .ZN(n20073) );
  AOI211_X1 U23013 ( .C1(n20076), .C2(n20075), .A(n20074), .B(n20073), .ZN(
        n20086) );
  INV_X1 U23014 ( .A(n20077), .ZN(n20078) );
  AOI22_X1 U23015 ( .A1(n20080), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20079), .B2(n20078), .ZN(n20085) );
  NAND2_X1 U23016 ( .A1(n20099), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n20084) );
  NAND3_X1 U23017 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20082), .A3(
        n20081), .ZN(n20083) );
  NAND4_X1 U23018 ( .A1(n20086), .A2(n20085), .A3(n20084), .A4(n20083), .ZN(
        P1_U3029) );
  NOR2_X1 U23019 ( .A1(n20088), .A2(n20087), .ZN(n20098) );
  INV_X1 U23020 ( .A(n20089), .ZN(n20091) );
  AOI21_X1 U23021 ( .B1(n20092), .B2(n20091), .A(n20090), .ZN(n20097) );
  AOI211_X1 U23022 ( .C1(n20095), .C2(n20094), .A(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n20093), .ZN(n20096) );
  AOI211_X1 U23023 ( .C1(n20098), .C2(n13300), .A(n20097), .B(n20096), .ZN(
        n20101) );
  NAND2_X1 U23024 ( .A1(n20099), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20100) );
  OAI211_X1 U23025 ( .C1(n20103), .C2(n20102), .A(n20101), .B(n20100), .ZN(
        P1_U3030) );
  NOR2_X1 U23026 ( .A1(n20105), .A2(n20104), .ZN(P1_U3032) );
  NAND2_X1 U23027 ( .A1(n20417), .A2(n20472), .ZN(n20296) );
  NAND2_X1 U23028 ( .A1(n20123), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20641) );
  NAND2_X1 U23029 ( .A1(n20299), .A2(n20641), .ZN(n20419) );
  INV_X1 U23030 ( .A(n13420), .ZN(n20106) );
  INV_X1 U23031 ( .A(n20548), .ZN(n20108) );
  OAI21_X1 U23032 ( .B1(n20205), .B2(n20717), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20110) );
  NAND2_X1 U23033 ( .A1(n20110), .A2(n20613), .ZN(n20126) );
  OR2_X1 U23034 ( .A1(n20416), .A2(n20111), .ZN(n20220) );
  NAND2_X1 U23035 ( .A1(n20260), .A2(n20642), .ZN(n20125) );
  INV_X1 U23036 ( .A(n20125), .ZN(n20112) );
  NAND3_X1 U23037 ( .A1(n20515), .A2(n11766), .A3(n20555), .ZN(n20189) );
  NOR2_X1 U23038 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20189), .ZN(
        n20120) );
  OAI22_X1 U23039 ( .A1(n20126), .A2(n20112), .B1(n20120), .B2(n21100), .ZN(
        n20113) );
  INV_X1 U23040 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n20130) );
  INV_X1 U23041 ( .A(n20172), .ZN(n20175) );
  INV_X1 U23042 ( .A(DATAI_24_), .ZN(n20117) );
  OAI22_X2 U23043 ( .A1(n20118), .A2(n20175), .B1(n20117), .B2(n20174), .ZN(
        n20686) );
  INV_X1 U23044 ( .A(n20686), .ZN(n20255) );
  NAND2_X1 U23045 ( .A1(n20177), .A2(n11464), .ZN(n20556) );
  INV_X1 U23046 ( .A(n20120), .ZN(n20178) );
  OAI22_X1 U23047 ( .A1(n20737), .A2(n20255), .B1(n20556), .B2(n20178), .ZN(
        n20121) );
  INV_X1 U23048 ( .A(n20121), .ZN(n20129) );
  NOR2_X2 U23049 ( .A1(n20122), .A2(n20182), .ZN(n20677) );
  INV_X1 U23050 ( .A(n20123), .ZN(n20124) );
  NAND2_X1 U23051 ( .A1(n20124), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20471) );
  AOI22_X2 U23052 ( .A1(DATAI_16_), .A2(n20173), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n20172), .ZN(n20689) );
  INV_X1 U23053 ( .A(n20689), .ZN(n20127) );
  AOI22_X1 U23054 ( .A1(n20677), .A2(n20183), .B1(n20205), .B2(n20127), .ZN(
        n20128) );
  OAI211_X1 U23055 ( .C1(n20180), .C2(n20130), .A(n20129), .B(n20128), .ZN(
        P1_U3033) );
  INV_X1 U23056 ( .A(DATAI_25_), .ZN(n20131) );
  OAI22_X2 U23057 ( .A1(n14943), .A2(n20175), .B1(n20131), .B2(n20174), .ZN(
        n20692) );
  INV_X1 U23058 ( .A(n20692), .ZN(n20485) );
  NAND2_X1 U23059 ( .A1(n20177), .A2(n12355), .ZN(n20567) );
  OAI22_X1 U23060 ( .A1(n20737), .A2(n20485), .B1(n20567), .B2(n20178), .ZN(
        n20132) );
  INV_X1 U23061 ( .A(n20132), .ZN(n20135) );
  NOR2_X2 U23062 ( .A1(n20133), .A2(n20182), .ZN(n20690) );
  AOI22_X2 U23063 ( .A1(DATAI_17_), .A2(n20173), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n20172), .ZN(n20695) );
  INV_X1 U23064 ( .A(n20695), .ZN(n20487) );
  AOI22_X1 U23065 ( .A1(n20690), .A2(n20183), .B1(n20205), .B2(n20487), .ZN(
        n20134) );
  OAI211_X1 U23066 ( .C1(n20180), .C2(n11543), .A(n20135), .B(n20134), .ZN(
        P1_U3034) );
  AOI22_X2 U23067 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20172), .B1(DATAI_26_), 
        .B2(n20173), .ZN(n20701) );
  NAND2_X1 U23068 ( .A1(n20177), .A2(n20136), .ZN(n20572) );
  OAI22_X1 U23069 ( .A1(n20737), .A2(n20701), .B1(n20572), .B2(n20178), .ZN(
        n20137) );
  INV_X1 U23070 ( .A(n20137), .ZN(n20142) );
  NOR2_X2 U23071 ( .A1(n20138), .A2(n20182), .ZN(n20696) );
  INV_X1 U23072 ( .A(DATAI_18_), .ZN(n20140) );
  OAI22_X2 U23073 ( .A1(n20140), .A2(n20174), .B1(n20139), .B2(n20175), .ZN(
        n20698) );
  AOI22_X1 U23074 ( .A1(n20696), .A2(n20183), .B1(n20205), .B2(n20698), .ZN(
        n20141) );
  OAI211_X1 U23075 ( .C1(n20180), .C2(n20143), .A(n20142), .B(n20141), .ZN(
        P1_U3035) );
  INV_X1 U23076 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n20151) );
  INV_X1 U23077 ( .A(DATAI_27_), .ZN(n20144) );
  OAI22_X2 U23078 ( .A1(n21078), .A2(n20175), .B1(n20144), .B2(n20174), .ZN(
        n20704) );
  INV_X1 U23079 ( .A(n20704), .ZN(n20275) );
  NAND2_X1 U23080 ( .A1(n20177), .A2(n20145), .ZN(n20579) );
  OAI22_X1 U23081 ( .A1(n20737), .A2(n20275), .B1(n20579), .B2(n20178), .ZN(
        n20146) );
  INV_X1 U23082 ( .A(n20146), .ZN(n20150) );
  NOR2_X2 U23083 ( .A1(n20147), .A2(n20182), .ZN(n20702) );
  AOI22_X2 U23084 ( .A1(DATAI_19_), .A2(n20173), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n20172), .ZN(n20707) );
  INV_X1 U23085 ( .A(n20707), .ZN(n20148) );
  AOI22_X1 U23086 ( .A1(n20702), .A2(n20183), .B1(n20205), .B2(n20148), .ZN(
        n20149) );
  OAI211_X1 U23087 ( .C1(n20180), .C2(n20151), .A(n20150), .B(n20149), .ZN(
        P1_U3036) );
  AOI22_X2 U23088 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20172), .B1(DATAI_28_), 
        .B2(n20173), .ZN(n20713) );
  NAND2_X1 U23089 ( .A1(n20177), .A2(n20152), .ZN(n20584) );
  OAI22_X1 U23090 ( .A1(n20737), .A2(n20713), .B1(n20584), .B2(n20178), .ZN(
        n20153) );
  INV_X1 U23091 ( .A(n20153), .ZN(n20158) );
  NOR2_X2 U23092 ( .A1(n20154), .A2(n20182), .ZN(n20708) );
  INV_X1 U23093 ( .A(DATAI_20_), .ZN(n20156) );
  OAI22_X2 U23094 ( .A1(n20156), .A2(n20174), .B1(n20155), .B2(n20175), .ZN(
        n20710) );
  AOI22_X1 U23095 ( .A1(n20708), .A2(n20183), .B1(n20205), .B2(n20710), .ZN(
        n20157) );
  OAI211_X1 U23096 ( .C1(n20180), .C2(n20159), .A(n20158), .B(n20157), .ZN(
        P1_U3037) );
  AOI22_X1 U23097 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20172), .B1(DATAI_29_), 
        .B2(n20173), .ZN(n20721) );
  NAND2_X1 U23098 ( .A1(n20177), .A2(n20160), .ZN(n20591) );
  OAI22_X1 U23099 ( .A1(n20737), .A2(n20721), .B1(n20591), .B2(n20178), .ZN(
        n20161) );
  INV_X1 U23100 ( .A(n20161), .ZN(n20164) );
  NOR2_X2 U23101 ( .A1(n20162), .A2(n20182), .ZN(n20714) );
  AOI22_X2 U23102 ( .A1(DATAI_21_), .A2(n20173), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n20172), .ZN(n20665) );
  INV_X1 U23103 ( .A(n20665), .ZN(n20716) );
  AOI22_X1 U23104 ( .A1(n20714), .A2(n20183), .B1(n20205), .B2(n20716), .ZN(
        n20163) );
  OAI211_X1 U23105 ( .C1(n20180), .C2(n11623), .A(n20164), .B(n20163), .ZN(
        P1_U3038) );
  INV_X1 U23106 ( .A(DATAI_30_), .ZN(n20165) );
  OAI22_X2 U23107 ( .A1(n20166), .A2(n20175), .B1(n20165), .B2(n20174), .ZN(
        n20724) );
  INV_X1 U23108 ( .A(n20724), .ZN(n20377) );
  NAND2_X1 U23109 ( .A1(n20177), .A2(n11473), .ZN(n20596) );
  OAI22_X1 U23110 ( .A1(n20737), .A2(n20377), .B1(n20596), .B2(n20178), .ZN(
        n20167) );
  INV_X1 U23111 ( .A(n20167), .ZN(n20170) );
  NOR2_X2 U23112 ( .A1(n20168), .A2(n20182), .ZN(n20722) );
  AOI22_X2 U23113 ( .A1(DATAI_22_), .A2(n20173), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n20172), .ZN(n20727) );
  INV_X1 U23114 ( .A(n20727), .ZN(n20379) );
  AOI22_X1 U23115 ( .A1(n20722), .A2(n20183), .B1(n20205), .B2(n20379), .ZN(
        n20169) );
  OAI211_X1 U23116 ( .C1(n20180), .C2(n20171), .A(n20170), .B(n20169), .ZN(
        P1_U3039) );
  AOI22_X1 U23117 ( .A1(DATAI_23_), .A2(n20173), .B1(BUF1_REG_23__SCAN_IN), 
        .B2(n20172), .ZN(n20738) );
  INV_X1 U23118 ( .A(DATAI_31_), .ZN(n20864) );
  OAI22_X1 U23119 ( .A1(n20176), .A2(n20175), .B1(n20864), .B2(n20174), .ZN(
        n20732) );
  INV_X1 U23120 ( .A(n20732), .ZN(n20547) );
  NAND2_X1 U23121 ( .A1(n20177), .A2(n11456), .ZN(n20602) );
  OAI22_X1 U23122 ( .A1(n20737), .A2(n20547), .B1(n20602), .B2(n20178), .ZN(
        n20179) );
  INV_X1 U23123 ( .A(n20179), .ZN(n20186) );
  INV_X1 U23124 ( .A(n20180), .ZN(n20184) );
  NOR2_X2 U23125 ( .A1(n20182), .A2(n20181), .ZN(n20729) );
  AOI22_X1 U23126 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20184), .B1(
        n20729), .B2(n20183), .ZN(n20185) );
  OAI211_X1 U23127 ( .C1(n20738), .C2(n20213), .A(n20186), .B(n20185), .ZN(
        P1_U3040) );
  INV_X1 U23128 ( .A(n20610), .ZN(n20187) );
  NOR2_X1 U23129 ( .A1(n20611), .A2(n20189), .ZN(n20209) );
  INV_X1 U23130 ( .A(n20188), .ZN(n20444) );
  AOI21_X1 U23131 ( .B1(n20260), .B2(n20444), .A(n20209), .ZN(n20190) );
  OAI22_X1 U23132 ( .A1(n20190), .A2(n20836), .B1(n20189), .B2(n20742), .ZN(
        n20208) );
  AOI22_X1 U23133 ( .A1(n20678), .A2(n20209), .B1(n20677), .B2(n20208), .ZN(
        n20194) );
  INV_X1 U23134 ( .A(n20189), .ZN(n20192) );
  OAI21_X1 U23135 ( .B1(n20257), .B2(n20643), .A(n20190), .ZN(n20191) );
  OAI221_X1 U23136 ( .B1(n20613), .B2(n20192), .C1(n20836), .C2(n20191), .A(
        n20684), .ZN(n20210) );
  AOI22_X1 U23137 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20210), .B1(
        n20205), .B2(n20686), .ZN(n20193) );
  OAI211_X1 U23138 ( .C1(n20689), .C2(n20247), .A(n20194), .B(n20193), .ZN(
        P1_U3041) );
  AOI22_X1 U23139 ( .A1(n20691), .A2(n20209), .B1(n20690), .B2(n20208), .ZN(
        n20196) );
  AOI22_X1 U23140 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20210), .B1(
        n20205), .B2(n20692), .ZN(n20195) );
  OAI211_X1 U23141 ( .C1(n20695), .C2(n20247), .A(n20196), .B(n20195), .ZN(
        P1_U3042) );
  AOI22_X1 U23142 ( .A1(n20697), .A2(n20209), .B1(n20696), .B2(n20208), .ZN(
        n20198) );
  AOI22_X1 U23143 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20210), .B1(
        n20217), .B2(n20698), .ZN(n20197) );
  OAI211_X1 U23144 ( .C1(n20701), .C2(n20213), .A(n20198), .B(n20197), .ZN(
        P1_U3043) );
  AOI22_X1 U23145 ( .A1(n20703), .A2(n20209), .B1(n20702), .B2(n20208), .ZN(
        n20200) );
  AOI22_X1 U23146 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20210), .B1(
        n20205), .B2(n20704), .ZN(n20199) );
  OAI211_X1 U23147 ( .C1(n20707), .C2(n20247), .A(n20200), .B(n20199), .ZN(
        P1_U3044) );
  AOI22_X1 U23148 ( .A1(n20709), .A2(n20209), .B1(n20708), .B2(n20208), .ZN(
        n20202) );
  AOI22_X1 U23149 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20210), .B1(
        n20217), .B2(n20710), .ZN(n20201) );
  OAI211_X1 U23150 ( .C1(n20713), .C2(n20213), .A(n20202), .B(n20201), .ZN(
        P1_U3045) );
  AOI22_X1 U23151 ( .A1(n20715), .A2(n20209), .B1(n20714), .B2(n20208), .ZN(
        n20204) );
  INV_X1 U23152 ( .A(n20721), .ZN(n20662) );
  AOI22_X1 U23153 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20210), .B1(
        n20205), .B2(n20662), .ZN(n20203) );
  OAI211_X1 U23154 ( .C1(n20665), .C2(n20247), .A(n20204), .B(n20203), .ZN(
        P1_U3046) );
  AOI22_X1 U23155 ( .A1(n20723), .A2(n20209), .B1(n20722), .B2(n20208), .ZN(
        n20207) );
  AOI22_X1 U23156 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20210), .B1(
        n20205), .B2(n20724), .ZN(n20206) );
  OAI211_X1 U23157 ( .C1(n20727), .C2(n20247), .A(n20207), .B(n20206), .ZN(
        P1_U3047) );
  AOI22_X1 U23158 ( .A1(n20731), .A2(n20209), .B1(n20729), .B2(n20208), .ZN(
        n20212) );
  INV_X1 U23159 ( .A(n20738), .ZN(n20542) );
  AOI22_X1 U23160 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20210), .B1(
        n20217), .B2(n20542), .ZN(n20211) );
  OAI211_X1 U23161 ( .C1(n20547), .C2(n20213), .A(n20212), .B(n20211), .ZN(
        P1_U3048) );
  INV_X1 U23162 ( .A(n20639), .ZN(n20215) );
  NAND3_X1 U23163 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20515), .A3(
        n11766), .ZN(n20264) );
  OR2_X1 U23164 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20264), .ZN(
        n20246) );
  OAI22_X1 U23165 ( .A1(n20247), .A2(n20255), .B1(n20556), .B2(n20246), .ZN(
        n20216) );
  INV_X1 U23166 ( .A(n20216), .ZN(n20227) );
  INV_X1 U23167 ( .A(n20294), .ZN(n20218) );
  OAI21_X1 U23168 ( .B1(n20218), .B2(n20217), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20219) );
  NAND2_X1 U23169 ( .A1(n20219), .A2(n20613), .ZN(n20225) );
  NOR2_X1 U23170 ( .A1(n20220), .A2(n20642), .ZN(n20222) );
  OR2_X1 U23171 ( .A1(n20472), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20223) );
  INV_X1 U23172 ( .A(n20223), .ZN(n20351) );
  NOR2_X1 U23173 ( .A1(n20351), .A2(n20742), .ZN(n20354) );
  AOI211_X1 U23174 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n20246), .A(n20354), 
        .B(n20419), .ZN(n20221) );
  INV_X1 U23175 ( .A(n20222), .ZN(n20224) );
  AOI22_X1 U23176 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20250), .B1(
        n20677), .B2(n20249), .ZN(n20226) );
  OAI211_X1 U23177 ( .C1(n20689), .C2(n20294), .A(n20227), .B(n20226), .ZN(
        P1_U3049) );
  OAI22_X1 U23178 ( .A1(n20247), .A2(n20485), .B1(n20567), .B2(n20246), .ZN(
        n20228) );
  INV_X1 U23179 ( .A(n20228), .ZN(n20230) );
  AOI22_X1 U23180 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20250), .B1(
        n20690), .B2(n20249), .ZN(n20229) );
  OAI211_X1 U23181 ( .C1(n20695), .C2(n20294), .A(n20230), .B(n20229), .ZN(
        P1_U3050) );
  INV_X1 U23182 ( .A(n20698), .ZN(n20573) );
  OAI22_X1 U23183 ( .A1(n20294), .A2(n20573), .B1(n20572), .B2(n20246), .ZN(
        n20231) );
  INV_X1 U23184 ( .A(n20231), .ZN(n20233) );
  AOI22_X1 U23185 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20250), .B1(
        n20696), .B2(n20249), .ZN(n20232) );
  OAI211_X1 U23186 ( .C1(n20701), .C2(n20247), .A(n20233), .B(n20232), .ZN(
        P1_U3051) );
  OAI22_X1 U23187 ( .A1(n20247), .A2(n20275), .B1(n20579), .B2(n20246), .ZN(
        n20234) );
  INV_X1 U23188 ( .A(n20234), .ZN(n20236) );
  AOI22_X1 U23189 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20250), .B1(
        n20702), .B2(n20249), .ZN(n20235) );
  OAI211_X1 U23190 ( .C1(n20707), .C2(n20294), .A(n20236), .B(n20235), .ZN(
        P1_U3052) );
  INV_X1 U23191 ( .A(n20710), .ZN(n20585) );
  OAI22_X1 U23192 ( .A1(n20294), .A2(n20585), .B1(n20584), .B2(n20246), .ZN(
        n20237) );
  INV_X1 U23193 ( .A(n20237), .ZN(n20239) );
  AOI22_X1 U23194 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20250), .B1(
        n20708), .B2(n20249), .ZN(n20238) );
  OAI211_X1 U23195 ( .C1(n20713), .C2(n20247), .A(n20239), .B(n20238), .ZN(
        P1_U3053) );
  OAI22_X1 U23196 ( .A1(n20247), .A2(n20721), .B1(n20591), .B2(n20246), .ZN(
        n20240) );
  INV_X1 U23197 ( .A(n20240), .ZN(n20242) );
  AOI22_X1 U23198 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20250), .B1(
        n20714), .B2(n20249), .ZN(n20241) );
  OAI211_X1 U23199 ( .C1(n20665), .C2(n20294), .A(n20242), .B(n20241), .ZN(
        P1_U3054) );
  OAI22_X1 U23200 ( .A1(n20247), .A2(n20377), .B1(n20596), .B2(n20246), .ZN(
        n20243) );
  INV_X1 U23201 ( .A(n20243), .ZN(n20245) );
  AOI22_X1 U23202 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20250), .B1(
        n20722), .B2(n20249), .ZN(n20244) );
  OAI211_X1 U23203 ( .C1(n20727), .C2(n20294), .A(n20245), .B(n20244), .ZN(
        P1_U3055) );
  OAI22_X1 U23204 ( .A1(n20247), .A2(n20547), .B1(n20602), .B2(n20246), .ZN(
        n20248) );
  INV_X1 U23205 ( .A(n20248), .ZN(n20252) );
  AOI22_X1 U23206 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20250), .B1(
        n20729), .B2(n20249), .ZN(n20251) );
  OAI211_X1 U23207 ( .C1(n20738), .C2(n20294), .A(n20252), .B(n20251), .ZN(
        P1_U3056) );
  INV_X1 U23208 ( .A(n20513), .ZN(n20253) );
  INV_X1 U23209 ( .A(n20516), .ZN(n20254) );
  NAND2_X1 U23210 ( .A1(n20254), .A2(n20515), .ZN(n20288) );
  OAI22_X1 U23211 ( .A1(n20294), .A2(n20255), .B1(n20556), .B2(n20288), .ZN(
        n20256) );
  INV_X1 U23212 ( .A(n20256), .ZN(n20268) );
  OAI21_X1 U23213 ( .B1(n20257), .B2(n20521), .A(n20613), .ZN(n20265) );
  AND2_X1 U23214 ( .A1(n20258), .A2(n11849), .ZN(n20517) );
  INV_X1 U23215 ( .A(n20288), .ZN(n20259) );
  AOI21_X1 U23216 ( .B1(n20260), .B2(n20517), .A(n20259), .ZN(n20266) );
  INV_X1 U23217 ( .A(n20266), .ZN(n20263) );
  AOI21_X1 U23218 ( .B1(n20836), .B2(n20264), .A(n20261), .ZN(n20262) );
  OAI22_X1 U23219 ( .A1(n20266), .A2(n20265), .B1(n20742), .B2(n20264), .ZN(
        n20290) );
  AOI22_X1 U23220 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20291), .B1(
        n20677), .B2(n20290), .ZN(n20267) );
  OAI211_X1 U23221 ( .C1(n20689), .C2(n20311), .A(n20268), .B(n20267), .ZN(
        P1_U3057) );
  OAI22_X1 U23222 ( .A1(n20294), .A2(n20485), .B1(n20567), .B2(n20288), .ZN(
        n20269) );
  INV_X1 U23223 ( .A(n20269), .ZN(n20271) );
  AOI22_X1 U23224 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20291), .B1(
        n20690), .B2(n20290), .ZN(n20270) );
  OAI211_X1 U23225 ( .C1(n20695), .C2(n20311), .A(n20271), .B(n20270), .ZN(
        P1_U3058) );
  OAI22_X1 U23226 ( .A1(n20311), .A2(n20573), .B1(n20572), .B2(n20288), .ZN(
        n20272) );
  INV_X1 U23227 ( .A(n20272), .ZN(n20274) );
  AOI22_X1 U23228 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20291), .B1(
        n20696), .B2(n20290), .ZN(n20273) );
  OAI211_X1 U23229 ( .C1(n20701), .C2(n20294), .A(n20274), .B(n20273), .ZN(
        P1_U3059) );
  OAI22_X1 U23230 ( .A1(n20294), .A2(n20275), .B1(n20579), .B2(n20288), .ZN(
        n20276) );
  INV_X1 U23231 ( .A(n20276), .ZN(n20278) );
  AOI22_X1 U23232 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20291), .B1(
        n20702), .B2(n20290), .ZN(n20277) );
  OAI211_X1 U23233 ( .C1(n20707), .C2(n20311), .A(n20278), .B(n20277), .ZN(
        P1_U3060) );
  OAI22_X1 U23234 ( .A1(n20311), .A2(n20585), .B1(n20584), .B2(n20288), .ZN(
        n20279) );
  INV_X1 U23235 ( .A(n20279), .ZN(n20281) );
  AOI22_X1 U23236 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20291), .B1(
        n20708), .B2(n20290), .ZN(n20280) );
  OAI211_X1 U23237 ( .C1(n20713), .C2(n20294), .A(n20281), .B(n20280), .ZN(
        P1_U3061) );
  OAI22_X1 U23238 ( .A1(n20311), .A2(n20665), .B1(n20591), .B2(n20288), .ZN(
        n20282) );
  INV_X1 U23239 ( .A(n20282), .ZN(n20284) );
  AOI22_X1 U23240 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20291), .B1(
        n20714), .B2(n20290), .ZN(n20283) );
  OAI211_X1 U23241 ( .C1(n20721), .C2(n20294), .A(n20284), .B(n20283), .ZN(
        P1_U3062) );
  OAI22_X1 U23242 ( .A1(n20294), .A2(n20377), .B1(n20596), .B2(n20288), .ZN(
        n20285) );
  INV_X1 U23243 ( .A(n20285), .ZN(n20287) );
  AOI22_X1 U23244 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20291), .B1(
        n20722), .B2(n20290), .ZN(n20286) );
  OAI211_X1 U23245 ( .C1(n20727), .C2(n20311), .A(n20287), .B(n20286), .ZN(
        P1_U3063) );
  OAI22_X1 U23246 ( .A1(n20311), .A2(n20738), .B1(n20602), .B2(n20288), .ZN(
        n20289) );
  INV_X1 U23247 ( .A(n20289), .ZN(n20293) );
  AOI22_X1 U23248 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20291), .B1(
        n20729), .B2(n20290), .ZN(n20292) );
  OAI211_X1 U23249 ( .C1(n20547), .C2(n20294), .A(n20293), .B(n20292), .ZN(
        P1_U3064) );
  NAND3_X1 U23250 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20515), .A3(
        n20555), .ZN(n20324) );
  NOR2_X1 U23251 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20324), .ZN(
        n20317) );
  NOR2_X1 U23252 ( .A1(n20552), .A2(n20295), .ZN(n20350) );
  NAND2_X1 U23253 ( .A1(n20350), .A2(n20613), .ZN(n20390) );
  OAI22_X1 U23254 ( .A1(n20390), .A2(n20645), .B1(n20296), .B2(n20641), .ZN(
        n20316) );
  AOI22_X1 U23255 ( .A1(n20678), .A2(n20317), .B1(n20677), .B2(n20316), .ZN(
        n20302) );
  INV_X1 U23256 ( .A(n20350), .ZN(n20298) );
  OAI21_X1 U23257 ( .B1(n20318), .B2(n20340), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20297) );
  OAI21_X1 U23258 ( .B1(n20645), .B2(n20298), .A(n20297), .ZN(n20300) );
  AOI22_X1 U23259 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20319), .B1(
        n20318), .B2(n20686), .ZN(n20301) );
  OAI211_X1 U23260 ( .C1(n20689), .C2(n20348), .A(n20302), .B(n20301), .ZN(
        P1_U3065) );
  AOI22_X1 U23261 ( .A1(n20691), .A2(n20317), .B1(n20690), .B2(n20316), .ZN(
        n20304) );
  AOI22_X1 U23262 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20319), .B1(
        n20318), .B2(n20692), .ZN(n20303) );
  OAI211_X1 U23263 ( .C1(n20695), .C2(n20348), .A(n20304), .B(n20303), .ZN(
        P1_U3066) );
  AOI22_X1 U23264 ( .A1(n20697), .A2(n20317), .B1(n20696), .B2(n20316), .ZN(
        n20306) );
  AOI22_X1 U23265 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20319), .B1(
        n20340), .B2(n20698), .ZN(n20305) );
  OAI211_X1 U23266 ( .C1(n20701), .C2(n20311), .A(n20306), .B(n20305), .ZN(
        P1_U3067) );
  AOI22_X1 U23267 ( .A1(n20703), .A2(n20317), .B1(n20702), .B2(n20316), .ZN(
        n20308) );
  AOI22_X1 U23268 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20319), .B1(
        n20318), .B2(n20704), .ZN(n20307) );
  OAI211_X1 U23269 ( .C1(n20707), .C2(n20348), .A(n20308), .B(n20307), .ZN(
        P1_U3068) );
  AOI22_X1 U23270 ( .A1(n20709), .A2(n20317), .B1(n20708), .B2(n20316), .ZN(
        n20310) );
  AOI22_X1 U23271 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20319), .B1(
        n20340), .B2(n20710), .ZN(n20309) );
  OAI211_X1 U23272 ( .C1(n20713), .C2(n20311), .A(n20310), .B(n20309), .ZN(
        P1_U3069) );
  AOI22_X1 U23273 ( .A1(n20715), .A2(n20317), .B1(n20714), .B2(n20316), .ZN(
        n20313) );
  AOI22_X1 U23274 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20319), .B1(
        n20318), .B2(n20662), .ZN(n20312) );
  OAI211_X1 U23275 ( .C1(n20665), .C2(n20348), .A(n20313), .B(n20312), .ZN(
        P1_U3070) );
  AOI22_X1 U23276 ( .A1(n20723), .A2(n20317), .B1(n20722), .B2(n20316), .ZN(
        n20315) );
  AOI22_X1 U23277 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20319), .B1(
        n20318), .B2(n20724), .ZN(n20314) );
  OAI211_X1 U23278 ( .C1(n20727), .C2(n20348), .A(n20315), .B(n20314), .ZN(
        P1_U3071) );
  AOI22_X1 U23279 ( .A1(n20731), .A2(n20317), .B1(n20729), .B2(n20316), .ZN(
        n20321) );
  AOI22_X1 U23280 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20319), .B1(
        n20318), .B2(n20732), .ZN(n20320) );
  OAI211_X1 U23281 ( .C1(n20738), .C2(n20348), .A(n20321), .B(n20320), .ZN(
        P1_U3072) );
  NOR2_X1 U23282 ( .A1(n20611), .A2(n20324), .ZN(n20344) );
  INV_X1 U23283 ( .A(n20344), .ZN(n20322) );
  OAI222_X1 U23284 ( .A1(n20322), .A2(n20836), .B1(n20742), .B2(n20324), .C1(
        n20188), .C2(n20390), .ZN(n20343) );
  AOI22_X1 U23285 ( .A1(n20678), .A2(n20344), .B1(n20677), .B2(n20343), .ZN(
        n20329) );
  INV_X1 U23286 ( .A(n20389), .ZN(n20326) );
  INV_X1 U23287 ( .A(n20323), .ZN(n20325) );
  OAI21_X1 U23288 ( .B1(n20326), .B2(n20325), .A(n20324), .ZN(n20327) );
  NAND2_X1 U23289 ( .A1(n20327), .A2(n20684), .ZN(n20345) );
  AOI22_X1 U23290 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20345), .B1(
        n20340), .B2(n20686), .ZN(n20328) );
  OAI211_X1 U23291 ( .C1(n20689), .C2(n20383), .A(n20329), .B(n20328), .ZN(
        P1_U3073) );
  AOI22_X1 U23292 ( .A1(n20691), .A2(n20344), .B1(n20690), .B2(n20343), .ZN(
        n20331) );
  AOI22_X1 U23293 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20345), .B1(
        n20340), .B2(n20692), .ZN(n20330) );
  OAI211_X1 U23294 ( .C1(n20695), .C2(n20383), .A(n20331), .B(n20330), .ZN(
        P1_U3074) );
  AOI22_X1 U23295 ( .A1(n20697), .A2(n20344), .B1(n20696), .B2(n20343), .ZN(
        n20333) );
  AOI22_X1 U23296 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20345), .B1(
        n20371), .B2(n20698), .ZN(n20332) );
  OAI211_X1 U23297 ( .C1(n20701), .C2(n20348), .A(n20333), .B(n20332), .ZN(
        P1_U3075) );
  AOI22_X1 U23298 ( .A1(n20703), .A2(n20344), .B1(n20702), .B2(n20343), .ZN(
        n20335) );
  AOI22_X1 U23299 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20345), .B1(
        n20340), .B2(n20704), .ZN(n20334) );
  OAI211_X1 U23300 ( .C1(n20707), .C2(n20383), .A(n20335), .B(n20334), .ZN(
        P1_U3076) );
  AOI22_X1 U23301 ( .A1(n20709), .A2(n20344), .B1(n20708), .B2(n20343), .ZN(
        n20337) );
  AOI22_X1 U23302 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20345), .B1(
        n20371), .B2(n20710), .ZN(n20336) );
  OAI211_X1 U23303 ( .C1(n20713), .C2(n20348), .A(n20337), .B(n20336), .ZN(
        P1_U3077) );
  AOI22_X1 U23304 ( .A1(n20715), .A2(n20344), .B1(n20714), .B2(n20343), .ZN(
        n20339) );
  AOI22_X1 U23305 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20345), .B1(
        n20340), .B2(n20662), .ZN(n20338) );
  OAI211_X1 U23306 ( .C1(n20665), .C2(n20383), .A(n20339), .B(n20338), .ZN(
        P1_U3078) );
  AOI22_X1 U23307 ( .A1(n20723), .A2(n20344), .B1(n20722), .B2(n20343), .ZN(
        n20342) );
  AOI22_X1 U23308 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20345), .B1(
        n20340), .B2(n20724), .ZN(n20341) );
  OAI211_X1 U23309 ( .C1(n20727), .C2(n20383), .A(n20342), .B(n20341), .ZN(
        P1_U3079) );
  AOI22_X1 U23310 ( .A1(n20731), .A2(n20344), .B1(n20729), .B2(n20343), .ZN(
        n20347) );
  AOI22_X1 U23311 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20345), .B1(
        n20371), .B2(n20542), .ZN(n20346) );
  OAI211_X1 U23312 ( .C1(n20547), .C2(n20348), .A(n20347), .B(n20346), .ZN(
        P1_U3080) );
  NAND2_X1 U23313 ( .A1(n20415), .A2(n20383), .ZN(n20349) );
  AOI21_X1 U23314 ( .B1(n20349), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20836), 
        .ZN(n20356) );
  NAND2_X1 U23315 ( .A1(n20350), .A2(n20645), .ZN(n20355) );
  INV_X1 U23316 ( .A(n20355), .ZN(n20352) );
  INV_X1 U23317 ( .A(n20641), .ZN(n20554) );
  INV_X1 U23318 ( .A(n20677), .ZN(n20566) );
  INV_X1 U23319 ( .A(n20394), .ZN(n20391) );
  NOR2_X1 U23320 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20391), .ZN(
        n20358) );
  INV_X1 U23321 ( .A(n20358), .ZN(n20382) );
  OAI22_X1 U23322 ( .A1(n20415), .A2(n20689), .B1(n20556), .B2(n20382), .ZN(
        n20353) );
  INV_X1 U23323 ( .A(n20353), .ZN(n20360) );
  AOI21_X1 U23324 ( .B1(n20356), .B2(n20355), .A(n20354), .ZN(n20357) );
  OAI211_X1 U23325 ( .C1(n20358), .C2(n21100), .A(n20649), .B(n20357), .ZN(
        n20385) );
  AOI22_X1 U23326 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20385), .B1(
        n20371), .B2(n20686), .ZN(n20359) );
  OAI211_X1 U23327 ( .C1(n20388), .C2(n20566), .A(n20360), .B(n20359), .ZN(
        P1_U3081) );
  INV_X1 U23328 ( .A(n20690), .ZN(n20571) );
  OAI22_X1 U23329 ( .A1(n20383), .A2(n20485), .B1(n20567), .B2(n20382), .ZN(
        n20361) );
  INV_X1 U23330 ( .A(n20361), .ZN(n20363) );
  AOI22_X1 U23331 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20385), .B1(
        n20407), .B2(n20487), .ZN(n20362) );
  OAI211_X1 U23332 ( .C1(n20388), .C2(n20571), .A(n20363), .B(n20362), .ZN(
        P1_U3082) );
  INV_X1 U23333 ( .A(n20696), .ZN(n20578) );
  OAI22_X1 U23334 ( .A1(n20415), .A2(n20573), .B1(n20572), .B2(n20382), .ZN(
        n20364) );
  INV_X1 U23335 ( .A(n20364), .ZN(n20366) );
  INV_X1 U23336 ( .A(n20701), .ZN(n20575) );
  AOI22_X1 U23337 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20385), .B1(
        n20371), .B2(n20575), .ZN(n20365) );
  OAI211_X1 U23338 ( .C1(n20388), .C2(n20578), .A(n20366), .B(n20365), .ZN(
        P1_U3083) );
  INV_X1 U23339 ( .A(n20702), .ZN(n20583) );
  OAI22_X1 U23340 ( .A1(n20415), .A2(n20707), .B1(n20579), .B2(n20382), .ZN(
        n20367) );
  INV_X1 U23341 ( .A(n20367), .ZN(n20369) );
  AOI22_X1 U23342 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20385), .B1(
        n20371), .B2(n20704), .ZN(n20368) );
  OAI211_X1 U23343 ( .C1(n20388), .C2(n20583), .A(n20369), .B(n20368), .ZN(
        P1_U3084) );
  INV_X1 U23344 ( .A(n20708), .ZN(n20590) );
  OAI22_X1 U23345 ( .A1(n20415), .A2(n20585), .B1(n20584), .B2(n20382), .ZN(
        n20370) );
  INV_X1 U23346 ( .A(n20370), .ZN(n20373) );
  INV_X1 U23347 ( .A(n20713), .ZN(n20587) );
  AOI22_X1 U23348 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20385), .B1(
        n20371), .B2(n20587), .ZN(n20372) );
  OAI211_X1 U23349 ( .C1(n20388), .C2(n20590), .A(n20373), .B(n20372), .ZN(
        P1_U3085) );
  INV_X1 U23350 ( .A(n20714), .ZN(n20595) );
  OAI22_X1 U23351 ( .A1(n20383), .A2(n20721), .B1(n20591), .B2(n20382), .ZN(
        n20374) );
  INV_X1 U23352 ( .A(n20374), .ZN(n20376) );
  AOI22_X1 U23353 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20385), .B1(
        n20407), .B2(n20716), .ZN(n20375) );
  OAI211_X1 U23354 ( .C1(n20388), .C2(n20595), .A(n20376), .B(n20375), .ZN(
        P1_U3086) );
  INV_X1 U23355 ( .A(n20722), .ZN(n20600) );
  OAI22_X1 U23356 ( .A1(n20383), .A2(n20377), .B1(n20596), .B2(n20382), .ZN(
        n20378) );
  INV_X1 U23357 ( .A(n20378), .ZN(n20381) );
  AOI22_X1 U23358 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20385), .B1(
        n20407), .B2(n20379), .ZN(n20380) );
  OAI211_X1 U23359 ( .C1(n20388), .C2(n20600), .A(n20381), .B(n20380), .ZN(
        P1_U3087) );
  INV_X1 U23360 ( .A(n20729), .ZN(n20608) );
  OAI22_X1 U23361 ( .A1(n20383), .A2(n20547), .B1(n20602), .B2(n20382), .ZN(
        n20384) );
  INV_X1 U23362 ( .A(n20384), .ZN(n20387) );
  AOI22_X1 U23363 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20385), .B1(
        n20407), .B2(n20542), .ZN(n20386) );
  OAI211_X1 U23364 ( .C1(n20388), .C2(n20608), .A(n20387), .B(n20386), .ZN(
        P1_U3088) );
  INV_X1 U23365 ( .A(n20392), .ZN(n20411) );
  INV_X1 U23366 ( .A(n20517), .ZN(n20675) );
  OAI222_X1 U23367 ( .A1(n20836), .A2(n20392), .B1(n20391), .B2(n20742), .C1(
        n20675), .C2(n20390), .ZN(n20410) );
  AOI22_X1 U23368 ( .A1(n20678), .A2(n20411), .B1(n20677), .B2(n20410), .ZN(
        n20396) );
  AOI22_X1 U23369 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20412), .B1(
        n20407), .B2(n20686), .ZN(n20395) );
  OAI211_X1 U23370 ( .C1(n20689), .C2(n20433), .A(n20396), .B(n20395), .ZN(
        P1_U3089) );
  AOI22_X1 U23371 ( .A1(n20691), .A2(n20411), .B1(n20690), .B2(n20410), .ZN(
        n20398) );
  AOI22_X1 U23372 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20412), .B1(
        n20407), .B2(n20692), .ZN(n20397) );
  OAI211_X1 U23373 ( .C1(n20695), .C2(n20433), .A(n20398), .B(n20397), .ZN(
        P1_U3090) );
  AOI22_X1 U23374 ( .A1(n20697), .A2(n20411), .B1(n20696), .B2(n20410), .ZN(
        n20400) );
  AOI22_X1 U23375 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20412), .B1(
        n20440), .B2(n20698), .ZN(n20399) );
  OAI211_X1 U23376 ( .C1(n20701), .C2(n20415), .A(n20400), .B(n20399), .ZN(
        P1_U3091) );
  AOI22_X1 U23377 ( .A1(n20703), .A2(n20411), .B1(n20702), .B2(n20410), .ZN(
        n20402) );
  AOI22_X1 U23378 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20412), .B1(
        n20407), .B2(n20704), .ZN(n20401) );
  OAI211_X1 U23379 ( .C1(n20707), .C2(n20433), .A(n20402), .B(n20401), .ZN(
        P1_U3092) );
  AOI22_X1 U23380 ( .A1(n20709), .A2(n20411), .B1(n20708), .B2(n20410), .ZN(
        n20404) );
  AOI22_X1 U23381 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20412), .B1(
        n20440), .B2(n20710), .ZN(n20403) );
  OAI211_X1 U23382 ( .C1(n20713), .C2(n20415), .A(n20404), .B(n20403), .ZN(
        P1_U3093) );
  AOI22_X1 U23383 ( .A1(n20715), .A2(n20411), .B1(n20714), .B2(n20410), .ZN(
        n20406) );
  AOI22_X1 U23384 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20412), .B1(
        n20407), .B2(n20662), .ZN(n20405) );
  OAI211_X1 U23385 ( .C1(n20665), .C2(n20433), .A(n20406), .B(n20405), .ZN(
        P1_U3094) );
  AOI22_X1 U23386 ( .A1(n20723), .A2(n20411), .B1(n20722), .B2(n20410), .ZN(
        n20409) );
  AOI22_X1 U23387 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20412), .B1(
        n20407), .B2(n20724), .ZN(n20408) );
  OAI211_X1 U23388 ( .C1(n20727), .C2(n20433), .A(n20409), .B(n20408), .ZN(
        P1_U3095) );
  AOI22_X1 U23389 ( .A1(n20731), .A2(n20411), .B1(n20729), .B2(n20410), .ZN(
        n20414) );
  AOI22_X1 U23390 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20412), .B1(
        n20440), .B2(n20542), .ZN(n20413) );
  OAI211_X1 U23391 ( .C1(n20547), .C2(n20415), .A(n20414), .B(n20413), .ZN(
        P1_U3096) );
  NAND3_X1 U23392 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n11766), .A3(
        n20555), .ZN(n20445) );
  NOR2_X1 U23393 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20445), .ZN(
        n20439) );
  AND2_X1 U23394 ( .A1(n20416), .A2(n20552), .ZN(n20518) );
  AOI21_X1 U23395 ( .B1(n20518), .B2(n20642), .A(n20439), .ZN(n20420) );
  INV_X1 U23396 ( .A(n20472), .ZN(n20418) );
  NOR2_X1 U23397 ( .A1(n20418), .A2(n20417), .ZN(n20553) );
  INV_X1 U23398 ( .A(n20553), .ZN(n20559) );
  OAI22_X1 U23399 ( .A1(n20420), .A2(n20836), .B1(n20471), .B2(n20559), .ZN(
        n20438) );
  AOI22_X1 U23400 ( .A1(n20678), .A2(n20439), .B1(n20677), .B2(n20438), .ZN(
        n20424) );
  INV_X1 U23401 ( .A(n20419), .ZN(n20477) );
  OAI21_X1 U23402 ( .B1(n20466), .B2(n20440), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20421) );
  NAND2_X1 U23403 ( .A1(n20421), .A2(n20420), .ZN(n20422) );
  AOI22_X1 U23404 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20441), .B1(
        n20440), .B2(n20686), .ZN(n20423) );
  OAI211_X1 U23405 ( .C1(n20689), .C2(n20459), .A(n20424), .B(n20423), .ZN(
        P1_U3097) );
  AOI22_X1 U23406 ( .A1(n20691), .A2(n20439), .B1(n20690), .B2(n20438), .ZN(
        n20426) );
  AOI22_X1 U23407 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20441), .B1(
        n20440), .B2(n20692), .ZN(n20425) );
  OAI211_X1 U23408 ( .C1(n20695), .C2(n20459), .A(n20426), .B(n20425), .ZN(
        P1_U3098) );
  AOI22_X1 U23409 ( .A1(n20697), .A2(n20439), .B1(n20696), .B2(n20438), .ZN(
        n20428) );
  AOI22_X1 U23410 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20441), .B1(
        n20466), .B2(n20698), .ZN(n20427) );
  OAI211_X1 U23411 ( .C1(n20701), .C2(n20433), .A(n20428), .B(n20427), .ZN(
        P1_U3099) );
  AOI22_X1 U23412 ( .A1(n20703), .A2(n20439), .B1(n20702), .B2(n20438), .ZN(
        n20430) );
  AOI22_X1 U23413 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20441), .B1(
        n20440), .B2(n20704), .ZN(n20429) );
  OAI211_X1 U23414 ( .C1(n20707), .C2(n20459), .A(n20430), .B(n20429), .ZN(
        P1_U3100) );
  AOI22_X1 U23415 ( .A1(n20709), .A2(n20439), .B1(n20708), .B2(n20438), .ZN(
        n20432) );
  AOI22_X1 U23416 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20441), .B1(
        n20466), .B2(n20710), .ZN(n20431) );
  OAI211_X1 U23417 ( .C1(n20713), .C2(n20433), .A(n20432), .B(n20431), .ZN(
        P1_U3101) );
  AOI22_X1 U23418 ( .A1(n20715), .A2(n20439), .B1(n20714), .B2(n20438), .ZN(
        n20435) );
  AOI22_X1 U23419 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20441), .B1(
        n20440), .B2(n20662), .ZN(n20434) );
  OAI211_X1 U23420 ( .C1(n20665), .C2(n20459), .A(n20435), .B(n20434), .ZN(
        P1_U3102) );
  AOI22_X1 U23421 ( .A1(n20723), .A2(n20439), .B1(n20722), .B2(n20438), .ZN(
        n20437) );
  AOI22_X1 U23422 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20441), .B1(
        n20440), .B2(n20724), .ZN(n20436) );
  OAI211_X1 U23423 ( .C1(n20727), .C2(n20459), .A(n20437), .B(n20436), .ZN(
        P1_U3103) );
  AOI22_X1 U23424 ( .A1(n20731), .A2(n20439), .B1(n20729), .B2(n20438), .ZN(
        n20443) );
  AOI22_X1 U23425 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20441), .B1(
        n20440), .B2(n20732), .ZN(n20442) );
  OAI211_X1 U23426 ( .C1(n20738), .C2(n20459), .A(n20443), .B(n20442), .ZN(
        P1_U3104) );
  NOR2_X1 U23427 ( .A1(n20611), .A2(n20445), .ZN(n20465) );
  AOI21_X1 U23428 ( .B1(n20518), .B2(n20444), .A(n20465), .ZN(n20446) );
  OAI22_X1 U23429 ( .A1(n20446), .A2(n20836), .B1(n20445), .B2(n20742), .ZN(
        n20464) );
  AOI22_X1 U23430 ( .A1(n20678), .A2(n20465), .B1(n20677), .B2(n20464), .ZN(
        n20450) );
  INV_X1 U23431 ( .A(n20445), .ZN(n20448) );
  OAI21_X1 U23432 ( .B1(n20522), .B2(n20643), .A(n20446), .ZN(n20447) );
  OAI221_X1 U23433 ( .B1(n20613), .B2(n20448), .C1(n20836), .C2(n20447), .A(
        n20684), .ZN(n20467) );
  AOI22_X1 U23434 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20467), .B1(
        n20466), .B2(n20686), .ZN(n20449) );
  OAI211_X1 U23435 ( .C1(n20689), .C2(n20507), .A(n20450), .B(n20449), .ZN(
        P1_U3105) );
  AOI22_X1 U23436 ( .A1(n20691), .A2(n20465), .B1(n20690), .B2(n20464), .ZN(
        n20452) );
  AOI22_X1 U23437 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20467), .B1(
        n20466), .B2(n20692), .ZN(n20451) );
  OAI211_X1 U23438 ( .C1(n20695), .C2(n20507), .A(n20452), .B(n20451), .ZN(
        P1_U3106) );
  AOI22_X1 U23439 ( .A1(n20697), .A2(n20465), .B1(n20696), .B2(n20464), .ZN(
        n20454) );
  AOI22_X1 U23440 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20467), .B1(
        n20503), .B2(n20698), .ZN(n20453) );
  OAI211_X1 U23441 ( .C1(n20701), .C2(n20459), .A(n20454), .B(n20453), .ZN(
        P1_U3107) );
  AOI22_X1 U23442 ( .A1(n20703), .A2(n20465), .B1(n20702), .B2(n20464), .ZN(
        n20456) );
  AOI22_X1 U23443 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20467), .B1(
        n20466), .B2(n20704), .ZN(n20455) );
  OAI211_X1 U23444 ( .C1(n20707), .C2(n20507), .A(n20456), .B(n20455), .ZN(
        P1_U3108) );
  AOI22_X1 U23445 ( .A1(n20709), .A2(n20465), .B1(n20708), .B2(n20464), .ZN(
        n20458) );
  AOI22_X1 U23446 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20467), .B1(
        n20503), .B2(n20710), .ZN(n20457) );
  OAI211_X1 U23447 ( .C1(n20713), .C2(n20459), .A(n20458), .B(n20457), .ZN(
        P1_U3109) );
  AOI22_X1 U23448 ( .A1(n20715), .A2(n20465), .B1(n20714), .B2(n20464), .ZN(
        n20461) );
  AOI22_X1 U23449 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20467), .B1(
        n20466), .B2(n20662), .ZN(n20460) );
  OAI211_X1 U23450 ( .C1(n20665), .C2(n20507), .A(n20461), .B(n20460), .ZN(
        P1_U3110) );
  AOI22_X1 U23451 ( .A1(n20723), .A2(n20465), .B1(n20722), .B2(n20464), .ZN(
        n20463) );
  AOI22_X1 U23452 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20467), .B1(
        n20466), .B2(n20724), .ZN(n20462) );
  OAI211_X1 U23453 ( .C1(n20727), .C2(n20507), .A(n20463), .B(n20462), .ZN(
        P1_U3111) );
  AOI22_X1 U23454 ( .A1(n20731), .A2(n20465), .B1(n20729), .B2(n20464), .ZN(
        n20469) );
  AOI22_X1 U23455 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20467), .B1(
        n20466), .B2(n20732), .ZN(n20468) );
  OAI211_X1 U23456 ( .C1(n20738), .C2(n20507), .A(n20469), .B(n20468), .ZN(
        P1_U3112) );
  AOI21_X1 U23457 ( .B1(n20546), .B2(n20507), .A(n20643), .ZN(n20470) );
  NOR2_X1 U23458 ( .A1(n20470), .A2(n20836), .ZN(n20481) );
  AND2_X1 U23459 ( .A1(n20518), .A2(n20645), .ZN(n20476) );
  INV_X1 U23460 ( .A(n20471), .ZN(n20474) );
  OR2_X1 U23461 ( .A1(n20472), .A2(n20515), .ZN(n20640) );
  INV_X1 U23462 ( .A(n20640), .ZN(n20473) );
  NAND3_X1 U23463 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n11766), .ZN(n20519) );
  NOR2_X1 U23464 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20519), .ZN(
        n20478) );
  INV_X1 U23465 ( .A(n20478), .ZN(n20506) );
  OAI22_X1 U23466 ( .A1(n20546), .A2(n20689), .B1(n20556), .B2(n20506), .ZN(
        n20475) );
  INV_X1 U23467 ( .A(n20475), .ZN(n20484) );
  INV_X1 U23468 ( .A(n20476), .ZN(n20480) );
  NAND2_X1 U23469 ( .A1(n20640), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20648) );
  OAI211_X1 U23470 ( .C1(n21100), .C2(n20478), .A(n20648), .B(n20477), .ZN(
        n20479) );
  AOI21_X1 U23471 ( .B1(n20481), .B2(n20480), .A(n20479), .ZN(n20482) );
  AOI22_X1 U23472 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20509), .B1(
        n20503), .B2(n20686), .ZN(n20483) );
  OAI211_X1 U23473 ( .C1(n20512), .C2(n20566), .A(n20484), .B(n20483), .ZN(
        P1_U3113) );
  OAI22_X1 U23474 ( .A1(n20507), .A2(n20485), .B1(n20567), .B2(n20506), .ZN(
        n20486) );
  INV_X1 U23475 ( .A(n20486), .ZN(n20489) );
  AOI22_X1 U23476 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20509), .B1(
        n20537), .B2(n20487), .ZN(n20488) );
  OAI211_X1 U23477 ( .C1(n20512), .C2(n20571), .A(n20489), .B(n20488), .ZN(
        P1_U3114) );
  OAI22_X1 U23478 ( .A1(n20546), .A2(n20573), .B1(n20572), .B2(n20506), .ZN(
        n20490) );
  INV_X1 U23479 ( .A(n20490), .ZN(n20492) );
  AOI22_X1 U23480 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20509), .B1(
        n20503), .B2(n20575), .ZN(n20491) );
  OAI211_X1 U23481 ( .C1(n20512), .C2(n20578), .A(n20492), .B(n20491), .ZN(
        P1_U3115) );
  OAI22_X1 U23482 ( .A1(n20546), .A2(n20707), .B1(n20579), .B2(n20506), .ZN(
        n20493) );
  INV_X1 U23483 ( .A(n20493), .ZN(n20495) );
  AOI22_X1 U23484 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20509), .B1(
        n20503), .B2(n20704), .ZN(n20494) );
  OAI211_X1 U23485 ( .C1(n20512), .C2(n20583), .A(n20495), .B(n20494), .ZN(
        P1_U3116) );
  OAI22_X1 U23486 ( .A1(n20546), .A2(n20585), .B1(n20584), .B2(n20506), .ZN(
        n20496) );
  INV_X1 U23487 ( .A(n20496), .ZN(n20498) );
  AOI22_X1 U23488 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20509), .B1(
        n20503), .B2(n20587), .ZN(n20497) );
  OAI211_X1 U23489 ( .C1(n20512), .C2(n20590), .A(n20498), .B(n20497), .ZN(
        P1_U3117) );
  OAI22_X1 U23490 ( .A1(n20546), .A2(n20665), .B1(n20591), .B2(n20506), .ZN(
        n20499) );
  INV_X1 U23491 ( .A(n20499), .ZN(n20501) );
  AOI22_X1 U23492 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20509), .B1(
        n20503), .B2(n20662), .ZN(n20500) );
  OAI211_X1 U23493 ( .C1(n20512), .C2(n20595), .A(n20501), .B(n20500), .ZN(
        P1_U3118) );
  OAI22_X1 U23494 ( .A1(n20546), .A2(n20727), .B1(n20596), .B2(n20506), .ZN(
        n20502) );
  INV_X1 U23495 ( .A(n20502), .ZN(n20505) );
  AOI22_X1 U23496 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20509), .B1(
        n20503), .B2(n20724), .ZN(n20504) );
  OAI211_X1 U23497 ( .C1(n20512), .C2(n20600), .A(n20505), .B(n20504), .ZN(
        P1_U3119) );
  OAI22_X1 U23498 ( .A1(n20507), .A2(n20547), .B1(n20602), .B2(n20506), .ZN(
        n20508) );
  INV_X1 U23499 ( .A(n20508), .ZN(n20511) );
  AOI22_X1 U23500 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20509), .B1(
        n20537), .B2(n20542), .ZN(n20510) );
  OAI211_X1 U23501 ( .C1(n20512), .C2(n20608), .A(n20511), .B(n20510), .ZN(
        P1_U3120) );
  NOR2_X1 U23502 ( .A1(n20516), .A2(n20515), .ZN(n20541) );
  AOI21_X1 U23503 ( .B1(n20518), .B2(n20517), .A(n20541), .ZN(n20520) );
  OAI22_X1 U23504 ( .A1(n20520), .A2(n20836), .B1(n20519), .B2(n20742), .ZN(
        n20540) );
  AOI22_X1 U23505 ( .A1(n20678), .A2(n20541), .B1(n20677), .B2(n20540), .ZN(
        n20526) );
  INV_X1 U23506 ( .A(n20519), .ZN(n20524) );
  OAI21_X1 U23507 ( .B1(n20522), .B2(n20521), .A(n20520), .ZN(n20523) );
  OAI221_X1 U23508 ( .B1(n20613), .B2(n20524), .C1(n20836), .C2(n20523), .A(
        n20684), .ZN(n20543) );
  AOI22_X1 U23509 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20543), .B1(
        n20537), .B2(n20686), .ZN(n20525) );
  OAI211_X1 U23510 ( .C1(n20689), .C2(n20549), .A(n20526), .B(n20525), .ZN(
        P1_U3121) );
  AOI22_X1 U23511 ( .A1(n20691), .A2(n20541), .B1(n20690), .B2(n20540), .ZN(
        n20528) );
  AOI22_X1 U23512 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20543), .B1(
        n20537), .B2(n20692), .ZN(n20527) );
  OAI211_X1 U23513 ( .C1(n20695), .C2(n20549), .A(n20528), .B(n20527), .ZN(
        P1_U3122) );
  AOI22_X1 U23514 ( .A1(n20697), .A2(n20541), .B1(n20696), .B2(n20540), .ZN(
        n20530) );
  AOI22_X1 U23515 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20543), .B1(
        n20604), .B2(n20698), .ZN(n20529) );
  OAI211_X1 U23516 ( .C1(n20701), .C2(n20546), .A(n20530), .B(n20529), .ZN(
        P1_U3123) );
  AOI22_X1 U23517 ( .A1(n20703), .A2(n20541), .B1(n20702), .B2(n20540), .ZN(
        n20532) );
  AOI22_X1 U23518 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20543), .B1(
        n20537), .B2(n20704), .ZN(n20531) );
  OAI211_X1 U23519 ( .C1(n20707), .C2(n20549), .A(n20532), .B(n20531), .ZN(
        P1_U3124) );
  AOI22_X1 U23520 ( .A1(n20709), .A2(n20541), .B1(n20708), .B2(n20540), .ZN(
        n20534) );
  AOI22_X1 U23521 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20543), .B1(
        n20604), .B2(n20710), .ZN(n20533) );
  OAI211_X1 U23522 ( .C1(n20713), .C2(n20546), .A(n20534), .B(n20533), .ZN(
        P1_U3125) );
  AOI22_X1 U23523 ( .A1(n20715), .A2(n20541), .B1(n20714), .B2(n20540), .ZN(
        n20536) );
  AOI22_X1 U23524 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20543), .B1(
        n20537), .B2(n20662), .ZN(n20535) );
  OAI211_X1 U23525 ( .C1(n20665), .C2(n20549), .A(n20536), .B(n20535), .ZN(
        P1_U3126) );
  AOI22_X1 U23526 ( .A1(n20723), .A2(n20541), .B1(n20722), .B2(n20540), .ZN(
        n20539) );
  AOI22_X1 U23527 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20543), .B1(
        n20537), .B2(n20724), .ZN(n20538) );
  OAI211_X1 U23528 ( .C1(n20727), .C2(n20549), .A(n20539), .B(n20538), .ZN(
        P1_U3127) );
  AOI22_X1 U23529 ( .A1(n20731), .A2(n20541), .B1(n20729), .B2(n20540), .ZN(
        n20545) );
  AOI22_X1 U23530 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20543), .B1(
        n20604), .B2(n20542), .ZN(n20544) );
  OAI211_X1 U23531 ( .C1(n20547), .C2(n20546), .A(n20545), .B(n20544), .ZN(
        P1_U3128) );
  AOI21_X1 U23532 ( .B1(n20549), .B2(n20630), .A(n20643), .ZN(n20550) );
  NOR2_X1 U23533 ( .A1(n20550), .A2(n20836), .ZN(n20561) );
  OR2_X1 U23534 ( .A1(n20552), .A2(n20551), .ZN(n20612) );
  NOR2_X1 U23535 ( .A1(n20612), .A2(n20645), .ZN(n20558) );
  NAND3_X1 U23536 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20555), .ZN(n20615) );
  NOR2_X1 U23537 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20615), .ZN(
        n20563) );
  INV_X1 U23538 ( .A(n20563), .ZN(n20601) );
  OAI22_X1 U23539 ( .A1(n20630), .A2(n20689), .B1(n20556), .B2(n20601), .ZN(
        n20557) );
  INV_X1 U23540 ( .A(n20557), .ZN(n20565) );
  INV_X1 U23541 ( .A(n20558), .ZN(n20560) );
  AOI22_X1 U23542 ( .A1(n20561), .A2(n20560), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20559), .ZN(n20562) );
  AOI22_X1 U23543 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20605), .B1(
        n20604), .B2(n20686), .ZN(n20564) );
  OAI211_X1 U23544 ( .C1(n20609), .C2(n20566), .A(n20565), .B(n20564), .ZN(
        P1_U3129) );
  OAI22_X1 U23545 ( .A1(n20630), .A2(n20695), .B1(n20567), .B2(n20601), .ZN(
        n20568) );
  INV_X1 U23546 ( .A(n20568), .ZN(n20570) );
  AOI22_X1 U23547 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20605), .B1(
        n20604), .B2(n20692), .ZN(n20569) );
  OAI211_X1 U23548 ( .C1(n20609), .C2(n20571), .A(n20570), .B(n20569), .ZN(
        P1_U3130) );
  OAI22_X1 U23549 ( .A1(n20630), .A2(n20573), .B1(n20572), .B2(n20601), .ZN(
        n20574) );
  INV_X1 U23550 ( .A(n20574), .ZN(n20577) );
  AOI22_X1 U23551 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20605), .B1(
        n20604), .B2(n20575), .ZN(n20576) );
  OAI211_X1 U23552 ( .C1(n20609), .C2(n20578), .A(n20577), .B(n20576), .ZN(
        P1_U3131) );
  OAI22_X1 U23553 ( .A1(n20630), .A2(n20707), .B1(n20579), .B2(n20601), .ZN(
        n20580) );
  INV_X1 U23554 ( .A(n20580), .ZN(n20582) );
  AOI22_X1 U23555 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20605), .B1(
        n20604), .B2(n20704), .ZN(n20581) );
  OAI211_X1 U23556 ( .C1(n20609), .C2(n20583), .A(n20582), .B(n20581), .ZN(
        P1_U3132) );
  OAI22_X1 U23557 ( .A1(n20630), .A2(n20585), .B1(n20584), .B2(n20601), .ZN(
        n20586) );
  INV_X1 U23558 ( .A(n20586), .ZN(n20589) );
  AOI22_X1 U23559 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20605), .B1(
        n20604), .B2(n20587), .ZN(n20588) );
  OAI211_X1 U23560 ( .C1(n20609), .C2(n20590), .A(n20589), .B(n20588), .ZN(
        P1_U3133) );
  OAI22_X1 U23561 ( .A1(n20630), .A2(n20665), .B1(n20591), .B2(n20601), .ZN(
        n20592) );
  INV_X1 U23562 ( .A(n20592), .ZN(n20594) );
  AOI22_X1 U23563 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20605), .B1(
        n20604), .B2(n20662), .ZN(n20593) );
  OAI211_X1 U23564 ( .C1(n20609), .C2(n20595), .A(n20594), .B(n20593), .ZN(
        P1_U3134) );
  OAI22_X1 U23565 ( .A1(n20630), .A2(n20727), .B1(n20596), .B2(n20601), .ZN(
        n20597) );
  INV_X1 U23566 ( .A(n20597), .ZN(n20599) );
  AOI22_X1 U23567 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20605), .B1(
        n20604), .B2(n20724), .ZN(n20598) );
  OAI211_X1 U23568 ( .C1(n20609), .C2(n20600), .A(n20599), .B(n20598), .ZN(
        P1_U3135) );
  OAI22_X1 U23569 ( .A1(n20630), .A2(n20738), .B1(n20602), .B2(n20601), .ZN(
        n20603) );
  INV_X1 U23570 ( .A(n20603), .ZN(n20607) );
  AOI22_X1 U23571 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20605), .B1(
        n20604), .B2(n20732), .ZN(n20606) );
  OAI211_X1 U23572 ( .C1(n20609), .C2(n20608), .A(n20607), .B(n20606), .ZN(
        P1_U3136) );
  NOR2_X1 U23573 ( .A1(n20611), .A2(n20615), .ZN(n20634) );
  INV_X1 U23574 ( .A(n20634), .ZN(n20614) );
  INV_X1 U23575 ( .A(n20612), .ZN(n20646) );
  NAND2_X1 U23576 ( .A1(n20646), .A2(n20613), .ZN(n20676) );
  OAI222_X1 U23577 ( .A1(n20614), .A2(n20836), .B1(n20742), .B2(n20615), .C1(
        n20188), .C2(n20676), .ZN(n20633) );
  AOI22_X1 U23578 ( .A1(n20678), .A2(n20634), .B1(n20677), .B2(n20633), .ZN(
        n20619) );
  INV_X1 U23579 ( .A(n20615), .ZN(n20617) );
  INV_X1 U23580 ( .A(n20630), .ZN(n20635) );
  AOI22_X1 U23581 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20636), .B1(
        n20635), .B2(n20686), .ZN(n20618) );
  OAI211_X1 U23582 ( .C1(n20689), .C2(n20661), .A(n20619), .B(n20618), .ZN(
        P1_U3137) );
  AOI22_X1 U23583 ( .A1(n20691), .A2(n20634), .B1(n20690), .B2(n20633), .ZN(
        n20621) );
  AOI22_X1 U23584 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20636), .B1(
        n20635), .B2(n20692), .ZN(n20620) );
  OAI211_X1 U23585 ( .C1(n20695), .C2(n20661), .A(n20621), .B(n20620), .ZN(
        P1_U3138) );
  AOI22_X1 U23586 ( .A1(n20697), .A2(n20634), .B1(n20696), .B2(n20633), .ZN(
        n20623) );
  AOI22_X1 U23587 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20636), .B1(
        n20670), .B2(n20698), .ZN(n20622) );
  OAI211_X1 U23588 ( .C1(n20701), .C2(n20630), .A(n20623), .B(n20622), .ZN(
        P1_U3139) );
  AOI22_X1 U23589 ( .A1(n20703), .A2(n20634), .B1(n20702), .B2(n20633), .ZN(
        n20625) );
  AOI22_X1 U23590 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20636), .B1(
        n20635), .B2(n20704), .ZN(n20624) );
  OAI211_X1 U23591 ( .C1(n20707), .C2(n20661), .A(n20625), .B(n20624), .ZN(
        P1_U3140) );
  AOI22_X1 U23592 ( .A1(n20709), .A2(n20634), .B1(n20708), .B2(n20633), .ZN(
        n20627) );
  AOI22_X1 U23593 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20636), .B1(
        n20670), .B2(n20710), .ZN(n20626) );
  OAI211_X1 U23594 ( .C1(n20713), .C2(n20630), .A(n20627), .B(n20626), .ZN(
        P1_U3141) );
  AOI22_X1 U23595 ( .A1(n20715), .A2(n20634), .B1(n20714), .B2(n20633), .ZN(
        n20629) );
  AOI22_X1 U23596 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20636), .B1(
        n20670), .B2(n20716), .ZN(n20628) );
  OAI211_X1 U23597 ( .C1(n20721), .C2(n20630), .A(n20629), .B(n20628), .ZN(
        P1_U3142) );
  AOI22_X1 U23598 ( .A1(n20723), .A2(n20634), .B1(n20722), .B2(n20633), .ZN(
        n20632) );
  AOI22_X1 U23599 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20636), .B1(
        n20635), .B2(n20724), .ZN(n20631) );
  OAI211_X1 U23600 ( .C1(n20727), .C2(n20661), .A(n20632), .B(n20631), .ZN(
        P1_U3143) );
  AOI22_X1 U23601 ( .A1(n20731), .A2(n20634), .B1(n20729), .B2(n20633), .ZN(
        n20638) );
  AOI22_X1 U23602 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20636), .B1(
        n20635), .B2(n20732), .ZN(n20637) );
  OAI211_X1 U23603 ( .C1(n20738), .C2(n20661), .A(n20638), .B(n20637), .ZN(
        P1_U3144) );
  NOR2_X1 U23604 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20681), .ZN(
        n20669) );
  OAI22_X1 U23605 ( .A1(n20676), .A2(n20642), .B1(n20641), .B2(n20640), .ZN(
        n20668) );
  AOI22_X1 U23606 ( .A1(n20678), .A2(n20669), .B1(n20677), .B2(n20668), .ZN(
        n20652) );
  AOI21_X1 U23607 ( .B1(n20720), .B2(n20661), .A(n20643), .ZN(n20644) );
  AOI21_X1 U23608 ( .B1(n20646), .B2(n20645), .A(n20644), .ZN(n20647) );
  NOR2_X1 U23609 ( .A1(n20647), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20650) );
  AOI22_X1 U23610 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20671), .B1(
        n20670), .B2(n20686), .ZN(n20651) );
  OAI211_X1 U23611 ( .C1(n20689), .C2(n20720), .A(n20652), .B(n20651), .ZN(
        P1_U3145) );
  AOI22_X1 U23612 ( .A1(n20691), .A2(n20669), .B1(n20690), .B2(n20668), .ZN(
        n20654) );
  AOI22_X1 U23613 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20671), .B1(
        n20670), .B2(n20692), .ZN(n20653) );
  OAI211_X1 U23614 ( .C1(n20695), .C2(n20720), .A(n20654), .B(n20653), .ZN(
        P1_U3146) );
  AOI22_X1 U23615 ( .A1(n20697), .A2(n20669), .B1(n20696), .B2(n20668), .ZN(
        n20656) );
  AOI22_X1 U23616 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20671), .B1(
        n20733), .B2(n20698), .ZN(n20655) );
  OAI211_X1 U23617 ( .C1(n20701), .C2(n20661), .A(n20656), .B(n20655), .ZN(
        P1_U3147) );
  AOI22_X1 U23618 ( .A1(n20703), .A2(n20669), .B1(n20702), .B2(n20668), .ZN(
        n20658) );
  AOI22_X1 U23619 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20671), .B1(
        n20670), .B2(n20704), .ZN(n20657) );
  OAI211_X1 U23620 ( .C1(n20707), .C2(n20720), .A(n20658), .B(n20657), .ZN(
        P1_U3148) );
  AOI22_X1 U23621 ( .A1(n20709), .A2(n20669), .B1(n20708), .B2(n20668), .ZN(
        n20660) );
  AOI22_X1 U23622 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20671), .B1(
        n20733), .B2(n20710), .ZN(n20659) );
  OAI211_X1 U23623 ( .C1(n20713), .C2(n20661), .A(n20660), .B(n20659), .ZN(
        P1_U3149) );
  AOI22_X1 U23624 ( .A1(n20715), .A2(n20669), .B1(n20714), .B2(n20668), .ZN(
        n20664) );
  AOI22_X1 U23625 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20671), .B1(
        n20670), .B2(n20662), .ZN(n20663) );
  OAI211_X1 U23626 ( .C1(n20665), .C2(n20720), .A(n20664), .B(n20663), .ZN(
        P1_U3150) );
  AOI22_X1 U23627 ( .A1(n20723), .A2(n20669), .B1(n20722), .B2(n20668), .ZN(
        n20667) );
  AOI22_X1 U23628 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20671), .B1(
        n20670), .B2(n20724), .ZN(n20666) );
  OAI211_X1 U23629 ( .C1(n20727), .C2(n20720), .A(n20667), .B(n20666), .ZN(
        P1_U3151) );
  AOI22_X1 U23630 ( .A1(n20731), .A2(n20669), .B1(n20729), .B2(n20668), .ZN(
        n20673) );
  AOI22_X1 U23631 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20671), .B1(
        n20670), .B2(n20732), .ZN(n20672) );
  OAI211_X1 U23632 ( .C1(n20738), .C2(n20720), .A(n20673), .B(n20672), .ZN(
        P1_U3152) );
  INV_X1 U23633 ( .A(n20674), .ZN(n20730) );
  OAI222_X1 U23634 ( .A1(n20676), .A2(n20675), .B1(n20742), .B2(n20681), .C1(
        n20836), .C2(n20674), .ZN(n20728) );
  AOI22_X1 U23635 ( .A1(n20678), .A2(n20730), .B1(n20677), .B2(n20728), .ZN(
        n20688) );
  INV_X1 U23636 ( .A(n20679), .ZN(n20683) );
  INV_X1 U23637 ( .A(n20680), .ZN(n20682) );
  OAI21_X1 U23638 ( .B1(n20683), .B2(n20682), .A(n20681), .ZN(n20685) );
  NAND2_X1 U23639 ( .A1(n20685), .A2(n20684), .ZN(n20734) );
  AOI22_X1 U23640 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20734), .B1(
        n20733), .B2(n20686), .ZN(n20687) );
  OAI211_X1 U23641 ( .C1(n20689), .C2(n20737), .A(n20688), .B(n20687), .ZN(
        P1_U3153) );
  AOI22_X1 U23642 ( .A1(n20691), .A2(n20730), .B1(n20690), .B2(n20728), .ZN(
        n20694) );
  AOI22_X1 U23643 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20734), .B1(
        n20733), .B2(n20692), .ZN(n20693) );
  OAI211_X1 U23644 ( .C1(n20695), .C2(n20737), .A(n20694), .B(n20693), .ZN(
        P1_U3154) );
  AOI22_X1 U23645 ( .A1(n20697), .A2(n20730), .B1(n20696), .B2(n20728), .ZN(
        n20700) );
  AOI22_X1 U23646 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20734), .B1(
        n20717), .B2(n20698), .ZN(n20699) );
  OAI211_X1 U23647 ( .C1(n20701), .C2(n20720), .A(n20700), .B(n20699), .ZN(
        P1_U3155) );
  AOI22_X1 U23648 ( .A1(n20703), .A2(n20730), .B1(n20702), .B2(n20728), .ZN(
        n20706) );
  AOI22_X1 U23649 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20734), .B1(
        n20733), .B2(n20704), .ZN(n20705) );
  OAI211_X1 U23650 ( .C1(n20707), .C2(n20737), .A(n20706), .B(n20705), .ZN(
        P1_U3156) );
  AOI22_X1 U23651 ( .A1(n20709), .A2(n20730), .B1(n20708), .B2(n20728), .ZN(
        n20712) );
  AOI22_X1 U23652 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20734), .B1(
        n20717), .B2(n20710), .ZN(n20711) );
  OAI211_X1 U23653 ( .C1(n20713), .C2(n20720), .A(n20712), .B(n20711), .ZN(
        P1_U3157) );
  AOI22_X1 U23654 ( .A1(n20715), .A2(n20730), .B1(n20714), .B2(n20728), .ZN(
        n20719) );
  AOI22_X1 U23655 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20734), .B1(
        n20717), .B2(n20716), .ZN(n20718) );
  OAI211_X1 U23656 ( .C1(n20721), .C2(n20720), .A(n20719), .B(n20718), .ZN(
        P1_U3158) );
  AOI22_X1 U23657 ( .A1(n20723), .A2(n20730), .B1(n20722), .B2(n20728), .ZN(
        n20726) );
  AOI22_X1 U23658 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20734), .B1(
        n20733), .B2(n20724), .ZN(n20725) );
  OAI211_X1 U23659 ( .C1(n20727), .C2(n20737), .A(n20726), .B(n20725), .ZN(
        P1_U3159) );
  AOI22_X1 U23660 ( .A1(n20731), .A2(n20730), .B1(n20729), .B2(n20728), .ZN(
        n20736) );
  AOI22_X1 U23661 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20734), .B1(
        n20733), .B2(n20732), .ZN(n20735) );
  OAI211_X1 U23662 ( .C1(n20738), .C2(n20737), .A(n20736), .B(n20735), .ZN(
        P1_U3160) );
  NOR2_X1 U23663 ( .A1(n11495), .A2(n20739), .ZN(n20743) );
  INV_X1 U23664 ( .A(n20740), .ZN(n20741) );
  OAI21_X1 U23665 ( .B1(n20743), .B2(n20742), .A(n20741), .ZN(P1_U3163) );
  AND2_X1 U23666 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20814), .ZN(
        P1_U3164) );
  AND2_X1 U23667 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20814), .ZN(
        P1_U3165) );
  AND2_X1 U23668 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20814), .ZN(
        P1_U3166) );
  AND2_X1 U23669 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20814), .ZN(
        P1_U3167) );
  AND2_X1 U23670 ( .A1(n20814), .A2(P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(
        P1_U3168) );
  AND2_X1 U23671 ( .A1(n20814), .A2(P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(
        P1_U3169) );
  AND2_X1 U23672 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20814), .ZN(
        P1_U3170) );
  AND2_X1 U23673 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20814), .ZN(
        P1_U3171) );
  AND2_X1 U23674 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20814), .ZN(
        P1_U3172) );
  AND2_X1 U23675 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20814), .ZN(
        P1_U3173) );
  AND2_X1 U23676 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20814), .ZN(
        P1_U3174) );
  AND2_X1 U23677 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20814), .ZN(
        P1_U3175) );
  AND2_X1 U23678 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20814), .ZN(
        P1_U3176) );
  AND2_X1 U23679 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20814), .ZN(
        P1_U3177) );
  AND2_X1 U23680 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20814), .ZN(
        P1_U3178) );
  AND2_X1 U23681 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20814), .ZN(
        P1_U3179) );
  AND2_X1 U23682 ( .A1(n20814), .A2(P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(
        P1_U3180) );
  AND2_X1 U23683 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20814), .ZN(
        P1_U3181) );
  AND2_X1 U23684 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20814), .ZN(
        P1_U3182) );
  AND2_X1 U23685 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20814), .ZN(
        P1_U3183) );
  AND2_X1 U23686 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20814), .ZN(
        P1_U3184) );
  AND2_X1 U23687 ( .A1(n20814), .A2(P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(
        P1_U3185) );
  AND2_X1 U23688 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20814), .ZN(P1_U3186) );
  AND2_X1 U23689 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20814), .ZN(P1_U3187) );
  AND2_X1 U23690 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20814), .ZN(P1_U3188) );
  AND2_X1 U23691 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20814), .ZN(P1_U3189) );
  AND2_X1 U23692 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20814), .ZN(P1_U3190) );
  AND2_X1 U23693 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20814), .ZN(P1_U3191) );
  AND2_X1 U23694 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20814), .ZN(P1_U3192) );
  AND2_X1 U23695 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20814), .ZN(P1_U3193) );
  AOI21_X1 U23696 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20838), .A(n20746), 
        .ZN(n20755) );
  NOR2_X1 U23697 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20744) );
  NOR2_X1 U23698 ( .A1(n20744), .A2(n21002), .ZN(n20745) );
  AOI211_X1 U23699 ( .C1(NA), .C2(n20746), .A(n20745), .B(n20749), .ZN(n20747)
         );
  OAI22_X1 U23700 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20755), .B1(n20800), 
        .B2(n20747), .ZN(P1_U3194) );
  AOI21_X1 U23701 ( .B1(n20838), .B2(n20753), .A(n20748), .ZN(n20757) );
  OAI211_X1 U23702 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20749), .A(
        P1_STATE_REG_0__SCAN_IN), .B(HOLD), .ZN(n20756) );
  INV_X1 U23703 ( .A(n20750), .ZN(n20751) );
  AOI221_X1 U23704 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n20753), .C1(n20752), 
        .C2(n20753), .A(n20751), .ZN(n20754) );
  OAI22_X1 U23705 ( .A1(n20757), .A2(n20756), .B1(n20755), .B2(n20754), .ZN(
        P1_U3196) );
  NOR2_X1 U23706 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20833), .ZN(n20805) );
  AOI22_X1 U23707 ( .A1(P1_ADDRESS_REG_0__SCAN_IN), .A2(n20833), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n20805), .ZN(n20758) );
  OAI21_X1 U23708 ( .B1(n13735), .B2(n20803), .A(n20758), .ZN(P1_U3197) );
  AOI22_X1 U23709 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(n20833), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n20806), .ZN(n20759) );
  OAI21_X1 U23710 ( .B1(n13563), .B2(n20798), .A(n20759), .ZN(P1_U3198) );
  OAI222_X1 U23711 ( .A1(n20803), .A2(n13563), .B1(n20760), .B2(n20800), .C1(
        n20761), .C2(n20798), .ZN(P1_U3199) );
  INV_X1 U23712 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20876) );
  OAI222_X1 U23713 ( .A1(n20798), .A2(n20763), .B1(n20876), .B2(n20800), .C1(
        n20761), .C2(n20803), .ZN(P1_U3200) );
  AOI22_X1 U23714 ( .A1(P1_ADDRESS_REG_4__SCAN_IN), .A2(n20833), .B1(
        P1_REIP_REG_6__SCAN_IN), .B2(n20805), .ZN(n20762) );
  OAI21_X1 U23715 ( .B1(n20763), .B2(n20803), .A(n20762), .ZN(P1_U3201) );
  INV_X1 U23716 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20765) );
  AOI22_X1 U23717 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(n20833), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20805), .ZN(n20764) );
  OAI21_X1 U23718 ( .B1(n20765), .B2(n20803), .A(n20764), .ZN(P1_U3202) );
  AOI22_X1 U23719 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n20833), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20806), .ZN(n20766) );
  OAI21_X1 U23720 ( .B1(n21092), .B2(n20798), .A(n20766), .ZN(P1_U3203) );
  INV_X1 U23721 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20767) );
  OAI222_X1 U23722 ( .A1(n20798), .A2(n13899), .B1(n20767), .B2(n20800), .C1(
        n21092), .C2(n20803), .ZN(P1_U3204) );
  INV_X1 U23723 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n20911) );
  OAI222_X1 U23724 ( .A1(n20803), .A2(n13899), .B1(n20911), .B2(n20800), .C1(
        n20768), .C2(n20798), .ZN(P1_U3205) );
  INV_X1 U23725 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n20769) );
  OAI222_X1 U23726 ( .A1(n20798), .A2(n20771), .B1(n20769), .B2(n20800), .C1(
        n20768), .C2(n20803), .ZN(P1_U3206) );
  INV_X1 U23727 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n20770) );
  OAI222_X1 U23728 ( .A1(n20803), .A2(n20771), .B1(n20770), .B2(n20800), .C1(
        n20772), .C2(n20798), .ZN(P1_U3207) );
  INV_X1 U23729 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n20773) );
  OAI222_X1 U23730 ( .A1(n20798), .A2(n14017), .B1(n20773), .B2(n20800), .C1(
        n20772), .C2(n20803), .ZN(P1_U3208) );
  AOI22_X1 U23731 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n20833), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20805), .ZN(n20774) );
  OAI21_X1 U23732 ( .B1(n14017), .B2(n20803), .A(n20774), .ZN(P1_U3209) );
  INV_X1 U23733 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20777) );
  INV_X1 U23734 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n20974) );
  INV_X1 U23735 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n20775) );
  OAI222_X1 U23736 ( .A1(n20798), .A2(n20777), .B1(n20974), .B2(n20800), .C1(
        n20775), .C2(n20803), .ZN(P1_U3210) );
  AOI22_X1 U23737 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(n20833), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n20805), .ZN(n20776) );
  OAI21_X1 U23738 ( .B1(n20777), .B2(n20803), .A(n20776), .ZN(P1_U3211) );
  AOI22_X1 U23739 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20833), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n20806), .ZN(n20778) );
  OAI21_X1 U23740 ( .B1(n20780), .B2(n20798), .A(n20778), .ZN(P1_U3212) );
  INV_X1 U23741 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n20779) );
  INV_X1 U23742 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20943) );
  OAI222_X1 U23743 ( .A1(n20803), .A2(n20780), .B1(n20779), .B2(n20800), .C1(
        n20943), .C2(n20798), .ZN(P1_U3213) );
  INV_X1 U23744 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n20781) );
  OAI222_X1 U23745 ( .A1(n20798), .A2(n20783), .B1(n20781), .B2(n20800), .C1(
        n20943), .C2(n20803), .ZN(P1_U3214) );
  INV_X1 U23746 ( .A(P1_ADDRESS_REG_18__SCAN_IN), .ZN(n20782) );
  OAI222_X1 U23747 ( .A1(n20803), .A2(n20783), .B1(n20782), .B2(n20800), .C1(
        n20785), .C2(n20798), .ZN(P1_U3215) );
  INV_X1 U23748 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n20784) );
  OAI222_X1 U23749 ( .A1(n20803), .A2(n20785), .B1(n20784), .B2(n20800), .C1(
        n14514), .C2(n20798), .ZN(P1_U3216) );
  INV_X1 U23750 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20786) );
  OAI222_X1 U23751 ( .A1(n20803), .A2(n14514), .B1(n20786), .B2(n20800), .C1(
        n20788), .C2(n20798), .ZN(P1_U3217) );
  AOI22_X1 U23752 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n20833), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20805), .ZN(n20787) );
  OAI21_X1 U23753 ( .B1(n20788), .B2(n20803), .A(n20787), .ZN(P1_U3218) );
  AOI22_X1 U23754 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n20833), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20806), .ZN(n20789) );
  OAI21_X1 U23755 ( .B1(n20791), .B2(n20798), .A(n20789), .ZN(P1_U3219) );
  INV_X1 U23756 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n20790) );
  OAI222_X1 U23757 ( .A1(n20803), .A2(n20791), .B1(n20790), .B2(n20800), .C1(
        n20793), .C2(n20798), .ZN(P1_U3220) );
  INV_X1 U23758 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20792) );
  OAI222_X1 U23759 ( .A1(n20803), .A2(n20793), .B1(n20792), .B2(n20800), .C1(
        n20795), .C2(n20798), .ZN(P1_U3221) );
  INV_X1 U23760 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n20794) );
  OAI222_X1 U23761 ( .A1(n20803), .A2(n20795), .B1(n20794), .B2(n20800), .C1(
        n20797), .C2(n20798), .ZN(P1_U3222) );
  INV_X1 U23762 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n20796) );
  OAI222_X1 U23763 ( .A1(n20803), .A2(n20797), .B1(n20796), .B2(n20800), .C1(
        n20802), .C2(n20798), .ZN(P1_U3223) );
  INV_X1 U23764 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n20801) );
  OAI222_X1 U23765 ( .A1(n20803), .A2(n20802), .B1(n20801), .B2(n20800), .C1(
        n20799), .C2(n20798), .ZN(P1_U3224) );
  AOI222_X1 U23766 ( .A1(n20805), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20833), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20806), .ZN(n20804) );
  INV_X1 U23767 ( .A(n20804), .ZN(P1_U3225) );
  AOI222_X1 U23768 ( .A1(n20806), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20833), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20805), .ZN(n20807) );
  INV_X1 U23769 ( .A(n20807), .ZN(P1_U3226) );
  INV_X1 U23770 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20808) );
  AOI22_X1 U23771 ( .A1(n20800), .A2(n21081), .B1(n20808), .B2(n20833), .ZN(
        P1_U3458) );
  INV_X1 U23772 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20828) );
  INV_X1 U23773 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n20809) );
  AOI22_X1 U23774 ( .A1(n20800), .A2(n20828), .B1(n20809), .B2(n20833), .ZN(
        P1_U3459) );
  INV_X1 U23775 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20810) );
  AOI22_X1 U23776 ( .A1(n20800), .A2(n20811), .B1(n20810), .B2(n20833), .ZN(
        P1_U3460) );
  INV_X1 U23777 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20831) );
  INV_X1 U23778 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20812) );
  AOI22_X1 U23779 ( .A1(n20800), .A2(n20831), .B1(n20812), .B2(n20833), .ZN(
        P1_U3461) );
  INV_X1 U23780 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20815) );
  INV_X1 U23781 ( .A(n20816), .ZN(n20813) );
  AOI21_X1 U23782 ( .B1(n20815), .B2(n20814), .A(n20813), .ZN(P1_U3464) );
  OAI21_X1 U23783 ( .B1(n20818), .B2(n20817), .A(n20816), .ZN(P1_U3465) );
  INV_X1 U23784 ( .A(n20819), .ZN(n20823) );
  OAI22_X1 U23785 ( .A1(n20823), .A2(n20822), .B1(n20821), .B2(n20820), .ZN(
        n20825) );
  MUX2_X1 U23786 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n20825), .S(
        n20824), .Z(P1_U3469) );
  AOI21_X1 U23787 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20826) );
  AOI22_X1 U23788 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20826), .B2(n13735), .ZN(n20829) );
  AOI22_X1 U23789 ( .A1(n20832), .A2(n20829), .B1(n20828), .B2(n20827), .ZN(
        P1_U3481) );
  OAI21_X1 U23790 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20832), .ZN(n20830) );
  OAI21_X1 U23791 ( .B1(n20832), .B2(n20831), .A(n20830), .ZN(P1_U3482) );
  AOI22_X1 U23792 ( .A1(n20800), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20834), 
        .B2(n20833), .ZN(P1_U3483) );
  OAI211_X1 U23793 ( .C1(n20838), .C2(n20837), .A(n20836), .B(n20835), .ZN(
        n20839) );
  NOR2_X1 U23794 ( .A1(n20840), .A2(n20839), .ZN(n20847) );
  OAI211_X1 U23795 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20842), .A(n20841), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n20844) );
  AOI21_X1 U23796 ( .B1(n20844), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n20843), 
        .ZN(n20846) );
  NAND2_X1 U23797 ( .A1(n20847), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20845) );
  OAI21_X1 U23798 ( .B1(n20847), .B2(n20846), .A(n20845), .ZN(P1_U3485) );
  MUX2_X1 U23799 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(P1_MEMORYFETCH_REG_SCAN_IN), 
        .S(n20800), .Z(P1_U3486) );
  OAI21_X1 U23800 ( .B1(n20850), .B2(n20849), .A(n20848), .ZN(n20853) );
  NAND4_X1 U23801 ( .A1(P3_REQUESTPENDING_REG_SCAN_IN), .A2(n20853), .A3(
        n20852), .A4(n20851), .ZN(n20854) );
  AOI22_X1 U23802 ( .A1(NA), .A2(n20855), .B1(n18801), .B2(n20854), .ZN(n21167) );
  INV_X1 U23803 ( .A(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n20857) );
  AOI22_X1 U23804 ( .A1(n20858), .A2(keyinput85), .B1(n20857), .B2(keyinput108), .ZN(n20856) );
  OAI221_X1 U23805 ( .B1(n20858), .B2(keyinput85), .C1(n20857), .C2(
        keyinput108), .A(n20856), .ZN(n20871) );
  INV_X1 U23806 ( .A(keyinput16), .ZN(n20860) );
  AOI22_X1 U23807 ( .A1(n20861), .A2(keyinput93), .B1(P3_DATAO_REG_19__SCAN_IN), .B2(n20860), .ZN(n20859) );
  OAI221_X1 U23808 ( .B1(n20861), .B2(keyinput93), .C1(n20860), .C2(
        P3_DATAO_REG_19__SCAN_IN), .A(n20859), .ZN(n20870) );
  AOI22_X1 U23809 ( .A1(n20864), .A2(keyinput124), .B1(n20863), .B2(
        keyinput103), .ZN(n20862) );
  OAI221_X1 U23810 ( .B1(n20864), .B2(keyinput124), .C1(n20863), .C2(
        keyinput103), .A(n20862), .ZN(n20869) );
  AOI22_X1 U23811 ( .A1(n20867), .A2(keyinput125), .B1(n20866), .B2(keyinput56), .ZN(n20865) );
  OAI221_X1 U23812 ( .B1(n20867), .B2(keyinput125), .C1(n20866), .C2(
        keyinput56), .A(n20865), .ZN(n20868) );
  NOR4_X1 U23813 ( .A1(n20871), .A2(n20870), .A3(n20869), .A4(n20868), .ZN(
        n20922) );
  INV_X1 U23814 ( .A(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n20874) );
  INV_X1 U23815 ( .A(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n20873) );
  AOI22_X1 U23816 ( .A1(n20874), .A2(keyinput104), .B1(keyinput3), .B2(n20873), 
        .ZN(n20872) );
  OAI221_X1 U23817 ( .B1(n20874), .B2(keyinput104), .C1(n20873), .C2(keyinput3), .A(n20872), .ZN(n20886) );
  AOI22_X1 U23818 ( .A1(n20877), .A2(keyinput119), .B1(n20876), .B2(keyinput63), .ZN(n20875) );
  OAI221_X1 U23819 ( .B1(n20877), .B2(keyinput119), .C1(n20876), .C2(
        keyinput63), .A(n20875), .ZN(n20885) );
  INV_X1 U23820 ( .A(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n20879) );
  AOI22_X1 U23821 ( .A1(n20880), .A2(keyinput26), .B1(keyinput8), .B2(n20879), 
        .ZN(n20878) );
  OAI221_X1 U23822 ( .B1(n20880), .B2(keyinput26), .C1(n20879), .C2(keyinput8), 
        .A(n20878), .ZN(n20884) );
  INV_X1 U23823 ( .A(P3_LWORD_REG_10__SCAN_IN), .ZN(n20882) );
  AOI22_X1 U23824 ( .A1(n12653), .A2(keyinput43), .B1(keyinput120), .B2(n20882), .ZN(n20881) );
  OAI221_X1 U23825 ( .B1(n12653), .B2(keyinput43), .C1(n20882), .C2(
        keyinput120), .A(n20881), .ZN(n20883) );
  NOR4_X1 U23826 ( .A1(n20886), .A2(n20885), .A3(n20884), .A4(n20883), .ZN(
        n20921) );
  INV_X1 U23827 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n20888) );
  AOI22_X1 U23828 ( .A1(n20889), .A2(keyinput126), .B1(n20888), .B2(keyinput58), .ZN(n20887) );
  OAI221_X1 U23829 ( .B1(n20889), .B2(keyinput126), .C1(n20888), .C2(
        keyinput58), .A(n20887), .ZN(n20890) );
  INV_X1 U23830 ( .A(n20890), .ZN(n20894) );
  XOR2_X1 U23831 ( .A(keyinput61), .B(n20891), .Z(n20893) );
  XNOR2_X1 U23832 ( .A(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B(keyinput80), .ZN(
        n20892) );
  NAND3_X1 U23833 ( .A1(n20894), .A2(n20893), .A3(n20892), .ZN(n20903) );
  AOI22_X1 U23834 ( .A1(n20897), .A2(keyinput87), .B1(n20896), .B2(keyinput46), 
        .ZN(n20895) );
  OAI221_X1 U23835 ( .B1(n20897), .B2(keyinput87), .C1(n20896), .C2(keyinput46), .A(n20895), .ZN(n20902) );
  INV_X1 U23836 ( .A(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n20900) );
  INV_X1 U23837 ( .A(keyinput74), .ZN(n20899) );
  AOI22_X1 U23838 ( .A1(n20900), .A2(keyinput70), .B1(
        P3_DATAWIDTH_REG_2__SCAN_IN), .B2(n20899), .ZN(n20898) );
  OAI221_X1 U23839 ( .B1(n20900), .B2(keyinput70), .C1(n20899), .C2(
        P3_DATAWIDTH_REG_2__SCAN_IN), .A(n20898), .ZN(n20901) );
  NOR3_X1 U23840 ( .A1(n20903), .A2(n20902), .A3(n20901), .ZN(n20920) );
  INV_X1 U23841 ( .A(keyinput117), .ZN(n20905) );
  AOI22_X1 U23842 ( .A1(n19544), .A2(keyinput66), .B1(
        P1_DATAWIDTH_REG_27__SCAN_IN), .B2(n20905), .ZN(n20904) );
  OAI221_X1 U23843 ( .B1(n19544), .B2(keyinput66), .C1(n20905), .C2(
        P1_DATAWIDTH_REG_27__SCAN_IN), .A(n20904), .ZN(n20918) );
  INV_X1 U23844 ( .A(P2_UWORD_REG_6__SCAN_IN), .ZN(n20908) );
  AOI22_X1 U23845 ( .A1(n20908), .A2(keyinput4), .B1(n20907), .B2(keyinput111), 
        .ZN(n20906) );
  OAI221_X1 U23846 ( .B1(n20908), .B2(keyinput4), .C1(n20907), .C2(keyinput111), .A(n20906), .ZN(n20917) );
  INV_X1 U23847 ( .A(READY2), .ZN(n20910) );
  AOI22_X1 U23848 ( .A1(n20911), .A2(keyinput65), .B1(keyinput22), .B2(n20910), 
        .ZN(n20909) );
  OAI221_X1 U23849 ( .B1(n20911), .B2(keyinput65), .C1(n20910), .C2(keyinput22), .A(n20909), .ZN(n20916) );
  INV_X1 U23850 ( .A(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n20912) );
  XOR2_X1 U23851 ( .A(n20912), .B(keyinput123), .Z(n20914) );
  XNOR2_X1 U23852 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B(keyinput78), .ZN(
        n20913) );
  NAND2_X1 U23853 ( .A1(n20914), .A2(n20913), .ZN(n20915) );
  NOR4_X1 U23854 ( .A1(n20918), .A2(n20917), .A3(n20916), .A4(n20915), .ZN(
        n20919) );
  NAND4_X1 U23855 ( .A1(n20922), .A2(n20921), .A3(n20920), .A4(n20919), .ZN(
        n21165) );
  INV_X1 U23856 ( .A(P3_LWORD_REG_2__SCAN_IN), .ZN(n20925) );
  INV_X1 U23857 ( .A(keyinput114), .ZN(n20924) );
  AOI22_X1 U23858 ( .A1(n20925), .A2(keyinput105), .B1(
        P3_DATAWIDTH_REG_11__SCAN_IN), .B2(n20924), .ZN(n20923) );
  OAI221_X1 U23859 ( .B1(n20925), .B2(keyinput105), .C1(n20924), .C2(
        P3_DATAWIDTH_REG_11__SCAN_IN), .A(n20923), .ZN(n20937) );
  INV_X1 U23860 ( .A(keyinput12), .ZN(n20927) );
  AOI22_X1 U23861 ( .A1(n20928), .A2(keyinput29), .B1(
        P3_ADDRESS_REG_8__SCAN_IN), .B2(n20927), .ZN(n20926) );
  OAI221_X1 U23862 ( .B1(n20928), .B2(keyinput29), .C1(n20927), .C2(
        P3_ADDRESS_REG_8__SCAN_IN), .A(n20926), .ZN(n20936) );
  INV_X1 U23863 ( .A(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n20930) );
  AOI22_X1 U23864 ( .A1(n20931), .A2(keyinput106), .B1(n20930), .B2(keyinput48), .ZN(n20929) );
  OAI221_X1 U23865 ( .B1(n20931), .B2(keyinput106), .C1(n20930), .C2(
        keyinput48), .A(n20929), .ZN(n20935) );
  XNOR2_X1 U23866 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B(keyinput0), .ZN(
        n20933) );
  XNOR2_X1 U23867 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B(keyinput72), .ZN(
        n20932) );
  NAND2_X1 U23868 ( .A1(n20933), .A2(n20932), .ZN(n20934) );
  NOR4_X1 U23869 ( .A1(n20937), .A2(n20936), .A3(n20935), .A4(n20934), .ZN(
        n20982) );
  INV_X1 U23870 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n20940) );
  INV_X1 U23871 ( .A(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n20939) );
  AOI22_X1 U23872 ( .A1(n20940), .A2(keyinput18), .B1(keyinput42), .B2(n20939), 
        .ZN(n20938) );
  OAI221_X1 U23873 ( .B1(n20940), .B2(keyinput18), .C1(n20939), .C2(keyinput42), .A(n20938), .ZN(n20951) );
  AOI22_X1 U23874 ( .A1(n20943), .A2(keyinput97), .B1(keyinput92), .B2(n20942), 
        .ZN(n20941) );
  OAI221_X1 U23875 ( .B1(n20943), .B2(keyinput97), .C1(n20942), .C2(keyinput92), .A(n20941), .ZN(n20950) );
  INV_X1 U23876 ( .A(keyinput45), .ZN(n20945) );
  AOI22_X1 U23877 ( .A1(n13292), .A2(keyinput121), .B1(
        P3_DATAWIDTH_REG_30__SCAN_IN), .B2(n20945), .ZN(n20944) );
  OAI221_X1 U23878 ( .B1(n13292), .B2(keyinput121), .C1(n20945), .C2(
        P3_DATAWIDTH_REG_30__SCAN_IN), .A(n20944), .ZN(n20949) );
  XNOR2_X1 U23879 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(keyinput76), 
        .ZN(n20947) );
  XNOR2_X1 U23880 ( .A(P1_EAX_REG_4__SCAN_IN), .B(keyinput57), .ZN(n20946) );
  NAND2_X1 U23881 ( .A1(n20947), .A2(n20946), .ZN(n20948) );
  NOR4_X1 U23882 ( .A1(n20951), .A2(n20950), .A3(n20949), .A4(n20948), .ZN(
        n20981) );
  AOI22_X1 U23883 ( .A1(n20954), .A2(keyinput7), .B1(n20953), .B2(keyinput68), 
        .ZN(n20952) );
  OAI221_X1 U23884 ( .B1(n20954), .B2(keyinput7), .C1(n20953), .C2(keyinput68), 
        .A(n20952), .ZN(n20964) );
  AOI22_X1 U23885 ( .A1(n12832), .A2(keyinput15), .B1(keyinput118), .B2(n10840), .ZN(n20955) );
  OAI221_X1 U23886 ( .B1(n12832), .B2(keyinput15), .C1(n10840), .C2(
        keyinput118), .A(n20955), .ZN(n20963) );
  INV_X1 U23887 ( .A(DATAI_19_), .ZN(n20957) );
  AOI22_X1 U23888 ( .A1(n20958), .A2(keyinput35), .B1(keyinput95), .B2(n20957), 
        .ZN(n20956) );
  OAI221_X1 U23889 ( .B1(n20958), .B2(keyinput35), .C1(n20957), .C2(keyinput95), .A(n20956), .ZN(n20962) );
  INV_X1 U23890 ( .A(keyinput62), .ZN(n20960) );
  AOI22_X1 U23891 ( .A1(n10855), .A2(keyinput81), .B1(
        P3_DATAWIDTH_REG_14__SCAN_IN), .B2(n20960), .ZN(n20959) );
  OAI221_X1 U23892 ( .B1(n10855), .B2(keyinput81), .C1(n20960), .C2(
        P3_DATAWIDTH_REG_14__SCAN_IN), .A(n20959), .ZN(n20961) );
  NOR4_X1 U23893 ( .A1(n20964), .A2(n20963), .A3(n20962), .A4(n20961), .ZN(
        n20980) );
  INV_X1 U23894 ( .A(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n20966) );
  AOI22_X1 U23895 ( .A1(n20966), .A2(keyinput73), .B1(n11841), .B2(keyinput32), 
        .ZN(n20965) );
  OAI221_X1 U23896 ( .B1(n20966), .B2(keyinput73), .C1(n11841), .C2(keyinput32), .A(n20965), .ZN(n20978) );
  AOI22_X1 U23897 ( .A1(n20968), .A2(keyinput64), .B1(n11114), .B2(keyinput1), 
        .ZN(n20967) );
  OAI221_X1 U23898 ( .B1(n20968), .B2(keyinput64), .C1(n11114), .C2(keyinput1), 
        .A(n20967), .ZN(n20977) );
  AOI22_X1 U23899 ( .A1(n20971), .A2(keyinput33), .B1(n20970), .B2(keyinput47), 
        .ZN(n20969) );
  OAI221_X1 U23900 ( .B1(n20971), .B2(keyinput33), .C1(n20970), .C2(keyinput47), .A(n20969), .ZN(n20976) );
  AOI22_X1 U23901 ( .A1(n20974), .A2(keyinput77), .B1(n20973), .B2(keyinput89), 
        .ZN(n20972) );
  OAI221_X1 U23902 ( .B1(n20974), .B2(keyinput77), .C1(n20973), .C2(keyinput89), .A(n20972), .ZN(n20975) );
  NOR4_X1 U23903 ( .A1(n20978), .A2(n20977), .A3(n20976), .A4(n20975), .ZN(
        n20979) );
  NAND4_X1 U23904 ( .A1(n20982), .A2(n20981), .A3(n20980), .A4(n20979), .ZN(
        n21164) );
  AOI22_X1 U23905 ( .A1(n20984), .A2(keyinput91), .B1(n15001), .B2(keyinput99), 
        .ZN(n20983) );
  OAI221_X1 U23906 ( .B1(n20984), .B2(keyinput91), .C1(n15001), .C2(keyinput99), .A(n20983), .ZN(n20997) );
  AOI22_X1 U23907 ( .A1(n20987), .A2(keyinput101), .B1(keyinput82), .B2(n20986), .ZN(n20985) );
  OAI221_X1 U23908 ( .B1(n20987), .B2(keyinput101), .C1(n20986), .C2(
        keyinput82), .A(n20985), .ZN(n20996) );
  AOI22_X1 U23909 ( .A1(n20990), .A2(keyinput25), .B1(n20989), .B2(keyinput59), 
        .ZN(n20988) );
  OAI221_X1 U23910 ( .B1(n20990), .B2(keyinput25), .C1(n20989), .C2(keyinput59), .A(n20988), .ZN(n20995) );
  INV_X1 U23911 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n20993) );
  INV_X1 U23912 ( .A(keyinput30), .ZN(n20992) );
  AOI22_X1 U23913 ( .A1(n20993), .A2(keyinput20), .B1(
        P1_DATAWIDTH_REG_10__SCAN_IN), .B2(n20992), .ZN(n20991) );
  OAI221_X1 U23914 ( .B1(n20993), .B2(keyinput20), .C1(n20992), .C2(
        P1_DATAWIDTH_REG_10__SCAN_IN), .A(n20991), .ZN(n20994) );
  NOR4_X1 U23915 ( .A1(n20997), .A2(n20996), .A3(n20995), .A4(n20994), .ZN(
        n21044) );
  INV_X1 U23916 ( .A(P3_DATAO_REG_27__SCAN_IN), .ZN(n21000) );
  INV_X1 U23917 ( .A(keyinput102), .ZN(n20999) );
  AOI22_X1 U23918 ( .A1(n21000), .A2(keyinput79), .B1(
        P1_DATAWIDTH_REG_26__SCAN_IN), .B2(n20999), .ZN(n20998) );
  OAI221_X1 U23919 ( .B1(n21000), .B2(keyinput79), .C1(n20999), .C2(
        P1_DATAWIDTH_REG_26__SCAN_IN), .A(n20998), .ZN(n21013) );
  AOI22_X1 U23920 ( .A1(n21003), .A2(keyinput17), .B1(keyinput49), .B2(n21002), 
        .ZN(n21001) );
  OAI221_X1 U23921 ( .B1(n21003), .B2(keyinput17), .C1(n21002), .C2(keyinput49), .A(n21001), .ZN(n21012) );
  INV_X1 U23922 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n21006) );
  AOI22_X1 U23923 ( .A1(n21006), .A2(keyinput14), .B1(keyinput10), .B2(n21005), 
        .ZN(n21004) );
  OAI221_X1 U23924 ( .B1(n21006), .B2(keyinput14), .C1(n21005), .C2(keyinput10), .A(n21004), .ZN(n21011) );
  INV_X1 U23925 ( .A(P1_EAX_REG_31__SCAN_IN), .ZN(n21009) );
  AOI22_X1 U23926 ( .A1(n21009), .A2(keyinput13), .B1(n21008), .B2(keyinput52), 
        .ZN(n21007) );
  OAI221_X1 U23927 ( .B1(n21009), .B2(keyinput13), .C1(n21008), .C2(keyinput52), .A(n21007), .ZN(n21010) );
  NOR4_X1 U23928 ( .A1(n21013), .A2(n21012), .A3(n21011), .A4(n21010), .ZN(
        n21043) );
  AOI22_X1 U23929 ( .A1(n21016), .A2(keyinput11), .B1(keyinput23), .B2(n21015), 
        .ZN(n21014) );
  OAI221_X1 U23930 ( .B1(n21016), .B2(keyinput11), .C1(n21015), .C2(keyinput23), .A(n21014), .ZN(n21027) );
  INV_X1 U23931 ( .A(P2_UWORD_REG_11__SCAN_IN), .ZN(n21018) );
  AOI22_X1 U23932 ( .A1(n21019), .A2(keyinput83), .B1(keyinput88), .B2(n21018), 
        .ZN(n21017) );
  OAI221_X1 U23933 ( .B1(n21019), .B2(keyinput83), .C1(n21018), .C2(keyinput88), .A(n21017), .ZN(n21026) );
  INV_X1 U23934 ( .A(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n21020) );
  XOR2_X1 U23935 ( .A(n21020), .B(keyinput94), .Z(n21024) );
  XNOR2_X1 U23936 ( .A(keyinput115), .B(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n21023) );
  XNOR2_X1 U23937 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(keyinput84), 
        .ZN(n21022) );
  XNOR2_X1 U23938 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B(keyinput6), .ZN(
        n21021) );
  NAND4_X1 U23939 ( .A1(n21024), .A2(n21023), .A3(n21022), .A4(n21021), .ZN(
        n21025) );
  NOR3_X1 U23940 ( .A1(n21027), .A2(n21026), .A3(n21025), .ZN(n21042) );
  AOI22_X1 U23941 ( .A1(n21030), .A2(keyinput31), .B1(keyinput28), .B2(n21029), 
        .ZN(n21028) );
  OAI221_X1 U23942 ( .B1(n21030), .B2(keyinput31), .C1(n21029), .C2(keyinput28), .A(n21028), .ZN(n21040) );
  INV_X1 U23943 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n21032) );
  AOI22_X1 U23944 ( .A1(n13542), .A2(keyinput50), .B1(n21032), .B2(keyinput55), 
        .ZN(n21031) );
  OAI221_X1 U23945 ( .B1(n13542), .B2(keyinput50), .C1(n21032), .C2(keyinput55), .A(n21031), .ZN(n21039) );
  AOI22_X1 U23946 ( .A1(n21034), .A2(keyinput109), .B1(keyinput98), .B2(n14179), .ZN(n21033) );
  OAI221_X1 U23947 ( .B1(n21034), .B2(keyinput109), .C1(n14179), .C2(
        keyinput98), .A(n21033), .ZN(n21038) );
  INV_X1 U23948 ( .A(keyinput75), .ZN(n21036) );
  AOI22_X1 U23949 ( .A1(n11208), .A2(keyinput5), .B1(P3_ADDRESS_REG_0__SCAN_IN), .B2(n21036), .ZN(n21035) );
  OAI221_X1 U23950 ( .B1(n11208), .B2(keyinput5), .C1(n21036), .C2(
        P3_ADDRESS_REG_0__SCAN_IN), .A(n21035), .ZN(n21037) );
  NOR4_X1 U23951 ( .A1(n21040), .A2(n21039), .A3(n21038), .A4(n21037), .ZN(
        n21041) );
  NAND4_X1 U23952 ( .A1(n21044), .A2(n21043), .A3(n21042), .A4(n21041), .ZN(
        n21163) );
  AOI22_X1 U23953 ( .A1(n21046), .A2(keyinput34), .B1(n11740), .B2(keyinput51), 
        .ZN(n21045) );
  OAI221_X1 U23954 ( .B1(n21046), .B2(keyinput34), .C1(n11740), .C2(keyinput51), .A(n21045), .ZN(n21058) );
  INV_X1 U23955 ( .A(DATAI_0_), .ZN(n21049) );
  AOI22_X1 U23956 ( .A1(n21049), .A2(keyinput122), .B1(n21048), .B2(keyinput60), .ZN(n21047) );
  OAI221_X1 U23957 ( .B1(n21049), .B2(keyinput122), .C1(n21048), .C2(
        keyinput60), .A(n21047), .ZN(n21057) );
  XOR2_X1 U23958 ( .A(n21050), .B(keyinput19), .Z(n21055) );
  XOR2_X1 U23959 ( .A(n21051), .B(keyinput37), .Z(n21054) );
  XNOR2_X1 U23960 ( .A(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B(keyinput86), .ZN(
        n21053) );
  XNOR2_X1 U23961 ( .A(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B(keyinput127), .ZN(
        n21052) );
  NAND4_X1 U23962 ( .A1(n21055), .A2(n21054), .A3(n21053), .A4(n21052), .ZN(
        n21056) );
  NOR3_X1 U23963 ( .A1(n21058), .A2(n21057), .A3(n21056), .ZN(n21161) );
  INV_X1 U23964 ( .A(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n21061) );
  INV_X1 U23965 ( .A(keyinput36), .ZN(n21060) );
  AOI22_X1 U23966 ( .A1(n21061), .A2(keyinput54), .B1(
        P3_BYTEENABLE_REG_0__SCAN_IN), .B2(n21060), .ZN(n21059) );
  OAI221_X1 U23967 ( .B1(n21061), .B2(keyinput54), .C1(n21060), .C2(
        P3_BYTEENABLE_REG_0__SCAN_IN), .A(n21059), .ZN(n21073) );
  INV_X1 U23968 ( .A(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n21064) );
  AOI22_X1 U23969 ( .A1(n21064), .A2(keyinput107), .B1(keyinput90), .B2(n21063), .ZN(n21062) );
  OAI221_X1 U23970 ( .B1(n21064), .B2(keyinput107), .C1(n21063), .C2(
        keyinput90), .A(n21062), .ZN(n21072) );
  AOI22_X1 U23971 ( .A1(n21066), .A2(keyinput2), .B1(n10495), .B2(keyinput113), 
        .ZN(n21065) );
  OAI221_X1 U23972 ( .B1(n21066), .B2(keyinput2), .C1(n10495), .C2(keyinput113), .A(n21065), .ZN(n21071) );
  INV_X1 U23973 ( .A(keyinput69), .ZN(n21067) );
  XOR2_X1 U23974 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n21067), .Z(n21069) );
  XNOR2_X1 U23975 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B(keyinput27), .ZN(
        n21068) );
  NAND2_X1 U23976 ( .A1(n21069), .A2(n21068), .ZN(n21070) );
  NOR4_X1 U23977 ( .A1(n21073), .A2(n21072), .A3(n21071), .A4(n21070), .ZN(
        n21160) );
  INV_X1 U23978 ( .A(keyinput44), .ZN(n21075) );
  OAI22_X1 U23979 ( .A1(n21076), .A2(keyinput112), .B1(n21075), .B2(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n21074) );
  AOI221_X1 U23980 ( .B1(n21076), .B2(keyinput112), .C1(
        P2_DATAWIDTH_REG_31__SCAN_IN), .C2(n21075), .A(n21074), .ZN(n21089) );
  OAI22_X1 U23981 ( .A1(n21079), .A2(keyinput67), .B1(n21078), .B2(keyinput71), 
        .ZN(n21077) );
  AOI221_X1 U23982 ( .B1(n21079), .B2(keyinput67), .C1(keyinput71), .C2(n21078), .A(n21077), .ZN(n21088) );
  OAI22_X1 U23983 ( .A1(keyinput110), .A2(n21082), .B1(n21081), .B2(keyinput41), .ZN(n21080) );
  AOI221_X1 U23984 ( .B1(n21082), .B2(keyinput110), .C1(n21081), .C2(
        keyinput41), .A(n21080), .ZN(n21087) );
  INV_X1 U23985 ( .A(keyinput38), .ZN(n21084) );
  OAI22_X1 U23986 ( .A1(n21085), .A2(keyinput96), .B1(n21084), .B2(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n21083) );
  AOI221_X1 U23987 ( .B1(n21085), .B2(keyinput96), .C1(
        P1_DATAWIDTH_REG_15__SCAN_IN), .C2(n21084), .A(n21083), .ZN(n21086) );
  NAND4_X1 U23988 ( .A1(n21089), .A2(n21088), .A3(n21087), .A4(n21086), .ZN(
        n21104) );
  AOI22_X1 U23989 ( .A1(n21092), .A2(keyinput9), .B1(n21091), .B2(keyinput116), 
        .ZN(n21090) );
  OAI221_X1 U23990 ( .B1(n21092), .B2(keyinput9), .C1(n21091), .C2(keyinput116), .A(n21090), .ZN(n21103) );
  AOI22_X1 U23991 ( .A1(n12111), .A2(keyinput53), .B1(keyinput40), .B2(n21094), 
        .ZN(n21093) );
  OAI221_X1 U23992 ( .B1(n12111), .B2(keyinput53), .C1(n21094), .C2(keyinput40), .A(n21093), .ZN(n21097) );
  XOR2_X1 U23993 ( .A(keyinput21), .B(P3_ADDRESS_REG_16__SCAN_IN), .Z(n21096)
         );
  XNOR2_X1 U23994 ( .A(n11566), .B(keyinput39), .ZN(n21095) );
  OR3_X1 U23995 ( .A1(n21097), .A2(n21096), .A3(n21095), .ZN(n21102) );
  INV_X1 U23996 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n21099) );
  AOI22_X1 U23997 ( .A1(n21100), .A2(keyinput100), .B1(n21099), .B2(keyinput24), .ZN(n21098) );
  OAI221_X1 U23998 ( .B1(n21100), .B2(keyinput100), .C1(n21099), .C2(
        keyinput24), .A(n21098), .ZN(n21101) );
  NOR4_X1 U23999 ( .A1(n21104), .A2(n21103), .A3(n21102), .A4(n21101), .ZN(
        n21159) );
  NAND2_X1 U24000 ( .A1(keyinput25), .A2(keyinput101), .ZN(n21105) );
  NOR3_X1 U24001 ( .A1(keyinput82), .A2(keyinput59), .A3(n21105), .ZN(n21106)
         );
  NAND3_X1 U24002 ( .A1(keyinput20), .A2(keyinput30), .A3(n21106), .ZN(n21118)
         );
  NAND4_X1 U24003 ( .A1(keyinput115), .A2(keyinput84), .A3(keyinput94), .A4(
        keyinput6), .ZN(n21107) );
  NOR3_X1 U24004 ( .A1(keyinput11), .A2(keyinput23), .A3(n21107), .ZN(n21116)
         );
  INV_X1 U24005 ( .A(keyinput52), .ZN(n21108) );
  NAND4_X1 U24006 ( .A1(keyinput13), .A2(keyinput14), .A3(keyinput10), .A4(
        n21108), .ZN(n21114) );
  NOR2_X1 U24007 ( .A1(keyinput49), .A2(keyinput102), .ZN(n21109) );
  NAND3_X1 U24008 ( .A1(keyinput17), .A2(keyinput79), .A3(n21109), .ZN(n21113)
         );
  NOR3_X1 U24009 ( .A1(keyinput31), .A2(keyinput5), .A3(keyinput28), .ZN(
        n21110) );
  NAND2_X1 U24010 ( .A1(keyinput75), .A2(n21110), .ZN(n21112) );
  NAND4_X1 U24011 ( .A1(keyinput50), .A2(keyinput55), .A3(keyinput109), .A4(
        keyinput98), .ZN(n21111) );
  NOR4_X1 U24012 ( .A1(n21114), .A2(n21113), .A3(n21112), .A4(n21111), .ZN(
        n21115) );
  NAND4_X1 U24013 ( .A1(keyinput83), .A2(keyinput88), .A3(n21116), .A4(n21115), 
        .ZN(n21117) );
  NOR4_X1 U24014 ( .A1(keyinput91), .A2(keyinput99), .A3(n21118), .A4(n21117), 
        .ZN(n21157) );
  NAND4_X1 U24015 ( .A1(keyinput56), .A2(keyinput60), .A3(keyinput22), .A4(
        keyinput61), .ZN(n21122) );
  NAND4_X1 U24016 ( .A1(keyinput80), .A2(keyinput96), .A3(keyinput93), .A4(
        keyinput69), .ZN(n21121) );
  NAND4_X1 U24017 ( .A1(keyinput63), .A2(keyinput46), .A3(keyinput108), .A4(
        keyinput116), .ZN(n21120) );
  NAND4_X1 U24018 ( .A1(keyinput27), .A2(keyinput3), .A3(keyinput51), .A4(
        keyinput54), .ZN(n21119) );
  NOR4_X1 U24019 ( .A1(n21122), .A2(n21121), .A3(n21120), .A4(n21119), .ZN(
        n21156) );
  NAND4_X1 U24020 ( .A1(keyinput70), .A2(keyinput71), .A3(keyinput74), .A4(
        keyinput103), .ZN(n21127) );
  INV_X1 U24021 ( .A(keyinput104), .ZN(n21123) );
  NAND4_X1 U24022 ( .A1(keyinput122), .A2(keyinput119), .A3(keyinput127), .A4(
        n21123), .ZN(n21126) );
  NAND4_X1 U24023 ( .A1(keyinput8), .A2(keyinput9), .A3(keyinput24), .A4(
        keyinput16), .ZN(n21125) );
  NAND4_X1 U24024 ( .A1(keyinput111), .A2(keyinput41), .A3(keyinput37), .A4(
        keyinput40), .ZN(n21124) );
  NOR4_X1 U24025 ( .A1(n21127), .A2(n21126), .A3(n21125), .A4(n21124), .ZN(
        n21155) );
  INV_X1 U24026 ( .A(keyinput72), .ZN(n21128) );
  NAND4_X1 U24027 ( .A1(keyinput0), .A2(keyinput106), .A3(keyinput48), .A4(
        n21128), .ZN(n21129) );
  NOR3_X1 U24028 ( .A1(keyinput105), .A2(keyinput114), .A3(n21129), .ZN(n21142) );
  NAND2_X1 U24029 ( .A1(keyinput42), .A2(keyinput92), .ZN(n21130) );
  NOR3_X1 U24030 ( .A1(keyinput97), .A2(keyinput18), .A3(n21130), .ZN(n21131)
         );
  NAND3_X1 U24031 ( .A1(keyinput76), .A2(keyinput57), .A3(n21131), .ZN(n21140)
         );
  INV_X1 U24032 ( .A(keyinput33), .ZN(n21132) );
  NOR4_X1 U24033 ( .A1(keyinput77), .A2(keyinput89), .A3(keyinput47), .A4(
        n21132), .ZN(n21138) );
  NAND2_X1 U24034 ( .A1(keyinput32), .A2(keyinput64), .ZN(n21133) );
  NOR3_X1 U24035 ( .A1(keyinput73), .A2(keyinput1), .A3(n21133), .ZN(n21137)
         );
  NAND2_X1 U24036 ( .A1(keyinput35), .A2(keyinput68), .ZN(n21134) );
  NOR3_X1 U24037 ( .A1(keyinput7), .A2(keyinput95), .A3(n21134), .ZN(n21136)
         );
  NOR4_X1 U24038 ( .A1(keyinput15), .A2(keyinput118), .A3(keyinput81), .A4(
        keyinput62), .ZN(n21135) );
  NAND4_X1 U24039 ( .A1(n21138), .A2(n21137), .A3(n21136), .A4(n21135), .ZN(
        n21139) );
  NOR4_X1 U24040 ( .A1(keyinput121), .A2(keyinput45), .A3(n21140), .A4(n21139), 
        .ZN(n21141) );
  NAND4_X1 U24041 ( .A1(keyinput29), .A2(keyinput12), .A3(n21142), .A4(n21141), 
        .ZN(n21153) );
  NOR4_X1 U24042 ( .A1(keyinput53), .A2(keyinput65), .A3(keyinput4), .A4(
        keyinput21), .ZN(n21146) );
  NOR4_X1 U24043 ( .A1(keyinput38), .A2(keyinput43), .A3(keyinput36), .A4(
        keyinput44), .ZN(n21145) );
  NOR4_X1 U24044 ( .A1(keyinput124), .A2(keyinput125), .A3(keyinput85), .A4(
        keyinput100), .ZN(n21144) );
  NOR4_X1 U24045 ( .A1(keyinput112), .A2(keyinput113), .A3(keyinput117), .A4(
        keyinput120), .ZN(n21143) );
  NAND4_X1 U24046 ( .A1(n21146), .A2(n21145), .A3(n21144), .A4(n21143), .ZN(
        n21152) );
  NOR4_X1 U24047 ( .A1(keyinput78), .A2(keyinput107), .A3(keyinput110), .A4(
        keyinput87), .ZN(n21150) );
  NOR4_X1 U24048 ( .A1(keyinput123), .A2(keyinput126), .A3(keyinput67), .A4(
        keyinput66), .ZN(n21149) );
  NOR4_X1 U24049 ( .A1(keyinput2), .A2(keyinput58), .A3(keyinput34), .A4(
        keyinput39), .ZN(n21148) );
  NOR4_X1 U24050 ( .A1(keyinput86), .A2(keyinput90), .A3(keyinput19), .A4(
        keyinput26), .ZN(n21147) );
  NAND4_X1 U24051 ( .A1(n21150), .A2(n21149), .A3(n21148), .A4(n21147), .ZN(
        n21151) );
  NOR3_X1 U24052 ( .A1(n21153), .A2(n21152), .A3(n21151), .ZN(n21154) );
  NAND4_X1 U24053 ( .A1(n21157), .A2(n21156), .A3(n21155), .A4(n21154), .ZN(
        n21158) );
  NAND4_X1 U24054 ( .A1(n21161), .A2(n21160), .A3(n21159), .A4(n21158), .ZN(
        n21162) );
  NOR4_X1 U24055 ( .A1(n21165), .A2(n21164), .A3(n21163), .A4(n21162), .ZN(
        n21166) );
  XNOR2_X1 U24056 ( .A(n21167), .B(n21166), .ZN(P3_U3029) );
  XNOR2_X1 U13341 ( .A(n10352), .B(n10348), .ZN(n12528) );
  INV_X1 U11196 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19680) );
  INV_X1 U11301 ( .A(n14126), .ZN(n13216) );
  CLKBUF_X1 U11195 ( .A(n12318), .Z(n12248) );
  CLKBUF_X1 U11237 ( .A(n11099), .Z(n12696) );
  AND2_X1 U11250 ( .A1(n10268), .A2(n10267), .ZN(n10958) );
  CLKBUF_X1 U11252 ( .A(n10252), .Z(n12509) );
  NOR2_X1 U11266 ( .A1(n10353), .A2(n10360), .ZN(n10363) );
  CLKBUF_X1 U11268 ( .A(n11477), .Z(n9786) );
  CLKBUF_X1 U11302 ( .A(n11461), .Z(n11466) );
  CLKBUF_X1 U11341 ( .A(n11476), .Z(n14652) );
  OAI221_X2 U11343 ( .B1(n14670), .B2(n16368), .C1(n15363), .C2(n16368), .A(
        n18894), .ZN(n19424) );
  CLKBUF_X1 U11493 ( .A(n17463), .Z(n9783) );
  CLKBUF_X1 U11564 ( .A(n12528), .Z(n9792) );
  INV_X1 U11580 ( .A(n14704), .ZN(n19032) );
  CLKBUF_X2 U11600 ( .A(n11013), .Z(n9788) );
  CLKBUF_X1 U11605 ( .A(n15006), .Z(n16215) );
  CLKBUF_X1 U11849 ( .A(n17775), .Z(n9754) );
  CLKBUF_X1 U11970 ( .A(n17256), .Z(n9756) );
endmodule

