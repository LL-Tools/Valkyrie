

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
         n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
         n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
         n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
         n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
         n12125, n12126, n12127, n12128, n12129, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
         n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
         n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
         n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
         n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
         n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
         n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
         n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
         n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
         n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
         n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
         n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
         n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
         n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
         n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
         n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
         n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325,
         n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333,
         n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
         n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
         n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
         n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
         n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
         n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
         n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
         n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
         n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
         n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429,
         n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
         n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
         n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
         n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
         n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
         n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477,
         n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
         n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
         n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501,
         n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
         n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
         n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
         n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533,
         n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
         n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549,
         n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
         n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565,
         n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573,
         n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
         n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
         n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
         n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621,
         n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
         n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
         n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
         n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
         n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
         n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
         n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
         n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
         n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
         n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
         n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
         n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
         n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
         n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
         n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
         n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
         n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
         n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
         n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
         n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
         n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541,
         n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549,
         n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
         n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
         n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
         n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
         n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669,
         n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
         n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
         n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
         n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
         n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
         n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
         n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
         n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
         n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
         n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
         n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
         n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
         n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
         n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
         n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
         n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
         n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
         n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
         n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
         n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885,
         n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
         n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901,
         n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909,
         n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
         n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
         n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
         n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957,
         n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
         n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973,
         n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981,
         n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989,
         n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
         n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005,
         n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
         n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
         n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
         n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
         n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
         n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
         n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
         n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
         n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
         n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
         n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125,
         n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
         n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
         n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
         n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
         n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
         n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173,
         n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
         n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189,
         n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197,
         n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
         n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
         n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221,
         n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
         n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
         n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245,
         n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
         n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261,
         n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
         n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
         n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
         n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293,
         n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
         n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
         n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317,
         n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
         n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333,
         n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341,
         n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349,
         n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
         n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365,
         n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373,
         n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381,
         n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389,
         n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397,
         n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405,
         n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413,
         n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421,
         n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429,
         n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437,
         n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445,
         n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453,
         n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461,
         n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469,
         n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477,
         n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485,
         n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493,
         n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501,
         n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509,
         n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517,
         n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525,
         n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533,
         n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541,
         n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549,
         n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557,
         n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565,
         n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573,
         n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581,
         n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589,
         n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597,
         n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605,
         n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613,
         n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621,
         n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629,
         n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637,
         n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645,
         n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653,
         n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661,
         n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669,
         n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677,
         n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685,
         n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693,
         n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701,
         n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709,
         n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717,
         n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725,
         n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733,
         n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741,
         n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749,
         n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757,
         n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765,
         n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773,
         n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781,
         n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789,
         n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797,
         n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805,
         n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813,
         n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821,
         n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829,
         n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837,
         n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845,
         n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853,
         n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861,
         n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869,
         n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877,
         n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885,
         n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893,
         n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901,
         n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909,
         n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917,
         n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925,
         n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933,
         n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941,
         n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949,
         n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957,
         n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965,
         n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973,
         n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981,
         n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989,
         n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997,
         n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005,
         n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013,
         n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021,
         n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029,
         n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037,
         n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045,
         n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053,
         n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061,
         n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069,
         n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077,
         n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085,
         n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093,
         n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101,
         n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109,
         n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117,
         n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125,
         n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133,
         n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141,
         n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149,
         n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157,
         n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165,
         n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173,
         n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181,
         n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189,
         n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197,
         n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205,
         n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213,
         n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221,
         n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229,
         n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237,
         n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245,
         n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253,
         n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261,
         n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269,
         n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277,
         n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285,
         n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293,
         n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301,
         n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309,
         n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317,
         n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325,
         n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333,
         n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341,
         n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349,
         n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357,
         n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365,
         n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373,
         n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381,
         n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389,
         n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397,
         n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405,
         n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413,
         n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421,
         n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429,
         n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437,
         n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445,
         n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453,
         n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461,
         n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469,
         n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
         n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485,
         n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493,
         n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501,
         n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509,
         n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517,
         n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525,
         n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533,
         n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541,
         n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549,
         n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557,
         n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565,
         n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573,
         n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581,
         n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589,
         n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597,
         n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605,
         n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613,
         n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
         n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629,
         n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637,
         n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645,
         n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653,
         n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661,
         n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669,
         n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677,
         n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685,
         n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693,
         n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701,
         n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709,
         n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717,
         n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725,
         n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733,
         n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741,
         n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749,
         n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757,
         n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765,
         n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773,
         n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781,
         n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789,
         n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797,
         n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805,
         n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813,
         n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821,
         n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829,
         n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837,
         n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845,
         n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853,
         n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861,
         n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869,
         n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877,
         n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885,
         n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893,
         n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901,
         n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909,
         n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917,
         n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925,
         n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933,
         n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941,
         n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949,
         n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957,
         n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965,
         n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973,
         n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981,
         n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989,
         n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997,
         n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005,
         n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013,
         n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021,
         n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029,
         n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037,
         n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045,
         n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053,
         n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061,
         n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069,
         n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077,
         n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085,
         n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093,
         n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101,
         n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109,
         n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117,
         n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125,
         n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133,
         n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141,
         n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149,
         n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157,
         n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165,
         n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173,
         n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181,
         n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189,
         n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197,
         n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205,
         n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213,
         n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221,
         n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229,
         n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237,
         n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245,
         n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253,
         n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261,
         n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269,
         n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277,
         n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285,
         n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293,
         n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301,
         n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309,
         n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317,
         n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325,
         n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333,
         n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341,
         n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349,
         n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357,
         n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365,
         n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373,
         n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381,
         n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389,
         n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397,
         n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405,
         n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413,
         n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421,
         n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429,
         n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437,
         n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445,
         n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453,
         n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461,
         n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469,
         n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477,
         n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485,
         n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493,
         n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501,
         n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509,
         n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517,
         n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525,
         n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533,
         n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541,
         n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549,
         n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557,
         n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565,
         n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573,
         n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581,
         n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589,
         n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597,
         n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605,
         n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613,
         n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621,
         n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629,
         n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637,
         n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645,
         n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653,
         n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661,
         n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669,
         n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677,
         n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685,
         n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693,
         n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701,
         n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709,
         n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717,
         n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725,
         n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733,
         n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741,
         n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749,
         n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757,
         n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765,
         n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773,
         n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781,
         n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789,
         n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797,
         n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805,
         n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813,
         n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821,
         n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829,
         n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837,
         n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845,
         n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853,
         n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861,
         n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869,
         n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877,
         n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885,
         n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893,
         n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901,
         n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909,
         n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917,
         n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925,
         n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933,
         n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941,
         n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949,
         n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957,
         n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965,
         n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973,
         n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981,
         n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989,
         n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997,
         n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005,
         n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013,
         n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021,
         n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029,
         n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037,
         n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045,
         n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053,
         n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061,
         n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069,
         n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077,
         n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085,
         n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093,
         n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101,
         n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109,
         n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117,
         n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125,
         n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133,
         n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141,
         n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149,
         n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157,
         n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165,
         n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173,
         n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181,
         n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189,
         n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197,
         n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205,
         n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213,
         n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221,
         n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229,
         n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237,
         n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245,
         n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253,
         n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261,
         n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269,
         n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277,
         n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285,
         n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293,
         n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301,
         n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309,
         n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317,
         n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325,
         n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333,
         n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341,
         n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349,
         n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357,
         n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365,
         n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373,
         n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381,
         n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389,
         n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397,
         n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405,
         n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413,
         n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421,
         n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429,
         n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437,
         n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445,
         n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453,
         n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461,
         n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469,
         n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477,
         n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485,
         n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493,
         n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501,
         n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509,
         n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517,
         n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525,
         n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533,
         n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541,
         n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549,
         n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557,
         n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565,
         n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573,
         n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581,
         n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589,
         n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597,
         n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605,
         n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613,
         n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621,
         n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629,
         n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637,
         n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645,
         n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653,
         n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661,
         n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669,
         n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677,
         n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685,
         n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693,
         n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701,
         n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709,
         n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717,
         n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725,
         n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733,
         n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741,
         n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749,
         n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757,
         n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765,
         n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773,
         n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781,
         n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789,
         n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797,
         n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805,
         n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813,
         n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821,
         n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829,
         n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837,
         n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845,
         n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853,
         n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861,
         n19862, n19863, n19864, n19865, n19866, n19867, n19869, n19870,
         n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878,
         n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886,
         n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894,
         n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902,
         n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910,
         n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918,
         n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926,
         n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934,
         n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942,
         n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950,
         n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958,
         n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966,
         n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974,
         n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982,
         n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990,
         n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998,
         n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006,
         n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014,
         n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022,
         n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030,
         n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038,
         n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046,
         n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054,
         n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062,
         n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070,
         n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078,
         n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086,
         n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094,
         n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102,
         n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110,
         n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118,
         n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126,
         n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134,
         n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142,
         n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150,
         n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158,
         n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166,
         n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174,
         n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182,
         n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190,
         n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198,
         n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206,
         n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214,
         n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222,
         n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230,
         n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238,
         n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246,
         n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254,
         n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262,
         n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270,
         n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278,
         n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286,
         n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294,
         n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302,
         n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310,
         n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318,
         n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326,
         n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334,
         n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342,
         n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350,
         n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358,
         n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366,
         n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374,
         n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382,
         n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390,
         n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398,
         n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406,
         n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414,
         n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422,
         n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430,
         n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438,
         n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446,
         n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454,
         n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462,
         n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470,
         n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478,
         n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486,
         n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494,
         n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502,
         n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510,
         n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518,
         n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526,
         n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534,
         n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542,
         n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550,
         n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558,
         n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566,
         n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574,
         n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582,
         n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590,
         n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598,
         n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606,
         n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614,
         n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622,
         n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630,
         n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638,
         n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646,
         n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654,
         n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662,
         n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670,
         n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678,
         n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686,
         n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694,
         n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702,
         n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710,
         n20711;

  NOR2_X1 U11046 ( .A1(n16277), .A2(n17191), .ZN(n16276) );
  OAI21_X1 U11047 ( .B1(n18216), .B2(n18215), .A(n16974), .ZN(n18384) );
  INV_X4 U11049 ( .A(n14368), .ZN(n15572) );
  OR2_X1 U11050 ( .A1(n13246), .A2(n15895), .ZN(n18933) );
  AND2_X1 U11051 ( .A1(n13262), .A2(n13225), .ZN(n19259) );
  BUF_X2 U11052 ( .A(n15226), .Z(n15219) );
  CLKBUF_X2 U11053 ( .A(n11573), .Z(n9604) );
  AND2_X2 U11054 ( .A1(n9625), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11629) );
  AND2_X2 U11055 ( .A1(n11654), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12032) );
  CLKBUF_X2 U11056 ( .A(n16624), .Z(n16733) );
  CLKBUF_X2 U11057 ( .A(n13606), .Z(n16668) );
  INV_X4 U11058 ( .A(n15218), .ZN(n16722) );
  CLKBUF_X2 U11059 ( .A(n10544), .Z(n10448) );
  CLKBUF_X2 U11060 ( .A(n10435), .Z(n11224) );
  CLKBUF_X2 U11061 ( .A(n10469), .Z(n11218) );
  INV_X1 U11062 ( .A(n12630), .ZN(n18926) );
  BUF_X1 U11063 ( .A(n15128), .Z(n9611) );
  INV_X1 U11064 ( .A(n18900), .ZN(n12549) );
  INV_X1 U11065 ( .A(n10396), .ZN(n12701) );
  AND4_X1 U11066 ( .A1(n10348), .A2(n10347), .A3(n10346), .A4(n10345), .ZN(
        n10364) );
  AND4_X1 U11067 ( .A1(n10352), .A2(n10351), .A3(n10350), .A4(n10349), .ZN(
        n10363) );
  AND4_X1 U11068 ( .A1(n10356), .A2(n10355), .A3(n10354), .A4(n10353), .ZN(
        n10362) );
  AND4_X1 U11069 ( .A1(n10386), .A2(n10385), .A3(n10384), .A4(n10383), .ZN(
        n10392) );
  AND2_X1 U11070 ( .A1(n10295), .A2(n12915), .ZN(n10470) );
  AND2_X1 U11071 ( .A1(n14427), .A2(n10297), .ZN(n10436) );
  AND2_X1 U11072 ( .A1(n10295), .A2(n10297), .ZN(n10435) );
  AND2_X1 U11073 ( .A1(n10290), .A2(n12915), .ZN(n10469) );
  AND2_X2 U11074 ( .A1(n12915), .A2(n14428), .ZN(n10570) );
  INV_X1 U11075 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11827) );
  BUF_X1 U11076 ( .A(n10403), .Z(n12500) );
  NOR2_X1 U11077 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11475) );
  CLKBUF_X3 U11078 ( .A(n10463), .Z(n11014) );
  BUF_X2 U11079 ( .A(n11470), .Z(n9606) );
  NAND2_X1 U11080 ( .A1(n13441), .A2(n13440), .ZN(n13860) );
  NAND2_X1 U11081 ( .A1(n18806), .A2(n18844), .ZN(n13363) );
  OR2_X1 U11082 ( .A1(n16465), .A2(n13573), .ZN(n15250) );
  INV_X1 U11083 ( .A(n12186), .ZN(n14826) );
  CLKBUF_X2 U11084 ( .A(n15269), .Z(n16716) );
  CLKBUF_X2 U11085 ( .A(n15128), .Z(n9612) );
  INV_X1 U11086 ( .A(n13715), .ZN(n13886) );
  NOR2_X1 U11087 ( .A1(n10535), .A2(n9844), .ZN(n10601) );
  INV_X1 U11088 ( .A(n12224), .ZN(n13327) );
  AND2_X1 U11089 ( .A1(n11395), .A2(n11394), .ZN(n11421) );
  NAND3_X1 U11090 ( .A1(n13642), .A2(n13641), .A3(n13640), .ZN(n15200) );
  NOR2_X1 U11091 ( .A1(n10093), .A2(n10092), .ZN(n16182) );
  NOR2_X1 U11092 ( .A1(n17101), .A2(n16209), .ZN(n16208) );
  OAI22_X1 U11093 ( .A1(n16256), .A2(n10076), .B1(n10073), .B2(n16247), .ZN(
        n16245) );
  NOR2_X1 U11094 ( .A1(n17152), .A2(n17153), .ZN(n17124) );
  INV_X1 U11095 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n17987) );
  AND2_X1 U11096 ( .A1(n13961), .A2(n12386), .ZN(n19644) );
  INV_X1 U11097 ( .A(n19798), .ZN(n19781) );
  AND2_X1 U11098 ( .A1(n10120), .A2(n15696), .ZN(n12264) );
  AND2_X1 U11099 ( .A1(n12769), .A2(n12768), .ZN(n12946) );
  CLKBUF_X2 U11100 ( .A(n12540), .Z(n18895) );
  NOR2_X2 U11101 ( .A1(n11997), .A2(n15853), .ZN(n11995) );
  INV_X1 U11102 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n15904) );
  NOR2_X2 U11103 ( .A1(n16141), .A2(n16200), .ZN(n16185) );
  INV_X2 U11104 ( .A(n17235), .ZN(n17318) );
  INV_X1 U11105 ( .A(n19644), .ZN(n19690) );
  INV_X2 U11106 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12617) );
  AOI21_X1 U11107 ( .B1(n16775), .B2(n16522), .A(n16535), .ZN(n16527) );
  OR3_X1 U11108 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18362), .A3(
        n13700), .ZN(n9602) );
  NAND2_X2 U11109 ( .A1(n10169), .A2(n9804), .ZN(n15060) );
  AND2_X1 U11110 ( .A1(n12921), .A2(n14428), .ZN(n10550) );
  NOR2_X2 U11111 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17253), .ZN(
        n17236) );
  NOR2_X2 U11112 ( .A1(n11982), .A2(n18456), .ZN(n11980) );
  INV_X1 U11113 ( .A(n9823), .ZN(n14368) );
  NAND4_X1 U11114 ( .A1(n18362), .A2(n18355), .A3(n18345), .A4(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15281) );
  NAND2_X2 U11115 ( .A1(n9777), .A2(n11081), .ZN(n11088) );
  AOI211_X2 U11116 ( .C1(n18875), .C2(n15702), .A(n14842), .B(n14841), .ZN(
        n14843) );
  NOR2_X2 U11117 ( .A1(n16604), .A2(n16631), .ZN(n16618) );
  MUX2_X2 U11118 ( .A(n13347), .B(n12216), .S(n11382), .Z(n12438) );
  AND2_X2 U11119 ( .A1(n13369), .A2(n12126), .ZN(n12625) );
  XNOR2_X2 U11120 ( .A(n11080), .B(n19831), .ZN(n12875) );
  AND2_X1 U11121 ( .A1(n9638), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11573) );
  NAND2_X2 U11122 ( .A1(n12888), .A2(n11072), .ZN(n11080) );
  BUF_X4 U11123 ( .A(n11470), .Z(n9605) );
  BUF_X4 U11124 ( .A(n11470), .Z(n9607) );
  INV_X1 U11125 ( .A(n9747), .ZN(n9608) );
  INV_X4 U11126 ( .A(n9608), .ZN(n9609) );
  XNOR2_X1 U11127 ( .A(n16133), .B(n15920), .ZN(n9747) );
  CLKBUF_X1 U11129 ( .A(n10545), .Z(n9610) );
  AND2_X1 U11130 ( .A1(n14428), .A2(n10297), .ZN(n10545) );
  CLKBUF_X1 U11131 ( .A(n10545), .Z(n11039) );
  XNOR2_X2 U11132 ( .A(n13359), .B(n13360), .ZN(n18806) );
  AND2_X4 U11133 ( .A1(n11475), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11804) );
  NOR2_X2 U11134 ( .A1(n20668), .A2(n15405), .ZN(n15927) );
  NAND2_X2 U11135 ( .A1(n11319), .A2(n9953), .ZN(n18919) );
  NAND2_X1 U11137 ( .A1(n14488), .A2(n11723), .ZN(n11745) );
  XNOR2_X1 U11138 ( .A(n11722), .B(n11718), .ZN(n14490) );
  AND2_X1 U11139 ( .A1(n10115), .A2(n9761), .ZN(n12001) );
  OR2_X1 U11140 ( .A1(n17093), .A2(n17435), .ZN(n10025) );
  NAND2_X1 U11141 ( .A1(n19783), .A2(n11096), .ZN(n15593) );
  NAND2_X1 U11142 ( .A1(n15356), .A2(n17144), .ZN(n17182) );
  XNOR2_X1 U11143 ( .A(n12658), .B(n12659), .ZN(n19540) );
  AND2_X1 U11144 ( .A1(n13802), .A2(n13779), .ZN(n13781) );
  NAND2_X1 U11145 ( .A1(n12740), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12888) );
  AND2_X1 U11146 ( .A1(n12734), .A2(n12733), .ZN(n12769) );
  NAND2_X1 U11147 ( .A1(n13235), .A2(n15895), .ZN(n19225) );
  OR2_X1 U11148 ( .A1(n13260), .A2(n13227), .ZN(n13246) );
  INV_X1 U11149 ( .A(n13187), .ZN(n15080) );
  CLKBUF_X2 U11150 ( .A(n18773), .Z(n18802) );
  AND2_X1 U11151 ( .A1(n9862), .A2(n12455), .ZN(n9861) );
  NOR2_X1 U11152 ( .A1(n11359), .A2(n11373), .ZN(n11370) );
  NAND2_X1 U11153 ( .A1(n11840), .A2(n11382), .ZN(n12626) );
  INV_X1 U11154 ( .A(n11382), .ZN(n12455) );
  INV_X2 U11155 ( .A(n16111), .ZN(n17736) );
  INV_X2 U11156 ( .A(n18895), .ZN(n9643) );
  INV_X1 U11157 ( .A(n11360), .ZN(n11832) );
  INV_X2 U11158 ( .A(n12003), .ZN(n9614) );
  NAND2_X1 U11159 ( .A1(n11990), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11987) );
  CLKBUF_X2 U11160 ( .A(n11360), .Z(n9634) );
  INV_X2 U11161 ( .A(n12581), .ZN(n9808) );
  INV_X1 U11162 ( .A(n12005), .ZN(n12540) );
  INV_X1 U11163 ( .A(n19858), .ZN(n9615) );
  CLKBUF_X2 U11164 ( .A(n15226), .Z(n16740) );
  CLKBUF_X2 U11165 ( .A(n16624), .Z(n16508) );
  CLKBUF_X2 U11166 ( .A(n10551), .Z(n10454) );
  AND2_X2 U11167 ( .A1(n11777), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11618) );
  BUF_X2 U11168 ( .A(n15097), .Z(n16738) );
  CLKBUF_X3 U11169 ( .A(n15140), .Z(n9621) );
  INV_X8 U11170 ( .A(n9679), .ZN(n9616) );
  AND2_X2 U11171 ( .A1(n11804), .A2(n9952), .ZN(n11533) );
  CLKBUF_X2 U11172 ( .A(n10575), .Z(n10453) );
  INV_X1 U11173 ( .A(n9635), .ZN(n9617) );
  AND2_X1 U11174 ( .A1(n12913), .A2(n10296), .ZN(n10552) );
  NOR2_X4 U11175 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10162) );
  NAND2_X1 U11176 ( .A1(n9687), .A2(n10145), .ZN(n14552) );
  NAND2_X1 U11177 ( .A1(n10253), .A2(n10252), .ZN(n10251) );
  AND2_X1 U11178 ( .A1(n9882), .A2(n9881), .ZN(n14996) );
  XNOR2_X1 U11179 ( .A(n10164), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14837) );
  OR2_X1 U11180 ( .A1(n13849), .A2(n14672), .ZN(n9935) );
  XNOR2_X1 U11181 ( .A(n14673), .B(n14675), .ZN(n14686) );
  AND2_X1 U11182 ( .A1(n9831), .A2(n9830), .ZN(n14673) );
  AND2_X1 U11183 ( .A1(n14720), .A2(n9812), .ZN(n14668) );
  OAI21_X1 U11184 ( .B1(n14772), .B2(n14739), .A(n9897), .ZN(n14752) );
  AOI21_X1 U11185 ( .B1(n14782), .B2(n14783), .A(n14737), .ZN(n14772) );
  NAND2_X1 U11186 ( .A1(n14716), .A2(n14721), .ZN(n10238) );
  NAND2_X1 U11187 ( .A1(n13831), .A2(n14714), .ZN(n10237) );
  OAI21_X1 U11188 ( .B1(n14917), .B2(n9939), .A(n9937), .ZN(n9936) );
  NAND2_X1 U11189 ( .A1(n14490), .A2(n14489), .ZN(n14488) );
  AOI21_X1 U11190 ( .B1(n9908), .B2(n9694), .A(n9900), .ZN(n14791) );
  OAI21_X1 U11191 ( .B1(n13864), .B2(n10170), .A(n13868), .ZN(n10166) );
  NOR2_X1 U11192 ( .A1(n9706), .A2(n9660), .ZN(n9969) );
  NAND2_X1 U11193 ( .A1(n14815), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9803) );
  NOR2_X1 U11194 ( .A1(n14652), .A2(n14651), .ZN(n10165) );
  OR2_X1 U11195 ( .A1(n11722), .A2(n11721), .ZN(n11723) );
  AOI21_X1 U11196 ( .B1(n9873), .B2(n9872), .A(n13821), .ZN(n14917) );
  NAND2_X1 U11197 ( .A1(n9834), .A2(n10243), .ZN(n9873) );
  OR2_X1 U11198 ( .A1(n14170), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14163) );
  NAND2_X1 U11199 ( .A1(n13755), .A2(n13754), .ZN(n15054) );
  NAND2_X1 U11200 ( .A1(n10225), .A2(n10223), .ZN(n13755) );
  NAND2_X1 U11201 ( .A1(n14508), .A2(n14507), .ZN(n14506) );
  XNOR2_X1 U11202 ( .A(n14514), .B(n11679), .ZN(n14508) );
  NOR2_X1 U11203 ( .A1(n18630), .A2(n15725), .ZN(n15716) );
  NAND2_X1 U11204 ( .A1(n9859), .A2(n9858), .ZN(n14514) );
  XNOR2_X1 U11205 ( .A(n14648), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10221) );
  NAND2_X1 U11206 ( .A1(n13481), .A2(n13480), .ZN(n13742) );
  AOI211_X1 U11207 ( .C1(n18875), .C2(n14553), .A(n14654), .B(n13880), .ZN(
        n13881) );
  AND2_X1 U11208 ( .A1(n9885), .A2(n13362), .ZN(n9964) );
  AND2_X1 U11209 ( .A1(n14830), .A2(n12203), .ZN(n14553) );
  NAND2_X1 U11210 ( .A1(n10265), .A2(n10268), .ZN(n15583) );
  AND2_X2 U11211 ( .A1(n13398), .A2(n13397), .ZN(n13501) );
  AND2_X1 U11212 ( .A1(n10650), .A2(n9668), .ZN(n13398) );
  OR2_X1 U11213 ( .A1(n13860), .A2(n13859), .ZN(n13865) );
  NAND2_X1 U11214 ( .A1(n9894), .A2(n18617), .ZN(n13479) );
  NAND2_X1 U11215 ( .A1(n11562), .A2(n10283), .ZN(n13195) );
  AND2_X1 U11216 ( .A1(n14893), .A2(n13878), .ZN(n14871) );
  NOR2_X1 U11217 ( .A1(n9928), .A2(n9875), .ZN(n9872) );
  XNOR2_X1 U11218 ( .A(n13439), .B(n13440), .ZN(n13364) );
  AND2_X1 U11219 ( .A1(n10263), .A2(n15580), .ZN(n9869) );
  NAND2_X1 U11220 ( .A1(n13330), .A2(n9811), .ZN(n13357) );
  AND2_X1 U11221 ( .A1(n11133), .A2(n9666), .ZN(n10263) );
  AND3_X1 U11222 ( .A1(n9847), .A2(n12990), .A3(n9846), .ZN(n13044) );
  NAND2_X1 U11223 ( .A1(n14644), .A2(n13738), .ZN(n13839) );
  AND2_X1 U11224 ( .A1(n10597), .A2(n12989), .ZN(n9847) );
  NAND2_X1 U11225 ( .A1(n11126), .A2(n11125), .ZN(n9823) );
  AOI21_X1 U11226 ( .B1(n10514), .B2(n10513), .A(n10512), .ZN(n12873) );
  OR2_X1 U11227 ( .A1(n18884), .A2(n13316), .ZN(n13317) );
  OR2_X1 U11228 ( .A1(n18962), .A2(n13460), .ZN(n13461) );
  CLKBUF_X1 U11229 ( .A(n11268), .Z(n14071) );
  AND2_X1 U11230 ( .A1(n9898), .A2(n15080), .ZN(n18887) );
  AND2_X1 U11231 ( .A1(n9898), .A2(n13263), .ZN(n13459) );
  OR2_X1 U11232 ( .A1(n19225), .A2(n13270), .ZN(n13271) );
  AND2_X1 U11233 ( .A1(n13262), .A2(n13223), .ZN(n19340) );
  NOR2_X2 U11234 ( .A1(n13264), .A2(n13263), .ZN(n19136) );
  XNOR2_X1 U11235 ( .A(n11462), .B(n11463), .ZN(n12659) );
  XNOR2_X1 U11236 ( .A(n11070), .B(n12680), .ZN(n12740) );
  CLKBUF_X1 U11237 ( .A(n12938), .Z(n9631) );
  AND2_X1 U11238 ( .A1(n13790), .A2(n10065), .ZN(n13802) );
  NAND2_X1 U11239 ( .A1(n13262), .A2(n13261), .ZN(n13264) );
  INV_X2 U11240 ( .A(n12957), .ZN(n19774) );
  NOR2_X1 U11241 ( .A1(n13257), .A2(n13222), .ZN(n13442) );
  NAND2_X1 U11242 ( .A1(n11461), .A2(n11460), .ZN(n11462) );
  NAND2_X1 U11243 ( .A1(n18864), .A2(n18870), .ZN(n14943) );
  NAND2_X1 U11244 ( .A1(n10507), .A2(n10506), .ZN(n10535) );
  OR2_X1 U11245 ( .A1(n12593), .A2(n12834), .ZN(n18864) );
  NAND2_X1 U11246 ( .A1(n11437), .A2(n11436), .ZN(n11438) );
  OR2_X1 U11247 ( .A1(n12593), .A2(n12592), .ZN(n18870) );
  OR2_X1 U11248 ( .A1(n13226), .A2(n14440), .ZN(n13257) );
  AND2_X1 U11249 ( .A1(n13226), .A2(n13221), .ZN(n13262) );
  NAND2_X1 U11250 ( .A1(n19710), .A2(n19886), .ZN(n14024) );
  NAND2_X1 U11251 ( .A1(n10515), .A2(n11062), .ZN(n10507) );
  AND2_X1 U11252 ( .A1(n11885), .A2(n12669), .ZN(n9652) );
  NAND2_X1 U11253 ( .A1(n9815), .A2(n10562), .ZN(n19837) );
  XNOR2_X1 U11254 ( .A(n9782), .B(n9813), .ZN(n9844) );
  NAND2_X1 U11255 ( .A1(n9955), .A2(n9731), .ZN(n11416) );
  AOI21_X1 U11256 ( .B1(n14440), .B2(n12461), .A(n11401), .ZN(n12664) );
  OAI21_X1 U11257 ( .B1(n11999), .B2(n18486), .A(n18485), .ZN(n18474) );
  XNOR2_X1 U11258 ( .A(n13231), .B(n11421), .ZN(n13187) );
  OR2_X1 U11259 ( .A1(n10505), .A2(n10504), .ZN(n10506) );
  XNOR2_X1 U11260 ( .A(n10505), .B(n10503), .ZN(n10515) );
  NAND2_X1 U11261 ( .A1(n10524), .A2(n9864), .ZN(n19922) );
  NAND2_X1 U11262 ( .A1(n11421), .A2(n11420), .ZN(n11424) );
  INV_X2 U11263 ( .A(n15696), .ZN(n18630) );
  NAND2_X1 U11264 ( .A1(n9916), .A2(n10429), .ZN(n12636) );
  NAND2_X1 U11265 ( .A1(n9887), .A2(n9886), .ZN(n10505) );
  NAND2_X1 U11266 ( .A1(n9888), .A2(n9697), .ZN(n9864) );
  AND2_X1 U11267 ( .A1(n11447), .A2(n11446), .ZN(n11452) );
  AND2_X1 U11268 ( .A1(n10074), .A2(n10073), .ZN(n16277) );
  OAI21_X1 U11269 ( .B1(n10526), .B2(n10477), .A(n9889), .ZN(n10524) );
  AND2_X1 U11270 ( .A1(n11409), .A2(n11408), .ZN(n11419) );
  CLKBUF_X1 U11271 ( .A(n10526), .Z(n19961) );
  AND2_X1 U11272 ( .A1(n9912), .A2(n10445), .ZN(n10497) );
  NOR2_X1 U11273 ( .A1(n12071), .A2(n12070), .ZN(n12085) );
  AND2_X1 U11274 ( .A1(n12530), .A2(n11853), .ZN(n12839) );
  NAND2_X1 U11275 ( .A1(n9911), .A2(n12578), .ZN(n11389) );
  AND2_X1 U11276 ( .A1(n12866), .A2(n12069), .ZN(n12070) );
  INV_X2 U11277 ( .A(n16977), .ZN(n17037) );
  NAND2_X2 U11278 ( .A1(n16974), .A2(n18234), .ZN(n17040) );
  AND2_X1 U11279 ( .A1(n12564), .A2(n12565), .ZN(n12563) );
  NAND3_X1 U11280 ( .A1(n9949), .A2(n12846), .A3(n9948), .ZN(n10037) );
  NAND2_X1 U11281 ( .A1(n9945), .A2(n9944), .ZN(n9949) );
  AND2_X1 U11282 ( .A1(n12859), .A2(n11379), .ZN(n11888) );
  AOI21_X1 U11283 ( .B1(n10478), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n9890), 
        .ZN(n9889) );
  AND2_X1 U11284 ( .A1(n11406), .A2(n9942), .ZN(n9948) );
  CLKBUF_X1 U11285 ( .A(n12443), .Z(n12848) );
  OR2_X1 U11286 ( .A1(n15917), .A2(n15193), .ZN(n15095) );
  INV_X2 U11287 ( .A(n14452), .ZN(n11957) );
  AND2_X1 U11288 ( .A1(n9947), .A2(n9946), .ZN(n9945) );
  AND2_X1 U11289 ( .A1(n11339), .A2(n11375), .ZN(n12859) );
  AND2_X1 U11290 ( .A1(n9820), .A2(n12715), .ZN(n9817) );
  NAND2_X1 U11291 ( .A1(n11370), .A2(n9634), .ZN(n12846) );
  AND3_X1 U11292 ( .A1(n11362), .A2(n12626), .A3(n9644), .ZN(n9944) );
  OR2_X1 U11293 ( .A1(n12045), .A2(n9808), .ZN(n9947) );
  AND2_X1 U11294 ( .A1(n9696), .A2(n9644), .ZN(n12576) );
  AND2_X1 U11295 ( .A1(n11338), .A2(n18900), .ZN(n11339) );
  NAND2_X1 U11296 ( .A1(n12706), .A2(n10401), .ZN(n12510) );
  NOR2_X1 U11297 ( .A1(n18907), .A2(n18926), .ZN(n11362) );
  OR2_X1 U11298 ( .A1(n12899), .A2(n10400), .ZN(n14422) );
  INV_X1 U11299 ( .A(n20541), .ZN(n11129) );
  NAND2_X1 U11300 ( .A1(n18919), .A2(n12003), .ZN(n12536) );
  AND2_X1 U11301 ( .A1(n9808), .A2(n18900), .ZN(n9644) );
  NAND2_X1 U11302 ( .A1(n9692), .A2(n11210), .ZN(n12706) );
  AND2_X1 U11303 ( .A1(n9615), .A2(n19863), .ZN(n11063) );
  NOR2_X2 U11304 ( .A1(n13652), .A2(n13651), .ZN(n17741) );
  NOR2_X2 U11305 ( .A1(n13612), .A2(n13611), .ZN(n17778) );
  AND2_X1 U11306 ( .A1(n19839), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11161) );
  OR2_X1 U11307 ( .A1(n10460), .A2(n10459), .ZN(n11128) );
  NAND2_X2 U11308 ( .A1(n9829), .A2(n9828), .ZN(n12630) );
  NOR2_X1 U11309 ( .A1(n19886), .A2(n20448), .ZN(n10508) );
  NAND2_X1 U11310 ( .A1(n11331), .A2(n9952), .ZN(n9807) );
  NAND2_X1 U11311 ( .A1(n9951), .A2(n9950), .ZN(n12003) );
  NAND2_X1 U11312 ( .A1(n11318), .A2(n9952), .ZN(n9953) );
  NAND2_X1 U11313 ( .A1(n11313), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11319) );
  OR2_X2 U11314 ( .A1(n10303), .A2(n10302), .ZN(n19858) );
  OR2_X2 U11315 ( .A1(n16045), .A2(n15991), .ZN(n16047) );
  INV_X2 U11316 ( .A(U212), .ZN(n16032) );
  NAND2_X1 U11317 ( .A1(n9810), .A2(n9809), .ZN(n12581) );
  INV_X2 U11318 ( .A(n12541), .ZN(n18907) );
  AND4_X1 U11319 ( .A1(n11330), .A2(n11329), .A3(n11328), .A4(n11327), .ZN(
        n11331) );
  AND4_X1 U11320 ( .A1(n11312), .A2(n11311), .A3(n11310), .A4(n11309), .ZN(
        n11313) );
  AND4_X1 U11321 ( .A1(n10378), .A2(n10377), .A3(n10376), .A4(n10375), .ZN(
        n10394) );
  OR2_X2 U11322 ( .A1(n10323), .A2(n10322), .ZN(n19878) );
  INV_X1 U11323 ( .A(n17244), .ZN(n17260) );
  MUX2_X1 U11324 ( .A(n11285), .B(n11284), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n12541) );
  INV_X1 U11325 ( .A(n16435), .ZN(n16610) );
  INV_X2 U11326 ( .A(n10462), .ZN(n9618) );
  INV_X2 U11327 ( .A(n11496), .ZN(n9639) );
  AND4_X1 U11328 ( .A1(n10360), .A2(n10359), .A3(n10358), .A4(n10357), .ZN(
        n10361) );
  AND2_X1 U11329 ( .A1(n11334), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11335) );
  NAND2_X2 U11330 ( .A1(n18270), .A2(n18380), .ZN(n18318) );
  INV_X2 U11331 ( .A(n9636), .ZN(n9638) );
  NAND2_X2 U11332 ( .A1(n18380), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18328) );
  INV_X1 U11334 ( .A(n9602), .ZN(n9640) );
  CLKBUF_X2 U11335 ( .A(n10334), .Z(n11037) );
  BUF_X2 U11336 ( .A(n10461), .Z(n11036) );
  BUF_X2 U11337 ( .A(n10461), .Z(n10903) );
  INV_X1 U11338 ( .A(n11298), .ZN(n9636) );
  INV_X2 U11339 ( .A(n16079), .ZN(U215) );
  NAND2_X2 U11340 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19509), .ZN(n19508) );
  NAND2_X2 U11341 ( .A1(n19509), .A2(n20627), .ZN(n19511) );
  INV_X2 U11342 ( .A(n9771), .ZN(n18251) );
  BUF_X2 U11343 ( .A(n10470), .Z(n10447) );
  BUF_X2 U11344 ( .A(n10971), .Z(n11038) );
  INV_X1 U11345 ( .A(n9680), .ZN(n16623) );
  BUF_X2 U11346 ( .A(n10464), .Z(n11226) );
  BUF_X4 U11347 ( .A(n15269), .Z(n9620) );
  INV_X2 U11348 ( .A(n16083), .ZN(n16085) );
  INV_X2 U11349 ( .A(n18401), .ZN(n18380) );
  INV_X2 U11350 ( .A(n15250), .ZN(n9622) );
  AND2_X1 U11351 ( .A1(n12796), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9623) );
  AND2_X2 U11352 ( .A1(n12795), .A2(n11827), .ZN(n9626) );
  AND2_X2 U11353 ( .A1(n12796), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11777) );
  INV_X2 U11354 ( .A(n11286), .ZN(n9627) );
  AND2_X2 U11355 ( .A1(n12796), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9624) );
  AND2_X1 U11356 ( .A1(n12921), .A2(n14427), .ZN(n10334) );
  BUF_X2 U11357 ( .A(n10463), .Z(n11044) );
  NAND2_X1 U11358 ( .A1(n11804), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11496) );
  NOR2_X1 U11359 ( .A1(n18348), .A2(n18255), .ZN(n18386) );
  BUF_X2 U11360 ( .A(n10552), .Z(n11225) );
  NAND2_X1 U11361 ( .A1(n18355), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13573) );
  NAND2_X1 U11362 ( .A1(n18369), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13574) );
  AND2_X1 U11363 ( .A1(n12617), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10290) );
  NAND2_X1 U11364 ( .A1(n18345), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13572) );
  AND2_X1 U11365 ( .A1(n9913), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12921) );
  AND2_X1 U11366 ( .A1(n11275), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12795) );
  AND2_X1 U11367 ( .A1(n9941), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12796) );
  AND2_X2 U11368 ( .A1(n10162), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11470) );
  AND2_X2 U11369 ( .A1(n12774), .A2(n11827), .ZN(n11654) );
  NAND2_X1 U11370 ( .A1(n12448), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12776) );
  NAND3_X1 U11371 ( .A1(n13713), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11286) );
  INV_X2 U11372 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18369) );
  INV_X2 U11373 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18362) );
  AND2_X1 U11374 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12774) );
  INV_X2 U11375 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18345) );
  AND2_X1 U11376 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12448) );
  INV_X2 U11377 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18355) );
  NAND2_X2 U11378 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18205) );
  NOR2_X1 U11379 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10296) );
  NAND2_X1 U11380 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13700) );
  AND2_X1 U11381 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12913) );
  AND2_X2 U11382 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14427) );
  NOR2_X2 U11383 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12915) );
  AND2_X1 U11384 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10297) );
  INV_X1 U11385 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9952) );
  NOR2_X2 U11386 ( .A1(n16480), .A2(n16772), .ZN(n16777) );
  NAND3_X1 U11387 ( .A1(n15420), .A2(n18391), .A3(n17736), .ZN(n16772) );
  OR2_X2 U11388 ( .A1(n13990), .A2(n13980), .ZN(n13982) );
  NAND2_X1 U11389 ( .A1(n18362), .A2(n18369), .ZN(n16465) );
  OAI21_X2 U11390 ( .B1(n13297), .B2(n13296), .A(n13295), .ZN(n13298) );
  NOR2_X2 U11391 ( .A1(n10399), .A2(n10396), .ZN(n10413) );
  NOR2_X2 U11392 ( .A1(n14642), .A2(n14661), .ZN(n10222) );
  INV_X1 U11393 ( .A(n9845), .ZN(n11062) );
  NOR2_X2 U11394 ( .A1(n13050), .A2(n13049), .ZN(n13119) );
  INV_X2 U11395 ( .A(n13682), .ZN(n18216) );
  AOI211_X2 U11396 ( .C1(n18830), .C2(n18459), .A(n14768), .B(n14767), .ZN(
        n14769) );
  NAND2_X1 U11397 ( .A1(n19960), .A2(n10497), .ZN(n10500) );
  NOR2_X1 U11398 ( .A1(n13572), .A2(n13574), .ZN(n15140) );
  NOR2_X2 U11399 ( .A1(n14011), .A2(n14012), .ZN(n13999) );
  OAI22_X2 U11400 ( .A1(n15904), .A2(n11967), .B1(n14650), .B2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n13164) );
  XNOR2_X2 U11401 ( .A(n11966), .B(n11965), .ZN(n14650) );
  NOR2_X2 U11402 ( .A1(n16759), .A2(n16763), .ZN(n16762) );
  AND2_X1 U11403 ( .A1(n12795), .A2(n11827), .ZN(n9625) );
  AND2_X2 U11404 ( .A1(n12795), .A2(n11827), .ZN(n11681) );
  INV_X1 U11405 ( .A(n11815), .ZN(n9628) );
  INV_X2 U11406 ( .A(n11286), .ZN(n11815) );
  BUF_X8 U11407 ( .A(n16663), .Z(n9629) );
  INV_X2 U11408 ( .A(n15151), .ZN(n16663) );
  INV_X2 U11409 ( .A(n9680), .ZN(n9630) );
  OR2_X1 U11410 ( .A1(n13571), .A2(n13573), .ZN(n9680) );
  NOR2_X2 U11411 ( .A1(n13622), .A2(n13621), .ZN(n17766) );
  INV_X1 U11412 ( .A(n9622), .ZN(n9633) );
  INV_X4 U11413 ( .A(n15250), .ZN(n15241) );
  NAND2_X1 U11414 ( .A1(n9856), .A2(n9855), .ZN(n11360) );
  INV_X1 U11415 ( .A(n12776), .ZN(n9635) );
  INV_X1 U11416 ( .A(n9636), .ZN(n9637) );
  AND2_X2 U11417 ( .A1(n9606), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12034) );
  NOR3_X2 U11418 ( .A1(n15096), .A2(n16756), .A3(n16753), .ZN(n16752) );
  NOR2_X4 U11419 ( .A1(n11981), .A2(n14742), .ZN(n11978) );
  NOR2_X1 U11420 ( .A1(n13575), .A2(n18205), .ZN(n15097) );
  INV_X1 U11421 ( .A(n9602), .ZN(n9641) );
  INV_X1 U11422 ( .A(n9602), .ZN(n9642) );
  BUF_X4 U11423 ( .A(n13164), .Z(n15696) );
  MUX2_X2 U11424 ( .A(n11358), .B(n11357), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n12005) );
  NOR2_X4 U11425 ( .A1(n11976), .A2(n14710), .ZN(n11974) );
  OR2_X2 U11426 ( .A1(n11214), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n19798) );
  NOR2_X1 U11427 ( .A1(n19994), .A2(n10599), .ZN(n10600) );
  AOI21_X1 U11428 ( .B1(n10243), .B2(n10242), .A(n9737), .ZN(n10241) );
  INV_X1 U11429 ( .A(n9686), .ZN(n10242) );
  INV_X1 U11430 ( .A(n17126), .ZN(n10105) );
  AND2_X1 U11431 ( .A1(n13469), .A2(n13468), .ZN(n13472) );
  OR2_X1 U11432 ( .A1(n13466), .A2(n13465), .ZN(n13469) );
  NAND2_X1 U11433 ( .A1(n9709), .A2(n10600), .ZN(n11126) );
  INV_X1 U11434 ( .A(n10443), .ZN(n11082) );
  AOI21_X1 U11435 ( .B1(n9889), .B2(n10477), .A(n11124), .ZN(n9886) );
  INV_X1 U11436 ( .A(n11187), .ZN(n11194) );
  NAND2_X1 U11437 ( .A1(n12701), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10543) );
  AND3_X1 U11438 ( .A1(n12003), .A2(n18907), .A3(n12631), .ZN(n9862) );
  AND2_X1 U11439 ( .A1(n15845), .A2(n10233), .ZN(n10232) );
  NAND2_X1 U11440 ( .A1(n13332), .A2(n10234), .ZN(n10233) );
  AND2_X1 U11441 ( .A1(n12224), .A2(n15903), .ZN(n10234) );
  NAND2_X1 U11442 ( .A1(n9711), .A2(n9808), .ZN(n9946) );
  NAND2_X1 U11443 ( .A1(n10600), .A2(n10601), .ZN(n10618) );
  AND2_X1 U11444 ( .A1(n11010), .A2(n10207), .ZN(n10206) );
  INV_X1 U11445 ( .A(n13917), .ZN(n10207) );
  AND2_X1 U11446 ( .A1(n14052), .A2(n14000), .ZN(n10202) );
  NAND2_X1 U11447 ( .A1(n12612), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11239) );
  NAND2_X1 U11448 ( .A1(n15583), .A2(n15581), .ZN(n9870) );
  INV_X1 U11449 ( .A(n10508), .ZN(n10999) );
  NAND2_X1 U11450 ( .A1(n14367), .A2(n9705), .ZN(n9914) );
  INV_X1 U11451 ( .A(n9994), .ZN(n9993) );
  OAI21_X1 U11452 ( .B1(n15572), .B2(n11140), .A(n9996), .ZN(n9994) );
  NAND2_X1 U11453 ( .A1(n9915), .A2(n9891), .ZN(n9868) );
  NOR2_X1 U11454 ( .A1(n14366), .A2(n9995), .ZN(n9891) );
  AND2_X1 U11455 ( .A1(n15572), .A2(n9996), .ZN(n9995) );
  NAND2_X1 U11456 ( .A1(n11161), .A2(n10396), .ZN(n11187) );
  NAND2_X1 U11457 ( .A1(n11158), .A2(n11157), .ZN(n11253) );
  NAND2_X1 U11458 ( .A1(n10541), .A2(n10540), .ZN(n19995) );
  AOI21_X1 U11459 ( .B1(n10406), .B2(n10195), .A(n10407), .ZN(n9781) );
  NAND2_X1 U11460 ( .A1(n10408), .A2(n10195), .ZN(n10194) );
  AND3_X2 U11461 ( .A1(n9816), .A2(n19839), .A3(n11063), .ZN(n12423) );
  AOI21_X1 U11462 ( .B1(n14467), .B2(n9760), .A(n10150), .ZN(n10148) );
  NAND2_X1 U11463 ( .A1(n9936), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13831) );
  INV_X1 U11464 ( .A(n10246), .ZN(n10244) );
  NOR2_X1 U11465 ( .A1(n10224), .A2(n9735), .ZN(n10223) );
  INV_X1 U11466 ( .A(n13744), .ZN(n10224) );
  AND4_X1 U11467 ( .A1(n12134), .A2(n12133), .A3(n12132), .A4(n12131), .ZN(
        n12152) );
  NAND2_X1 U11468 ( .A1(n11398), .A2(n19535), .ZN(n11459) );
  INV_X1 U11469 ( .A(n12536), .ZN(n11338) );
  NOR2_X1 U11470 ( .A1(n16465), .A2(n13575), .ZN(n13606) );
  NOR2_X1 U11471 ( .A1(n16910), .A2(n15293), .ZN(n15292) );
  NAND2_X1 U11472 ( .A1(n18176), .A2(n9787), .ZN(n13682) );
  INV_X1 U11473 ( .A(n15194), .ZN(n9787) );
  AND2_X1 U11474 ( .A1(n12691), .A2(n12705), .ZN(n12650) );
  AND2_X1 U11475 ( .A1(n20448), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11243) );
  AND2_X1 U11476 ( .A1(n11060), .A2(n10206), .ZN(n10205) );
  NAND2_X1 U11477 ( .A1(n9847), .A2(n12990), .ZN(n13006) );
  NAND2_X1 U11478 ( .A1(n12699), .A2(n12698), .ZN(n12717) );
  AND2_X1 U11479 ( .A1(n9670), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10134) );
  NAND2_X1 U11480 ( .A1(n11308), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9829) );
  NAND2_X1 U11481 ( .A1(n11307), .A2(n9952), .ZN(n9828) );
  NAND2_X1 U11482 ( .A1(n14809), .A2(n9907), .ZN(n9906) );
  INV_X1 U11483 ( .A(n14808), .ZN(n9907) );
  AND2_X1 U11484 ( .A1(n15904), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12461) );
  AND2_X1 U11485 ( .A1(n10171), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9812) );
  OAI21_X1 U11486 ( .B1(n9902), .B2(n9901), .A(n14801), .ZN(n9900) );
  INV_X1 U11487 ( .A(n14800), .ZN(n9901) );
  NOR2_X1 U11488 ( .A1(n10079), .A2(n10104), .ZN(n10103) );
  INV_X1 U11489 ( .A(n16902), .ZN(n15979) );
  INV_X1 U11490 ( .A(n19687), .ZN(n19662) );
  AND2_X1 U11491 ( .A1(n12906), .A2(n9863), .ZN(n11551) );
  NAND2_X1 U11492 ( .A1(n11830), .A2(n11829), .ZN(n11845) );
  AND2_X1 U11493 ( .A1(n11845), .A2(n11844), .ZN(n11847) );
  NOR2_X1 U11494 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n10532) );
  INV_X1 U11495 ( .A(n10409), .ZN(n10276) );
  OR2_X1 U11496 ( .A1(n10492), .A2(n10491), .ZN(n11073) );
  AOI21_X1 U11497 ( .B1(n11186), .B2(n11185), .A(n11155), .ZN(n11191) );
  NAND2_X1 U11498 ( .A1(n12899), .A2(n19863), .ZN(n10412) );
  NAND2_X1 U11499 ( .A1(n9710), .A2(n12701), .ZN(n10272) );
  NAND2_X2 U11500 ( .A1(n11247), .A2(n9817), .ZN(n10408) );
  NAND2_X1 U11501 ( .A1(n9992), .A2(n9662), .ZN(n9989) );
  NAND3_X1 U11502 ( .A1(n10405), .A2(n10404), .A3(n10410), .ZN(n10406) );
  AND2_X1 U11503 ( .A1(n11255), .A2(n10525), .ZN(n9816) );
  INV_X1 U11504 ( .A(n14498), .ZN(n10141) );
  INV_X1 U11505 ( .A(n14915), .ZN(n9940) );
  OR2_X1 U11506 ( .A1(n13322), .A2(n13321), .ZN(n13326) );
  AND2_X1 U11507 ( .A1(n13269), .A2(n9738), .ZN(n9827) );
  AOI21_X1 U11508 ( .B1(n11933), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n11451), .ZN(n11453) );
  AND2_X1 U11509 ( .A1(n11378), .A2(n12588), .ZN(n9911) );
  INV_X1 U11510 ( .A(n11419), .ZN(n11422) );
  AOI21_X1 U11511 ( .B1(n14452), .B2(P2_EBX_REG_2__SCAN_IN), .A(n9736), .ZN(
        n9917) );
  AOI21_X1 U11512 ( .B1(n12827), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11847), .ZN(n11843) );
  INV_X1 U11513 ( .A(n16923), .ZN(n15321) );
  INV_X1 U11514 ( .A(n17754), .ZN(n13663) );
  NAND2_X1 U11515 ( .A1(n9983), .A2(n14002), .ZN(n9982) );
  INV_X1 U11516 ( .A(n13964), .ZN(n9983) );
  AND2_X1 U11517 ( .A1(n9853), .A2(n13979), .ZN(n9852) );
  INV_X1 U11518 ( .A(n13931), .ZN(n9853) );
  INV_X1 U11519 ( .A(n13147), .ZN(n9849) );
  XNOR2_X1 U11520 ( .A(n11126), .B(n10644), .ZN(n11114) );
  INV_X1 U11521 ( .A(n13092), .ZN(n10649) );
  NAND2_X1 U11522 ( .A1(n9675), .A2(n12376), .ZN(n9976) );
  INV_X1 U11523 ( .A(n13933), .ZN(n9977) );
  NAND2_X1 U11524 ( .A1(n14153), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11145) );
  NAND2_X1 U11525 ( .A1(n9712), .A2(n9822), .ZN(n14182) );
  INV_X1 U11526 ( .A(n14207), .ZN(n9822) );
  AOI21_X1 U11527 ( .B1(n10263), .B2(n10262), .A(n9657), .ZN(n10261) );
  NOR2_X1 U11528 ( .A1(n13182), .A2(n9988), .ZN(n9987) );
  INV_X1 U11529 ( .A(n13148), .ZN(n9988) );
  NOR2_X1 U11530 ( .A1(n10270), .A2(n10267), .ZN(n10266) );
  INV_X1 U11531 ( .A(n11113), .ZN(n10270) );
  INV_X1 U11532 ( .A(n15592), .ZN(n10267) );
  INV_X1 U11533 ( .A(n11106), .ZN(n10269) );
  NAND2_X1 U11534 ( .A1(n13715), .A2(n12352), .ZN(n12365) );
  OR2_X1 U11535 ( .A1(n10476), .A2(n10475), .ZN(n11074) );
  INV_X1 U11536 ( .A(n10444), .ZN(n9813) );
  NAND2_X1 U11537 ( .A1(n9814), .A2(n9732), .ZN(n9782) );
  NAND2_X1 U11538 ( .A1(n10396), .A2(n19886), .ZN(n10400) );
  NAND2_X1 U11539 ( .A1(n20517), .A2(n20446), .ZN(n9815) );
  AND2_X1 U11540 ( .A1(n10069), .A2(n10068), .ZN(n10067) );
  INV_X1 U11541 ( .A(n13785), .ZN(n10068) );
  AND2_X1 U11542 ( .A1(n13788), .A2(n13783), .ZN(n10069) );
  AND2_X1 U11543 ( .A1(n13798), .A2(n13796), .ZN(n13790) );
  NOR2_X1 U11544 ( .A1(n13793), .A2(n13792), .ZN(n13798) );
  NOR2_X1 U11545 ( .A1(n13475), .A2(n13473), .ZN(n13750) );
  NAND2_X1 U11546 ( .A1(n13329), .A2(n13328), .ZN(n13475) );
  OR2_X1 U11547 ( .A1(n12064), .A2(n12063), .ZN(n13293) );
  NOR2_X1 U11548 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11656) );
  OR2_X1 U11549 ( .A1(n10160), .A2(n13420), .ZN(n10159) );
  NAND2_X1 U11550 ( .A1(n10161), .A2(n13385), .ZN(n10160) );
  INV_X1 U11551 ( .A(n13196), .ZN(n10161) );
  AND2_X1 U11552 ( .A1(n12017), .A2(n12634), .ZN(n10189) );
  AND2_X1 U11553 ( .A1(n10189), .A2(n12738), .ZN(n10188) );
  NAND2_X1 U11554 ( .A1(n11832), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11852) );
  OR2_X1 U11555 ( .A1(n10125), .A2(n20697), .ZN(n10124) );
  AND2_X1 U11556 ( .A1(n13120), .A2(n10053), .ZN(n10052) );
  INV_X1 U11557 ( .A(n13175), .ZN(n10053) );
  NAND2_X1 U11558 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10125) );
  NOR2_X1 U11559 ( .A1(n14818), .A2(n10129), .ZN(n10133) );
  INV_X1 U11560 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10129) );
  NAND2_X1 U11561 ( .A1(n10133), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10132) );
  NAND2_X1 U11562 ( .A1(n14483), .A2(n10042), .ZN(n10041) );
  NOR2_X1 U11563 ( .A1(n10043), .A2(n14492), .ZN(n10042) );
  INV_X1 U11564 ( .A(n14596), .ZN(n10186) );
  AOI21_X1 U11565 ( .B1(n10170), .B2(n13868), .A(n10168), .ZN(n10167) );
  INV_X1 U11566 ( .A(n14905), .ZN(n10168) );
  NAND2_X1 U11567 ( .A1(n10169), .A2(n9803), .ZN(n9968) );
  AND2_X1 U11568 ( .A1(n10052), .A2(n10051), .ZN(n10050) );
  INV_X1 U11569 ( .A(n13206), .ZN(n10051) );
  INV_X1 U11570 ( .A(n15056), .ZN(n10249) );
  NAND2_X1 U11571 ( .A1(n9871), .A2(n13858), .ZN(n13863) );
  NAND2_X1 U11572 ( .A1(n13471), .A2(n13438), .ZN(n13857) );
  INV_X1 U11573 ( .A(n13363), .ZN(n9806) );
  NOR2_X1 U11574 ( .A1(n13470), .A2(n9966), .ZN(n9965) );
  INV_X1 U11575 ( .A(n9964), .ZN(n9963) );
  NOR2_X1 U11576 ( .A1(n12087), .A2(n10178), .ZN(n10180) );
  NAND2_X1 U11577 ( .A1(n13017), .A2(n12031), .ZN(n10178) );
  AOI21_X1 U11578 ( .B1(n10232), .B2(n9733), .A(n10229), .ZN(n10228) );
  NOR2_X1 U11579 ( .A1(n13332), .A2(n10230), .ZN(n10229) );
  INV_X1 U11580 ( .A(n10235), .ZN(n10230) );
  NOR2_X1 U11581 ( .A1(n10232), .A2(n10235), .ZN(n10231) );
  NOR2_X1 U11582 ( .A1(n13074), .A2(n13073), .ZN(n13016) );
  NAND2_X1 U11583 ( .A1(n13016), .A2(n13015), .ZN(n13340) );
  INV_X1 U11584 ( .A(n9826), .ZN(n9811) );
  NAND2_X1 U11585 ( .A1(n12008), .A2(n9614), .ZN(n12169) );
  OR2_X1 U11586 ( .A1(n13233), .A2(n13240), .ZN(n13234) );
  OAI21_X1 U11587 ( .B1(n18228), .B2(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n13672), .ZN(n13680) );
  NOR2_X1 U11588 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18369), .ZN(
        n13693) );
  NOR2_X1 U11589 ( .A1(n10079), .A2(n10098), .ZN(n10097) );
  AND2_X1 U11590 ( .A1(n9609), .A2(n10099), .ZN(n10098) );
  INV_X1 U11591 ( .A(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n20650) );
  NOR2_X1 U11592 ( .A1(n13573), .A2(n13574), .ZN(n15128) );
  NOR2_X1 U11593 ( .A1(n13571), .A2(n13700), .ZN(n13570) );
  NAND2_X1 U11594 ( .A1(n16117), .A2(n15919), .ZN(n15945) );
  INV_X1 U11595 ( .A(n17043), .ZN(n15919) );
  NAND3_X1 U11596 ( .A1(n17260), .A2(n17250), .A3(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16128) );
  NAND2_X1 U11597 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10087) );
  OR2_X1 U11598 ( .A1(n15926), .A2(n17318), .ZN(n10015) );
  NAND2_X1 U11599 ( .A1(n17192), .A2(n17235), .ZN(n15356) );
  NAND2_X1 U11600 ( .A1(n9801), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15345) );
  INV_X1 U11601 ( .A(n17332), .ZN(n9801) );
  NAND2_X1 U11602 ( .A1(n17339), .A2(n15315), .ZN(n15316) );
  NAND2_X1 U11603 ( .A1(n17349), .A2(n15337), .ZN(n15339) );
  XNOR2_X1 U11604 ( .A(n16930), .B(n16923), .ZN(n15297) );
  XNOR2_X1 U11605 ( .A(n15329), .B(n16923), .ZN(n9799) );
  AND2_X1 U11606 ( .A1(n12504), .A2(n12690), .ZN(n12705) );
  INV_X1 U11607 ( .A(n13906), .ZN(n10204) );
  OR2_X1 U11608 ( .A1(n11009), .A2(n11008), .ZN(n12278) );
  NAND2_X1 U11609 ( .A1(n13977), .A2(n9851), .ZN(n13916) );
  AND2_X1 U11610 ( .A1(n11010), .A2(n9852), .ZN(n9851) );
  INV_X1 U11611 ( .A(n13997), .ZN(n10201) );
  INV_X1 U11612 ( .A(n9914), .ZN(n9867) );
  INV_X1 U11613 ( .A(n13528), .ZN(n10198) );
  NAND2_X1 U11614 ( .A1(n9870), .A2(n15580), .ZN(n13215) );
  NAND2_X1 U11615 ( .A1(n10569), .A2(n10568), .ZN(n12990) );
  NOR3_X1 U11616 ( .A1(n13982), .A2(n9979), .A3(n13933), .ZN(n13923) );
  NAND2_X1 U11617 ( .A1(n13215), .A2(n11132), .ZN(n10264) );
  NAND2_X1 U11618 ( .A1(n15593), .A2(n15592), .ZN(n15591) );
  NAND2_X1 U11619 ( .A1(n9972), .A2(n9971), .ZN(n12993) );
  INV_X1 U11620 ( .A(n12893), .ZN(n9971) );
  INV_X1 U11621 ( .A(n12894), .ZN(n9972) );
  NAND2_X1 U11622 ( .A1(n12302), .A2(n12372), .ZN(n13887) );
  NAND2_X1 U11623 ( .A1(n12717), .A2(n12705), .ZN(n19824) );
  INV_X1 U11624 ( .A(n10515), .ZN(n10517) );
  INV_X1 U11625 ( .A(n11062), .ZN(n10516) );
  OAI221_X1 U11626 ( .B1(n15684), .B2(n14426), .C1(n15683), .C2(n14426), .A(
        n20446), .ZN(n19897) );
  OAI21_X1 U11627 ( .B1(n11253), .B2(n11201), .A(n11200), .ZN(n11205) );
  INV_X1 U11628 ( .A(n19602), .ZN(n12696) );
  NAND2_X1 U11629 ( .A1(n10499), .A2(n10498), .ZN(n20317) );
  AND2_X1 U11630 ( .A1(n20000), .A2(n20172), .ZN(n20353) );
  NAND2_X1 U11631 ( .A1(n9631), .A2(n19838), .ZN(n20222) );
  XNOR2_X1 U11632 ( .A(n14645), .B(n12227), .ZN(n13853) );
  AND2_X1 U11633 ( .A1(n13781), .A2(n11922), .ZN(n12253) );
  NAND2_X1 U11634 ( .A1(n13790), .A2(n10067), .ZN(n13801) );
  NAND2_X1 U11635 ( .A1(n12225), .A2(n13770), .ZN(n13793) );
  OR2_X1 U11636 ( .A1(n13771), .A2(n13767), .ZN(n12225) );
  NAND2_X1 U11637 ( .A1(n13037), .A2(n13038), .ZN(n13049) );
  AND2_X1 U11638 ( .A1(n13745), .A2(n11874), .ZN(n10072) );
  AND2_X1 U11639 ( .A1(n13750), .A2(n13748), .ZN(n13746) );
  NOR2_X1 U11640 ( .A1(n9672), .A2(n12153), .ZN(n9863) );
  INV_X1 U11641 ( .A(n13031), .ZN(n10155) );
  INV_X1 U11642 ( .A(n11716), .ZN(n11762) );
  INV_X1 U11643 ( .A(n14516), .ZN(n9858) );
  INV_X1 U11644 ( .A(n14513), .ZN(n9859) );
  INV_X1 U11645 ( .A(n11852), .ZN(n18705) );
  NAND2_X1 U11646 ( .A1(n10032), .A2(n11886), .ZN(n10031) );
  AOI21_X1 U11647 ( .B1(n11886), .B2(n10026), .A(n12728), .ZN(n10030) );
  INV_X1 U11648 ( .A(n10219), .ZN(n10212) );
  NAND2_X1 U11649 ( .A1(n9935), .A2(n10216), .ZN(n9934) );
  INV_X1 U11650 ( .A(n14661), .ZN(n9933) );
  OAI21_X1 U11651 ( .B1(n13853), .B2(n13327), .A(n14832), .ZN(n14643) );
  NAND2_X1 U11652 ( .A1(n14720), .A2(n10171), .ZN(n14681) );
  AND3_X1 U11653 ( .A1(n15701), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n12224), .ZN(n14661) );
  INV_X1 U11654 ( .A(n14672), .ZN(n9830) );
  AND2_X1 U11655 ( .A1(n14720), .A2(n9678), .ZN(n14687) );
  NAND2_X1 U11656 ( .A1(n14720), .A2(n10172), .ZN(n14695) );
  NAND2_X1 U11657 ( .A1(n14720), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14702) );
  AND2_X1 U11658 ( .A1(n12189), .A2(n12188), .ZN(n12269) );
  NOR3_X1 U11659 ( .A1(n12268), .A2(n10186), .A3(n12269), .ZN(n14895) );
  NAND2_X1 U11660 ( .A1(n14621), .A2(n12258), .ZN(n12268) );
  NOR2_X1 U11661 ( .A1(n13423), .A2(n12184), .ZN(n14629) );
  AND2_X1 U11662 ( .A1(n14629), .A2(n14619), .ZN(n14621) );
  AND2_X1 U11663 ( .A1(n14762), .A2(n14771), .ZN(n9897) );
  OR2_X1 U11664 ( .A1(n18445), .A2(n13819), .ZN(n14750) );
  NAND2_X1 U11665 ( .A1(n15793), .A2(n9903), .ZN(n9902) );
  INV_X1 U11666 ( .A(n15794), .ZN(n9903) );
  NOR2_X1 U11667 ( .A1(n9905), .A2(n14733), .ZN(n9904) );
  INV_X1 U11668 ( .A(n9906), .ZN(n9905) );
  NAND2_X1 U11669 ( .A1(n15054), .A2(n10243), .ZN(n9931) );
  NAND2_X1 U11670 ( .A1(n10243), .A2(n9877), .ZN(n9876) );
  INV_X1 U11671 ( .A(n13754), .ZN(n9877) );
  INV_X1 U11672 ( .A(n13755), .ZN(n9834) );
  NAND2_X1 U11673 ( .A1(n9714), .A2(n9656), .ZN(n10246) );
  NAND2_X1 U11674 ( .A1(n10248), .A2(n9685), .ZN(n10247) );
  INV_X1 U11675 ( .A(n12087), .ZN(n10177) );
  AND4_X1 U11676 ( .A1(n12142), .A2(n12141), .A3(n12140), .A4(n12139), .ZN(
        n12151) );
  AND4_X1 U11677 ( .A1(n12146), .A2(n12145), .A3(n12144), .A4(n12143), .ZN(
        n12150) );
  INV_X1 U11678 ( .A(n11400), .ZN(n11401) );
  NAND2_X1 U11679 ( .A1(n9857), .A2(n10137), .ZN(n11440) );
  OAI22_X2 U11680 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19525), .B1(n12863), 
        .B2(n19585), .ZN(n19377) );
  OR2_X1 U11681 ( .A1(n16160), .A2(n16161), .ZN(n10085) );
  NOR2_X1 U11682 ( .A1(n17047), .A2(n16170), .ZN(n16169) );
  INV_X1 U11683 ( .A(n10097), .ZN(n10096) );
  AND2_X1 U11684 ( .A1(n16122), .A2(n10105), .ZN(n10102) );
  INV_X1 U11685 ( .A(n17170), .ZN(n10077) );
  NOR2_X1 U11686 ( .A1(n16266), .A2(n9609), .ZN(n16256) );
  NAND2_X1 U11687 ( .A1(n10078), .A2(n10077), .ZN(n10080) );
  INV_X1 U11688 ( .A(n16256), .ZN(n10078) );
  NOR2_X1 U11689 ( .A1(n17178), .A2(n16267), .ZN(n16266) );
  AND2_X1 U11690 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10018) );
  INV_X1 U11691 ( .A(n15257), .ZN(n10019) );
  INV_X1 U11692 ( .A(n15258), .ZN(n10021) );
  AOI21_X1 U11693 ( .B1(n13682), .B2(n9693), .A(n13696), .ZN(n15422) );
  NOR2_X1 U11694 ( .A1(n15945), .A2(n16167), .ZN(n15944) );
  AND2_X1 U11695 ( .A1(n17124), .A2(n10106), .ZN(n16117) );
  AND2_X1 U11696 ( .A1(n10107), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10106) );
  AND2_X1 U11697 ( .A1(n17186), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10281) );
  NAND2_X1 U11698 ( .A1(n17232), .A2(n9802), .ZN(n17131) );
  INV_X1 U11699 ( .A(n17232), .ZN(n17576) );
  NAND2_X1 U11700 ( .A1(n17061), .A2(n15969), .ZN(n15406) );
  OAI21_X1 U11701 ( .B1(n15359), .B2(n17235), .A(n17076), .ZN(n15360) );
  INV_X1 U11702 ( .A(n10025), .ZN(n15359) );
  NAND2_X1 U11703 ( .A1(n17090), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17415) );
  INV_X1 U11704 ( .A(n17092), .ZN(n10023) );
  NAND2_X1 U11705 ( .A1(n17235), .A2(n17435), .ZN(n10024) );
  NAND2_X1 U11706 ( .A1(n9842), .A2(n9841), .ZN(n17076) );
  AND2_X1 U11707 ( .A1(n10023), .A2(n17418), .ZN(n9842) );
  AND2_X1 U11708 ( .A1(n17235), .A2(n17102), .ZN(n17092) );
  NOR2_X1 U11709 ( .A1(n17091), .A2(n17435), .ZN(n17090) );
  NOR2_X1 U11710 ( .A1(n17131), .A2(n15348), .ZN(n17450) );
  NAND2_X1 U11711 ( .A1(n17616), .A2(n17609), .ZN(n10004) );
  NAND2_X1 U11712 ( .A1(n17327), .A2(n17235), .ZN(n17300) );
  NAND2_X1 U11713 ( .A1(n17355), .A2(n17667), .ZN(n9835) );
  NAND2_X1 U11714 ( .A1(n15313), .A2(n17368), .ZN(n17357) );
  NAND2_X1 U11715 ( .A1(n17741), .A2(n17630), .ZN(n17468) );
  AND2_X1 U11716 ( .A1(n13961), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19675) );
  AND2_X1 U11717 ( .A1(n13063), .A2(n12383), .ZN(n19687) );
  INV_X1 U11718 ( .A(n14118), .ZN(n14036) );
  NAND2_X1 U11719 ( .A1(n13905), .A2(n11061), .ZN(n13737) );
  AND2_X1 U11720 ( .A1(n14190), .A2(n11213), .ZN(n15566) );
  INV_X1 U11721 ( .A(n19787), .ZN(n19835) );
  NAND2_X1 U11722 ( .A1(n10259), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10257) );
  AND2_X1 U11723 ( .A1(n10258), .A2(n14238), .ZN(n10256) );
  NAND2_X1 U11724 ( .A1(n9974), .A2(n19807), .ZN(n9973) );
  INV_X1 U11725 ( .A(n14220), .ZN(n9974) );
  XNOR2_X1 U11726 ( .A(n11150), .B(n14247), .ZN(n14267) );
  XNOR2_X1 U11727 ( .A(n14114), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14283) );
  INV_X1 U11728 ( .A(n11148), .ZN(n14112) );
  NAND2_X1 U11729 ( .A1(n9990), .A2(n11247), .ZN(n12703) );
  XNOR2_X1 U11730 ( .A(n19994), .B(n10601), .ZN(n20524) );
  INV_X1 U11731 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19586) );
  INV_X1 U11732 ( .A(n18540), .ZN(n18639) );
  XNOR2_X1 U11733 ( .A(n14457), .B(n14456), .ZN(n15700) );
  NAND2_X1 U11734 ( .A1(n10146), .A2(n9695), .ZN(n10145) );
  AND2_X1 U11735 ( .A1(n10153), .A2(n10152), .ZN(n10151) );
  INV_X1 U11736 ( .A(n12947), .ZN(n10152) );
  AND2_X1 U11737 ( .A1(n14540), .A2(n12630), .ZN(n14522) );
  AND2_X1 U11738 ( .A1(n10210), .A2(n18808), .ZN(n10055) );
  NAND2_X1 U11739 ( .A1(n19552), .A2(n19377), .ZN(n18811) );
  NAND2_X1 U11740 ( .A1(n14668), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10164) );
  AND2_X1 U11741 ( .A1(n10210), .A2(n18846), .ZN(n10209) );
  AND2_X1 U11742 ( .A1(n10213), .A2(n10056), .ZN(n10211) );
  INV_X1 U11743 ( .A(n10214), .ZN(n10213) );
  NAND2_X1 U11744 ( .A1(n9935), .A2(n9690), .ZN(n10056) );
  OAI21_X1 U11745 ( .B1(n10219), .B2(n10216), .A(n10217), .ZN(n10214) );
  INV_X1 U11746 ( .A(n14836), .ZN(n10035) );
  AOI21_X1 U11747 ( .B1(n15004), .B2(n18856), .A(n15006), .ZN(n9881) );
  NAND2_X1 U11748 ( .A1(n9884), .A2(n9883), .ZN(n9882) );
  NAND2_X1 U11749 ( .A1(n18861), .A2(n18864), .ZN(n9883) );
  OR2_X1 U11750 ( .A1(n12593), .A2(n12559), .ZN(n18839) );
  OR2_X1 U11751 ( .A1(n12593), .A2(n12562), .ZN(n15898) );
  INV_X1 U11752 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19571) );
  INV_X1 U11753 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19535) );
  NOR2_X1 U11754 ( .A1(n19373), .A2(n19019), .ZN(n19089) );
  NOR2_X1 U11755 ( .A1(n19108), .A2(n19297), .ZN(n19095) );
  INV_X1 U11756 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18394) );
  NOR2_X2 U11757 ( .A1(n17778), .A2(n16772), .ZN(n16765) );
  NAND2_X1 U11758 ( .A1(n16791), .A2(P3_EAX_REG_29__SCAN_IN), .ZN(n16790) );
  NAND2_X1 U11759 ( .A1(n16818), .A2(n17778), .ZN(n16812) );
  NOR2_X1 U11760 ( .A1(n16819), .A2(n16993), .ZN(n16818) );
  NOR2_X1 U11761 ( .A1(n15225), .A2(n15224), .ZN(n16902) );
  NOR2_X1 U11762 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n15351), .ZN(
        n17327) );
  NAND2_X1 U11763 ( .A1(n15351), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17310) );
  NOR2_X1 U11764 ( .A1(n15979), .A2(n17411), .ZN(n17309) );
  NOR2_X1 U11765 ( .A1(n18391), .A2(n16095), .ZN(n17401) );
  INV_X1 U11766 ( .A(n17401), .ZN(n17412) );
  NAND2_X1 U11767 ( .A1(n10009), .A2(n10005), .ZN(n15965) );
  NAND2_X1 U11768 ( .A1(n10007), .A2(n10006), .ZN(n10005) );
  NAND2_X1 U11769 ( .A1(n10010), .A2(n15928), .ZN(n10009) );
  INV_X1 U11770 ( .A(n15928), .ZN(n10006) );
  NAND2_X1 U11771 ( .A1(n17419), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9794) );
  INV_X1 U11772 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17616) );
  NOR2_X1 U11773 ( .A1(n11201), .A2(n11250), .ZN(n11179) );
  AOI21_X1 U11774 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n18209), .A(
        n13670), .ZN(n13671) );
  NAND2_X1 U11775 ( .A1(n11154), .A2(n11153), .ZN(n11186) );
  CLKBUF_X1 U11776 ( .A(n10570), .Z(n11219) );
  INV_X1 U11777 ( .A(n11132), .ZN(n10262) );
  AND3_X1 U11778 ( .A1(n10496), .A2(n10495), .A3(n10494), .ZN(n10503) );
  OR2_X1 U11779 ( .A1(n10442), .A2(n10441), .ZN(n10443) );
  OR2_X1 U11780 ( .A1(n19839), .A2(n20446), .ZN(n10542) );
  OAI21_X1 U11781 ( .B1(n10408), .B2(n10406), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n10536) );
  NOR2_X1 U11782 ( .A1(n12517), .A2(n20446), .ZN(n10195) );
  INV_X1 U11783 ( .A(n13472), .ZN(n13859) );
  OR2_X1 U11784 ( .A1(n12027), .A2(n12026), .ZN(n13299) );
  NAND2_X1 U11785 ( .A1(n13269), .A2(n13268), .ZN(n9826) );
  OR2_X1 U11786 ( .A1(n12099), .A2(n12098), .ZN(n12221) );
  NOR2_X1 U11787 ( .A1(n10038), .A2(n15904), .ZN(n10036) );
  AND2_X1 U11788 ( .A1(n12455), .A2(n9644), .ZN(n11388) );
  NOR2_X1 U11789 ( .A1(n12792), .A2(n15904), .ZN(n9910) );
  INV_X1 U11790 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9878) );
  INV_X1 U11791 ( .A(n11363), .ZN(n12584) );
  XNOR2_X1 U11792 ( .A(n11827), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11833) );
  OR2_X1 U11793 ( .A1(n11847), .A2(n11846), .ZN(n12219) );
  AND3_X1 U11794 ( .A1(n15192), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(
        n11843), .ZN(n12214) );
  AOI21_X1 U11795 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n17987), .A(
        n13669), .ZN(n13677) );
  AND2_X1 U11796 ( .A1(n13695), .A2(n13693), .ZN(n13669) );
  NAND2_X1 U11797 ( .A1(n18355), .A2(n18345), .ZN(n13575) );
  NAND2_X1 U11798 ( .A1(n18362), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13571) );
  NOR2_X1 U11799 ( .A1(n16918), .A2(n15311), .ZN(n15294) );
  AOI21_X1 U11800 ( .B1(n17748), .B2(n16111), .A(n15423), .ZN(n13653) );
  NAND2_X1 U11801 ( .A1(n16890), .A2(n13663), .ZN(n13683) );
  OR2_X1 U11802 ( .A1(n11055), .A2(n14107), .ZN(n11056) );
  INV_X1 U11803 ( .A(n12278), .ZN(n11010) );
  NAND2_X1 U11804 ( .A1(n13957), .A2(n10197), .ZN(n10196) );
  INV_X1 U11805 ( .A(n14022), .ZN(n10197) );
  AND2_X1 U11806 ( .A1(n10746), .A2(n10200), .ZN(n10199) );
  OR2_X1 U11807 ( .A1(n15528), .A2(n13500), .ZN(n10200) );
  AND2_X1 U11808 ( .A1(n13505), .A2(n13520), .ZN(n10746) );
  NAND2_X1 U11809 ( .A1(n13501), .A2(n13500), .ZN(n13503) );
  AND3_X1 U11810 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A3(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10589) );
  NAND2_X1 U11811 ( .A1(n9708), .A2(n10600), .ZN(n10641) );
  NAND2_X1 U11812 ( .A1(n10275), .A2(n10277), .ZN(n9912) );
  NAND2_X1 U11813 ( .A1(n10408), .A2(n10278), .ZN(n10277) );
  NOR2_X1 U11814 ( .A1(n12617), .A2(n20446), .ZN(n10278) );
  OAI21_X1 U11815 ( .B1(n12952), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n10502), 
        .ZN(n9845) );
  AOI21_X1 U11816 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20446), .A(
        n11199), .ZN(n11200) );
  OAI21_X1 U11817 ( .B1(n11198), .B2(n11197), .A(n11196), .ZN(n11199) );
  AND2_X1 U11818 ( .A1(n10543), .A2(n10542), .ZN(n11201) );
  NAND2_X1 U11819 ( .A1(n9816), .A2(n11063), .ZN(n12686) );
  NAND2_X1 U11820 ( .A1(n10397), .A2(n9615), .ZN(n10274) );
  INV_X1 U11821 ( .A(n11210), .ZN(n12420) );
  INV_X1 U11822 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12926) );
  NAND2_X1 U11823 ( .A1(n10062), .A2(n10061), .ZN(n14645) );
  INV_X1 U11824 ( .A(n13851), .ZN(n10061) );
  NOR2_X1 U11825 ( .A1(n13839), .A2(n13840), .ZN(n10062) );
  AND2_X1 U11826 ( .A1(n9674), .A2(n10064), .ZN(n10063) );
  AND2_X1 U11827 ( .A1(n11402), .A2(n18919), .ZN(n11716) );
  AND2_X1 U11828 ( .A1(n9643), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11402) );
  INV_X1 U11829 ( .A(n14565), .ZN(n10175) );
  OAI21_X1 U11830 ( .B1(n11745), .B2(n9755), .A(n9860), .ZN(n11768) );
  NAND2_X1 U11831 ( .A1(n11745), .A2(n9757), .ZN(n9860) );
  NAND2_X1 U11832 ( .A1(n10139), .A2(n10140), .ZN(n11722) );
  NAND2_X1 U11833 ( .A1(n10141), .A2(n9673), .ZN(n10140) );
  OR2_X1 U11834 ( .A1(n12113), .A2(n12112), .ZN(n13323) );
  NAND2_X1 U11835 ( .A1(n9614), .A2(n18919), .ZN(n12065) );
  NOR2_X1 U11836 ( .A1(n14688), .A2(n10136), .ZN(n10135) );
  INV_X1 U11837 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10136) );
  AND2_X1 U11838 ( .A1(n10112), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10111) );
  NOR2_X1 U11839 ( .A1(n10114), .A2(n10113), .ZN(n10112) );
  NAND2_X1 U11840 ( .A1(n10218), .A2(n10222), .ZN(n10060) );
  INV_X1 U11841 ( .A(n14643), .ZN(n10218) );
  AND2_X1 U11842 ( .A1(n10239), .A2(n9716), .ZN(n10236) );
  AND2_X1 U11843 ( .A1(n9678), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10171) );
  NOR2_X1 U11844 ( .A1(n14694), .A2(n10240), .ZN(n10239) );
  INV_X1 U11845 ( .A(n14705), .ZN(n10240) );
  NAND2_X1 U11846 ( .A1(n10185), .A2(n14894), .ZN(n10184) );
  INV_X1 U11847 ( .A(n12269), .ZN(n10185) );
  NOR2_X1 U11848 ( .A1(n14877), .A2(n14886), .ZN(n10172) );
  AND2_X1 U11849 ( .A1(n15737), .A2(n12224), .ZN(n13838) );
  AOI21_X1 U11850 ( .B1(n14724), .B2(n9938), .A(n9664), .ZN(n9937) );
  NAND2_X1 U11851 ( .A1(n14724), .A2(n9940), .ZN(n9939) );
  NAND2_X1 U11852 ( .A1(n12270), .A2(n10046), .ZN(n10045) );
  INV_X1 U11853 ( .A(n14528), .ZN(n10046) );
  NOR2_X1 U11854 ( .A1(n12630), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12004) );
  NOR2_X1 U11855 ( .A1(n13760), .A2(n15061), .ZN(n9918) );
  NAND2_X1 U11856 ( .A1(n10169), .A2(n10170), .ZN(n9919) );
  NAND2_X1 U11857 ( .A1(n9927), .A2(n13476), .ZN(n13743) );
  NAND2_X1 U11858 ( .A1(n13856), .A2(n13327), .ZN(n9927) );
  NAND2_X1 U11859 ( .A1(n15848), .A2(n13355), .ZN(n13359) );
  INV_X1 U11860 ( .A(n13299), .ZN(n13356) );
  INV_X1 U11861 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11275) );
  NAND2_X1 U11862 ( .A1(n9945), .A2(n9943), .ZN(n12794) );
  AND2_X1 U11863 ( .A1(n11362), .A2(n12626), .ZN(n9943) );
  NAND2_X1 U11864 ( .A1(n12576), .A2(n11361), .ZN(n11406) );
  INV_X1 U11865 ( .A(n10138), .ZN(n9857) );
  CLKBUF_X1 U11866 ( .A(n12448), .Z(n12815) );
  NAND2_X1 U11867 ( .A1(n11296), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9809) );
  NAND2_X1 U11868 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19571), .ZN(
        n11837) );
  NOR4_X1 U11869 ( .A1(n13663), .A2(n15093), .A3(n13662), .A4(n13656), .ZN(
        n13665) );
  OR2_X1 U11870 ( .A1(n13571), .A2(n13572), .ZN(n15151) );
  NOR2_X1 U11871 ( .A1(n15200), .A2(n13654), .ZN(n13664) );
  NOR2_X1 U11872 ( .A1(n10110), .A2(n10108), .ZN(n10107) );
  NAND2_X1 U11873 ( .A1(n9646), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10108) );
  INV_X1 U11874 ( .A(n17083), .ZN(n10110) );
  AND2_X1 U11875 ( .A1(n18349), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10014) );
  NAND2_X1 U11876 ( .A1(n10003), .A2(n10002), .ZN(n10001) );
  INV_X1 U11877 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10002) );
  INV_X1 U11878 ( .A(n10004), .ZN(n10003) );
  INV_X1 U11879 ( .A(n13683), .ZN(n15197) );
  INV_X1 U11880 ( .A(n16930), .ZN(n15320) );
  AOI21_X1 U11881 ( .B1(n13667), .B2(n17741), .A(n18215), .ZN(n18176) );
  NOR2_X1 U11882 ( .A1(n13663), .A2(n15200), .ZN(n18180) );
  INV_X1 U11883 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n20593) );
  AND2_X1 U11884 ( .A1(n12483), .A2(n12279), .ZN(n12414) );
  NAND2_X1 U11885 ( .A1(n13063), .A2(n12380), .ZN(n13963) );
  NAND2_X1 U11886 ( .A1(n12346), .A2(n9981), .ZN(n9980) );
  INV_X1 U11887 ( .A(n14335), .ZN(n9981) );
  NOR3_X1 U11888 ( .A1(n14021), .A2(n9985), .A3(n13964), .ZN(n14010) );
  AND2_X1 U11889 ( .A1(n15444), .A2(n12280), .ZN(n10937) );
  AND2_X1 U11890 ( .A1(n10877), .A2(n10876), .ZN(n14052) );
  AND2_X1 U11891 ( .A1(n12688), .A2(n12598), .ZN(n19716) );
  INV_X1 U11892 ( .A(n12959), .ZN(n19763) );
  AND2_X1 U11893 ( .A1(n11003), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11004) );
  NAND2_X1 U11894 ( .A1(n11004), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11055) );
  NAND2_X1 U11895 ( .A1(n13977), .A2(n13979), .ZN(n13978) );
  NAND2_X1 U11896 ( .A1(n10922), .A2(n10921), .ZN(n13943) );
  OR2_X1 U11897 ( .A1(n14149), .A2(n11028), .ZN(n10921) );
  NAND2_X1 U11898 ( .A1(n13999), .A2(n10202), .ZN(n14051) );
  AND2_X1 U11899 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n10874), .ZN(
        n10875) );
  INV_X1 U11900 ( .A(n10873), .ZN(n10874) );
  AND2_X1 U11901 ( .A1(n10858), .A2(n10857), .ZN(n14000) );
  AND2_X1 U11902 ( .A1(n13999), .A2(n14000), .ZN(n14053) );
  NOR2_X1 U11903 ( .A1(n10840), .A2(n15487), .ZN(n10841) );
  NAND2_X1 U11904 ( .A1(n10841), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10873) );
  NAND2_X1 U11905 ( .A1(n13526), .A2(n9854), .ZN(n14011) );
  NOR3_X1 U11906 ( .A1(n10196), .A2(n14014), .A3(n14077), .ZN(n9854) );
  NOR2_X1 U11907 ( .A1(n10797), .A2(n15498), .ZN(n10810) );
  NAND2_X1 U11908 ( .A1(n10794), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10797) );
  NAND2_X1 U11909 ( .A1(n13526), .A2(n10780), .ZN(n14074) );
  NOR2_X1 U11910 ( .A1(n20593), .A2(n10748), .ZN(n10794) );
  INV_X1 U11911 ( .A(n10747), .ZN(n10748) );
  NAND2_X1 U11912 ( .A1(n10731), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10715) );
  INV_X1 U11913 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n20629) );
  NAND2_X1 U11914 ( .A1(n13501), .A2(n10199), .ZN(n13527) );
  INV_X1 U11915 ( .A(n10714), .ZN(n10731) );
  NOR2_X1 U11916 ( .A1(n10699), .A2(n10698), .ZN(n10700) );
  NAND2_X1 U11917 ( .A1(n10682), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10699) );
  INV_X1 U11918 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10698) );
  INV_X1 U11919 ( .A(n13181), .ZN(n9848) );
  NOR2_X1 U11920 ( .A1(n10666), .A2(n10665), .ZN(n10682) );
  INV_X1 U11921 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10665) );
  AND3_X1 U11922 ( .A1(n10664), .A2(n10663), .A3(n10662), .ZN(n13147) );
  AOI21_X1 U11923 ( .B1(n11114), .B2(n10773), .A(n10648), .ZN(n13092) );
  NAND2_X1 U11924 ( .A1(n10650), .A2(n10649), .ZN(n13146) );
  NOR2_X1 U11925 ( .A1(n10632), .A2(n19654), .ZN(n10645) );
  INV_X1 U11926 ( .A(n13005), .ZN(n9846) );
  NAND2_X1 U11927 ( .A1(n10614), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10632) );
  NOR2_X1 U11928 ( .A1(n12691), .A2(n19602), .ZN(n12688) );
  AND2_X1 U11929 ( .A1(n12370), .A2(n12369), .ZN(n13933) );
  NOR2_X1 U11930 ( .A1(n13982), .A2(n13933), .ZN(n13932) );
  OR2_X1 U11931 ( .A1(n14334), .A2(n13992), .ZN(n13994) );
  NOR2_X1 U11932 ( .A1(n13994), .A2(n13944), .ZN(n13988) );
  NAND2_X1 U11933 ( .A1(n10280), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10279) );
  NOR2_X1 U11934 ( .A1(n9914), .A2(n9768), .ZN(n9866) );
  NOR2_X1 U11935 ( .A1(n14021), .A2(n13964), .ZN(n14016) );
  NOR2_X1 U11936 ( .A1(n14186), .A2(n14184), .ZN(n14367) );
  NAND2_X1 U11937 ( .A1(n9821), .A2(n11139), .ZN(n14366) );
  OAI21_X1 U11938 ( .B1(n14182), .B2(n14185), .A(n11141), .ZN(n9821) );
  AND3_X1 U11939 ( .A1(n12339), .A2(n12360), .A3(n12338), .ZN(n14019) );
  OR2_X1 U11940 ( .A1(n14401), .A2(n14019), .ZN(n14021) );
  NOR2_X1 U11941 ( .A1(n13534), .A2(n13533), .ZN(n14399) );
  AND3_X1 U11942 ( .A1(n12328), .A2(n12360), .A3(n12327), .ZN(n13524) );
  NAND2_X1 U11943 ( .A1(n13149), .A2(n9734), .ZN(n15520) );
  INV_X1 U11944 ( .A(n15523), .ZN(n9986) );
  NAND2_X1 U11945 ( .A1(n10264), .A2(n10263), .ZN(n15570) );
  CLKBUF_X1 U11946 ( .A(n13546), .Z(n15571) );
  NAND2_X1 U11947 ( .A1(n13149), .A2(n9655), .ZN(n15522) );
  NAND2_X1 U11948 ( .A1(n13149), .A2(n13148), .ZN(n13183) );
  NOR2_X1 U11949 ( .A1(n15669), .A2(n15667), .ZN(n13097) );
  AND2_X1 U11950 ( .A1(n12315), .A2(n12314), .ZN(n13096) );
  AND2_X1 U11951 ( .A1(n13097), .A2(n13096), .ZN(n13149) );
  AOI21_X1 U11952 ( .B1(n11113), .B2(n10269), .A(n9707), .ZN(n10268) );
  OR2_X1 U11953 ( .A1(n13009), .A2(n13010), .ZN(n15669) );
  NAND2_X1 U11954 ( .A1(n12995), .A2(n11089), .ZN(n19785) );
  NAND2_X1 U11955 ( .A1(n19785), .A2(n19784), .ZN(n19783) );
  NAND2_X1 U11956 ( .A1(n12991), .A2(n12974), .ZN(n13009) );
  NOR2_X1 U11957 ( .A1(n12993), .A2(n12992), .ZN(n12991) );
  AND2_X1 U11958 ( .A1(n13554), .A2(n15609), .ZN(n13559) );
  OAI21_X1 U11959 ( .B1(n19922), .B2(n11160), .A(n11069), .ZN(n12678) );
  NAND2_X1 U11960 ( .A1(n12678), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12680) );
  NAND2_X1 U11961 ( .A1(n9819), .A2(n9818), .ZN(n12715) );
  NAND2_X1 U11962 ( .A1(n12423), .A2(n9991), .ZN(n9990) );
  INV_X1 U11963 ( .A(n10535), .ZN(n9783) );
  INV_X1 U11964 ( .A(n10429), .ZN(n10190) );
  NAND2_X1 U11965 ( .A1(n10500), .A2(n10423), .ZN(n9916) );
  AND2_X1 U11966 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20000), .ZN(n19885) );
  INV_X1 U11967 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20315) );
  AND2_X1 U11968 ( .A1(n20445), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11206) );
  INV_X1 U11969 ( .A(n11206), .ZN(n15395) );
  OR2_X1 U11970 ( .A1(n12833), .A2(n12208), .ZN(n12843) );
  OR2_X1 U11971 ( .A1(n15696), .A2(n15705), .ZN(n10116) );
  OR2_X1 U11972 ( .A1(n15716), .A2(n9767), .ZN(n10115) );
  INV_X1 U11973 ( .A(n10062), .ZN(n13850) );
  INV_X1 U11974 ( .A(n15749), .ZN(n10127) );
  NAND2_X1 U11975 ( .A1(n12255), .A2(n9674), .ZN(n13828) );
  NAND2_X1 U11976 ( .A1(n12253), .A2(n12226), .ZN(n12265) );
  NAND2_X1 U11977 ( .A1(n12255), .A2(n12266), .ZN(n13824) );
  NAND2_X1 U11978 ( .A1(n10119), .A2(n10118), .ZN(n10120) );
  AOI21_X1 U11979 ( .B1(n15696), .B2(n18443), .A(n14746), .ZN(n10118) );
  OR2_X1 U11980 ( .A1(n18442), .A2(n18443), .ZN(n10121) );
  AND2_X1 U11981 ( .A1(n10067), .A2(n10066), .ZN(n10065) );
  INV_X1 U11982 ( .A(n13800), .ZN(n10066) );
  NAND2_X1 U11983 ( .A1(n13790), .A2(n10069), .ZN(n13786) );
  AND2_X1 U11984 ( .A1(n13790), .A2(n13788), .ZN(n13782) );
  NAND2_X1 U11985 ( .A1(n13119), .A2(n13120), .ZN(n13176) );
  AND2_X1 U11986 ( .A1(n10072), .A2(n10071), .ZN(n10070) );
  NAND2_X1 U11987 ( .A1(n13746), .A2(n13745), .ZN(n13757) );
  AND2_X1 U11988 ( .A1(n12218), .A2(n12217), .ZN(n13073) );
  INV_X1 U11989 ( .A(n14460), .ZN(n10149) );
  INV_X1 U11990 ( .A(n10148), .ZN(n10143) );
  INV_X1 U11991 ( .A(n11823), .ZN(n10147) );
  AND2_X1 U11992 ( .A1(n11468), .A2(n11469), .ZN(n10153) );
  AND2_X1 U11993 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n12724), .ZN(
        n11468) );
  AND2_X1 U11994 ( .A1(n9861), .A2(n9739), .ZN(n12775) );
  AND2_X1 U11995 ( .A1(n9751), .A2(n10174), .ZN(n10173) );
  INV_X1 U11996 ( .A(n14558), .ZN(n10174) );
  XNOR2_X1 U11997 ( .A(n11768), .B(n11767), .ZN(n14478) );
  NAND2_X1 U11998 ( .A1(n14581), .A2(n14573), .ZN(n14572) );
  NAND2_X1 U11999 ( .A1(n10158), .A2(n10157), .ZN(n10156) );
  INV_X1 U12000 ( .A(n14533), .ZN(n10157) );
  INV_X1 U12001 ( .A(n10159), .ZN(n10158) );
  OR2_X1 U12002 ( .A1(n13195), .A2(n10159), .ZN(n14534) );
  NOR2_X1 U12003 ( .A1(n13195), .A2(n13196), .ZN(n13386) );
  AND2_X1 U12004 ( .A1(n10188), .A2(n12160), .ZN(n10187) );
  AND2_X1 U12005 ( .A1(n12635), .A2(n10189), .ZN(n15884) );
  NAND2_X1 U12006 ( .A1(n12635), .A2(n10188), .ZN(n12746) );
  NAND2_X1 U12007 ( .A1(n12635), .A2(n12634), .ZN(n15885) );
  NOR2_X1 U12008 ( .A1(n18691), .A2(n12632), .ZN(n13199) );
  AND2_X1 U12009 ( .A1(n18704), .A2(n19582), .ZN(n18737) );
  AND2_X1 U12010 ( .A1(n12397), .A2(n9643), .ZN(n12401) );
  OAI21_X1 U12011 ( .B1(n12248), .B2(n12247), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n14610) );
  INV_X1 U12012 ( .A(n14610), .ZN(n14634) );
  NAND2_X1 U12013 ( .A1(n11974), .A2(n9670), .ZN(n11970) );
  NAND2_X1 U12014 ( .A1(n11974), .A2(n10135), .ZN(n11972) );
  NOR2_X1 U12015 ( .A1(n14537), .A2(n14528), .ZN(n14529) );
  NAND2_X1 U12016 ( .A1(n10123), .A2(n11964), .ZN(n10122) );
  INV_X1 U12017 ( .A(n10124), .ZN(n10123) );
  NAND2_X1 U12018 ( .A1(n13119), .A2(n10050), .ZN(n13416) );
  NAND2_X1 U12019 ( .A1(n13119), .A2(n10052), .ZN(n13207) );
  NOR2_X1 U12020 ( .A1(n13026), .A2(n13027), .ZN(n13037) );
  NOR2_X1 U12021 ( .A1(n10132), .A2(n15824), .ZN(n10131) );
  NAND2_X1 U12022 ( .A1(n12946), .A2(n12945), .ZN(n12944) );
  INV_X1 U12023 ( .A(n10132), .ZN(n10130) );
  NAND2_X1 U12024 ( .A1(n11443), .A2(n11441), .ZN(n10027) );
  AND2_X1 U12025 ( .A1(n11886), .A2(n10029), .ZN(n10028) );
  NAND2_X1 U12026 ( .A1(n11442), .A2(n11441), .ZN(n10029) );
  NAND2_X1 U12027 ( .A1(n10034), .A2(n9652), .ZN(n12727) );
  NAND3_X1 U12028 ( .A1(n13357), .A2(n15849), .A3(n13331), .ZN(n15848) );
  NAND2_X1 U12029 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11997) );
  INV_X1 U12030 ( .A(n10222), .ZN(n10220) );
  NAND2_X1 U12031 ( .A1(n10058), .A2(n10057), .ZN(n10217) );
  NAND2_X1 U12032 ( .A1(n10222), .A2(n10221), .ZN(n10057) );
  NAND2_X1 U12033 ( .A1(n10060), .A2(n10059), .ZN(n10058) );
  INV_X1 U12034 ( .A(n10221), .ZN(n10059) );
  AND2_X1 U12035 ( .A1(n14643), .A2(n10216), .ZN(n10215) );
  INV_X1 U12036 ( .A(n9935), .ZN(n14663) );
  NAND2_X1 U12037 ( .A1(n10040), .A2(n14470), .ZN(n10039) );
  INV_X1 U12038 ( .A(n10041), .ZN(n10040) );
  NOR2_X1 U12039 ( .A1(n15729), .A2(n13327), .ZN(n14675) );
  NOR2_X1 U12040 ( .A1(n14503), .A2(n10041), .ZN(n14475) );
  OR2_X1 U12041 ( .A1(n13847), .A2(n14886), .ZN(n14707) );
  AND2_X1 U12042 ( .A1(n10237), .A2(n10238), .ZN(n14704) );
  NAND2_X1 U12043 ( .A1(n14704), .A2(n14705), .ZN(n14703) );
  NOR2_X1 U12044 ( .A1(n14503), .A2(n14492), .ZN(n14491) );
  INV_X1 U12045 ( .A(n9936), .ZN(n14716) );
  AND2_X1 U12046 ( .A1(n10167), .A2(n14893), .ZN(n9967) );
  NOR3_X1 U12047 ( .A1(n14537), .A2(n10048), .A3(n14528), .ZN(n12271) );
  NAND2_X1 U12048 ( .A1(n9968), .A2(n10167), .ZN(n14919) );
  INV_X1 U12049 ( .A(n13415), .ZN(n10049) );
  INV_X1 U12050 ( .A(n13391), .ZN(n10182) );
  NOR2_X1 U12051 ( .A1(n15855), .A2(n9723), .ZN(n13392) );
  NOR2_X1 U12052 ( .A1(n12944), .A2(n12903), .ZN(n12966) );
  NAND2_X1 U12053 ( .A1(n12966), .A2(n12967), .ZN(n13026) );
  NOR2_X1 U12054 ( .A1(n15054), .A2(n15056), .ZN(n15053) );
  INV_X1 U12055 ( .A(n9803), .ZN(n9805) );
  NAND2_X1 U12056 ( .A1(n10225), .A2(n13744), .ZN(n15827) );
  XNOR2_X1 U12057 ( .A(n13743), .B(n13491), .ZN(n13741) );
  AOI21_X1 U12058 ( .B1(n9806), .B2(n9965), .A(n9661), .ZN(n9961) );
  AOI21_X1 U12059 ( .B1(n10228), .B2(n10231), .A(n9749), .ZN(n10226) );
  OR2_X1 U12060 ( .A1(n14943), .A2(n18855), .ZN(n18837) );
  AND2_X2 U12061 ( .A1(n11397), .A2(n11396), .ZN(n14440) );
  INV_X1 U12062 ( .A(n11421), .ZN(n11396) );
  NAND2_X1 U12063 ( .A1(n13187), .A2(n12461), .ZN(n9955) );
  INV_X1 U12064 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12792) );
  INV_X1 U12065 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9941) );
  XNOR2_X1 U12066 ( .A(n11438), .B(n9729), .ZN(n10138) );
  AND2_X1 U12067 ( .A1(n19546), .A2(n19557), .ZN(n19161) );
  AND2_X1 U12068 ( .A1(n19540), .A2(n19566), .ZN(n18959) );
  NAND2_X1 U12069 ( .A1(n19540), .A2(n19128), .ZN(n19108) );
  NAND2_X2 U12070 ( .A1(n9807), .A2(n11337), .ZN(n18900) );
  OR2_X1 U12071 ( .A1(n19540), .A2(n19566), .ZN(n19292) );
  INV_X1 U12072 ( .A(n18923), .ZN(n18915) );
  INV_X1 U12073 ( .A(n18924), .ZN(n18917) );
  OR2_X1 U12074 ( .A1(n19540), .A2(n19128), .ZN(n19331) );
  OR2_X1 U12075 ( .A1(n19546), .A2(n19557), .ZN(n19373) );
  OAI21_X1 U12076 ( .B1(n13681), .B2(n13680), .A(n13694), .ZN(n18222) );
  AND2_X1 U12077 ( .A1(n10085), .A2(n10073), .ZN(n16151) );
  INV_X1 U12078 ( .A(n10095), .ZN(n10092) );
  NOR2_X1 U12079 ( .A1(n16201), .A2(n10096), .ZN(n10093) );
  AOI21_X1 U12080 ( .B1(n10097), .B2(n17075), .A(n16183), .ZN(n10095) );
  NOR2_X1 U12081 ( .A1(n18311), .A2(n16223), .ZN(n16140) );
  OR2_X1 U12082 ( .A1(n16285), .A2(n17205), .ZN(n10074) );
  OR2_X1 U12083 ( .A1(n20706), .A2(n16327), .ZN(n16310) );
  NOR2_X1 U12084 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n16336), .ZN(n16320) );
  NAND2_X1 U12085 ( .A1(n16470), .A2(n16136), .ZN(n16353) );
  OR2_X1 U12086 ( .A1(n13700), .A2(n18205), .ZN(n9683) );
  NOR2_X1 U12087 ( .A1(n16111), .A2(n18384), .ZN(n16131) );
  NAND2_X1 U12088 ( .A1(n16784), .A2(n17772), .ZN(n18187) );
  INV_X1 U12089 ( .A(n18187), .ZN(n15423) );
  NOR2_X1 U12090 ( .A1(n16975), .A2(n16936), .ZN(n16953) );
  NAND2_X1 U12091 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17043) );
  NAND2_X1 U12092 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15918) );
  INV_X1 U12093 ( .A(n17228), .ZN(n17250) );
  NAND2_X1 U12094 ( .A1(n10089), .A2(n10088), .ZN(n17244) );
  AND2_X1 U12095 ( .A1(n10090), .A2(n10086), .ZN(n10088) );
  NOR2_X1 U12096 ( .A1(n10087), .A2(n17353), .ZN(n10086) );
  NAND2_X1 U12097 ( .A1(n17328), .A2(n15318), .ZN(n15351) );
  NAND2_X1 U12098 ( .A1(n10090), .A2(n10091), .ZN(n17313) );
  NOR2_X1 U12099 ( .A1(n17353), .A2(n16410), .ZN(n10091) );
  INV_X1 U12100 ( .A(n17741), .ZN(n18391) );
  INV_X1 U12101 ( .A(n15958), .ZN(n10011) );
  NAND2_X1 U12102 ( .A1(n10015), .A2(n10013), .ZN(n10012) );
  NAND2_X1 U12103 ( .A1(n10015), .A2(n10008), .ZN(n10007) );
  OAI21_X1 U12104 ( .B1(n15927), .B2(n17235), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10008) );
  NOR2_X1 U12105 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15406), .ZN(
        n15926) );
  AND2_X1 U12106 ( .A1(n15356), .A2(n9715), .ZN(n17104) );
  NOR2_X1 U12107 ( .A1(n17129), .A2(n17480), .ZN(n17109) );
  NAND2_X1 U12108 ( .A1(n17182), .A2(n10022), .ZN(n17129) );
  AND2_X1 U12109 ( .A1(n17475), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10022) );
  INV_X1 U12110 ( .A(n15356), .ZN(n17150) );
  OR3_X1 U12111 ( .A1(n17180), .A2(n17235), .A3(n17144), .ZN(n17163) );
  NOR2_X1 U12112 ( .A1(n17199), .A2(n15354), .ZN(n17193) );
  INV_X1 U12113 ( .A(n15353), .ZN(n15354) );
  AOI21_X1 U12114 ( .B1(n17200), .B2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n9843), .ZN(n15353) );
  AND2_X1 U12115 ( .A1(n17318), .A2(n17539), .ZN(n9843) );
  NAND2_X1 U12116 ( .A1(n17193), .A2(n17522), .ZN(n17192) );
  OR2_X1 U12117 ( .A1(n17310), .A2(n17507), .ZN(n17200) );
  INV_X1 U12118 ( .A(n17131), .ZN(n17548) );
  NOR2_X1 U12119 ( .A1(n17556), .A2(n17562), .ZN(n17533) );
  INV_X1 U12120 ( .A(n17239), .ZN(n17556) );
  OR2_X1 U12121 ( .A1(n17300), .A2(n9999), .ZN(n17253) );
  NAND2_X1 U12122 ( .A1(n10000), .A2(n17591), .ZN(n9999) );
  INV_X1 U12123 ( .A(n10001), .ZN(n10000) );
  NOR2_X1 U12124 ( .A1(n17300), .A2(n10001), .ZN(n17262) );
  NAND2_X1 U12125 ( .A1(n17320), .A2(n15347), .ZN(n17232) );
  INV_X1 U12126 ( .A(n15345), .ZN(n15342) );
  NAND2_X1 U12127 ( .A1(n17342), .A2(n15340), .ZN(n17333) );
  NOR2_X1 U12128 ( .A1(n17333), .A2(n17334), .ZN(n17332) );
  XNOR2_X1 U12129 ( .A(n15316), .B(n10016), .ZN(n17329) );
  INV_X1 U12130 ( .A(n15317), .ZN(n10016) );
  NAND2_X1 U12131 ( .A1(n17329), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17328) );
  XNOR2_X1 U12132 ( .A(n15339), .B(n9800), .ZN(n17343) );
  INV_X1 U12133 ( .A(n15338), .ZN(n9800) );
  NAND2_X1 U12134 ( .A1(n17364), .A2(n15336), .ZN(n17350) );
  NAND2_X1 U12135 ( .A1(n17350), .A2(n17351), .ZN(n17349) );
  NAND2_X1 U12136 ( .A1(n9798), .A2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n15332) );
  INV_X1 U12137 ( .A(n9799), .ZN(n9798) );
  NOR2_X1 U12138 ( .A1(n15212), .A2(n15211), .ZN(n15980) );
  XNOR2_X1 U12139 ( .A(n15297), .B(n15296), .ZN(n17391) );
  XNOR2_X1 U12140 ( .A(n9799), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n17388) );
  XNOR2_X1 U12141 ( .A(n16930), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17399) );
  NAND2_X1 U12142 ( .A1(n17406), .A2(n17399), .ZN(n17398) );
  INV_X1 U12143 ( .A(n18218), .ZN(n18185) );
  NOR2_X1 U12144 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n17734), .ZN(n18037) );
  NOR2_X1 U12145 ( .A1(n13581), .A2(n13580), .ZN(n17754) );
  NOR2_X1 U12146 ( .A1(n13591), .A2(n13590), .ZN(n17760) );
  INV_X1 U12147 ( .A(n15206), .ZN(n17772) );
  INV_X1 U12148 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18228) );
  CLKBUF_X1 U12149 ( .A(n14610), .Z(n14633) );
  NAND2_X1 U12150 ( .A1(n12642), .A2(n12412), .ZN(n20550) );
  INV_X1 U12151 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n19654) );
  INV_X1 U12152 ( .A(n19653), .ZN(n19678) );
  XNOR2_X1 U12153 ( .A(n13889), .B(n13888), .ZN(n14220) );
  NAND2_X2 U12154 ( .A1(n12653), .A2(n12652), .ZN(n19710) );
  OR2_X1 U12155 ( .A1(n12651), .A2(n13886), .ZN(n12652) );
  INV_X1 U12156 ( .A(n14025), .ZN(n19705) );
  INV_X1 U12157 ( .A(n19710), .ZN(n14004) );
  INV_X1 U12158 ( .A(n14097), .ZN(n14028) );
  INV_X1 U12159 ( .A(n14063), .ZN(n14069) );
  AND2_X1 U12160 ( .A1(n19713), .A2(n12901), .ZN(n15544) );
  INV_X1 U12161 ( .A(n15544), .ZN(n19712) );
  BUF_X1 U12162 ( .A(n19736), .Z(n19746) );
  OR2_X1 U12163 ( .A1(n19773), .A2(n19853), .ZN(n12957) );
  AND2_X1 U12164 ( .A1(n12276), .A2(n10203), .ZN(n11245) );
  AND2_X1 U12165 ( .A1(n10205), .A2(n10204), .ZN(n10203) );
  XOR2_X1 U12166 ( .A(n13906), .B(n13905), .Z(n14097) );
  INV_X1 U12167 ( .A(n13916), .ZN(n12277) );
  INV_X1 U12168 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14158) );
  INV_X1 U12169 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15487) );
  INV_X1 U12170 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15498) );
  NAND2_X1 U12171 ( .A1(n12989), .A2(n12990), .ZN(n12972) );
  AND2_X1 U12172 ( .A1(n12939), .A2(n20547), .ZN(n19787) );
  INV_X1 U12173 ( .A(n14190), .ZN(n19782) );
  NAND2_X1 U12174 ( .A1(n10264), .A2(n11133), .ZN(n13432) );
  NAND2_X1 U12175 ( .A1(n15591), .A2(n11106), .ZN(n15588) );
  NOR2_X1 U12176 ( .A1(n19827), .A2(n19828), .ZN(n9775) );
  NOR2_X1 U12177 ( .A1(n19795), .A2(n13559), .ZN(n19816) );
  NAND2_X1 U12178 ( .A1(n12717), .A2(n12712), .ZN(n15609) );
  INV_X1 U12179 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20262) );
  NOR2_X1 U12180 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12614) );
  OAI22_X1 U12181 ( .A1(n19930), .A2(n19929), .B1(n20172), .B2(n20055), .ZN(
        n19953) );
  NAND2_X1 U12182 ( .A1(n19958), .A2(n19894), .ZN(n19957) );
  OAI21_X1 U12183 ( .B1(n19969), .B2(n19968), .A(n19967), .ZN(n19990) );
  OAI21_X1 U12184 ( .B1(n20016), .B2(n20001), .A(n20353), .ZN(n20019) );
  OAI211_X1 U12185 ( .C1(n20140), .C2(n20270), .A(n20180), .B(n20125), .ZN(
        n20143) );
  OR2_X1 U12186 ( .A1(n20223), .A2(n20314), .ZN(n20198) );
  OAI211_X1 U12187 ( .C1(n20376), .C2(n20354), .A(n20353), .B(n20352), .ZN(
        n20379) );
  INV_X1 U12188 ( .A(n20263), .ZN(n20385) );
  INV_X1 U12189 ( .A(n20274), .ZN(n20386) );
  INV_X1 U12190 ( .A(n20275), .ZN(n20396) );
  INV_X1 U12191 ( .A(n20280), .ZN(n20402) );
  INV_X1 U12192 ( .A(n20284), .ZN(n20403) );
  INV_X1 U12193 ( .A(n20285), .ZN(n20408) );
  INV_X1 U12194 ( .A(n20289), .ZN(n20409) );
  INV_X1 U12195 ( .A(n20290), .ZN(n20414) );
  INV_X1 U12196 ( .A(n20295), .ZN(n20420) );
  INV_X1 U12197 ( .A(n20299), .ZN(n20421) );
  INV_X1 U12198 ( .A(n20300), .ZN(n20428) );
  INV_X1 U12199 ( .A(n20304), .ZN(n20429) );
  OR2_X1 U12200 ( .A1(n20389), .A2(n20222), .ZN(n20443) );
  INV_X1 U12201 ( .A(n20312), .ZN(n20436) );
  NAND2_X1 U12202 ( .A1(n11206), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n19602) );
  INV_X2 U12203 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20448) );
  INV_X1 U12204 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20445) );
  NOR2_X1 U12205 ( .A1(n15759), .A2(n15760), .ZN(n15758) );
  NOR2_X1 U12206 ( .A1(n15766), .A2(n18630), .ZN(n15759) );
  AND2_X1 U12207 ( .A1(n10121), .A2(n15696), .ZN(n12251) );
  NAND2_X1 U12208 ( .A1(n15690), .A2(n12213), .ZN(n18614) );
  NAND2_X1 U12209 ( .A1(n13746), .A2(n10072), .ZN(n13759) );
  INV_X1 U12210 ( .A(n18637), .ZN(n18616) );
  AND2_X1 U12211 ( .A1(n12401), .A2(n12211), .ZN(n18625) );
  OR2_X1 U12212 ( .A1(n11528), .A2(n11527), .ZN(n13036) );
  NOR2_X1 U12213 ( .A1(n11518), .A2(n11517), .ZN(n13031) );
  NAND2_X1 U12214 ( .A1(n11504), .A2(n11503), .ZN(n13030) );
  NOR2_X1 U12215 ( .A1(n11762), .A2(n11747), .ZN(n12724) );
  AOI21_X1 U12216 ( .B1(n11462), .B2(n11465), .A(n11464), .ZN(n11466) );
  INV_X1 U12217 ( .A(n14522), .ZN(n14550) );
  XNOR2_X1 U12218 ( .A(n9957), .B(n14460), .ZN(n14562) );
  OAI21_X1 U12219 ( .B1(n14476), .B2(n14467), .A(n14469), .ZN(n9957) );
  INV_X1 U12220 ( .A(n15778), .ZN(n14611) );
  NAND2_X1 U12221 ( .A1(n14506), .A2(n9645), .ZN(n14500) );
  AND2_X1 U12222 ( .A1(n13199), .A2(n14633), .ZN(n18651) );
  AND2_X1 U12223 ( .A1(n13199), .A2(n14634), .ZN(n18652) );
  INV_X1 U12224 ( .A(n18692), .ZN(n18687) );
  INV_X1 U12225 ( .A(n19566), .ZN(n19128) );
  NAND2_X1 U12226 ( .A1(n12628), .A2(n18699), .ZN(n18691) );
  OR2_X1 U12227 ( .A1(n12783), .A2(n12627), .ZN(n12628) );
  INV_X1 U12228 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14742) );
  INV_X1 U12229 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18456) );
  INV_X1 U12230 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n20697) );
  NAND2_X1 U12231 ( .A1(n9908), .A2(n9906), .ZN(n15796) );
  AOI21_X1 U12232 ( .B1(n18525), .B2(n18830), .A(n9924), .ZN(n9923) );
  OAI21_X1 U12233 ( .B1(n18816), .B2(n14813), .A(n9925), .ZN(n9924) );
  INV_X1 U12234 ( .A(n14814), .ZN(n9925) );
  INV_X1 U12235 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n18541) );
  INV_X1 U12236 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n15824) );
  INV_X1 U12237 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n15853) );
  NAND2_X1 U12238 ( .A1(n18418), .A2(n12460), .ZN(n15852) );
  AND2_X1 U12239 ( .A1(n15852), .A2(n12472), .ZN(n18829) );
  INV_X1 U12240 ( .A(n14440), .ZN(n13221) );
  XNOR2_X1 U12241 ( .A(n9932), .B(n9688), .ZN(n14660) );
  NAND2_X1 U12242 ( .A1(n9934), .A2(n9933), .ZN(n9932) );
  NOR2_X1 U12243 ( .A1(n12268), .A2(n12269), .ZN(n14595) );
  OAI21_X1 U12244 ( .B1(n14917), .B2(n14915), .A(n14914), .ZN(n14725) );
  XNOR2_X1 U12245 ( .A(n9895), .B(n9726), .ZN(n14931) );
  NAND2_X1 U12246 ( .A1(n9896), .A2(n9929), .ZN(n9895) );
  NAND2_X1 U12247 ( .A1(n14752), .A2(n14750), .ZN(n9896) );
  NAND2_X1 U12248 ( .A1(n9899), .A2(n9902), .ZN(n14803) );
  NAND2_X1 U12249 ( .A1(n9908), .A2(n9904), .ZN(n9899) );
  NAND2_X1 U12250 ( .A1(n9873), .A2(n9874), .ZN(n14811) );
  INV_X1 U12251 ( .A(n14812), .ZN(n15017) );
  NAND2_X1 U12252 ( .A1(n10245), .A2(n10246), .ZN(n15804) );
  NAND2_X1 U12253 ( .A1(n10248), .A2(n9686), .ZN(n10245) );
  AND2_X1 U12254 ( .A1(n10247), .A2(n10250), .ZN(n15027) );
  NAND2_X1 U12255 ( .A1(n13363), .A2(n13362), .ZN(n13365) );
  NAND2_X1 U12256 ( .A1(n10181), .A2(n9756), .ZN(n18632) );
  INV_X1 U12257 ( .A(n18839), .ZN(n18868) );
  OAI21_X1 U12258 ( .B1(n13345), .B2(n12224), .A(n13332), .ZN(n15847) );
  INV_X1 U12259 ( .A(n15898), .ZN(n18875) );
  INV_X1 U12260 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19560) );
  INV_X1 U12261 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19550) );
  NAND2_X1 U12262 ( .A1(n19586), .A2(n19535), .ZN(n19533) );
  NOR2_X1 U12263 ( .A1(n12980), .A2(n12087), .ZN(n13018) );
  INV_X1 U12264 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15419) );
  INV_X1 U12265 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13713) );
  INV_X1 U12266 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n13706) );
  XNOR2_X1 U12267 ( .A(n9954), .B(n12528), .ZN(n19557) );
  INV_X1 U12268 ( .A(n11416), .ZN(n9954) );
  AND2_X1 U12269 ( .A1(n18959), .A2(n19536), .ZN(n19007) );
  INV_X1 U12270 ( .A(n19007), .ZN(n19018) );
  OAI21_X1 U12271 ( .B1(n19028), .B2(n19043), .A(n19027), .ZN(n19046) );
  OR3_X1 U12272 ( .A1(n13188), .A2(n13189), .A3(n19104), .ZN(n19096) );
  AND2_X1 U12273 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n11457), .ZN(
        n19135) );
  OR2_X1 U12274 ( .A1(n19292), .A2(n19159), .ZN(n19190) );
  INV_X1 U12275 ( .A(n19383), .ZN(n19303) );
  INV_X1 U12276 ( .A(n19432), .ZN(n19325) );
  INV_X1 U12277 ( .A(n19366), .ZN(n19356) );
  OAI21_X1 U12278 ( .B1(n19343), .B2(n19342), .A(n19341), .ZN(n19362) );
  OR2_X1 U12279 ( .A1(n19292), .A2(n19297), .ZN(n19366) );
  OAI22_X1 U12280 ( .A1(n18894), .A2(n18917), .B1(n18893), .B2(n18915), .ZN(
        n19386) );
  OAI22_X1 U12281 ( .A1(n18899), .A2(n18917), .B1(n20604), .B2(n18915), .ZN(
        n19392) );
  INV_X1 U12282 ( .A(n19315), .ZN(n19398) );
  INV_X1 U12283 ( .A(n19431), .ZN(n19411) );
  INV_X1 U12284 ( .A(n19283), .ZN(n19410) );
  OR2_X1 U12285 ( .A1(n19331), .A2(n19373), .ZN(n19431) );
  INV_X1 U12286 ( .A(n19414), .ZN(n19427) );
  INV_X1 U12287 ( .A(n18416), .ZN(n18699) );
  NAND2_X1 U12288 ( .A1(n12434), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19525) );
  INV_X1 U12289 ( .A(n12839), .ZN(n12434) );
  NAND2_X1 U12290 ( .A1(n18231), .A2(n18235), .ZN(n16095) );
  XNOR2_X1 U12291 ( .A(n16151), .B(n10084), .ZN(n10083) );
  INV_X1 U12292 ( .A(n16152), .ZN(n10084) );
  OR2_X1 U12293 ( .A1(n16153), .A2(n10082), .ZN(n10081) );
  AND2_X1 U12294 ( .A1(n16163), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n10082) );
  INV_X1 U12295 ( .A(n10085), .ZN(n16159) );
  NOR2_X1 U12296 ( .A1(n16191), .A2(n17075), .ZN(n16190) );
  NOR2_X1 U12297 ( .A1(n16201), .A2(n10079), .ZN(n16191) );
  NAND2_X1 U12298 ( .A1(n16238), .A2(n10105), .ZN(n10101) );
  NOR2_X1 U12299 ( .A1(n18305), .A2(n16254), .ZN(n16241) );
  NAND2_X1 U12300 ( .A1(n17155), .A2(n10077), .ZN(n10076) );
  AND2_X1 U12301 ( .A1(n10080), .A2(n10073), .ZN(n16246) );
  INV_X1 U12302 ( .A(n10080), .ZN(n16255) );
  NOR2_X1 U12303 ( .A1(n16138), .A2(n16303), .ZN(n16269) );
  NOR2_X1 U12304 ( .A1(n9609), .A2(n10075), .ZN(n16285) );
  AND2_X1 U12305 ( .A1(n16294), .A2(n16478), .ZN(n10075) );
  INV_X1 U12306 ( .A(n10074), .ZN(n16284) );
  INV_X1 U12307 ( .A(n16291), .ZN(n16303) );
  NOR2_X1 U12308 ( .A1(n16137), .A2(n16353), .ZN(n16335) );
  NOR2_X1 U12309 ( .A1(n17226), .A2(n17313), .ZN(n16343) );
  NOR2_X1 U12310 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n16407), .ZN(n16387) );
  INV_X1 U12311 ( .A(n16482), .ZN(n16469) );
  INV_X1 U12312 ( .A(n16481), .ZN(n16466) );
  INV_X1 U12313 ( .A(n16477), .ZN(n16479) );
  NOR2_X1 U12314 ( .A1(n16577), .A2(n16578), .ZN(n16552) );
  NOR2_X1 U12315 ( .A1(n16890), .A2(n16602), .ZN(n16589) );
  NAND2_X1 U12316 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n16618), .ZN(n16602) );
  NOR2_X1 U12317 ( .A1(n16647), .A2(n16660), .ZN(n16632) );
  NAND2_X1 U12318 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n16632), .ZN(n16631) );
  NAND2_X1 U12319 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n16676), .ZN(n16660) );
  INV_X1 U12320 ( .A(n16748), .ZN(n16731) );
  NAND2_X1 U12321 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n16762), .ZN(n16753) );
  INV_X1 U12322 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n16756) );
  NAND2_X1 U12323 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n16770), .ZN(n16763) );
  NAND2_X1 U12324 ( .A1(P3_EBX_REG_1__SCAN_IN), .A2(n16777), .ZN(n16766) );
  NOR2_X2 U12325 ( .A1(n16767), .A2(n16766), .ZN(n16770) );
  INV_X1 U12326 ( .A(P3_EAX_REG_31__SCAN_IN), .ZN(n9785) );
  NAND2_X1 U12327 ( .A1(n16798), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n16795) );
  NOR2_X1 U12328 ( .A1(n16804), .A2(n17001), .ZN(n16798) );
  NAND2_X1 U12329 ( .A1(n16807), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n16804) );
  NOR2_X1 U12330 ( .A1(n16813), .A2(n16997), .ZN(n16807) );
  NAND2_X1 U12331 ( .A1(n16858), .A2(n9786), .ZN(n16819) );
  AND2_X1 U12332 ( .A1(n16781), .A2(n9770), .ZN(n9786) );
  NOR2_X1 U12333 ( .A1(n16985), .A2(n16845), .ZN(n16840) );
  NOR2_X1 U12334 ( .A1(n16863), .A2(n16979), .ZN(n16858) );
  NOR2_X1 U12335 ( .A1(n15236), .A2(n15235), .ZN(n16910) );
  NOR2_X1 U12336 ( .A1(n15256), .A2(n10021), .ZN(n10020) );
  NOR2_X1 U12337 ( .A1(n10019), .A2(n10018), .ZN(n10017) );
  INV_X1 U12338 ( .A(n16931), .ZN(n16924) );
  INV_X1 U12339 ( .A(n16932), .ZN(n16927) );
  AOI21_X1 U12340 ( .B1(n15422), .B2(n18235), .A(n15421), .ZN(n16929) );
  NOR2_X1 U12341 ( .A1(n18187), .A2(n16929), .ZN(n16931) );
  NOR2_X1 U12342 ( .A1(n18386), .A2(n16953), .ZN(n16963) );
  CLKBUF_X1 U12343 ( .A(n16963), .Z(n16970) );
  NOR2_X1 U12344 ( .A1(n17741), .A2(n17037), .ZN(n17030) );
  AOI21_X1 U12346 ( .B1(n15955), .B2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n9839), .ZN(n9838) );
  AOI21_X1 U12347 ( .B1(n15976), .B2(n20668), .A(n15956), .ZN(n9839) );
  INV_X1 U12348 ( .A(n17061), .ZN(n15977) );
  INV_X1 U12349 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17086) );
  NAND2_X1 U12350 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17228) );
  INV_X1 U12351 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17353) );
  NOR2_X1 U12352 ( .A1(n17396), .A2(n17044), .ZN(n17367) );
  NOR2_X1 U12353 ( .A1(n17352), .A2(n17353), .ZN(n17354) );
  NOR2_X2 U12354 ( .A1(n18035), .A2(n17896), .ZN(n18121) );
  OAI21_X1 U12355 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18388), .A(n16095), 
        .ZN(n17408) );
  NAND2_X1 U12356 ( .A1(n15405), .A2(n15406), .ZN(n15362) );
  AND2_X1 U12357 ( .A1(n15360), .A2(n15361), .ZN(n17061) );
  NOR2_X2 U12358 ( .A1(n15361), .A2(n15360), .ZN(n17060) );
  INV_X1 U12359 ( .A(n15291), .ZN(n15985) );
  OAI21_X1 U12360 ( .B1(n17420), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n17716), .ZN(n9793) );
  OAI21_X1 U12361 ( .B1(n17421), .B2(n17636), .A(n9790), .ZN(n9789) );
  AOI21_X1 U12362 ( .B1(n17699), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n9769), .ZN(n9790) );
  NAND2_X1 U12363 ( .A1(n9797), .A2(n9795), .ZN(n17424) );
  AOI21_X1 U12364 ( .B1(n17414), .B2(n17472), .A(n9796), .ZN(n9795) );
  NAND2_X1 U12365 ( .A1(n17415), .A2(n18217), .ZN(n9797) );
  AND2_X1 U12366 ( .A1(n9841), .A2(n10023), .ZN(n17077) );
  INV_X1 U12367 ( .A(n17200), .ZN(n17541) );
  INV_X1 U12368 ( .A(n17586), .ZN(n17597) );
  OR2_X1 U12369 ( .A1(n17300), .A2(n10004), .ZN(n17271) );
  NAND2_X1 U12370 ( .A1(n18185), .A2(n18202), .ZN(n17610) );
  NOR2_X1 U12371 ( .A1(n17300), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17283) );
  AND2_X1 U12372 ( .A1(n9691), .A2(n9835), .ZN(n17341) );
  NOR2_X1 U12373 ( .A1(n17710), .A2(n17716), .ZN(n17699) );
  INV_X1 U12374 ( .A(n15980), .ZN(n18224) );
  NOR2_X1 U12375 ( .A1(n18224), .A2(n17680), .ZN(n17721) );
  INV_X1 U12376 ( .A(n18190), .ZN(n18202) );
  INV_X1 U12377 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18209) );
  INV_X1 U12378 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18196) );
  INV_X1 U12379 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18339) );
  NAND2_X1 U12380 ( .A1(n20637), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18401) );
  AND2_X1 U12381 ( .A1(n11267), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n19836)
         );
  OR4_X1 U12383 ( .A1(n12393), .A2(n12392), .A3(n12391), .A4(n12390), .ZN(
        P1_U2813) );
  OAI21_X1 U12384 ( .B1(n14267), .B2(n19608), .A(n9824), .ZN(P1_U2970) );
  NOR2_X1 U12385 ( .A1(n9825), .A2(n9700), .ZN(n9824) );
  INV_X1 U12386 ( .A(n11217), .ZN(n9825) );
  NAND2_X1 U12387 ( .A1(n12876), .A2(n9774), .ZN(n12881) );
  AND2_X1 U12388 ( .A1(n9975), .A2(n9973), .ZN(n9892) );
  NOR3_X1 U12389 ( .A1(n14250), .A2(n14249), .A3(n14248), .ZN(n9975) );
  OAI21_X1 U12390 ( .B1(n14283), .B2(n19820), .A(n9997), .ZN(P1_U3004) );
  NOR2_X1 U12391 ( .A1(n14284), .A2(n9998), .ZN(n9997) );
  NOR2_X1 U12392 ( .A1(n14279), .A2(n14268), .ZN(n9998) );
  INV_X1 U12393 ( .A(n10193), .ZN(n20525) );
  AOI211_X1 U12394 ( .C1(n9772), .C2(P2_REIP_REG_0__SCAN_IN), .A(n14445), .B(
        n14444), .ZN(n14448) );
  OAI21_X1 U12395 ( .B1(n14656), .B2(n14548), .A(n11959), .ZN(n11960) );
  INV_X1 U12396 ( .A(n11551), .ZN(n13117) );
  NAND2_X1 U12397 ( .A1(n10211), .A2(n10055), .ZN(n10054) );
  NAND2_X1 U12398 ( .A1(n14837), .A2(n18821), .ZN(n10163) );
  NAND2_X1 U12399 ( .A1(n9926), .A2(n9921), .ZN(P2_U3001) );
  INV_X1 U12400 ( .A(n9922), .ZN(n9921) );
  NAND2_X1 U12401 ( .A1(n14812), .A2(n18821), .ZN(n9926) );
  OAI21_X1 U12402 ( .B1(n15022), .B2(n18833), .A(n9923), .ZN(n9922) );
  NAND2_X1 U12403 ( .A1(n10209), .A2(n10211), .ZN(n10208) );
  NAND2_X1 U12404 ( .A1(n14837), .A2(n18849), .ZN(n9970) );
  INV_X1 U12405 ( .A(n9879), .ZN(n15000) );
  OAI21_X1 U12406 ( .B1(n14996), .B2(n20666), .A(n9880), .ZN(n9879) );
  AOI21_X1 U12407 ( .B1(n14998), .B2(n14999), .A(n14997), .ZN(n9880) );
  AOI21_X1 U12408 ( .B1(n16782), .B2(P3_EAX_REG_30__SCAN_IN), .A(n9784), .ZN(
        n16783) );
  AOI21_X1 U12409 ( .B1(n16788), .B2(n9753), .A(n9785), .ZN(n9784) );
  AOI21_X1 U12410 ( .B1(n15965), .B2(n17293), .A(n9701), .ZN(n15929) );
  NAND2_X1 U12411 ( .A1(n9840), .A2(n9836), .ZN(P3_U2801) );
  NOR2_X1 U12412 ( .A1(n15954), .A2(n9837), .ZN(n9836) );
  NAND2_X1 U12413 ( .A1(n15951), .A2(n17293), .ZN(n9840) );
  OAI21_X1 U12414 ( .B1(n15952), .B2(n15953), .A(n9838), .ZN(n9837) );
  NAND2_X1 U12415 ( .A1(n17124), .A2(n10287), .ZN(n17115) );
  AOI21_X1 U12416 ( .B1(n15965), .B2(n17613), .A(n15964), .ZN(n15966) );
  NAND2_X1 U12417 ( .A1(n9791), .A2(n9788), .ZN(P3_U2835) );
  NAND2_X1 U12418 ( .A1(n9794), .A2(n9792), .ZN(n9791) );
  INV_X1 U12419 ( .A(n9789), .ZN(n9788) );
  INV_X1 U12420 ( .A(n9793), .ZN(n9792) );
  OR2_X2 U12421 ( .A1(n13574), .A2(n13575), .ZN(n9679) );
  CLKBUF_X3 U12422 ( .A(n15097), .Z(n16721) );
  NAND2_X1 U12423 ( .A1(n10162), .A2(n11275), .ZN(n11291) );
  OR2_X1 U12424 ( .A1(n14514), .A2(n11700), .ZN(n9645) );
  AND2_X1 U12425 ( .A1(n10287), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9646) );
  AND2_X2 U12426 ( .A1(n12915), .A2(n14427), .ZN(n10575) );
  NAND4_X2 U12427 ( .A1(n12152), .A2(n12151), .A3(n12150), .A4(n12149), .ZN(
        n12224) );
  AND2_X1 U12428 ( .A1(n11504), .A2(n9669), .ZN(n9647) );
  AND2_X1 U12429 ( .A1(n9669), .A2(n13036), .ZN(n9648) );
  INV_X1 U12430 ( .A(n9609), .ZN(n10073) );
  INV_X1 U12431 ( .A(n15054), .ZN(n10248) );
  OR2_X1 U12432 ( .A1(n12268), .A2(n9752), .ZN(n9649) );
  OR3_X2 U12433 ( .A1(n15855), .A2(n9723), .A3(n10182), .ZN(n9650) );
  AND2_X1 U12434 ( .A1(n19863), .A2(n19853), .ZN(n9692) );
  NAND2_X1 U12435 ( .A1(n11996), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11993) );
  NAND2_X1 U12436 ( .A1(n11996), .A2(n10130), .ZN(n11991) );
  NOR2_X1 U12437 ( .A1(n11987), .A2(n18518), .ZN(n11988) );
  OR2_X1 U12438 ( .A1(n14092), .A2(n10257), .ZN(n9651) );
  INV_X1 U12439 ( .A(n15834), .ZN(n10170) );
  NOR2_X1 U12440 ( .A1(n14074), .A2(n14022), .ZN(n13956) );
  OR2_X1 U12441 ( .A1(n13982), .A2(n9976), .ZN(n9653) );
  AND2_X1 U12442 ( .A1(n10649), .A2(n9849), .ZN(n9654) );
  AND2_X1 U12443 ( .A1(n9987), .A2(n13399), .ZN(n9655) );
  NAND2_X1 U12444 ( .A1(n15025), .A2(n15030), .ZN(n9656) );
  AND2_X1 U12445 ( .A1(n15572), .A2(n11134), .ZN(n9657) );
  AND4_X1 U12446 ( .A1(n14762), .A2(n14790), .A3(n13804), .A4(n14771), .ZN(
        n9658) );
  OR3_X1 U12447 ( .A1(n14537), .A2(n10045), .A3(n10048), .ZN(n9659) );
  NOR2_X1 U12448 ( .A1(n15700), .A2(n18839), .ZN(n9660) );
  AND2_X1 U12449 ( .A1(n13364), .A2(n9702), .ZN(n9661) );
  NAND2_X1 U12450 ( .A1(n19886), .A2(n10395), .ZN(n9662) );
  AND2_X1 U12451 ( .A1(n10180), .A2(n13370), .ZN(n9663) );
  NOR3_X1 U12452 ( .A1(n15770), .A2(n13327), .A3(n13827), .ZN(n9664) );
  AND2_X1 U12453 ( .A1(n18926), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9665) );
  OR2_X1 U12454 ( .A1(n15572), .A2(n11134), .ZN(n9666) );
  AND2_X1 U12455 ( .A1(n10619), .A2(n10640), .ZN(n9667) );
  AOI21_X1 U12456 ( .B1(n16201), .B2(n10099), .A(n10096), .ZN(n10094) );
  AND2_X1 U12457 ( .A1(n9654), .A2(n9848), .ZN(n9668) );
  AND2_X2 U12458 ( .A1(n12918), .A2(n14427), .ZN(n10551) );
  NAND2_X2 U12459 ( .A1(n12629), .A2(n12008), .ZN(n12103) );
  INV_X1 U12460 ( .A(n12980), .ZN(n10181) );
  NOR2_X1 U12461 ( .A1(n11987), .A2(n10124), .ZN(n11985) );
  INV_X1 U12462 ( .A(n14749), .ZN(n9929) );
  NAND2_X1 U12463 ( .A1(n11978), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11977) );
  NAND2_X1 U12464 ( .A1(n12667), .A2(n10153), .ZN(n12766) );
  INV_X1 U12465 ( .A(n10192), .ZN(n20117) );
  AND2_X1 U12466 ( .A1(n10155), .A2(n11503), .ZN(n9669) );
  AND2_X1 U12467 ( .A1(n10135), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9670) );
  NAND2_X1 U12468 ( .A1(n11983), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11982) );
  INV_X1 U12469 ( .A(n10154), .ZN(n13035) );
  OR3_X1 U12470 ( .A1(n14021), .A2(n9982), .A3(n9985), .ZN(n9671) );
  NAND2_X1 U12471 ( .A1(n9648), .A2(n13053), .ZN(n9672) );
  OR3_X1 U12472 ( .A1(n11700), .A2(n14496), .A3(n11699), .ZN(n9673) );
  AND2_X1 U12473 ( .A1(n9758), .A2(n12266), .ZN(n9674) );
  AND2_X1 U12474 ( .A1(n9977), .A2(n13922), .ZN(n9675) );
  AND2_X1 U12475 ( .A1(n10063), .A2(n14493), .ZN(n9676) );
  NAND2_X1 U12476 ( .A1(n11743), .A2(n14482), .ZN(n9677) );
  AND2_X1 U12477 ( .A1(n10172), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9678) );
  NOR2_X1 U12478 ( .A1(n16465), .A2(n13700), .ZN(n16624) );
  OR2_X1 U12479 ( .A1(n14503), .A2(n10039), .ZN(n9681) );
  OR2_X1 U12480 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n13836), .ZN(n9682) );
  AND2_X1 U12481 ( .A1(n12255), .A2(n10063), .ZN(n9684) );
  NOR2_X2 U12482 ( .A1(n16902), .A2(n17411), .ZN(n17293) );
  AND2_X1 U12483 ( .A1(n11996), .A2(n10133), .ZN(n11994) );
  INV_X1 U12484 ( .A(n13546), .ZN(n9915) );
  INV_X1 U12485 ( .A(n11291), .ZN(n11298) );
  AND2_X1 U12486 ( .A1(n15040), .A2(n10249), .ZN(n9685) );
  AND2_X1 U12487 ( .A1(n9656), .A2(n9685), .ZN(n9686) );
  INV_X1 U12488 ( .A(n10523), .ZN(n9890) );
  AND2_X1 U12489 ( .A1(n13942), .A2(n13985), .ZN(n13977) );
  AND2_X1 U12490 ( .A1(n10144), .A2(n10142), .ZN(n9687) );
  INV_X1 U12491 ( .A(n19837), .ZN(n19994) );
  NOR2_X1 U12492 ( .A1(n14993), .A2(n14981), .ZN(n14987) );
  INV_X1 U12493 ( .A(n14987), .ZN(n9884) );
  AND2_X1 U12494 ( .A1(n13854), .A2(n14643), .ZN(n9688) );
  AND2_X1 U12495 ( .A1(n11995), .A2(n11963), .ZN(n11996) );
  OR3_X1 U12496 ( .A1(n12268), .A2(n10184), .A3(n10186), .ZN(n9689) );
  AND2_X1 U12497 ( .A1(n10221), .A2(n10215), .ZN(n9690) );
  OR2_X1 U12498 ( .A1(n17356), .A2(n17357), .ZN(n9691) );
  OR2_X1 U12499 ( .A1(n16976), .A2(n17741), .ZN(n9693) );
  AND2_X1 U12500 ( .A1(n9904), .A2(n14800), .ZN(n9694) );
  INV_X1 U12501 ( .A(n19839), .ZN(n12485) );
  AND2_X1 U12502 ( .A1(n10148), .A2(n10147), .ZN(n9695) );
  AND2_X1 U12503 ( .A1(n12631), .A2(n12540), .ZN(n9696) );
  AND2_X1 U12504 ( .A1(n10478), .A2(n9890), .ZN(n9697) );
  AND2_X1 U12505 ( .A1(n14825), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9698) );
  NOR3_X1 U12506 ( .A1(n13982), .A2(n13722), .A3(n9976), .ZN(n9978) );
  NOR3_X1 U12507 ( .A1(n14537), .A2(n10045), .A3(n9754), .ZN(n10047) );
  OR2_X1 U12508 ( .A1(n14074), .A2(n10196), .ZN(n9699) );
  NAND2_X1 U12509 ( .A1(n11440), .A2(n11439), .ZN(n12658) );
  NOR2_X1 U12510 ( .A1(n13737), .A2(n19835), .ZN(n9700) );
  AND2_X1 U12511 ( .A1(n15959), .A2(n17309), .ZN(n9701) );
  AND2_X1 U12512 ( .A1(n13859), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9702) );
  AND4_X1 U12513 ( .A1(n15255), .A2(n15254), .A3(n15253), .A4(n15252), .ZN(
        n9703) );
  NOR2_X1 U12514 ( .A1(n10244), .A2(n15802), .ZN(n10243) );
  NOR2_X1 U12515 ( .A1(n11768), .A2(n11767), .ZN(n14467) );
  AND2_X1 U12516 ( .A1(n13769), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9704) );
  AND2_X1 U12517 ( .A1(n13977), .A2(n9852), .ZN(n12276) );
  OR2_X1 U12518 ( .A1(n15572), .A2(n9993), .ZN(n9705) );
  OR2_X1 U12519 ( .A1(n9698), .A2(n10035), .ZN(n9706) );
  AND2_X1 U12520 ( .A1(n15586), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9707) );
  AND2_X1 U12521 ( .A1(n10601), .A2(n10619), .ZN(n9708) );
  AND2_X1 U12522 ( .A1(n10601), .A2(n9667), .ZN(n9709) );
  NOR2_X1 U12523 ( .A1(n13995), .A2(n13943), .ZN(n13942) );
  INV_X1 U12524 ( .A(n9875), .ZN(n9874) );
  NAND2_X1 U12525 ( .A1(n9876), .A2(n10241), .ZN(n9875) );
  AND2_X1 U12526 ( .A1(n19873), .A2(n19858), .ZN(n9710) );
  OR2_X1 U12527 ( .A1(n12536), .A2(n12005), .ZN(n9711) );
  AND2_X1 U12528 ( .A1(n14204), .A2(n13549), .ZN(n9712) );
  NAND2_X1 U12529 ( .A1(n14581), .A2(n10173), .ZN(n9713) );
  NOR2_X1 U12530 ( .A1(n10479), .A2(n20446), .ZN(n11124) );
  INV_X1 U12531 ( .A(n9992), .ZN(n9991) );
  NAND2_X1 U12532 ( .A1(n19886), .A2(n19853), .ZN(n9992) );
  INV_X1 U12533 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18518) );
  OR2_X1 U12534 ( .A1(n13764), .A2(n9704), .ZN(n9714) );
  OR2_X1 U12535 ( .A1(n15358), .A2(n10288), .ZN(n9715) );
  OR2_X1 U12537 ( .A1(n14675), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9716) );
  AND2_X1 U12538 ( .A1(n11342), .A2(n9952), .ZN(n9717) );
  AND2_X1 U12539 ( .A1(n11347), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9718) );
  AND2_X1 U12540 ( .A1(n11320), .A2(n9952), .ZN(n9719) );
  AND3_X1 U12541 ( .A1(n9833), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n9832), .ZN(n9720) );
  AND2_X1 U12542 ( .A1(n10117), .A2(n15696), .ZN(n9721) );
  AND2_X1 U12543 ( .A1(n12540), .A2(n11832), .ZN(n9722) );
  AND2_X2 U12544 ( .A1(n12918), .A2(n10290), .ZN(n10544) );
  XNOR2_X1 U12545 ( .A(n10517), .B(n10516), .ZN(n12938) );
  OR2_X1 U12546 ( .A1(n13195), .A2(n10160), .ZN(n13384) );
  NOR2_X1 U12547 ( .A1(n11989), .A2(n18541), .ZN(n11990) );
  AND2_X1 U12548 ( .A1(n11996), .A2(n10131), .ZN(n11992) );
  OR3_X1 U12549 ( .A1(n10183), .A2(n15856), .A3(n13198), .ZN(n9723) );
  AND2_X1 U12550 ( .A1(n15848), .A2(n9958), .ZN(n9724) );
  NAND2_X1 U12551 ( .A1(n14519), .A2(n14520), .ZN(n14513) );
  NOR2_X1 U12552 ( .A1(n11987), .A2(n10122), .ZN(n11983) );
  NAND2_X1 U12553 ( .A1(n13044), .A2(n13043), .ZN(n13042) );
  INV_X1 U12554 ( .A(n14740), .ZN(n9930) );
  NOR2_X1 U12555 ( .A1(n14621), .A2(n14620), .ZN(n9725) );
  INV_X1 U12556 ( .A(n13438), .ZN(n9966) );
  AND2_X1 U12557 ( .A1(n14535), .A2(n14526), .ZN(n14519) );
  AND2_X1 U12558 ( .A1(n9930), .A2(n14741), .ZN(n9726) );
  INV_X1 U12559 ( .A(n14914), .ZN(n9938) );
  NAND2_X2 U12560 ( .A1(n12287), .A2(n19839), .ZN(n12302) );
  OR2_X1 U12561 ( .A1(n11987), .A2(n10125), .ZN(n9727) );
  INV_X1 U12562 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17402) );
  NAND2_X1 U12563 ( .A1(n13331), .A2(n13357), .ZN(n13345) );
  OR3_X1 U12564 ( .A1(n15855), .A2(n10183), .A3(n15856), .ZN(n9728) );
  AND2_X1 U12565 ( .A1(n11716), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n9729) );
  NAND2_X1 U12566 ( .A1(n19878), .A2(n19886), .ZN(n12684) );
  INV_X1 U12567 ( .A(n12684), .ZN(n9818) );
  AND2_X1 U12568 ( .A1(n9863), .A2(n11550), .ZN(n9730) );
  NOR3_X1 U12569 ( .A1(n14021), .A2(n9982), .A3(n9980), .ZN(n9984) );
  NAND2_X1 U12570 ( .A1(n10650), .A2(n9654), .ZN(n9850) );
  AND2_X1 U12571 ( .A1(n11414), .A2(n19194), .ZN(n9731) );
  INV_X1 U12572 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20446) );
  OR2_X1 U12573 ( .A1(n11082), .A2(n10543), .ZN(n9732) );
  NAND2_X1 U12574 ( .A1(n13332), .A2(n15903), .ZN(n9733) );
  AND2_X1 U12575 ( .A1(n9655), .A2(n9986), .ZN(n9734) );
  NAND2_X1 U12576 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n16731), .ZN(n16730) );
  NAND2_X1 U12577 ( .A1(n11504), .A2(n9648), .ZN(n10154) );
  AND2_X1 U12578 ( .A1(n13501), .A2(n9741), .ZN(n13526) );
  INV_X1 U12579 ( .A(n14077), .ZN(n10780) );
  AND3_X1 U12580 ( .A1(n10779), .A2(n10778), .A3(n10777), .ZN(n14077) );
  OR2_X1 U12581 ( .A1(n15829), .A2(n15825), .ZN(n9735) );
  AND2_X1 U12582 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n9736) );
  OR2_X1 U12583 ( .A1(n11491), .A2(n11490), .ZN(n12907) );
  AND2_X1 U12584 ( .A1(n13775), .A2(n13774), .ZN(n9737) );
  AND2_X1 U12585 ( .A1(n13268), .A2(n13299), .ZN(n9738) );
  AND2_X1 U12586 ( .A1(n9644), .A2(n18926), .ZN(n9739) );
  AND2_X1 U12587 ( .A1(n10050), .A2(n10049), .ZN(n9740) );
  AND2_X1 U12588 ( .A1(n10199), .A2(n10198), .ZN(n9741) );
  AND2_X1 U12589 ( .A1(n10101), .A2(n10103), .ZN(n9742) );
  AND2_X1 U12590 ( .A1(n9776), .A2(n9775), .ZN(n9743) );
  AND2_X1 U12591 ( .A1(n10202), .A2(n10201), .ZN(n9744) );
  OR2_X1 U12592 ( .A1(n10103), .A2(n17112), .ZN(n9745) );
  INV_X1 U12593 ( .A(n13764), .ZN(n10250) );
  INV_X1 U12594 ( .A(n19820), .ZN(n19810) );
  OR3_X2 U12595 ( .A1(n18343), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(
        P3_STATE2_REG_0__SCAN_IN), .ZN(n9746) );
  INV_X1 U12596 ( .A(n18833), .ZN(n18808) );
  INV_X1 U12597 ( .A(n17075), .ZN(n10099) );
  NAND2_X1 U12598 ( .A1(n12667), .A2(n11468), .ZN(n12725) );
  NAND2_X1 U12599 ( .A1(n10028), .A2(n10027), .ZN(n10034) );
  AND2_X1 U12600 ( .A1(n12688), .A2(n15381), .ZN(n19788) );
  AND2_X1 U12601 ( .A1(n12667), .A2(n10151), .ZN(n12906) );
  NAND2_X1 U12602 ( .A1(n11974), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11971) );
  OR2_X1 U12603 ( .A1(n12593), .A2(n19573), .ZN(n18859) );
  AND2_X1 U12604 ( .A1(n11978), .A2(n10112), .ZN(n9748) );
  INV_X1 U12605 ( .A(n9949), .ZN(n12558) );
  XOR2_X1 U12606 ( .A(n18638), .B(n18844), .Z(n9749) );
  AND2_X1 U12607 ( .A1(n13149), .A2(n9987), .ZN(n9750) );
  NAND2_X1 U12608 ( .A1(n12871), .A2(n10534), .ZN(n12989) );
  AND2_X1 U12609 ( .A1(n10175), .A2(n14573), .ZN(n9751) );
  OR3_X1 U12610 ( .A1(n10184), .A2(n10186), .A3(n14586), .ZN(n9752) );
  OR2_X1 U12611 ( .A1(n16928), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n9753) );
  OR2_X1 U12612 ( .A1(n10048), .A2(n14510), .ZN(n9754) );
  AND2_X1 U12613 ( .A1(n11744), .A2(n14482), .ZN(n9755) );
  NAND2_X1 U12614 ( .A1(n12906), .A2(n12907), .ZN(n12964) );
  INV_X1 U12615 ( .A(n12964), .ZN(n11504) );
  NAND2_X1 U12616 ( .A1(n12906), .A2(n9730), .ZN(n13178) );
  INV_X1 U12617 ( .A(n13178), .ZN(n11562) );
  INV_X1 U12618 ( .A(n13767), .ZN(n13834) );
  AND2_X1 U12619 ( .A1(n13746), .A2(n9614), .ZN(n13767) );
  AND2_X1 U12620 ( .A1(n10177), .A2(n13017), .ZN(n9756) );
  AND2_X1 U12621 ( .A1(n9677), .A2(n11743), .ZN(n9757) );
  INV_X1 U12622 ( .A(n14483), .ZN(n10044) );
  NAND2_X2 U12623 ( .A1(n15979), .A2(n15985), .ZN(n17235) );
  NAND2_X1 U12624 ( .A1(n18911), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n9758) );
  INV_X1 U12625 ( .A(n10259), .ZN(n10258) );
  NOR2_X1 U12626 ( .A1(n9823), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10259) );
  AND2_X1 U12627 ( .A1(n9760), .A2(n11823), .ZN(n9759) );
  AND2_X1 U12628 ( .A1(n10149), .A2(n14469), .ZN(n9760) );
  INV_X1 U12629 ( .A(n10033), .ZN(n12733) );
  OAI211_X1 U12630 ( .C1(n10031), .C2(n11443), .A(n9652), .B(n10030), .ZN(
        n10033) );
  INV_X1 U12631 ( .A(n10179), .ZN(n18634) );
  AND2_X1 U12632 ( .A1(n10116), .A2(n15696), .ZN(n9761) );
  AND2_X1 U12633 ( .A1(n10127), .A2(n14718), .ZN(n9762) );
  AND2_X1 U12634 ( .A1(n10173), .A2(n12202), .ZN(n9763) );
  AND2_X1 U12635 ( .A1(n10034), .A2(n11885), .ZN(n9764) );
  AND2_X1 U12636 ( .A1(n11857), .A2(n18699), .ZN(n14540) );
  INV_X2 U12637 ( .A(n14540), .ZN(n14548) );
  INV_X1 U12638 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10109) );
  AND2_X1 U12639 ( .A1(n17124), .A2(n9646), .ZN(n9765) );
  INV_X1 U12640 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n10071) );
  AND2_X1 U12641 ( .A1(n17124), .A2(n10107), .ZN(n9766) );
  INV_X1 U12642 ( .A(n12202), .ZN(n10176) );
  OR2_X1 U12643 ( .A1(n18418), .A2(n12005), .ZN(n15838) );
  INV_X1 U12644 ( .A(n15838), .ZN(n18821) );
  INV_X1 U12645 ( .A(n12376), .ZN(n9979) );
  OR2_X1 U12646 ( .A1(n15705), .A2(n15715), .ZN(n9767) );
  INV_X1 U12647 ( .A(n19437), .ZN(n18623) );
  INV_X1 U12648 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n10064) );
  INV_X1 U12649 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10114) );
  OR2_X1 U12650 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n9768) );
  INV_X1 U12651 ( .A(n20316), .ZN(n20516) );
  AND2_X1 U12652 ( .A1(n17710), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n9769) );
  NAND3_X1 U12653 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17352) );
  INV_X1 U12654 ( .A(n17352), .ZN(n10090) );
  NAND2_X1 U12655 ( .A1(n17533), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17507) );
  INV_X1 U12656 ( .A(n17507), .ZN(n9802) );
  AND2_X1 U12657 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_21__SCAN_IN), 
        .ZN(n9770) );
  INV_X1 U12658 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n10038) );
  INV_X1 U12659 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n9996) );
  INV_X1 U12660 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10113) );
  INV_X1 U12661 ( .A(n14329), .ZN(n10280) );
  CLKBUF_X1 U12662 ( .A(n16459), .Z(n9771) );
  NOR4_X1 U12663 ( .A1(n18348), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(
        P3_STATE2_REG_2__SCAN_IN), .A4(P3_STATEBS16_REG_SCAN_IN), .ZN(n16459)
         );
  AOI22_X2 U12664 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19883), .B1(DATAI_19_), 
        .B2(n19884), .ZN(n20413) );
  AOI22_X2 U12665 ( .A1(DATAI_17_), .A2(n19884), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n19883), .ZN(n20401) );
  AOI22_X2 U12666 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19883), .B1(DATAI_20_), 
        .B2(n19884), .ZN(n20369) );
  AOI22_X2 U12667 ( .A1(DATAI_23_), .A2(n19884), .B1(BUF1_REG_23__SCAN_IN), 
        .B2(n19883), .ZN(n20444) );
  NOR2_X2 U12668 ( .A1(n18926), .A2(n18925), .ZN(n19423) );
  AOI22_X2 U12669 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n18924), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n18923), .ZN(n19401) );
  NOR2_X2 U12670 ( .A1(n14634), .A2(n18811), .ZN(n18923) );
  NAND2_X1 U12671 ( .A1(n16790), .A2(n16922), .ZN(n16788) );
  INV_X1 U12672 ( .A(n16922), .ZN(n16868) );
  NOR2_X1 U12673 ( .A1(n16922), .A2(n17772), .ZN(n16856) );
  AOI22_X2 U12674 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19883), .B1(DATAI_16_), 
        .B2(n19884), .ZN(n20395) );
  CLKBUF_X1 U12675 ( .A(n18636), .Z(n9772) );
  INV_X1 U12676 ( .A(n9772), .ZN(n18601) );
  NOR4_X1 U12677 ( .A1(n18850), .A2(n18414), .A3(n18623), .A4(n15907), .ZN(
        n18636) );
  NOR2_X1 U12678 ( .A1(n18919), .A2(n18925), .ZN(n9773) );
  AND2_X1 U12679 ( .A1(n9777), .A2(n19788), .ZN(n9774) );
  NAND2_X1 U12680 ( .A1(n19829), .A2(n9777), .ZN(n9776) );
  NAND2_X1 U12681 ( .A1(n12874), .A2(n12875), .ZN(n9777) );
  NAND2_X1 U12682 ( .A1(n9778), .A2(n9892), .ZN(P1_U3000) );
  NAND4_X1 U12683 ( .A1(n10251), .A2(n10254), .A3(n9651), .A4(n19810), .ZN(
        n9778) );
  NAND2_X1 U12684 ( .A1(n9779), .A2(n14090), .ZN(P1_U2968) );
  NAND4_X1 U12685 ( .A1(n10251), .A2(n10254), .A3(n9651), .A4(n19788), .ZN(
        n9779) );
  NAND2_X1 U12686 ( .A1(n12997), .A2(n12996), .ZN(n12995) );
  OAI21_X2 U12687 ( .B1(n14353), .B2(n10279), .A(n15572), .ZN(n14153) );
  NAND2_X2 U12688 ( .A1(n14177), .A2(n14176), .ZN(n14353) );
  NAND2_X2 U12689 ( .A1(n9868), .A2(n9867), .ZN(n14177) );
  XNOR2_X2 U12690 ( .A(n9780), .B(n10419), .ZN(n19960) );
  NAND2_X1 U12691 ( .A1(n10194), .A2(n9781), .ZN(n9780) );
  OR2_X2 U12692 ( .A1(n14085), .A2(n10256), .ZN(n10253) );
  AND2_X2 U12693 ( .A1(n14084), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14085) );
  NOR2_X2 U12694 ( .A1(n14082), .A2(n14081), .ZN(n14084) );
  NAND2_X2 U12695 ( .A1(n11148), .A2(n14245), .ZN(n14082) );
  XNOR2_X1 U12696 ( .A(n9783), .B(n9844), .ZN(n10192) );
  NAND3_X1 U12697 ( .A1(n17429), .A2(n17416), .A3(n17417), .ZN(n9796) );
  NAND2_X1 U12698 ( .A1(n9803), .A2(n13864), .ZN(n15833) );
  NAND2_X1 U12699 ( .A1(n9803), .A2(n10169), .ZN(n9920) );
  NAND2_X1 U12700 ( .A1(n9805), .A2(n15834), .ZN(n9804) );
  NAND2_X1 U12701 ( .A1(n11297), .A2(n9952), .ZN(n9810) );
  NAND2_X1 U12702 ( .A1(n13298), .A2(n9826), .ZN(n13331) );
  INV_X1 U12703 ( .A(n13298), .ZN(n13330) );
  NOR2_X2 U12704 ( .A1(n14729), .A2(n14721), .ZN(n14720) );
  INV_X2 U12705 ( .A(n14452), .ZN(n11949) );
  AND3_X2 U12706 ( .A1(n9644), .A2(n9861), .A3(n9665), .ZN(n14452) );
  NAND3_X1 U12707 ( .A1(n12636), .A2(n20446), .A3(n10430), .ZN(n9814) );
  OR2_X2 U12708 ( .A1(n14146), .A2(n14099), .ZN(n11144) );
  NAND2_X2 U12709 ( .A1(n11145), .A2(n14154), .ZN(n14146) );
  XNOR2_X2 U12710 ( .A(n12636), .B(n19995), .ZN(n20517) );
  INV_X1 U12711 ( .A(n12511), .ZN(n9819) );
  NAND2_X1 U12712 ( .A1(n12423), .A2(n9989), .ZN(n9820) );
  NAND2_X1 U12713 ( .A1(n13364), .A2(n13327), .ZN(n9894) );
  NAND2_X2 U12714 ( .A1(n9827), .A2(n13330), .ZN(n13439) );
  NAND2_X1 U12715 ( .A1(n9862), .A2(n18926), .ZN(n11363) );
  NAND3_X1 U12716 ( .A1(n10237), .A2(n10238), .A3(n10239), .ZN(n9831) );
  INV_X2 U12717 ( .A(n12776), .ZN(n11348) );
  NAND2_X1 U12718 ( .A1(n9627), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n9832) );
  NAND2_X1 U12719 ( .A1(n11348), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n9833) );
  OR2_X2 U12720 ( .A1(n15268), .A2(n15267), .ZN(n16930) );
  NAND3_X1 U12721 ( .A1(n9691), .A2(n17340), .A3(n9835), .ZN(n17339) );
  NAND2_X1 U12722 ( .A1(n10025), .A2(n10024), .ZN(n9841) );
  INV_X4 U12723 ( .A(n15281), .ZN(n15217) );
  NAND2_X2 U12724 ( .A1(n20317), .A2(n10500), .ZN(n12952) );
  INV_X1 U12725 ( .A(n9850), .ZN(n13145) );
  NAND2_X1 U12726 ( .A1(n10012), .A2(n10011), .ZN(n10010) );
  NAND2_X1 U12727 ( .A1(n17104), .A2(n17103), .ZN(n17102) );
  NOR2_X1 U12728 ( .A1(n15927), .A2(n10014), .ZN(n10013) );
  AOI21_X1 U12729 ( .B1(n15352), .B2(n17236), .A(n17318), .ZN(n17199) );
  NAND4_X1 U12730 ( .A1(n9717), .A2(n11340), .A3(n11341), .A4(n11343), .ZN(
        n9855) );
  NAND4_X1 U12731 ( .A1(n9718), .A2(n11344), .A3(n11345), .A4(n11346), .ZN(
        n9856) );
  NOR2_X2 U12732 ( .A1(n13195), .A2(n10156), .ZN(n14535) );
  XNOR2_X1 U12733 ( .A(n11745), .B(n11743), .ZN(n14481) );
  NOR2_X2 U12734 ( .A1(n14478), .A2(n14477), .ZN(n14476) );
  AND2_X2 U12735 ( .A1(n12918), .A2(n10295), .ZN(n10461) );
  AND2_X2 U12736 ( .A1(n12517), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10295) );
  INV_X2 U12737 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12517) );
  AND2_X2 U12738 ( .A1(n12516), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12918) );
  INV_X2 U12739 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12516) );
  NOR2_X2 U12740 ( .A1(n14083), .A2(n14084), .ZN(n14092) );
  NAND2_X2 U12741 ( .A1(n14121), .A2(n14111), .ZN(n11148) );
  NOR2_X2 U12742 ( .A1(n9865), .A2(n10396), .ZN(n11210) );
  INV_X1 U12743 ( .A(n19873), .ZN(n9865) );
  OR2_X4 U12744 ( .A1(n10333), .A2(n10332), .ZN(n19873) );
  NAND2_X1 U12745 ( .A1(n9868), .A2(n9866), .ZN(n14170) );
  NAND2_X1 U12746 ( .A1(n9870), .A2(n9869), .ZN(n10260) );
  NAND2_X1 U12747 ( .A1(n9603), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11138) );
  XNOR2_X2 U12748 ( .A(n13863), .B(n13861), .ZN(n14815) );
  NAND2_X1 U12749 ( .A1(n13855), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9871) );
  NAND3_X1 U12750 ( .A1(n9962), .A2(n9961), .A3(n9960), .ZN(n13855) );
  OAI21_X2 U12751 ( .B1(n11444), .B2(n9878), .A(n11425), .ZN(n11430) );
  NAND2_X2 U12752 ( .A1(n11389), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11444) );
  INV_X1 U12753 ( .A(n13366), .ZN(n9885) );
  NOR2_X1 U12754 ( .A1(n13364), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13366) );
  NAND3_X1 U12755 ( .A1(n10238), .A2(n10237), .A3(n10236), .ZN(n13845) );
  NAND2_X1 U12756 ( .A1(n10526), .A2(n9889), .ZN(n9887) );
  NAND2_X1 U12757 ( .A1(n10526), .A2(n20446), .ZN(n9888) );
  INV_X1 U12758 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9893) );
  AND4_X2 U12759 ( .A1(n9893), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A4(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10463) );
  NOR2_X1 U12760 ( .A1(n13257), .A2(n13260), .ZN(n9898) );
  NAND2_X1 U12761 ( .A1(n9931), .A2(n9909), .ZN(n9908) );
  AND2_X1 U12762 ( .A1(n10241), .A2(n14809), .ZN(n9909) );
  NAND2_X1 U12763 ( .A1(n11389), .A2(n9910), .ZN(n11409) );
  OAI22_X2 U12764 ( .A1(n11366), .A2(n9634), .B1(n12584), .B2(n12583), .ZN(
        n12578) );
  XNOR2_X2 U12765 ( .A(n9912), .B(n10446), .ZN(n10526) );
  INV_X1 U12766 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9913) );
  NAND2_X1 U12767 ( .A1(n12636), .A2(n10430), .ZN(n20259) );
  NAND2_X1 U12768 ( .A1(n9603), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14194) );
  NAND2_X1 U12769 ( .A1(n9917), .A2(n11426), .ZN(n11428) );
  NAND2_X1 U12770 ( .A1(n13364), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13438) );
  NAND3_X1 U12771 ( .A1(n9920), .A2(n9919), .A3(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15059) );
  NAND3_X1 U12772 ( .A1(n9920), .A2(n9919), .A3(n9918), .ZN(n15023) );
  NOR2_X2 U12773 ( .A1(n15023), .A2(n15030), .ZN(n15799) );
  NAND3_X1 U12774 ( .A1(n9930), .A2(n9658), .A3(n9929), .ZN(n9928) );
  NAND3_X1 U12775 ( .A1(n11375), .A2(n11339), .A3(n9722), .ZN(n9942) );
  NAND3_X1 U12776 ( .A1(n11375), .A2(n11339), .A3(n11832), .ZN(n12209) );
  NAND4_X1 U12777 ( .A1(n9720), .A2(n11325), .A3(n11326), .A4(n11324), .ZN(
        n9950) );
  NAND4_X1 U12778 ( .A1(n9719), .A2(n11321), .A3(n11323), .A4(n11322), .ZN(
        n9951) );
  NAND2_X1 U12779 ( .A1(n9956), .A2(n11422), .ZN(n11423) );
  XNOR2_X2 U12780 ( .A(n9956), .B(n11422), .ZN(n13231) );
  INV_X1 U12781 ( .A(n11418), .ZN(n9956) );
  NAND3_X1 U12782 ( .A1(n14506), .A2(n9673), .A3(n9645), .ZN(n10139) );
  NAND2_X1 U12783 ( .A1(n13345), .A2(n9959), .ZN(n9958) );
  INV_X1 U12784 ( .A(n15849), .ZN(n9959) );
  NAND3_X1 U12785 ( .A1(n13363), .A2(n13470), .A3(n9964), .ZN(n9960) );
  NAND2_X1 U12786 ( .A1(n9963), .A2(n9965), .ZN(n9962) );
  NAND2_X1 U12787 ( .A1(n13363), .A2(n9964), .ZN(n13471) );
  NAND2_X1 U12788 ( .A1(n9968), .A2(n9967), .ZN(n14729) );
  INV_X1 U12789 ( .A(n10166), .ZN(n10169) );
  NAND3_X1 U12790 ( .A1(n9970), .A2(n10208), .A3(n9969), .ZN(P2_U3015) );
  NAND2_X1 U12791 ( .A1(n12296), .A2(n12295), .ZN(n12894) );
  INV_X1 U12792 ( .A(n9978), .ZN(n13898) );
  INV_X1 U12793 ( .A(n9984), .ZN(n14334) );
  INV_X1 U12794 ( .A(n12346), .ZN(n9985) );
  AND2_X1 U12795 ( .A1(n12423), .A2(n19886), .ZN(n11246) );
  OAI21_X2 U12796 ( .B1(n14163), .B2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n9603), .ZN(n14154) );
  AND3_X2 U12797 ( .A1(n9703), .A2(n10020), .A3(n10017), .ZN(n16923) );
  INV_X1 U12798 ( .A(n11441), .ZN(n10026) );
  INV_X1 U12799 ( .A(n11442), .ZN(n10032) );
  OAI21_X2 U12800 ( .B1(n11443), .B2(n11442), .A(n11441), .ZN(n11887) );
  NAND2_X2 U12801 ( .A1(n10037), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11895) );
  NAND2_X1 U12802 ( .A1(n10037), .A2(n10036), .ZN(n11385) );
  NAND2_X1 U12803 ( .A1(n12558), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11391) );
  NOR3_X2 U12804 ( .A1(n14503), .A2(n10044), .A3(n14492), .ZN(n14485) );
  INV_X1 U12805 ( .A(n14473), .ZN(n10043) );
  INV_X1 U12806 ( .A(n10047), .ZN(n14509) );
  INV_X1 U12807 ( .A(n12256), .ZN(n10048) );
  AND2_X2 U12808 ( .A1(n13119), .A2(n9740), .ZN(n14544) );
  NAND3_X1 U12809 ( .A1(n10054), .A2(n10165), .A3(n10163), .ZN(P2_U2983) );
  NAND2_X1 U12810 ( .A1(n12255), .A2(n9676), .ZN(n13836) );
  NAND2_X1 U12811 ( .A1(n13746), .A2(n10070), .ZN(n13765) );
  CLKBUF_X1 U12812 ( .A(n9609), .Z(n10079) );
  AOI21_X1 U12813 ( .B1(n10083), .B2(n9771), .A(n10081), .ZN(n16154) );
  INV_X1 U12814 ( .A(n17226), .ZN(n10089) );
  NAND2_X1 U12815 ( .A1(n10100), .A2(n9745), .ZN(n16216) );
  NAND2_X1 U12816 ( .A1(n16238), .A2(n10102), .ZN(n10100) );
  AND2_X1 U12817 ( .A1(n9609), .A2(n10105), .ZN(n10104) );
  NOR2_X1 U12818 ( .A1(n16227), .A2(n17126), .ZN(n16226) );
  NOR2_X1 U12819 ( .A1(n16238), .A2(n9609), .ZN(n16227) );
  NAND2_X1 U12820 ( .A1(n11978), .A2(n10111), .ZN(n11976) );
  NAND2_X1 U12821 ( .A1(n10115), .A2(n10116), .ZN(n15704) );
  OR2_X1 U12822 ( .A1(n15716), .A2(n15715), .ZN(n10117) );
  INV_X1 U12823 ( .A(n10117), .ZN(n15714) );
  NAND2_X1 U12824 ( .A1(n18442), .A2(n15696), .ZN(n10119) );
  INV_X1 U12825 ( .A(n10121), .ZN(n18441) );
  INV_X1 U12826 ( .A(n10120), .ZN(n12250) );
  AOI21_X1 U12827 ( .B1(n15766), .B2(n14718), .A(n18630), .ZN(n10128) );
  INV_X1 U12828 ( .A(n10126), .ZN(n15748) );
  AOI22_X1 U12829 ( .A1(n15766), .A2(n9762), .B1(n18630), .B2(n10127), .ZN(
        n10126) );
  AND2_X2 U12830 ( .A1(n11974), .A2(n10134), .ZN(n12000) );
  INV_X1 U12831 ( .A(n11417), .ZN(n10137) );
  XNOR2_X1 U12832 ( .A(n11417), .B(n10138), .ZN(n19546) );
  NAND2_X1 U12833 ( .A1(n10143), .A2(n11823), .ZN(n10142) );
  NAND2_X1 U12834 ( .A1(n14476), .A2(n9759), .ZN(n10144) );
  NAND2_X1 U12835 ( .A1(n14552), .A2(n18694), .ZN(n14557) );
  NAND2_X1 U12836 ( .A1(n14476), .A2(n9760), .ZN(n10146) );
  NOR2_X1 U12837 ( .A1(n11800), .A2(n11799), .ZN(n10150) );
  NOR2_X1 U12838 ( .A1(n12815), .A2(n10162), .ZN(n12779) );
  NAND2_X1 U12839 ( .A1(n14581), .A2(n9763), .ZN(n14830) );
  NAND2_X1 U12840 ( .A1(n14581), .A2(n9751), .ZN(n14563) );
  NAND2_X1 U12841 ( .A1(n10181), .A2(n10180), .ZN(n10179) );
  NAND2_X1 U12842 ( .A1(n9663), .A2(n10181), .ZN(n13369) );
  NOR2_X1 U12843 ( .A1(n15855), .A2(n15856), .ZN(n15854) );
  INV_X1 U12844 ( .A(n13048), .ZN(n10183) );
  AND2_X2 U12845 ( .A1(n12635), .A2(n10187), .ZN(n12911) );
  NAND3_X1 U12846 ( .A1(n10500), .A2(n10190), .A3(n10423), .ZN(n10430) );
  NAND2_X1 U12847 ( .A1(n10192), .A2(n10773), .ZN(n10514) );
  CLKBUF_X1 U12848 ( .A(n10192), .Z(n10191) );
  NAND2_X1 U12849 ( .A1(n10192), .A2(n11123), .ZN(n11079) );
  NOR2_X1 U12850 ( .A1(n20524), .A2(n10191), .ZN(n19958) );
  NAND2_X1 U12851 ( .A1(n10191), .A2(n19994), .ZN(n20521) );
  NAND2_X1 U12852 ( .A1(n10191), .A2(n19837), .ZN(n20389) );
  OAI21_X1 U12853 ( .B1(n20117), .B2(n20347), .A(n20316), .ZN(n10193) );
  NAND2_X1 U12854 ( .A1(n13999), .A2(n9744), .ZN(n13995) );
  NAND2_X1 U12855 ( .A1(n12276), .A2(n10205), .ZN(n13905) );
  AND2_X1 U12856 ( .A1(n12276), .A2(n10206), .ZN(n13915) );
  NAND2_X1 U12857 ( .A1(n14663), .A2(n10212), .ZN(n10210) );
  INV_X1 U12858 ( .A(n14662), .ZN(n10216) );
  OR2_X2 U12859 ( .A1(n10221), .A2(n10220), .ZN(n10219) );
  NAND2_X1 U12860 ( .A1(n13742), .A2(n13741), .ZN(n10225) );
  OAI21_X1 U12861 ( .B1(n13345), .B2(n10231), .A(n10228), .ZN(n18807) );
  NAND2_X1 U12862 ( .A1(n10227), .A2(n10226), .ZN(n13344) );
  NAND2_X1 U12863 ( .A1(n13345), .A2(n10228), .ZN(n10227) );
  AOI21_X1 U12864 ( .B1(n13332), .B2(n12224), .A(n15903), .ZN(n10235) );
  NOR2_X4 U12865 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14428) );
  NAND2_X1 U12866 ( .A1(n14085), .A2(n14238), .ZN(n10252) );
  NAND3_X1 U12867 ( .A1(n14092), .A2(n10255), .A3(n14238), .ZN(n10254) );
  INV_X1 U12868 ( .A(n14085), .ZN(n10255) );
  NOR2_X1 U12869 ( .A1(n14092), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14091) );
  NAND2_X1 U12870 ( .A1(n10260), .A2(n10261), .ZN(n13546) );
  NAND2_X1 U12871 ( .A1(n15593), .A2(n10266), .ZN(n10265) );
  NAND3_X1 U12872 ( .A1(n10273), .A2(n10412), .A3(n10271), .ZN(n10403) );
  NAND2_X1 U12873 ( .A1(n10272), .A2(n10274), .ZN(n10271) );
  NAND2_X1 U12874 ( .A1(n10400), .A2(n12684), .ZN(n10273) );
  NOR2_X2 U12875 ( .A1(n10403), .A2(n12420), .ZN(n12478) );
  NAND3_X1 U12876 ( .A1(n14121), .A2(n14111), .A3(n11149), .ZN(n14080) );
  NAND2_X2 U12877 ( .A1(n11147), .A2(n11146), .ZN(n14111) );
  NAND2_X2 U12878 ( .A1(n11144), .A2(n9603), .ZN(n14121) );
  AOI21_X1 U12879 ( .B1(n10406), .B2(n10278), .A(n10276), .ZN(n10275) );
  MUX2_X1 U12880 ( .A(n20216), .B(n20387), .S(n20117), .Z(n12941) );
  NAND2_X1 U12881 ( .A1(n11467), .A2(n11466), .ZN(n12667) );
  NAND2_X1 U12882 ( .A1(n11992), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11989) );
  NOR2_X1 U12883 ( .A1(n12394), .A2(n12209), .ZN(n12397) );
  OR2_X1 U12884 ( .A1(n11444), .A2(n9952), .ZN(n11447) );
  NAND2_X1 U12885 ( .A1(n11980), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11981) );
  NOR2_X1 U12886 ( .A1(n18919), .A2(n18925), .ZN(n19416) );
  AND2_X1 U12887 ( .A1(n18686), .A2(n18926), .ZN(n18692) );
  NAND2_X1 U12888 ( .A1(n12664), .A2(n12663), .ZN(n19566) );
  NAND2_X1 U12889 ( .A1(n10408), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10419) );
  NOR2_X2 U12890 ( .A1(n19878), .A2(n20448), .ZN(n10773) );
  INV_X1 U12891 ( .A(n11895), .ZN(n11448) );
  INV_X1 U12892 ( .A(n10532), .ZN(n11028) );
  INV_X1 U12893 ( .A(n13570), .ZN(n15218) );
  INV_X1 U12894 ( .A(n12004), .ZN(n12187) );
  NOR2_X1 U12895 ( .A1(n13771), .A2(n13768), .ZN(n10282) );
  OR2_X1 U12896 ( .A1(n11561), .A2(n11560), .ZN(n10283) );
  CLKBUF_X3 U12897 ( .A(n11888), .Z(n14451) );
  INV_X1 U12898 ( .A(n17310), .ZN(n17574) );
  INV_X2 U12899 ( .A(n16765), .ZN(n16774) );
  AND2_X1 U12900 ( .A1(n12396), .A2(n15904), .ZN(n13482) );
  NAND2_X1 U12901 ( .A1(n11405), .A2(n11415), .ZN(n12528) );
  AND2_X1 U12902 ( .A1(n19195), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10284) );
  AND2_X1 U12903 ( .A1(n11333), .A2(n11332), .ZN(n10285) );
  INV_X1 U12904 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17207) );
  AND2_X1 U12905 ( .A1(n19136), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n10286) );
  INV_X1 U12906 ( .A(n12006), .ZN(n12186) );
  NOR2_X1 U12907 ( .A1(n18255), .A2(n17396), .ZN(n17154) );
  INV_X4 U12908 ( .A(n9614), .ZN(n18911) );
  NOR2_X1 U12909 ( .A1(n13572), .A2(n18205), .ZN(n15251) );
  NOR2_X1 U12910 ( .A1(n13572), .A2(n16465), .ZN(n15226) );
  AND2_X1 U12911 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10287) );
  AND3_X1 U12912 ( .A1(n17127), .A2(n17451), .A3(n17480), .ZN(n10288) );
  INV_X1 U12913 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17214) );
  INV_X1 U12914 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17187) );
  INV_X1 U12915 ( .A(n12965), .ZN(n11503) );
  INV_X1 U12916 ( .A(n13118), .ZN(n11550) );
  AND4_X1 U12917 ( .A1(n13256), .A2(n13255), .A3(n13254), .A4(n13253), .ZN(
        n10289) );
  AOI22_X1 U12918 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19023), .B1(
        n13442), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13292) );
  INV_X1 U12919 ( .A(n11159), .ZN(n11167) );
  OR2_X1 U12920 ( .A1(n10581), .A2(n10580), .ZN(n11098) );
  XNOR2_X1 U12921 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11185) );
  AND2_X1 U12922 ( .A1(n11191), .A2(n11190), .ZN(n11251) );
  OR2_X1 U12923 ( .A1(n10611), .A2(n10610), .ZN(n11116) );
  OR2_X1 U12924 ( .A1(n10629), .A2(n10628), .ZN(n11115) );
  NOR2_X1 U12925 ( .A1(n11194), .A2(n11192), .ZN(n11197) );
  NAND2_X1 U12926 ( .A1(n11363), .A2(n9808), .ZN(n11364) );
  INV_X1 U12927 ( .A(n12857), .ZN(n11445) );
  OR2_X1 U12928 ( .A1(n10559), .A2(n10558), .ZN(n11099) );
  XNOR2_X1 U12929 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12435) );
  AND2_X1 U12930 ( .A1(n13326), .A2(n13325), .ZN(n13440) );
  INV_X1 U12931 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12827) );
  AND2_X1 U12932 ( .A1(n12334), .A2(n12333), .ZN(n13533) );
  OR2_X1 U12933 ( .A1(n11056), .A2(n11215), .ZN(n12284) );
  AND2_X1 U12934 ( .A1(n10957), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10958) );
  NOR2_X1 U12935 ( .A1(n20629), .A2(n10715), .ZN(n10747) );
  INV_X1 U12936 ( .A(n11099), .ZN(n11084) );
  INV_X1 U12937 ( .A(n9692), .ZN(n12352) );
  NOR2_X1 U12938 ( .A1(n11187), .A2(n11160), .ZN(n11203) );
  NAND2_X1 U12939 ( .A1(n10428), .A2(n10427), .ZN(n10429) );
  OR2_X2 U12940 ( .A1(n10344), .A2(n10343), .ZN(n10396) );
  NOR2_X1 U12941 ( .A1(n12214), .A2(n12219), .ZN(n12440) );
  AND2_X1 U12942 ( .A1(n18911), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n13792) );
  INV_X1 U12943 ( .A(n11655), .ZN(n11801) );
  OR2_X1 U12944 ( .A1(n11740), .A2(n11742), .ZN(n11763) );
  NOR2_X1 U12945 ( .A1(n11373), .A2(n12549), .ZN(n11374) );
  AND4_X1 U12946 ( .A1(n11317), .A2(n11316), .A3(n11315), .A4(n11314), .ZN(
        n11318) );
  INV_X1 U12947 ( .A(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n20658) );
  INV_X1 U12948 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n15296) );
  NOR2_X1 U12949 ( .A1(n10917), .A2(n14158), .ZN(n10918) );
  AND2_X1 U12950 ( .A1(n12337), .A2(n12336), .ZN(n14398) );
  INV_X1 U12951 ( .A(n10999), .ZN(n11237) );
  INV_X1 U12952 ( .A(n11239), .ZN(n11051) );
  NOR2_X1 U12953 ( .A1(n12284), .A2(n14095), .ZN(n12285) );
  AND2_X1 U12954 ( .A1(n12284), .A2(n11057), .ZN(n13731) );
  NAND2_X1 U12955 ( .A1(n10958), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11002) );
  INV_X1 U12956 ( .A(n11028), .ZN(n12280) );
  INV_X1 U12957 ( .A(n12971), .ZN(n10597) );
  AND3_X1 U12958 ( .A1(n12502), .A2(n11063), .A3(n11209), .ZN(n12484) );
  AND2_X1 U12959 ( .A1(n12312), .A2(n12311), .ZN(n15667) );
  AND2_X1 U12960 ( .A1(n10538), .A2(n20384), .ZN(n19844) );
  AOI221_X1 U12961 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n11843), 
        .C1(n15192), .C2(n11843), .A(n11831), .ZN(n12442) );
  NOR2_X1 U12962 ( .A1(n12765), .A2(n11809), .ZN(n11469) );
  OR2_X1 U12963 ( .A1(n11763), .A2(n11765), .ZN(n11786) );
  NOR2_X1 U12964 ( .A1(n12125), .A2(n12124), .ZN(n13467) );
  INV_X1 U12965 ( .A(n18837), .ZN(n15028) );
  AND2_X1 U12966 ( .A1(n12548), .A2(n12547), .ZN(n12784) );
  OR2_X1 U12967 ( .A1(n12575), .A2(n12574), .ZN(n12834) );
  INV_X1 U12968 ( .A(n17760), .ZN(n15093) );
  OR3_X1 U12969 ( .A1(n16890), .A2(n15093), .A3(n15092), .ZN(n15094) );
  INV_X1 U12970 ( .A(n17627), .ZN(n17671) );
  NOR2_X1 U12971 ( .A1(n17580), .A2(n17559), .ZN(n17239) );
  INV_X1 U12972 ( .A(n18188), .ZN(n17602) );
  NAND2_X1 U12973 ( .A1(n17391), .A2(n17390), .ZN(n17389) );
  NOR2_X1 U12974 ( .A1(n17766), .A2(n15200), .ZN(n15205) );
  INV_X1 U12975 ( .A(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n20623) );
  NAND2_X1 U12976 ( .A1(n10918), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10956) );
  AND2_X1 U12977 ( .A1(n13961), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13063) );
  OR3_X1 U12978 ( .A1(n20550), .A2(n12283), .A3(n12282), .ZN(n13961) );
  NAND2_X1 U12979 ( .A1(n14399), .A2(n14398), .ZN(n14401) );
  AOI21_X1 U12980 ( .B1(n11097), .B2(n10773), .A(n10617), .ZN(n13005) );
  AND4_X1 U12981 ( .A1(n10390), .A2(n10389), .A3(n10388), .A4(n10387), .ZN(
        n10391) );
  AOI21_X1 U12982 ( .B1(n15566), .B2(n13731), .A(n11216), .ZN(n11217) );
  INV_X1 U12983 ( .A(n12276), .ZN(n13930) );
  NAND2_X1 U12984 ( .A1(n10810), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10840) );
  INV_X1 U12985 ( .A(n13526), .ZN(n14076) );
  OR2_X1 U12986 ( .A1(n19788), .A2(n11211), .ZN(n14190) );
  OR2_X1 U12987 ( .A1(n14303), .A2(n14243), .ZN(n14289) );
  OR2_X1 U12988 ( .A1(n19824), .A2(n14240), .ZN(n14324) );
  AND2_X1 U12989 ( .A1(n15609), .A2(n14326), .ZN(n19795) );
  AND2_X1 U12990 ( .A1(n12478), .A2(n13062), .ZN(n12712) );
  AND2_X1 U12991 ( .A1(n11205), .A2(n11204), .ZN(n12691) );
  AND2_X1 U12992 ( .A1(n19959), .A2(n20089), .ZN(n19969) );
  INV_X1 U12993 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19923) );
  OR2_X1 U12994 ( .A1(n20223), .A2(n20222), .ZN(n20255) );
  OR2_X1 U12995 ( .A1(n20389), .A2(n20254), .ZN(n20322) );
  INV_X1 U12996 ( .A(n19922), .ZN(n19838) );
  NOR2_X1 U12997 ( .A1(n18630), .A2(n15748), .ZN(n15735) );
  NOR2_X1 U12998 ( .A1(n18630), .A2(n18473), .ZN(n18463) );
  OAI21_X1 U12999 ( .B1(n12528), .B2(n11416), .A(n11415), .ZN(n11417) );
  INV_X1 U13000 ( .A(n11700), .ZN(n11679) );
  OR2_X1 U13001 ( .A1(n11584), .A2(n11583), .ZN(n13385) );
  OR2_X1 U13002 ( .A1(n14960), .A2(n13876), .ZN(n14935) );
  OR2_X1 U13003 ( .A1(n14992), .A2(n14732), .ZN(n14960) );
  INV_X1 U13004 ( .A(n13482), .ZN(n18600) );
  AND2_X1 U13005 ( .A1(n15894), .A2(n13870), .ZN(n15029) );
  INV_X1 U13006 ( .A(n13482), .ZN(n18496) );
  INV_X1 U13007 ( .A(n18959), .ZN(n19019) );
  OR2_X1 U13008 ( .A1(n19108), .A2(n19373), .ZN(n19129) );
  INV_X1 U13009 ( .A(n19557), .ZN(n19538) );
  NAND2_X1 U13010 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19377), .ZN(n18925) );
  OAI21_X1 U13011 ( .B1(n13692), .B2(n13679), .A(n13678), .ZN(n13694) );
  NOR2_X1 U13012 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n16230), .ZN(n16217) );
  NOR2_X1 U13013 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n16270), .ZN(n16257) );
  NOR2_X1 U13014 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n16306), .ZN(n16297) );
  INV_X1 U13015 ( .A(n16131), .ZN(n16112) );
  NAND2_X1 U13016 ( .A1(n16976), .A2(n13691), .ZN(n18215) );
  INV_X1 U13017 ( .A(n16730), .ZN(n16646) );
  INV_X1 U13018 ( .A(n17766), .ZN(n16784) );
  INV_X1 U13019 ( .A(n17154), .ZN(n17070) );
  NOR3_X1 U13020 ( .A1(n17140), .A2(n17138), .A3(n16125), .ZN(n17084) );
  INV_X1 U13021 ( .A(n17186), .ZN(n17188) );
  NOR2_X1 U13022 ( .A1(n17610), .A2(n17602), .ZN(n17630) );
  AOI21_X1 U13023 ( .B1(n18180), .B2(n18176), .A(n18179), .ZN(n18188) );
  NOR2_X1 U13024 ( .A1(n18364), .A2(n18253), .ZN(n17734) );
  INV_X1 U13025 ( .A(n18121), .ZN(n18090) );
  INV_X1 U13026 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18348) );
  NAND2_X1 U13027 ( .A1(n10875), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10917) );
  NOR2_X1 U13028 ( .A1(n13963), .A2(n13508), .ZN(n15525) );
  AND2_X1 U13029 ( .A1(n13961), .A2(n12286), .ZN(n19659) );
  AND2_X1 U13030 ( .A1(n13063), .A2(n12378), .ZN(n19686) );
  NAND2_X1 U13031 ( .A1(n13988), .A2(n13987), .ZN(n13990) );
  INV_X1 U13032 ( .A(n14024), .ZN(n19706) );
  NAND2_X1 U13033 ( .A1(n12650), .A2(n12696), .ZN(n12653) );
  INV_X1 U13034 ( .A(n19713), .ZN(n15545) );
  NAND2_X1 U13035 ( .A1(n10700), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10714) );
  NAND2_X1 U13036 ( .A1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n10645), .ZN(
        n10666) );
  AND2_X1 U13037 ( .A1(n10589), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10614) );
  NAND2_X1 U13038 ( .A1(n12717), .A2(n12716), .ZN(n19823) );
  AND2_X1 U13039 ( .A1(n19826), .A2(n15623), .ZN(n19809) );
  INV_X1 U13040 ( .A(n19795), .ZN(n19818) );
  INV_X1 U13041 ( .A(n19823), .ZN(n19807) );
  NOR2_X1 U13042 ( .A1(n20270), .A2(n12691), .ZN(n14426) );
  OAI22_X1 U13043 ( .A1(n19850), .A2(n19849), .B1(n20172), .B2(n19997), .ZN(
        n19890) );
  INV_X1 U13044 ( .A(n19915), .ZN(n19918) );
  AND2_X1 U13045 ( .A1(n9631), .A2(n19922), .ZN(n20048) );
  INV_X1 U13046 ( .A(n19988), .ZN(n19984) );
  NOR2_X2 U13047 ( .A1(n19964), .A2(n20222), .ZN(n20018) );
  OR2_X1 U13048 ( .A1(n9631), .A2(n19838), .ZN(n20254) );
  INV_X1 U13049 ( .A(n20116), .ZN(n20142) );
  INV_X1 U13050 ( .A(n20254), .ZN(n20118) );
  INV_X1 U13051 ( .A(n20198), .ZN(n20205) );
  NAND2_X1 U13052 ( .A1(n20117), .A2(n20524), .ZN(n20223) );
  INV_X1 U13053 ( .A(n20255), .ZN(n20308) );
  INV_X1 U13054 ( .A(n19897), .ZN(n20000) );
  OR2_X1 U13055 ( .A1(n9631), .A2(n19922), .ZN(n20314) );
  INV_X1 U13056 ( .A(n20355), .ZN(n20378) );
  INV_X1 U13057 ( .A(n20279), .ZN(n20397) );
  INV_X1 U13058 ( .A(n20294), .ZN(n20415) );
  INV_X1 U13059 ( .A(n20306), .ZN(n20434) );
  AND2_X1 U13060 ( .A1(n20446), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20547) );
  INV_X1 U13061 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20451) );
  NAND2_X1 U13062 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n11856), .ZN(n18416) );
  NAND2_X1 U13063 ( .A1(n18601), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n18540) );
  NAND2_X1 U13064 ( .A1(n14544), .A2(n14543), .ZN(n14546) );
  AND2_X1 U13065 ( .A1(n12401), .A2(n12229), .ZN(n18637) );
  OR2_X1 U13066 ( .A1(n11539), .A2(n11538), .ZN(n13053) );
  AND2_X1 U13067 ( .A1(n18686), .A2(n12045), .ZN(n18694) );
  NOR2_X1 U13068 ( .A1(n12410), .A2(n18801), .ZN(n18773) );
  INV_X1 U13069 ( .A(n18804), .ZN(n12410) );
  AOI21_X1 U13070 ( .B1(n14463), .B2(n9681), .A(n14462), .ZN(n15703) );
  INV_X1 U13071 ( .A(n18811), .ZN(n18830) );
  INV_X1 U13072 ( .A(n15852), .ZN(n18820) );
  NOR2_X1 U13073 ( .A1(n15881), .A2(n15880), .ZN(n15862) );
  INV_X1 U13074 ( .A(n15029), .ZN(n15068) );
  OR2_X1 U13075 ( .A1(n12848), .A2(n12444), .ZN(n19575) );
  NAND2_X1 U13076 ( .A1(n12557), .A2(n18699), .ZN(n12593) );
  INV_X1 U13077 ( .A(n18859), .ZN(n18846) );
  INV_X1 U13078 ( .A(n18861), .ZN(n18849) );
  INV_X1 U13079 ( .A(n19377), .ZN(n19104) );
  OAI21_X1 U13080 ( .B1(n18890), .B2(n18889), .A(n18888), .ZN(n18929) );
  INV_X1 U13081 ( .A(n19536), .ZN(n19191) );
  INV_X1 U13082 ( .A(n19010), .ZN(n19045) );
  NOR2_X1 U13083 ( .A1(n19019), .A2(n19297), .ZN(n19068) );
  INV_X1 U13084 ( .A(n19129), .ZN(n19154) );
  INV_X1 U13085 ( .A(n19161), .ZN(n19159) );
  INV_X1 U13086 ( .A(n19190), .ZN(n19217) );
  NOR2_X1 U13087 ( .A1(n19331), .A2(n19191), .ZN(n19254) );
  AND2_X1 U13088 ( .A1(n19546), .A2(n19538), .ZN(n19536) );
  OR2_X1 U13089 ( .A1(n19546), .A2(n19538), .ZN(n19297) );
  OAI22_X1 U13090 ( .A1(n18918), .A2(n18917), .B1(n18916), .B2(n18915), .ZN(
        n19418) );
  NOR2_X2 U13091 ( .A1(n14633), .A2(n18811), .ZN(n18924) );
  INV_X1 U13092 ( .A(n19563), .ZN(n12863) );
  INV_X1 U13093 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20627) );
  NOR2_X1 U13094 ( .A1(n13601), .A2(n13600), .ZN(n16111) );
  NOR2_X1 U13095 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n16210), .ZN(n16198) );
  NOR2_X1 U13096 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16248), .ZN(n16236) );
  NOR2_X1 U13097 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n16286), .ZN(n16274) );
  NOR2_X1 U13098 ( .A1(n20705), .A2(n16310), .ZN(n16291) );
  NOR2_X1 U13099 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n16360), .ZN(n16345) );
  NOR2_X1 U13100 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n16382), .ZN(n16367) );
  NOR2_X1 U13101 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n16430), .ZN(n16411) );
  NOR2_X2 U13102 ( .A1(n18339), .A2(n16479), .ZN(n16443) );
  NAND2_X1 U13103 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16552), .ZN(n16546) );
  NAND2_X1 U13104 ( .A1(n16646), .A2(n16645), .ZN(n15183) );
  INV_X1 U13105 ( .A(n16795), .ZN(n16791) );
  OR2_X1 U13106 ( .A1(n16995), .A2(n16812), .ZN(n16813) );
  NOR2_X1 U13107 ( .A1(n16981), .A2(n16849), .ZN(n16850) );
  NOR4_X1 U13108 ( .A1(n16896), .A2(n17032), .A3(n17029), .A4(n16780), .ZN(
        n16867) );
  INV_X2 U13109 ( .A(n17778), .ZN(n16890) );
  NAND2_X1 U13110 ( .A1(n16890), .A2(n15426), .ZN(n16922) );
  NOR2_X1 U13111 ( .A1(n17418), .A2(n17081), .ZN(n17042) );
  INV_X1 U13112 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17152) );
  INV_X1 U13113 ( .A(n17247), .ZN(n17258) );
  INV_X1 U13114 ( .A(n17408), .ZN(n17396) );
  NOR2_X1 U13115 ( .A1(n15307), .A2(n15306), .ZN(n17407) );
  INV_X1 U13116 ( .A(n17573), .ZN(n17472) );
  INV_X1 U13117 ( .A(n17636), .ZN(n17613) );
  INV_X1 U13118 ( .A(n9746), .ZN(n17715) );
  INV_X1 U13119 ( .A(n18037), .ZN(n17896) );
  NOR2_X1 U13120 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18339), .ZN(
        n18364) );
  INV_X1 U13121 ( .A(n17836), .ZN(n17846) );
  INV_X1 U13122 ( .A(n17881), .ZN(n17891) );
  INV_X1 U13123 ( .A(n17905), .ZN(n17937) );
  INV_X1 U13124 ( .A(n17980), .ZN(n17982) );
  INV_X1 U13125 ( .A(n18029), .ZN(n18031) );
  INV_X1 U13126 ( .A(n18081), .ZN(n18083) );
  INV_X1 U13127 ( .A(n18115), .ZN(n18106) );
  OAI22_X1 U13128 ( .A1(n15917), .A2(n17468), .B1(n15916), .B2(n18224), .ZN(
        n18231) );
  NOR3_X1 U13129 ( .A1(n18403), .A2(n18394), .A3(P3_STATE2_REG_1__SCAN_IN), 
        .ZN(n18235) );
  NOR2_X1 U13130 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12249), .ZN(n16072)
         );
  NAND2_X1 U13131 ( .A1(n12688), .A2(n11246), .ZN(n12642) );
  INV_X1 U13132 ( .A(n19675), .ZN(n19691) );
  INV_X1 U13133 ( .A(n19686), .ZN(n19681) );
  INV_X1 U13134 ( .A(n19659), .ZN(n15470) );
  INV_X1 U13135 ( .A(n19636), .ZN(n19669) );
  NAND2_X1 U13136 ( .A1(n19710), .A2(n13724), .ZN(n14025) );
  OR2_X1 U13137 ( .A1(n13523), .A2(n13522), .ZN(n15543) );
  NAND2_X1 U13138 ( .A1(n12959), .A2(n11257), .ZN(n19713) );
  INV_X1 U13139 ( .A(n19716), .ZN(n19748) );
  OR3_X1 U13140 ( .A1(n12642), .A2(n12597), .A3(n20457), .ZN(n12959) );
  INV_X1 U13141 ( .A(n15566), .ZN(n19793) );
  INV_X1 U13142 ( .A(n19788), .ZN(n19608) );
  NAND2_X1 U13143 ( .A1(n12717), .A2(n12704), .ZN(n19820) );
  INV_X1 U13144 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20528) );
  NAND2_X1 U13145 ( .A1(n19958), .A2(n20118), .ZN(n19915) );
  NAND2_X1 U13146 ( .A1(n19958), .A2(n20048), .ZN(n19988) );
  AOI22_X1 U13147 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n19965), .B1(n19963), 
        .B2(n19968), .ZN(n19993) );
  OR2_X1 U13148 ( .A1(n20521), .A2(n20254), .ZN(n20047) );
  OR2_X1 U13149 ( .A1(n20521), .A2(n20314), .ZN(n20084) );
  OR2_X1 U13150 ( .A1(n20521), .A2(n20343), .ZN(n20109) );
  OR2_X1 U13151 ( .A1(n20521), .A2(n20222), .ZN(n20116) );
  NAND2_X1 U13152 ( .A1(n20119), .A2(n20118), .ZN(n20170) );
  AOI22_X1 U13153 ( .A1(n20177), .A2(n20175), .B1(n20344), .B2(n20173), .ZN(
        n20209) );
  OR2_X1 U13154 ( .A1(n20223), .A2(n20343), .ZN(n20252) );
  AOI22_X1 U13155 ( .A1(n20268), .A2(n20265), .B1(n20261), .B2(n20260), .ZN(
        n20313) );
  OR2_X1 U13156 ( .A1(n20389), .A2(n20314), .ZN(n20355) );
  OR2_X1 U13157 ( .A1(n20389), .A2(n20343), .ZN(n20426) );
  INV_X1 U13158 ( .A(n20503), .ZN(n20540) );
  NOR2_X1 U13159 ( .A1(n12843), .A2(n18416), .ZN(n18414) );
  AOI21_X1 U13160 ( .B1(n14553), .B2(n18647), .A(n12233), .ZN(n12234) );
  INV_X1 U13161 ( .A(n18625), .ZN(n18643) );
  INV_X1 U13162 ( .A(n18503), .ZN(n15002) );
  INV_X1 U13163 ( .A(n18694), .ZN(n18671) );
  INV_X1 U13164 ( .A(n18691), .ZN(n18686) );
  NOR2_X1 U13165 ( .A1(n18694), .A2(n18692), .ZN(n18675) );
  AND2_X1 U13166 ( .A1(n14611), .A2(n12633), .ZN(n18698) );
  NAND2_X1 U13167 ( .A1(n18737), .A2(n18705), .ZN(n18735) );
  INV_X1 U13168 ( .A(n18737), .ZN(n18769) );
  NAND2_X1 U13169 ( .A1(n12397), .A2(n18895), .ZN(n18702) );
  OR2_X1 U13170 ( .A1(n18418), .A2(n18895), .ZN(n18833) );
  INV_X1 U13171 ( .A(n18829), .ZN(n18816) );
  OR2_X1 U13172 ( .A1(n12593), .A2(n19575), .ZN(n18861) );
  INV_X1 U13173 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15192) );
  NAND2_X1 U13174 ( .A1(n19161), .A2(n18959), .ZN(n18958) );
  OR2_X1 U13175 ( .A1(n19108), .A2(n19191), .ZN(n19010) );
  INV_X1 U13176 ( .A(n19068), .ZN(n19078) );
  INV_X1 U13177 ( .A(n19095), .ZN(n19092) );
  INV_X1 U13178 ( .A(n19089), .ZN(n19127) );
  OR2_X1 U13179 ( .A1(n19331), .A2(n19159), .ZN(n19182) );
  INV_X1 U13180 ( .A(n19254), .ZN(n19221) );
  INV_X1 U13181 ( .A(n19386), .ZN(n19239) );
  NAND2_X1 U13182 ( .A1(n19222), .A2(n19536), .ZN(n19291) );
  INV_X1 U13183 ( .A(n19418), .ZN(n19360) );
  OR2_X1 U13184 ( .A1(n19292), .A2(n19373), .ZN(n19414) );
  INV_X1 U13185 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19263) );
  INV_X1 U13186 ( .A(n19518), .ZN(n19441) );
  INV_X1 U13187 ( .A(n16975), .ZN(n16974) );
  NAND4_X1 U13188 ( .A1(n16131), .A2(P3_EBX_REG_31__SCAN_IN), .A3(n18391), 
        .A4(n16114), .ZN(n16481) );
  INV_X1 U13189 ( .A(n16443), .ZN(n16467) );
  AND2_X1 U13190 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16551), .ZN(n16545) );
  NOR2_X2 U13191 ( .A1(n16308), .A2(n15183), .ZN(n16676) );
  INV_X1 U13192 ( .A(n16856), .ZN(n16825) );
  NOR2_X1 U13193 ( .A1(n15247), .A2(n15246), .ZN(n16918) );
  INV_X1 U13194 ( .A(n16929), .ZN(n15426) );
  INV_X1 U13195 ( .A(n16953), .ZN(n16973) );
  NAND2_X1 U13196 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17367), .ZN(n17247) );
  INV_X1 U13197 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17559) );
  INV_X1 U13198 ( .A(n17293), .ZN(n17322) );
  OR2_X1 U13199 ( .A1(n16095), .A2(n17741), .ZN(n17411) );
  INV_X1 U13200 ( .A(n17699), .ZN(n17705) );
  INV_X1 U13201 ( .A(n17716), .ZN(n17680) );
  INV_X1 U13202 ( .A(n9746), .ZN(n17710) );
  NAND2_X1 U13203 ( .A1(n15979), .A2(n17721), .ZN(n17636) );
  INV_X1 U13204 ( .A(n17719), .ZN(n17703) );
  INV_X1 U13205 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n17988) );
  INV_X1 U13206 ( .A(n17788), .ZN(n18131) );
  INV_X1 U13207 ( .A(n17797), .ZN(n18156) );
  INV_X1 U13208 ( .A(n18336), .ZN(n18256) );
  INV_X1 U13209 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n20637) );
  BUF_X2 U13210 ( .A(n10461), .Z(n11013) );
  AOI22_X1 U13211 ( .A1(n11013), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10469), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10294) );
  AOI22_X1 U13212 ( .A1(n10334), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10470), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10293) );
  AND2_X2 U13213 ( .A1(n10295), .A2(n12921), .ZN(n10971) );
  AOI22_X1 U13214 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10570), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10292) );
  AOI22_X1 U13215 ( .A1(n10544), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10545), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10291) );
  NAND4_X1 U13216 ( .A1(n10294), .A2(n10293), .A3(n10292), .A4(n10291), .ZN(
        n10303) );
  AOI22_X1 U13217 ( .A1(n10550), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10435), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10301) );
  AOI22_X1 U13218 ( .A1(n10551), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10575), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10300) );
  AOI22_X1 U13219 ( .A1(n11014), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10552), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10299) );
  AOI22_X1 U13221 ( .A1(n10464), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10436), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10298) );
  NAND4_X1 U13222 ( .A1(n10301), .A2(n10300), .A3(n10299), .A4(n10298), .ZN(
        n10302) );
  AOI22_X1 U13223 ( .A1(n10469), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10435), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10307) );
  AOI22_X1 U13224 ( .A1(n10334), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10470), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10306) );
  AOI22_X1 U13225 ( .A1(n10544), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10436), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10305) );
  AOI22_X1 U13226 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10545), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10304) );
  NAND4_X1 U13227 ( .A1(n10307), .A2(n10306), .A3(n10305), .A4(n10304), .ZN(
        n10313) );
  INV_X1 U13228 ( .A(n10550), .ZN(n10462) );
  AOI22_X1 U13229 ( .A1(n11013), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10550), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10311) );
  AOI22_X1 U13230 ( .A1(n10551), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10575), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10310) );
  AOI22_X1 U13231 ( .A1(n10464), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10570), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10309) );
  AOI22_X1 U13232 ( .A1(n11014), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10552), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10308) );
  NAND4_X1 U13233 ( .A1(n10311), .A2(n10310), .A3(n10309), .A4(n10308), .ZN(
        n10312) );
  AOI22_X1 U13235 ( .A1(n11013), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10469), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10317) );
  AOI22_X1 U13236 ( .A1(n10334), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10470), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10316) );
  AOI22_X1 U13237 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10570), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10315) );
  AOI22_X1 U13238 ( .A1(n10544), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10545), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10314) );
  NAND4_X1 U13239 ( .A1(n10317), .A2(n10316), .A3(n10315), .A4(n10314), .ZN(
        n10323) );
  AOI22_X1 U13240 ( .A1(n10550), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10435), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10321) );
  AOI22_X1 U13241 ( .A1(n10551), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10575), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10320) );
  AOI22_X1 U13242 ( .A1(n11014), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10552), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10319) );
  AOI22_X1 U13243 ( .A1(n10464), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10436), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10318) );
  NAND4_X1 U13244 ( .A1(n10321), .A2(n10320), .A3(n10319), .A4(n10318), .ZN(
        n10322) );
  INV_X2 U13245 ( .A(n19878), .ZN(n10525) );
  AOI22_X1 U13246 ( .A1(n10334), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10544), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10327) );
  AOI22_X1 U13247 ( .A1(n10469), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10470), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10326) );
  AOI22_X1 U13248 ( .A1(n10550), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10570), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10325) );
  AOI22_X1 U13249 ( .A1(n10551), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10436), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10324) );
  NAND4_X1 U13250 ( .A1(n10327), .A2(n10326), .A3(n10325), .A4(n10324), .ZN(
        n10333) );
  AOI22_X1 U13251 ( .A1(n10903), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10971), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10331) );
  AOI22_X1 U13252 ( .A1(n10435), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10575), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10330) );
  AOI22_X1 U13253 ( .A1(n10464), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10545), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10329) );
  AOI22_X1 U13254 ( .A1(n10463), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10552), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10328) );
  NAND4_X1 U13255 ( .A1(n10331), .A2(n10330), .A3(n10329), .A4(n10328), .ZN(
        n10332) );
  AOI22_X1 U13256 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10469), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10338) );
  AOI22_X1 U13257 ( .A1(n10334), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10470), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10337) );
  AOI22_X1 U13258 ( .A1(n11044), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10552), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10336) );
  AOI22_X1 U13259 ( .A1(n10544), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10545), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10335) );
  NAND4_X1 U13260 ( .A1(n10338), .A2(n10337), .A3(n10336), .A4(n10335), .ZN(
        n10344) );
  AOI22_X1 U13261 ( .A1(n10550), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10435), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10342) );
  AOI22_X1 U13262 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10570), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10341) );
  AOI22_X1 U13263 ( .A1(n10551), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10575), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10340) );
  AOI22_X1 U13264 ( .A1(n10464), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10436), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10339) );
  NAND4_X1 U13265 ( .A1(n10342), .A2(n10341), .A3(n10340), .A4(n10339), .ZN(
        n10343) );
  NOR2_X1 U13266 ( .A1(n19873), .A2(n10396), .ZN(n11255) );
  NAND2_X1 U13267 ( .A1(n10550), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n10348) );
  NAND2_X1 U13268 ( .A1(n10464), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10347) );
  NAND2_X1 U13269 ( .A1(n10435), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10346) );
  NAND2_X1 U13270 ( .A1(n10436), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10345) );
  NAND2_X1 U13271 ( .A1(n10903), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10352) );
  NAND2_X1 U13272 ( .A1(n10334), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10351) );
  NAND2_X1 U13273 ( .A1(n10469), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10350) );
  NAND2_X1 U13274 ( .A1(n10470), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n10349) );
  NAND2_X1 U13275 ( .A1(n10544), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10356) );
  NAND2_X1 U13276 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n10355) );
  NAND2_X1 U13277 ( .A1(n10545), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n10354) );
  NAND2_X1 U13278 ( .A1(n10570), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10353) );
  NAND2_X1 U13279 ( .A1(n10551), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10360) );
  NAND2_X1 U13280 ( .A1(n10552), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n10359) );
  NAND2_X1 U13281 ( .A1(n10575), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n10358) );
  NAND2_X1 U13282 ( .A1(n10463), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n10357) );
  NAND4_X4 U13283 ( .A1(n10364), .A2(n10363), .A3(n10362), .A4(n10361), .ZN(
        n19839) );
  AOI22_X1 U13284 ( .A1(n11013), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10469), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10368) );
  AOI22_X1 U13285 ( .A1(n10334), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10470), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10367) );
  AOI22_X1 U13286 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10570), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10366) );
  AOI22_X1 U13287 ( .A1(n10544), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10545), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10365) );
  NAND4_X1 U13288 ( .A1(n10368), .A2(n10367), .A3(n10366), .A4(n10365), .ZN(
        n10374) );
  AOI22_X1 U13289 ( .A1(n10550), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10435), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10372) );
  AOI22_X1 U13290 ( .A1(n10551), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10575), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10371) );
  AOI22_X1 U13291 ( .A1(n11014), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10552), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10370) );
  AOI22_X1 U13292 ( .A1(n10464), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10436), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10369) );
  NAND4_X1 U13293 ( .A1(n10372), .A2(n10371), .A3(n10370), .A4(n10369), .ZN(
        n10373) );
  OR2_X4 U13294 ( .A1(n10374), .A2(n10373), .ZN(n19886) );
  NAND2_X1 U13295 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20465) );
  OAI21_X1 U13296 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(P1_STATE_REG_2__SCAN_IN), 
        .A(n20465), .ZN(n12379) );
  INV_X1 U13297 ( .A(n12379), .ZN(n10395) );
  NOR2_X2 U13298 ( .A1(n19863), .A2(n19858), .ZN(n12520) );
  NAND2_X1 U13299 ( .A1(n10464), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10378) );
  NAND2_X1 U13300 ( .A1(n10550), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10377) );
  NAND2_X1 U13301 ( .A1(n10469), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10376) );
  NAND2_X1 U13302 ( .A1(n10470), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10375) );
  NAND2_X1 U13303 ( .A1(n10334), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10382) );
  NAND2_X1 U13304 ( .A1(n10903), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10381) );
  NAND2_X1 U13305 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10380) );
  NAND2_X1 U13306 ( .A1(n10570), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10379) );
  AND4_X2 U13307 ( .A1(n10382), .A2(n10381), .A3(n10380), .A4(n10379), .ZN(
        n10393) );
  NAND2_X1 U13308 ( .A1(n10544), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10386) );
  NAND2_X1 U13309 ( .A1(n10551), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10385) );
  NAND2_X1 U13310 ( .A1(n10545), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10384) );
  NAND2_X1 U13311 ( .A1(n10436), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10383) );
  NAND2_X1 U13312 ( .A1(n10435), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10390) );
  NAND2_X1 U13313 ( .A1(n10575), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10389) );
  NAND2_X1 U13314 ( .A1(n11044), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10388) );
  NAND2_X1 U13315 ( .A1(n10552), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10387) );
  NAND4_X4 U13316 ( .A1(n10394), .A2(n10393), .A3(n10392), .A4(n10391), .ZN(
        n19853) );
  NOR2_X4 U13317 ( .A1(n19853), .A2(n19839), .ZN(n13056) );
  NAND3_X1 U13318 ( .A1(n12520), .A2(n13056), .A3(n9865), .ZN(n12511) );
  NAND2_X2 U13319 ( .A1(n10525), .A2(n19873), .ZN(n12899) );
  NAND2_X1 U13320 ( .A1(n19873), .A2(n19878), .ZN(n10397) );
  NAND2_X1 U13322 ( .A1(n9865), .A2(n19878), .ZN(n10398) );
  AND2_X1 U13323 ( .A1(n10398), .A2(n19886), .ZN(n11207) );
  INV_X1 U13324 ( .A(n11207), .ZN(n10399) );
  NAND2_X1 U13325 ( .A1(n10413), .A2(n12899), .ZN(n12488) );
  NAND2_X1 U13326 ( .A1(n12488), .A2(n14422), .ZN(n10410) );
  NAND2_X1 U13327 ( .A1(n19858), .A2(n19839), .ZN(n10401) );
  INV_X2 U13328 ( .A(n19853), .ZN(n12597) );
  NAND2_X1 U13329 ( .A1(n12597), .A2(n19839), .ZN(n20541) );
  NAND2_X1 U13330 ( .A1(n12485), .A2(n19853), .ZN(n12492) );
  INV_X1 U13331 ( .A(n12520), .ZN(n12917) );
  OAI211_X1 U13332 ( .C1(n20541), .C2(n12701), .A(n12492), .B(n12917), .ZN(
        n10402) );
  NOR2_X1 U13333 ( .A1(n12510), .A2(n10402), .ZN(n10405) );
  NAND2_X1 U13334 ( .A1(n12500), .A2(n12485), .ZN(n10404) );
  NAND2_X1 U13335 ( .A1(n12614), .A2(n20446), .ZN(n11214) );
  NAND2_X1 U13336 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10425) );
  OAI21_X1 U13337 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n10425), .ZN(n20178) );
  NAND2_X1 U13338 ( .A1(n15395), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10420) );
  OAI21_X1 U13339 ( .B1(n11214), .B2(n20178), .A(n10420), .ZN(n10407) );
  MUX2_X1 U13340 ( .A(n11214), .B(n11206), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n10409) );
  OR2_X1 U13341 ( .A1(n10410), .A2(n12597), .ZN(n10418) );
  NAND2_X1 U13342 ( .A1(n12520), .A2(n10525), .ZN(n12707) );
  NAND4_X1 U13343 ( .A1(n12707), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n12614), 
        .A4(n12492), .ZN(n10411) );
  NOR2_X1 U13344 ( .A1(n10411), .A2(n12510), .ZN(n10417) );
  OAI21_X1 U13345 ( .B1(n13056), .B2(n10412), .A(n12500), .ZN(n10416) );
  INV_X1 U13346 ( .A(n10413), .ZN(n10414) );
  NAND2_X1 U13347 ( .A1(n10414), .A2(n11129), .ZN(n10415) );
  NAND4_X1 U13348 ( .A1(n10418), .A2(n10417), .A3(n10416), .A4(n10415), .ZN(
        n10445) );
  INV_X1 U13349 ( .A(n10419), .ZN(n10422) );
  NAND2_X1 U13350 ( .A1(n10420), .A2(n12517), .ZN(n10421) );
  NAND2_X1 U13351 ( .A1(n10422), .A2(n10421), .ZN(n10423) );
  OR2_X1 U13352 ( .A1(n10536), .A2(n12516), .ZN(n10428) );
  INV_X1 U13353 ( .A(n10425), .ZN(n10424) );
  NAND2_X1 U13354 ( .A1(n10424), .A2(n20262), .ZN(n20211) );
  NAND2_X1 U13355 ( .A1(n10425), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10426) );
  NAND2_X1 U13356 ( .A1(n20211), .A2(n10426), .ZN(n19848) );
  INV_X1 U13357 ( .A(n11214), .ZN(n10539) );
  AOI22_X1 U13358 ( .A1(n19848), .A2(n10539), .B1(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15395), .ZN(n10427) );
  AOI22_X1 U13359 ( .A1(n11013), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11218), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10434) );
  AOI22_X1 U13360 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10433) );
  AOI22_X1 U13361 ( .A1(n11038), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10570), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10432) );
  AOI22_X1 U13362 ( .A1(n10448), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11039), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10431) );
  NAND4_X1 U13363 ( .A1(n10434), .A2(n10433), .A3(n10432), .A4(n10431), .ZN(
        n10442) );
  AOI22_X1 U13364 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10440) );
  AOI22_X1 U13365 ( .A1(n10454), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10453), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10439) );
  AOI22_X1 U13366 ( .A1(n11014), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10438) );
  INV_X1 U13367 ( .A(n10436), .ZN(n10553) );
  AOI22_X1 U13368 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10437) );
  NAND4_X1 U13369 ( .A1(n10440), .A2(n10439), .A3(n10438), .A4(n10437), .ZN(
        n10441) );
  INV_X1 U13370 ( .A(n10542), .ZN(n10493) );
  AOI22_X1 U13371 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10493), .B2(n10443), .ZN(n10444) );
  INV_X1 U13372 ( .A(n10445), .ZN(n10446) );
  AOI22_X1 U13373 ( .A1(n11013), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11218), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10452) );
  AOI22_X1 U13374 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10451) );
  AOI22_X1 U13375 ( .A1(n11038), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10570), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10450) );
  AOI22_X1 U13376 ( .A1(n10448), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9610), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10449) );
  NAND4_X1 U13377 ( .A1(n10452), .A2(n10451), .A3(n10450), .A4(n10449), .ZN(
        n10460) );
  AOI22_X1 U13378 ( .A1(n10550), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10458) );
  AOI22_X1 U13379 ( .A1(n10454), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10453), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10457) );
  AOI22_X1 U13380 ( .A1(n11014), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10456) );
  AOI22_X1 U13381 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10455) );
  NAND4_X1 U13382 ( .A1(n10458), .A2(n10457), .A3(n10456), .A4(n10455), .ZN(
        n10459) );
  NAND2_X1 U13383 ( .A1(n12701), .A2(n11128), .ZN(n10479) );
  NOR2_X1 U13384 ( .A1(n10543), .A2(n11128), .ZN(n10482) );
  AOI22_X1 U13385 ( .A1(n10903), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9618), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10468) );
  AOI22_X1 U13386 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10467) );
  AOI22_X1 U13387 ( .A1(n11014), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10466) );
  AOI22_X1 U13388 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11039), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10465) );
  NAND4_X1 U13389 ( .A1(n10468), .A2(n10467), .A3(n10466), .A4(n10465), .ZN(
        n10476) );
  AOI22_X1 U13390 ( .A1(n10448), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10454), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10474) );
  AOI22_X1 U13391 ( .A1(n11218), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10473) );
  AOI22_X1 U13392 ( .A1(n10447), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10570), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10472) );
  AOI22_X1 U13393 ( .A1(n10453), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10471) );
  NAND4_X1 U13394 ( .A1(n10474), .A2(n10473), .A3(n10472), .A4(n10471), .ZN(
        n10475) );
  MUX2_X1 U13395 ( .A(n11124), .B(n10482), .S(n11074), .Z(n10477) );
  INV_X1 U13396 ( .A(n10477), .ZN(n10478) );
  INV_X1 U13397 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10481) );
  AOI21_X1 U13398 ( .B1(n12485), .B2(n11074), .A(n20446), .ZN(n10480) );
  OAI211_X1 U13399 ( .C1(n11187), .C2(n10481), .A(n10480), .B(n10479), .ZN(
        n10523) );
  NAND2_X1 U13400 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10496) );
  INV_X1 U13401 ( .A(n10482), .ZN(n10495) );
  AOI22_X1 U13402 ( .A1(n10454), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U13403 ( .A1(n10448), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9618), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10485) );
  AOI22_X1 U13404 ( .A1(n11038), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10484) );
  AOI22_X1 U13405 ( .A1(n11014), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10483) );
  NAND4_X1 U13406 ( .A1(n10486), .A2(n10485), .A3(n10484), .A4(n10483), .ZN(
        n10492) );
  AOI22_X1 U13407 ( .A1(n10903), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11218), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10490) );
  AOI22_X1 U13408 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10453), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10489) );
  AOI22_X1 U13409 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11039), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10488) );
  AOI22_X1 U13410 ( .A1(n11219), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10487) );
  NAND4_X1 U13411 ( .A1(n10490), .A2(n10489), .A3(n10488), .A4(n10487), .ZN(
        n10491) );
  NAND2_X1 U13412 ( .A1(n10493), .A2(n11073), .ZN(n10494) );
  INV_X1 U13413 ( .A(n19960), .ZN(n10499) );
  INV_X1 U13414 ( .A(n10497), .ZN(n10498) );
  INV_X1 U13415 ( .A(n11073), .ZN(n10501) );
  OR2_X1 U13416 ( .A1(n10543), .A2(n10501), .ZN(n10502) );
  INV_X1 U13417 ( .A(n10503), .ZN(n10504) );
  NAND2_X1 U13418 ( .A1(n9818), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10587) );
  XNOR2_X1 U13419 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12877) );
  AOI21_X1 U13420 ( .B1(n10532), .B2(n12877), .A(n11243), .ZN(n10510) );
  NAND2_X1 U13421 ( .A1(n10508), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n10509) );
  OAI211_X1 U13422 ( .C1(n10587), .C2(n12516), .A(n10510), .B(n10509), .ZN(
        n10511) );
  INV_X1 U13423 ( .A(n10511), .ZN(n10513) );
  NAND2_X1 U13424 ( .A1(n11243), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10534) );
  INV_X1 U13425 ( .A(n10534), .ZN(n10512) );
  NAND2_X1 U13426 ( .A1(n12938), .A2(n10773), .ZN(n10522) );
  AOI22_X1 U13427 ( .A1(n10508), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20448), .ZN(n10520) );
  INV_X1 U13428 ( .A(n10587), .ZN(n10518) );
  NAND2_X1 U13429 ( .A1(n10518), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10519) );
  AND2_X1 U13430 ( .A1(n10520), .A2(n10519), .ZN(n10521) );
  NAND2_X1 U13431 ( .A1(n10522), .A2(n10521), .ZN(n12649) );
  AOI21_X1 U13432 ( .B1(n19922), .B2(n10525), .A(n20448), .ZN(n12674) );
  NAND2_X1 U13433 ( .A1(n19961), .A2(n10773), .ZN(n10531) );
  NAND2_X1 U13434 ( .A1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20448), .ZN(
        n10528) );
  NAND2_X1 U13435 ( .A1(n10508), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n10527) );
  OAI211_X1 U13436 ( .C1(n10587), .C2(n12617), .A(n10528), .B(n10527), .ZN(
        n10529) );
  INV_X1 U13437 ( .A(n10529), .ZN(n10530) );
  NAND2_X1 U13438 ( .A1(n10531), .A2(n10530), .ZN(n12673) );
  NAND2_X1 U13439 ( .A1(n12674), .A2(n12673), .ZN(n12676) );
  OR2_X1 U13440 ( .A1(n12673), .A2(n11028), .ZN(n10533) );
  NAND2_X1 U13441 ( .A1(n12676), .A2(n10533), .ZN(n12648) );
  NAND2_X1 U13442 ( .A1(n12649), .A2(n12648), .ZN(n12647) );
  INV_X1 U13443 ( .A(n12647), .ZN(n12872) );
  NAND2_X1 U13444 ( .A1(n12873), .A2(n12872), .ZN(n12871) );
  OR2_X1 U13445 ( .A1(n10536), .A2(n12926), .ZN(n10541) );
  NAND3_X1 U13446 ( .A1(n20528), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20088) );
  INV_X1 U13447 ( .A(n20088), .ZN(n20094) );
  NAND2_X1 U13448 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20094), .ZN(
        n20085) );
  NAND2_X1 U13449 ( .A1(n20528), .A2(n20085), .ZN(n10538) );
  NAND3_X1 U13450 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20388) );
  INV_X1 U13451 ( .A(n20388), .ZN(n10537) );
  NAND2_X1 U13452 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n10537), .ZN(
        n20384) );
  AOI22_X1 U13453 ( .A1(n10539), .A2(n19844), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15395), .ZN(n10540) );
  AOI22_X1 U13454 ( .A1(n10903), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11218), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10549) );
  AOI22_X1 U13455 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10548) );
  AOI22_X1 U13456 ( .A1(n11038), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10570), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10547) );
  AOI22_X1 U13457 ( .A1(n10448), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11039), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10546) );
  NAND4_X1 U13458 ( .A1(n10549), .A2(n10548), .A3(n10547), .A4(n10546), .ZN(
        n10559) );
  AOI22_X1 U13459 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10557) );
  AOI22_X1 U13460 ( .A1(n10454), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10453), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10556) );
  AOI22_X1 U13461 ( .A1(n11014), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10555) );
  INV_X2 U13462 ( .A(n10553), .ZN(n12914) );
  AOI22_X1 U13463 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10554) );
  NAND4_X1 U13464 ( .A1(n10557), .A2(n10556), .A3(n10555), .A4(n10554), .ZN(
        n10558) );
  INV_X1 U13465 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10560) );
  OAI22_X1 U13466 ( .A1(n11201), .A2(n11084), .B1(n10560), .B2(n11187), .ZN(
        n10561) );
  INV_X1 U13467 ( .A(n10561), .ZN(n10562) );
  NAND2_X1 U13468 ( .A1(n20524), .A2(n10773), .ZN(n10569) );
  INV_X1 U13469 ( .A(n10589), .ZN(n10591) );
  INV_X1 U13470 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n19692) );
  NAND2_X1 U13471 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10563) );
  NAND2_X1 U13472 ( .A1(n19692), .A2(n10563), .ZN(n10564) );
  NAND2_X1 U13473 ( .A1(n10591), .A2(n10564), .ZN(n19689) );
  AOI22_X1 U13474 ( .A1(n19689), .A2(n12280), .B1(n11243), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10566) );
  NAND2_X1 U13475 ( .A1(n11237), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n10565) );
  OAI211_X1 U13476 ( .C1(n10587), .C2(n12926), .A(n10566), .B(n10565), .ZN(
        n10567) );
  INV_X1 U13477 ( .A(n10567), .ZN(n10568) );
  NAND2_X1 U13478 ( .A1(n10601), .A2(n19837), .ZN(n10584) );
  AOI22_X1 U13479 ( .A1(n10903), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11218), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10574) );
  AOI22_X1 U13480 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10573) );
  AOI22_X1 U13481 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n11038), .B1(
        n11219), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10572) );
  AOI22_X1 U13482 ( .A1(n10448), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11039), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10571) );
  NAND4_X1 U13483 ( .A1(n10574), .A2(n10573), .A3(n10572), .A4(n10571), .ZN(
        n10581) );
  AOI22_X1 U13484 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n9618), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10579) );
  AOI22_X1 U13485 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n10454), .B1(
        n10453), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10578) );
  AOI22_X1 U13486 ( .A1(n11014), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10577) );
  AOI22_X1 U13487 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10576) );
  NAND4_X1 U13488 ( .A1(n10579), .A2(n10578), .A3(n10577), .A4(n10576), .ZN(
        n10580) );
  INV_X1 U13489 ( .A(n11098), .ZN(n10583) );
  INV_X1 U13490 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10582) );
  OAI22_X1 U13491 ( .A1(n11201), .A2(n10583), .B1(n10582), .B2(n11187), .ZN(
        n10598) );
  XNOR2_X1 U13492 ( .A(n10584), .B(n10598), .ZN(n11090) );
  INV_X1 U13493 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12637) );
  NAND2_X1 U13494 ( .A1(n20448), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10586) );
  NAND2_X1 U13495 ( .A1(n10508), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n10585) );
  OAI211_X1 U13496 ( .C1(n10587), .C2(n12637), .A(n10586), .B(n10585), .ZN(
        n10588) );
  NAND2_X1 U13497 ( .A1(n10588), .A2(n11028), .ZN(n10595) );
  INV_X1 U13498 ( .A(n10614), .ZN(n10593) );
  INV_X1 U13499 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10590) );
  NAND2_X1 U13500 ( .A1(n10591), .A2(n10590), .ZN(n10592) );
  NAND2_X1 U13501 ( .A1(n10593), .A2(n10592), .ZN(n19792) );
  NAND2_X1 U13502 ( .A1(n19792), .A2(n12280), .ZN(n10594) );
  NAND2_X1 U13503 ( .A1(n10595), .A2(n10594), .ZN(n10596) );
  AOI21_X1 U13504 ( .B1(n11090), .B2(n10773), .A(n10596), .ZN(n12971) );
  INV_X1 U13505 ( .A(n10598), .ZN(n10599) );
  AOI22_X1 U13506 ( .A1(n10903), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11218), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10605) );
  AOI22_X1 U13507 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10604) );
  AOI22_X1 U13508 ( .A1(n11038), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11219), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10603) );
  AOI22_X1 U13509 ( .A1(n10448), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11039), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10602) );
  NAND4_X1 U13510 ( .A1(n10605), .A2(n10604), .A3(n10603), .A4(n10602), .ZN(
        n10611) );
  AOI22_X1 U13511 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10609) );
  AOI22_X1 U13512 ( .A1(n10454), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10453), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10608) );
  AOI22_X1 U13513 ( .A1(n11014), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10607) );
  AOI22_X1 U13514 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10606) );
  NAND4_X1 U13515 ( .A1(n10609), .A2(n10608), .A3(n10607), .A4(n10606), .ZN(
        n10610) );
  INV_X1 U13516 ( .A(n11116), .ZN(n10613) );
  INV_X1 U13517 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10612) );
  OAI22_X1 U13518 ( .A1(n11201), .A2(n10613), .B1(n10612), .B2(n11187), .ZN(
        n10619) );
  XNOR2_X1 U13519 ( .A(n10618), .B(n10619), .ZN(n11097) );
  INV_X1 U13520 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n10616) );
  OAI21_X1 U13521 ( .B1(n10614), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n10632), .ZN(n19673) );
  AOI22_X1 U13522 ( .A1(n19673), .A2(n12280), .B1(n11243), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10615) );
  OAI21_X1 U13523 ( .B1(n10999), .B2(n10616), .A(n10615), .ZN(n10617) );
  AOI22_X1 U13524 ( .A1(n10903), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11218), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10623) );
  AOI22_X1 U13525 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10622) );
  AOI22_X1 U13526 ( .A1(n11038), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11219), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10621) );
  AOI22_X1 U13527 ( .A1(n10448), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11039), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10620) );
  NAND4_X1 U13528 ( .A1(n10623), .A2(n10622), .A3(n10621), .A4(n10620), .ZN(
        n10629) );
  AOI22_X1 U13529 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10627) );
  AOI22_X1 U13530 ( .A1(n10454), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10453), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10626) );
  AOI22_X1 U13531 ( .A1(n11014), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10625) );
  AOI22_X1 U13532 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10624) );
  NAND4_X1 U13533 ( .A1(n10627), .A2(n10626), .A3(n10625), .A4(n10624), .ZN(
        n10628) );
  INV_X1 U13534 ( .A(n11115), .ZN(n10631) );
  INV_X1 U13535 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10630) );
  OAI22_X1 U13536 ( .A1(n11201), .A2(n10631), .B1(n11187), .B2(n10630), .ZN(
        n10640) );
  XNOR2_X1 U13537 ( .A(n10641), .B(n10640), .ZN(n11107) );
  NAND2_X1 U13538 ( .A1(n11107), .A2(n10773), .ZN(n10639) );
  INV_X1 U13539 ( .A(n11243), .ZN(n10636) );
  NAND2_X1 U13540 ( .A1(n10632), .A2(n19654), .ZN(n10634) );
  INV_X1 U13541 ( .A(n10645), .ZN(n10633) );
  NAND2_X1 U13542 ( .A1(n10634), .A2(n10633), .ZN(n19656) );
  NAND2_X1 U13543 ( .A1(n19656), .A2(n12280), .ZN(n10635) );
  OAI21_X1 U13544 ( .B1(n19654), .B2(n10636), .A(n10635), .ZN(n10637) );
  AOI21_X1 U13545 ( .B1(n11237), .B2(P1_EAX_REG_6__SCAN_IN), .A(n10637), .ZN(
        n10638) );
  NAND2_X1 U13546 ( .A1(n10639), .A2(n10638), .ZN(n13043) );
  INV_X1 U13547 ( .A(n13042), .ZN(n10650) );
  INV_X1 U13548 ( .A(n11128), .ZN(n10643) );
  INV_X1 U13549 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10642) );
  OAI22_X1 U13550 ( .A1(n11201), .A2(n10643), .B1(n10642), .B2(n11187), .ZN(
        n10644) );
  INV_X1 U13551 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n10647) );
  OAI21_X1 U13552 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n10645), .A(
        n10666), .ZN(n19642) );
  AOI22_X1 U13553 ( .A1(n12280), .A2(n19642), .B1(n11243), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10646) );
  OAI21_X1 U13554 ( .B1(n10999), .B2(n10647), .A(n10646), .ZN(n10648) );
  AOI22_X1 U13555 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11218), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10654) );
  AOI22_X1 U13556 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10653) );
  AOI22_X1 U13557 ( .A1(n11014), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10652) );
  AOI22_X1 U13558 ( .A1(n10454), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10453), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10651) );
  NAND4_X1 U13559 ( .A1(n10654), .A2(n10653), .A3(n10652), .A4(n10651), .ZN(
        n10660) );
  AOI22_X1 U13560 ( .A1(n10448), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10658) );
  AOI22_X1 U13561 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11219), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10657) );
  AOI22_X1 U13562 ( .A1(n10447), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11039), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10656) );
  AOI22_X1 U13563 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10655) );
  NAND4_X1 U13564 ( .A1(n10658), .A2(n10657), .A3(n10656), .A4(n10655), .ZN(
        n10659) );
  OAI21_X1 U13565 ( .B1(n10660), .B2(n10659), .A(n10773), .ZN(n10664) );
  INV_X1 U13566 ( .A(n10666), .ZN(n10661) );
  XNOR2_X1 U13567 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n10661), .ZN(
        n13217) );
  AOI22_X1 U13568 ( .A1(n12280), .A2(n13217), .B1(n11243), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10663) );
  NAND2_X1 U13569 ( .A1(n10508), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n10662) );
  XOR2_X1 U13570 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n10682), .Z(n19631) );
  INV_X1 U13571 ( .A(n19631), .ZN(n10681) );
  AOI22_X1 U13572 ( .A1(n10903), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10670) );
  AOI22_X1 U13573 ( .A1(n11224), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10453), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10669) );
  AOI22_X1 U13574 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11039), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10668) );
  AOI22_X1 U13575 ( .A1(n11014), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10667) );
  NAND4_X1 U13576 ( .A1(n10670), .A2(n10669), .A3(n10668), .A4(n10667), .ZN(
        n10676) );
  AOI22_X1 U13577 ( .A1(n10454), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9618), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10674) );
  AOI22_X1 U13578 ( .A1(n11038), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11218), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10673) );
  AOI22_X1 U13579 ( .A1(n10448), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11219), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10672) );
  AOI22_X1 U13580 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10671) );
  NAND4_X1 U13581 ( .A1(n10674), .A2(n10673), .A3(n10672), .A4(n10671), .ZN(
        n10675) );
  OAI21_X1 U13582 ( .B1(n10676), .B2(n10675), .A(n10773), .ZN(n10679) );
  NAND2_X1 U13583 ( .A1(n10508), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n10678) );
  NAND2_X1 U13584 ( .A1(n11243), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10677) );
  NAND3_X1 U13585 ( .A1(n10679), .A2(n10678), .A3(n10677), .ZN(n10680) );
  AOI21_X1 U13586 ( .B1(n10681), .B2(n12280), .A(n10680), .ZN(n13181) );
  XNOR2_X1 U13587 ( .A(n10699), .B(n10698), .ZN(n14215) );
  NAND2_X1 U13588 ( .A1(n14215), .A2(n12280), .ZN(n10697) );
  AOI22_X1 U13589 ( .A1(n10448), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11218), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10686) );
  AOI22_X1 U13590 ( .A1(n10447), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10685) );
  AOI22_X1 U13591 ( .A1(n10463), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10684) );
  AOI22_X1 U13592 ( .A1(n10454), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10453), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10683) );
  NAND4_X1 U13593 ( .A1(n10686), .A2(n10685), .A3(n10684), .A4(n10683), .ZN(
        n10692) );
  AOI22_X1 U13594 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11226), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10690) );
  AOI22_X1 U13595 ( .A1(n10461), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9610), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10689) );
  AOI22_X1 U13596 ( .A1(n11038), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11219), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10688) );
  AOI22_X1 U13597 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10687) );
  NAND4_X1 U13598 ( .A1(n10690), .A2(n10689), .A3(n10688), .A4(n10687), .ZN(
        n10691) );
  OAI21_X1 U13599 ( .B1(n10692), .B2(n10691), .A(n10773), .ZN(n10695) );
  NAND2_X1 U13600 ( .A1(n10508), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n10694) );
  NAND2_X1 U13601 ( .A1(n11243), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10693) );
  AND3_X1 U13602 ( .A1(n10695), .A2(n10694), .A3(n10693), .ZN(n10696) );
  NAND2_X1 U13603 ( .A1(n10697), .A2(n10696), .ZN(n13397) );
  NAND2_X1 U13604 ( .A1(n10508), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n10702) );
  OAI21_X1 U13605 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n10700), .A(
        n10714), .ZN(n15579) );
  AOI22_X1 U13606 ( .A1(n12280), .A2(n15579), .B1(n11243), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10701) );
  NAND2_X1 U13607 ( .A1(n10702), .A2(n10701), .ZN(n13500) );
  AOI22_X1 U13608 ( .A1(n10461), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11226), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10706) );
  AOI22_X1 U13609 ( .A1(n10448), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11218), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10705) );
  AOI22_X1 U13610 ( .A1(n11014), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10704) );
  AOI22_X1 U13611 ( .A1(n11224), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10453), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10703) );
  NAND4_X1 U13612 ( .A1(n10706), .A2(n10705), .A3(n10704), .A4(n10703), .ZN(
        n10712) );
  AOI22_X1 U13613 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10710) );
  AOI22_X1 U13614 ( .A1(n11038), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11219), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10709) );
  AOI22_X1 U13615 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(n9610), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10708) );
  AOI22_X1 U13616 ( .A1(n10454), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10707) );
  NAND4_X1 U13617 ( .A1(n10710), .A2(n10709), .A3(n10708), .A4(n10707), .ZN(
        n10711) );
  OR2_X1 U13618 ( .A1(n10712), .A2(n10711), .ZN(n10713) );
  AND2_X1 U13619 ( .A1(n10773), .A2(n10713), .ZN(n15528) );
  AOI21_X1 U13620 ( .B1(n20629), .B2(n10715), .A(n10747), .ZN(n14208) );
  OR2_X1 U13621 ( .A1(n14208), .A2(n11028), .ZN(n10730) );
  AOI22_X1 U13622 ( .A1(n11013), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9618), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10719) );
  AOI22_X1 U13623 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10718) );
  AOI22_X1 U13624 ( .A1(n10448), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11218), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10717) );
  AOI22_X1 U13625 ( .A1(n11014), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10716) );
  NAND4_X1 U13626 ( .A1(n10719), .A2(n10718), .A3(n10717), .A4(n10716), .ZN(
        n10725) );
  AOI22_X1 U13627 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10723) );
  AOI22_X1 U13628 ( .A1(n10454), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11219), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10722) );
  AOI22_X1 U13629 ( .A1(n10447), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11039), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10721) );
  AOI22_X1 U13630 ( .A1(n10453), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10720) );
  NAND4_X1 U13631 ( .A1(n10723), .A2(n10722), .A3(n10721), .A4(n10720), .ZN(
        n10724) );
  OAI21_X1 U13632 ( .B1(n10725), .B2(n10724), .A(n10773), .ZN(n10728) );
  NAND2_X1 U13633 ( .A1(n10508), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n10727) );
  NAND2_X1 U13634 ( .A1(n11243), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10726) );
  AND3_X1 U13635 ( .A1(n10728), .A2(n10727), .A3(n10726), .ZN(n10729) );
  NAND2_X1 U13636 ( .A1(n10730), .A2(n10729), .ZN(n13505) );
  XOR2_X1 U13637 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n10731), .Z(
        n15565) );
  AOI22_X1 U13638 ( .A1(n10454), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10453), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10735) );
  AOI22_X1 U13639 ( .A1(n10447), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11219), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10734) );
  AOI22_X1 U13640 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11039), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10733) );
  AOI22_X1 U13641 ( .A1(n11044), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10732) );
  NAND4_X1 U13642 ( .A1(n10735), .A2(n10734), .A3(n10733), .A4(n10732), .ZN(
        n10741) );
  AOI22_X1 U13643 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n9618), .B1(
        n10448), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10739) );
  AOI22_X1 U13644 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11037), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10738) );
  AOI22_X1 U13645 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n11226), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10737) );
  AOI22_X1 U13646 ( .A1(n11218), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10736) );
  NAND4_X1 U13647 ( .A1(n10739), .A2(n10738), .A3(n10737), .A4(n10736), .ZN(
        n10740) );
  OAI21_X1 U13648 ( .B1(n10741), .B2(n10740), .A(n10773), .ZN(n10744) );
  NAND2_X1 U13649 ( .A1(n11237), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n10743) );
  NAND2_X1 U13650 ( .A1(n11243), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10742) );
  AND3_X1 U13651 ( .A1(n10744), .A2(n10743), .A3(n10742), .ZN(n10745) );
  OAI21_X1 U13652 ( .B1(n15565), .B2(n11028), .A(n10745), .ZN(n13520) );
  OR2_X1 U13653 ( .A1(n10747), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10750) );
  INV_X1 U13654 ( .A(n10794), .ZN(n10749) );
  NAND2_X1 U13655 ( .A1(n10750), .A2(n10749), .ZN(n14199) );
  AOI22_X1 U13656 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11226), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10754) );
  AOI22_X1 U13657 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10448), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10753) );
  AOI22_X1 U13658 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11218), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10752) );
  AOI22_X1 U13659 ( .A1(n11044), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10751) );
  NAND4_X1 U13660 ( .A1(n10754), .A2(n10753), .A3(n10752), .A4(n10751), .ZN(
        n10760) );
  AOI22_X1 U13661 ( .A1(n11038), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11219), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10758) );
  AOI22_X1 U13662 ( .A1(n10454), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10453), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10757) );
  AOI22_X1 U13663 ( .A1(n10447), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11039), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10756) );
  AOI22_X1 U13664 ( .A1(n11224), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10755) );
  NAND4_X1 U13665 ( .A1(n10758), .A2(n10757), .A3(n10756), .A4(n10755), .ZN(
        n10759) );
  OAI21_X1 U13666 ( .B1(n10760), .B2(n10759), .A(n10773), .ZN(n10763) );
  NAND2_X1 U13667 ( .A1(n11237), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n10762) );
  NAND2_X1 U13668 ( .A1(n11243), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10761) );
  NAND3_X1 U13669 ( .A1(n10763), .A2(n10762), .A3(n10761), .ZN(n10764) );
  AOI21_X1 U13670 ( .B1(n14199), .B2(n12280), .A(n10764), .ZN(n13528) );
  AOI22_X1 U13671 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11226), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10768) );
  AOI22_X1 U13672 ( .A1(n10454), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10453), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10767) );
  AOI22_X1 U13673 ( .A1(n10447), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11219), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10766) );
  AOI22_X1 U13674 ( .A1(n11044), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10765) );
  NAND4_X1 U13675 ( .A1(n10768), .A2(n10767), .A3(n10766), .A4(n10765), .ZN(
        n10775) );
  AOI22_X1 U13676 ( .A1(n10448), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10772) );
  AOI22_X1 U13677 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11218), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10771) );
  AOI22_X1 U13678 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(n9610), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10770) );
  AOI22_X1 U13679 ( .A1(n11224), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10769) );
  NAND4_X1 U13680 ( .A1(n10772), .A2(n10771), .A3(n10770), .A4(n10769), .ZN(
        n10774) );
  OAI21_X1 U13681 ( .B1(n10775), .B2(n10774), .A(n10773), .ZN(n10779) );
  NAND2_X1 U13682 ( .A1(n11237), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n10778) );
  XOR2_X1 U13683 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n10794), .Z(
        n15559) );
  INV_X1 U13684 ( .A(n15559), .ZN(n10776) );
  AOI22_X1 U13685 ( .A1(n11243), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n12280), .B2(n10776), .ZN(n10777) );
  INV_X1 U13686 ( .A(n14422), .ZN(n12612) );
  AOI22_X1 U13687 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11218), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10784) );
  AOI22_X1 U13688 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10783) );
  AOI22_X1 U13689 ( .A1(n11044), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10782) );
  AOI22_X1 U13690 ( .A1(n10454), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10453), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10781) );
  NAND4_X1 U13691 ( .A1(n10784), .A2(n10783), .A3(n10782), .A4(n10781), .ZN(
        n10790) );
  AOI22_X1 U13692 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10788) );
  AOI22_X1 U13693 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10787) );
  AOI22_X1 U13694 ( .A1(n10448), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11219), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10786) );
  AOI22_X1 U13695 ( .A1(n11039), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10785) );
  NAND4_X1 U13696 ( .A1(n10788), .A2(n10787), .A3(n10786), .A4(n10785), .ZN(
        n10789) );
  NOR2_X1 U13697 ( .A1(n10790), .A2(n10789), .ZN(n10793) );
  OAI21_X1 U13698 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n15498), .A(n11028), 
        .ZN(n10791) );
  AOI21_X1 U13699 ( .B1(n11237), .B2(P1_EAX_REG_16__SCAN_IN), .A(n10791), .ZN(
        n10792) );
  OAI21_X1 U13700 ( .B1(n11239), .B2(n10793), .A(n10792), .ZN(n10796) );
  XNOR2_X1 U13701 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B(n10797), .ZN(
        n15496) );
  NAND2_X1 U13702 ( .A1(n15496), .A2(n12280), .ZN(n10795) );
  NAND2_X1 U13703 ( .A1(n10796), .A2(n10795), .ZN(n14022) );
  XOR2_X1 U13704 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n10810), .Z(
        n15554) );
  AOI22_X1 U13705 ( .A1(n10508), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n11243), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10809) );
  AOI22_X1 U13706 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11226), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10801) );
  AOI22_X1 U13707 ( .A1(n10454), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10800) );
  AOI22_X1 U13708 ( .A1(n11044), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10799) );
  AOI22_X1 U13709 ( .A1(n10544), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11039), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10798) );
  NAND4_X1 U13710 ( .A1(n10801), .A2(n10800), .A3(n10799), .A4(n10798), .ZN(
        n10807) );
  AOI22_X1 U13711 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10805) );
  AOI22_X1 U13712 ( .A1(n11038), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11219), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10804) );
  AOI22_X1 U13713 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10453), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10803) );
  AOI22_X1 U13714 ( .A1(n11218), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10802) );
  NAND4_X1 U13715 ( .A1(n10805), .A2(n10804), .A3(n10803), .A4(n10802), .ZN(
        n10806) );
  OAI21_X1 U13716 ( .B1(n10807), .B2(n10806), .A(n11051), .ZN(n10808) );
  OAI211_X1 U13717 ( .C1(n15554), .C2(n11028), .A(n10809), .B(n10808), .ZN(
        n13957) );
  XNOR2_X1 U13718 ( .A(n10840), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15490) );
  NAND2_X1 U13719 ( .A1(n15490), .A2(n12280), .ZN(n10825) );
  AOI22_X1 U13720 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11218), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10814) );
  AOI22_X1 U13721 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10813) );
  AOI22_X1 U13722 ( .A1(n11038), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11219), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10812) );
  AOI22_X1 U13723 ( .A1(n10544), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11039), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10811) );
  NAND4_X1 U13724 ( .A1(n10814), .A2(n10813), .A3(n10812), .A4(n10811), .ZN(
        n10820) );
  AOI22_X1 U13725 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10818) );
  AOI22_X1 U13726 ( .A1(n10454), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10453), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10817) );
  AOI22_X1 U13727 ( .A1(n11044), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10816) );
  AOI22_X1 U13728 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10815) );
  NAND4_X1 U13729 ( .A1(n10818), .A2(n10817), .A3(n10816), .A4(n10815), .ZN(
        n10819) );
  NOR2_X1 U13730 ( .A1(n10820), .A2(n10819), .ZN(n10823) );
  AOI21_X1 U13731 ( .B1(n15487), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10821) );
  AOI21_X1 U13732 ( .B1(n11237), .B2(P1_EAX_REG_18__SCAN_IN), .A(n10821), .ZN(
        n10822) );
  OAI21_X1 U13733 ( .B1(n11239), .B2(n10823), .A(n10822), .ZN(n10824) );
  NAND2_X1 U13734 ( .A1(n10825), .A2(n10824), .ZN(n14014) );
  AOI22_X1 U13735 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11218), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10829) );
  AOI22_X1 U13736 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10828) );
  AOI22_X1 U13737 ( .A1(n11044), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10827) );
  AOI22_X1 U13738 ( .A1(n10551), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10575), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10826) );
  NAND4_X1 U13739 ( .A1(n10829), .A2(n10828), .A3(n10827), .A4(n10826), .ZN(
        n10835) );
  AOI22_X1 U13740 ( .A1(n10544), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10833) );
  AOI22_X1 U13741 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10832) );
  AOI22_X1 U13742 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10831) );
  AOI22_X1 U13743 ( .A1(n11219), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9610), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10830) );
  NAND4_X1 U13744 ( .A1(n10833), .A2(n10832), .A3(n10831), .A4(n10830), .ZN(
        n10834) );
  NOR2_X1 U13745 ( .A1(n10835), .A2(n10834), .ZN(n10839) );
  NAND2_X1 U13746 ( .A1(n20448), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10836) );
  NAND2_X1 U13747 ( .A1(n11028), .A2(n10836), .ZN(n10837) );
  AOI21_X1 U13748 ( .B1(n11237), .B2(P1_EAX_REG_19__SCAN_IN), .A(n10837), .ZN(
        n10838) );
  OAI21_X1 U13749 ( .B1(n11239), .B2(n10839), .A(n10838), .ZN(n10843) );
  OAI21_X1 U13750 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n10841), .A(
        n10873), .ZN(n15552) );
  OR2_X1 U13751 ( .A1(n11028), .A2(n15552), .ZN(n10842) );
  NAND2_X1 U13752 ( .A1(n10843), .A2(n10842), .ZN(n14012) );
  AOI22_X1 U13753 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11218), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10847) );
  AOI22_X1 U13754 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10846) );
  AOI22_X1 U13755 ( .A1(n11038), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11219), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10845) );
  AOI22_X1 U13756 ( .A1(n10448), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11039), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10844) );
  NAND4_X1 U13757 ( .A1(n10847), .A2(n10846), .A3(n10845), .A4(n10844), .ZN(
        n10853) );
  AOI22_X1 U13758 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n9618), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10851) );
  AOI22_X1 U13759 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n10551), .B1(
        n10453), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10850) );
  AOI22_X1 U13760 ( .A1(n11044), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10849) );
  AOI22_X1 U13761 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10848) );
  NAND4_X1 U13762 ( .A1(n10851), .A2(n10850), .A3(n10849), .A4(n10848), .ZN(
        n10852) );
  NOR2_X1 U13763 ( .A1(n10853), .A2(n10852), .ZN(n10856) );
  INV_X1 U13764 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15476) );
  AOI21_X1 U13765 ( .B1(n15476), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10854) );
  AOI21_X1 U13766 ( .B1(n11237), .B2(P1_EAX_REG_20__SCAN_IN), .A(n10854), .ZN(
        n10855) );
  OAI21_X1 U13767 ( .B1(n11239), .B2(n10856), .A(n10855), .ZN(n10858) );
  XNOR2_X1 U13768 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n10873), .ZN(
        n15467) );
  NAND2_X1 U13769 ( .A1(n15467), .A2(n12280), .ZN(n10857) );
  AOI22_X1 U13770 ( .A1(n10551), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10862) );
  AOI22_X1 U13771 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10861) );
  AOI22_X1 U13772 ( .A1(n11044), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10860) );
  AOI22_X1 U13773 ( .A1(n10544), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11039), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10859) );
  NAND4_X1 U13774 ( .A1(n10862), .A2(n10861), .A3(n10860), .A4(n10859), .ZN(
        n10868) );
  AOI22_X1 U13775 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11218), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10866) );
  AOI22_X1 U13776 ( .A1(n11038), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11219), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10865) );
  AOI22_X1 U13777 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10575), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10864) );
  AOI22_X1 U13778 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10863) );
  NAND4_X1 U13779 ( .A1(n10866), .A2(n10865), .A3(n10864), .A4(n10863), .ZN(
        n10867) );
  NOR2_X1 U13780 ( .A1(n10868), .A2(n10867), .ZN(n10872) );
  NAND2_X1 U13781 ( .A1(n20448), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10869) );
  NAND2_X1 U13782 ( .A1(n11028), .A2(n10869), .ZN(n10870) );
  AOI21_X1 U13783 ( .B1(n11237), .B2(P1_EAX_REG_21__SCAN_IN), .A(n10870), .ZN(
        n10871) );
  OAI21_X1 U13784 ( .B1(n11239), .B2(n10872), .A(n10871), .ZN(n10877) );
  OAI21_X1 U13785 ( .B1(n10875), .B2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n10917), .ZN(n15466) );
  OR2_X1 U13786 ( .A1(n15466), .A2(n11028), .ZN(n10876) );
  AOI22_X1 U13787 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11218), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10881) );
  AOI22_X1 U13788 ( .A1(n11038), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10880) );
  AOI22_X1 U13789 ( .A1(n11044), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10879) );
  AOI22_X1 U13790 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10575), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10878) );
  NAND4_X1 U13791 ( .A1(n10881), .A2(n10880), .A3(n10879), .A4(n10878), .ZN(
        n10887) );
  AOI22_X1 U13792 ( .A1(n10551), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11226), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10885) );
  AOI22_X1 U13793 ( .A1(n10544), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10884) );
  AOI22_X1 U13794 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10883) );
  AOI22_X1 U13795 ( .A1(n11219), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9610), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10882) );
  NAND4_X1 U13796 ( .A1(n10885), .A2(n10884), .A3(n10883), .A4(n10882), .ZN(
        n10886) );
  NOR2_X1 U13797 ( .A1(n10887), .A2(n10886), .ZN(n10890) );
  AOI21_X1 U13798 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14158), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10888) );
  AOI21_X1 U13799 ( .B1(n11237), .B2(P1_EAX_REG_22__SCAN_IN), .A(n10888), .ZN(
        n10889) );
  OAI21_X1 U13800 ( .B1(n11239), .B2(n10890), .A(n10889), .ZN(n10892) );
  XNOR2_X1 U13801 ( .A(n10917), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15451) );
  NAND2_X1 U13802 ( .A1(n15451), .A2(n12280), .ZN(n10891) );
  NAND2_X1 U13803 ( .A1(n10892), .A2(n10891), .ZN(n13997) );
  AOI22_X1 U13804 ( .A1(n11013), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11218), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10896) );
  AOI22_X1 U13805 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10895) );
  AOI22_X1 U13806 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11219), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10894) );
  AOI22_X1 U13807 ( .A1(n10448), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9610), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10893) );
  NAND4_X1 U13808 ( .A1(n10896), .A2(n10895), .A3(n10894), .A4(n10893), .ZN(
        n10902) );
  AOI22_X1 U13809 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10900) );
  AOI22_X1 U13810 ( .A1(n10454), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10453), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10899) );
  AOI22_X1 U13811 ( .A1(n11014), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10898) );
  AOI22_X1 U13812 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10897) );
  NAND4_X1 U13813 ( .A1(n10900), .A2(n10899), .A3(n10898), .A4(n10897), .ZN(
        n10901) );
  OR2_X1 U13814 ( .A1(n10902), .A2(n10901), .ZN(n10923) );
  AOI22_X1 U13815 ( .A1(n10903), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11218), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10907) );
  AOI22_X1 U13816 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10906) );
  AOI22_X1 U13817 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11219), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10905) );
  AOI22_X1 U13818 ( .A1(n10448), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9610), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10904) );
  NAND4_X1 U13819 ( .A1(n10907), .A2(n10906), .A3(n10905), .A4(n10904), .ZN(
        n10913) );
  AOI22_X1 U13820 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10911) );
  AOI22_X1 U13821 ( .A1(n10551), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10453), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10910) );
  AOI22_X1 U13822 ( .A1(n10463), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10909) );
  AOI22_X1 U13823 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10908) );
  NAND4_X1 U13824 ( .A1(n10911), .A2(n10910), .A3(n10909), .A4(n10908), .ZN(
        n10912) );
  OR2_X1 U13825 ( .A1(n10913), .A2(n10912), .ZN(n10924) );
  XNOR2_X1 U13826 ( .A(n10923), .B(n10924), .ZN(n10916) );
  INV_X1 U13827 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n13947) );
  AOI21_X1 U13828 ( .B1(n13947), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10914) );
  AOI21_X1 U13829 ( .B1(n11237), .B2(P1_EAX_REG_23__SCAN_IN), .A(n10914), .ZN(
        n10915) );
  OAI21_X1 U13830 ( .B1(n11239), .B2(n10916), .A(n10915), .ZN(n10922) );
  INV_X1 U13831 ( .A(n10918), .ZN(n10919) );
  NAND2_X1 U13832 ( .A1(n10919), .A2(n13947), .ZN(n10920) );
  NAND2_X1 U13833 ( .A1(n10956), .A2(n10920), .ZN(n14149) );
  NAND2_X1 U13834 ( .A1(n10924), .A2(n10923), .ZN(n10940) );
  AOI22_X1 U13835 ( .A1(n10544), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10928) );
  AOI22_X1 U13836 ( .A1(n11013), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10927) );
  AOI22_X1 U13837 ( .A1(n11014), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10926) );
  AOI22_X1 U13838 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9610), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10925) );
  NAND4_X1 U13839 ( .A1(n10928), .A2(n10927), .A3(n10926), .A4(n10925), .ZN(
        n10934) );
  AOI22_X1 U13840 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10932) );
  AOI22_X1 U13841 ( .A1(n11218), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11219), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10931) );
  AOI22_X1 U13842 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10453), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10930) );
  AOI22_X1 U13843 ( .A1(n10454), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10929) );
  NAND4_X1 U13844 ( .A1(n10932), .A2(n10931), .A3(n10930), .A4(n10929), .ZN(
        n10933) );
  NOR2_X1 U13845 ( .A1(n10934), .A2(n10933), .ZN(n10941) );
  XOR2_X1 U13846 ( .A(n10940), .B(n10941), .Z(n10935) );
  NAND2_X1 U13847 ( .A1(n10935), .A2(n11051), .ZN(n10939) );
  INV_X1 U13848 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15439) );
  AOI21_X1 U13849 ( .B1(n15439), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10936) );
  AOI21_X1 U13850 ( .B1(n11237), .B2(P1_EAX_REG_24__SCAN_IN), .A(n10936), .ZN(
        n10938) );
  XNOR2_X1 U13851 ( .A(n10956), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15444) );
  AOI21_X1 U13852 ( .B1(n10939), .B2(n10938), .A(n10937), .ZN(n13985) );
  NOR2_X1 U13853 ( .A1(n10941), .A2(n10940), .ZN(n10966) );
  AOI22_X1 U13854 ( .A1(n11013), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11218), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10945) );
  AOI22_X1 U13855 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10944) );
  AOI22_X1 U13856 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10570), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10943) );
  AOI22_X1 U13857 ( .A1(n10448), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9610), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10942) );
  NAND4_X1 U13858 ( .A1(n10945), .A2(n10944), .A3(n10943), .A4(n10942), .ZN(
        n10951) );
  AOI22_X1 U13859 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10949) );
  AOI22_X1 U13860 ( .A1(n10454), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10575), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10948) );
  AOI22_X1 U13861 ( .A1(n11014), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10947) );
  AOI22_X1 U13862 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10946) );
  NAND4_X1 U13863 ( .A1(n10949), .A2(n10948), .A3(n10947), .A4(n10946), .ZN(
        n10950) );
  OR2_X1 U13864 ( .A1(n10951), .A2(n10950), .ZN(n10965) );
  INV_X1 U13865 ( .A(n10965), .ZN(n10952) );
  XNOR2_X1 U13866 ( .A(n10966), .B(n10952), .ZN(n10953) );
  NAND2_X1 U13867 ( .A1(n10953), .A2(n11051), .ZN(n10964) );
  NAND2_X1 U13868 ( .A1(n20448), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10954) );
  NAND2_X1 U13869 ( .A1(n11028), .A2(n10954), .ZN(n10955) );
  AOI21_X1 U13870 ( .B1(n11237), .B2(P1_EAX_REG_25__SCAN_IN), .A(n10955), .ZN(
        n10963) );
  INV_X1 U13871 ( .A(n10956), .ZN(n10957) );
  INV_X1 U13872 ( .A(n10958), .ZN(n10960) );
  INV_X1 U13873 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n10959) );
  NAND2_X1 U13874 ( .A1(n10960), .A2(n10959), .ZN(n10961) );
  NAND2_X1 U13875 ( .A1(n11002), .A2(n10961), .ZN(n15432) );
  NOR2_X1 U13876 ( .A1(n15432), .A2(n11028), .ZN(n10962) );
  AOI21_X1 U13877 ( .B1(n10964), .B2(n10963), .A(n10962), .ZN(n13979) );
  NAND2_X1 U13878 ( .A1(n10966), .A2(n10965), .ZN(n10985) );
  AOI22_X1 U13879 ( .A1(n11013), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11037), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10970) );
  AOI22_X1 U13880 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10969) );
  AOI22_X1 U13881 ( .A1(n11014), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10968) );
  AOI22_X1 U13882 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10967) );
  NAND4_X1 U13883 ( .A1(n10970), .A2(n10969), .A3(n10968), .A4(n10967), .ZN(
        n10977) );
  AOI22_X1 U13884 ( .A1(n11218), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10975) );
  AOI22_X1 U13885 ( .A1(n10551), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10575), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10974) );
  AOI22_X1 U13886 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10570), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10973) );
  AOI22_X1 U13887 ( .A1(n10448), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11039), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10972) );
  NAND4_X1 U13888 ( .A1(n10975), .A2(n10974), .A3(n10973), .A4(n10972), .ZN(
        n10976) );
  NOR2_X1 U13889 ( .A1(n10977), .A2(n10976), .ZN(n10986) );
  XOR2_X1 U13890 ( .A(n10985), .B(n10986), .Z(n10978) );
  NAND2_X1 U13891 ( .A1(n10978), .A2(n11051), .ZN(n10982) );
  NAND2_X1 U13892 ( .A1(n20448), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10979) );
  NAND2_X1 U13893 ( .A1(n11028), .A2(n10979), .ZN(n10980) );
  AOI21_X1 U13894 ( .B1(n11237), .B2(P1_EAX_REG_26__SCAN_IN), .A(n10980), .ZN(
        n10981) );
  NAND2_X1 U13895 ( .A1(n10982), .A2(n10981), .ZN(n10984) );
  XNOR2_X1 U13896 ( .A(n11002), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14123) );
  NAND2_X1 U13897 ( .A1(n14123), .A2(n12280), .ZN(n10983) );
  NAND2_X1 U13898 ( .A1(n10984), .A2(n10983), .ZN(n13931) );
  NOR2_X1 U13899 ( .A1(n10986), .A2(n10985), .ZN(n11012) );
  AOI22_X1 U13900 ( .A1(n11013), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11218), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10990) );
  AOI22_X1 U13901 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10989) );
  AOI22_X1 U13902 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11038), .B1(
        n10570), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10988) );
  AOI22_X1 U13903 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n10544), .B1(
        n9610), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10987) );
  NAND4_X1 U13904 ( .A1(n10990), .A2(n10989), .A3(n10988), .A4(n10987), .ZN(
        n10996) );
  AOI22_X1 U13905 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10994) );
  AOI22_X1 U13906 ( .A1(n10454), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10575), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10993) );
  AOI22_X1 U13907 ( .A1(n11014), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10992) );
  AOI22_X1 U13908 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10991) );
  NAND4_X1 U13909 ( .A1(n10994), .A2(n10993), .A3(n10992), .A4(n10991), .ZN(
        n10995) );
  OR2_X1 U13910 ( .A1(n10996), .A2(n10995), .ZN(n11011) );
  INV_X1 U13911 ( .A(n11011), .ZN(n10997) );
  XNOR2_X1 U13912 ( .A(n11012), .B(n10997), .ZN(n11001) );
  INV_X1 U13913 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n14032) );
  NAND2_X1 U13914 ( .A1(n20448), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10998) );
  OAI211_X1 U13915 ( .C1(n10999), .C2(n14032), .A(n11028), .B(n10998), .ZN(
        n11000) );
  AOI21_X1 U13916 ( .B1(n11001), .B2(n11051), .A(n11000), .ZN(n11009) );
  INV_X1 U13917 ( .A(n11002), .ZN(n11003) );
  INV_X1 U13918 ( .A(n11004), .ZN(n11006) );
  INV_X1 U13919 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11005) );
  NAND2_X1 U13920 ( .A1(n11006), .A2(n11005), .ZN(n11007) );
  NAND2_X1 U13921 ( .A1(n11055), .A2(n11007), .ZN(n14116) );
  NOR2_X1 U13922 ( .A1(n14116), .A2(n11028), .ZN(n11008) );
  NAND2_X1 U13923 ( .A1(n11012), .A2(n11011), .ZN(n11034) );
  AOI22_X1 U13924 ( .A1(n11013), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11018) );
  AOI22_X1 U13925 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11017) );
  AOI22_X1 U13926 ( .A1(n11014), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11016) );
  AOI22_X1 U13927 ( .A1(n11218), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11015) );
  NAND4_X1 U13928 ( .A1(n11018), .A2(n11017), .A3(n11016), .A4(n11015), .ZN(
        n11025) );
  AOI22_X1 U13929 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11023) );
  AOI22_X1 U13930 ( .A1(n10454), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10453), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11022) );
  AOI22_X1 U13931 ( .A1(n10448), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10570), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11021) );
  AOI22_X1 U13932 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11039), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11020) );
  NAND4_X1 U13933 ( .A1(n11023), .A2(n11022), .A3(n11021), .A4(n11020), .ZN(
        n11024) );
  NOR2_X1 U13934 ( .A1(n11025), .A2(n11024), .ZN(n11035) );
  XOR2_X1 U13935 ( .A(n11034), .B(n11035), .Z(n11026) );
  NAND2_X1 U13936 ( .A1(n11026), .A2(n11051), .ZN(n11031) );
  NAND2_X1 U13937 ( .A1(n20448), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11027) );
  NAND2_X1 U13938 ( .A1(n11028), .A2(n11027), .ZN(n11029) );
  AOI21_X1 U13939 ( .B1(n11237), .B2(P1_EAX_REG_28__SCAN_IN), .A(n11029), .ZN(
        n11030) );
  NAND2_X1 U13940 ( .A1(n11031), .A2(n11030), .ZN(n11033) );
  XNOR2_X1 U13941 ( .A(n11055), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14105) );
  NAND2_X1 U13942 ( .A1(n14105), .A2(n12280), .ZN(n11032) );
  NAND2_X1 U13943 ( .A1(n11033), .A2(n11032), .ZN(n13917) );
  NOR2_X1 U13944 ( .A1(n11035), .A2(n11034), .ZN(n11053) );
  AOI22_X1 U13945 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11218), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11043) );
  AOI22_X1 U13946 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11042) );
  AOI22_X1 U13947 ( .A1(n11038), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11219), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11041) );
  AOI22_X1 U13948 ( .A1(n10448), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9610), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11040) );
  NAND4_X1 U13949 ( .A1(n11043), .A2(n11042), .A3(n11041), .A4(n11040), .ZN(
        n11050) );
  AOI22_X1 U13950 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11048) );
  AOI22_X1 U13951 ( .A1(n10551), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10575), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11047) );
  AOI22_X1 U13952 ( .A1(n11044), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11046) );
  AOI22_X1 U13953 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11045) );
  NAND4_X1 U13954 ( .A1(n11048), .A2(n11047), .A3(n11046), .A4(n11045), .ZN(
        n11049) );
  OR2_X1 U13955 ( .A1(n11050), .A2(n11049), .ZN(n11052) );
  NAND2_X1 U13956 ( .A1(n11053), .A2(n11052), .ZN(n11234) );
  OAI211_X1 U13957 ( .C1(n11053), .C2(n11052), .A(n11234), .B(n11051), .ZN(
        n11059) );
  INV_X1 U13958 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11215) );
  NOR2_X1 U13959 ( .A1(n11215), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11054) );
  AOI211_X1 U13960 ( .C1(n11237), .C2(P1_EAX_REG_29__SCAN_IN), .A(n12280), .B(
        n11054), .ZN(n11058) );
  INV_X1 U13961 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14107) );
  NAND2_X1 U13962 ( .A1(n11056), .A2(n11215), .ZN(n11057) );
  AOI22_X1 U13963 ( .A1(n11059), .A2(n11058), .B1(n12280), .B2(n13731), .ZN(
        n11060) );
  OR2_X1 U13964 ( .A1(n13915), .A2(n11060), .ZN(n11061) );
  NOR2_X2 U13965 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20316) );
  AND2_X1 U13966 ( .A1(n20316), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12939) );
  NAND2_X1 U13967 ( .A1(n11062), .A2(n19853), .ZN(n11067) );
  XNOR2_X1 U13968 ( .A(n11073), .B(n11074), .ZN(n11064) );
  OAI211_X1 U13969 ( .C1(n11064), .C2(n20541), .A(n11063), .B(n19873), .ZN(
        n11065) );
  INV_X1 U13970 ( .A(n11065), .ZN(n11066) );
  NAND2_X1 U13971 ( .A1(n11067), .A2(n11066), .ZN(n11070) );
  NAND2_X1 U13972 ( .A1(n19873), .A2(n19853), .ZN(n11160) );
  NAND2_X1 U13973 ( .A1(n12485), .A2(n19863), .ZN(n11075) );
  OAI21_X1 U13974 ( .B1(n20541), .B2(n11074), .A(n11075), .ZN(n11068) );
  INV_X1 U13975 ( .A(n11068), .ZN(n11069) );
  INV_X1 U13976 ( .A(n11070), .ZN(n11071) );
  OR2_X1 U13977 ( .A1(n12680), .A2(n11071), .ZN(n11072) );
  INV_X1 U13978 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19831) );
  INV_X1 U13979 ( .A(n11160), .ZN(n11123) );
  NAND2_X1 U13980 ( .A1(n11074), .A2(n11073), .ZN(n11083) );
  XNOR2_X1 U13981 ( .A(n11083), .B(n11082), .ZN(n11077) );
  INV_X1 U13982 ( .A(n11075), .ZN(n11076) );
  AOI21_X1 U13983 ( .B1(n11077), .B2(n11129), .A(n11076), .ZN(n11078) );
  NAND2_X1 U13984 ( .A1(n11079), .A2(n11078), .ZN(n12874) );
  NAND2_X1 U13985 ( .A1(n11080), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11081) );
  INV_X1 U13986 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n19814) );
  XNOR2_X1 U13987 ( .A(n11088), .B(n19814), .ZN(n12997) );
  NAND2_X1 U13988 ( .A1(n20524), .A2(n11123), .ZN(n11087) );
  NAND2_X1 U13989 ( .A1(n11083), .A2(n11082), .ZN(n11101) );
  XNOR2_X1 U13990 ( .A(n11101), .B(n11084), .ZN(n11085) );
  NAND2_X1 U13991 ( .A1(n11085), .A2(n11129), .ZN(n11086) );
  NAND2_X1 U13992 ( .A1(n11087), .A2(n11086), .ZN(n12996) );
  NAND2_X1 U13993 ( .A1(n11088), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11089) );
  NAND2_X1 U13994 ( .A1(n11090), .A2(n11123), .ZN(n11094) );
  NAND2_X1 U13995 ( .A1(n11101), .A2(n11099), .ZN(n11091) );
  XNOR2_X1 U13996 ( .A(n11091), .B(n11098), .ZN(n11092) );
  NAND2_X1 U13997 ( .A1(n11092), .A2(n11129), .ZN(n11093) );
  NAND2_X1 U13998 ( .A1(n11094), .A2(n11093), .ZN(n11095) );
  INV_X1 U13999 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19804) );
  XNOR2_X1 U14000 ( .A(n11095), .B(n19804), .ZN(n19784) );
  NAND2_X1 U14001 ( .A1(n11095), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11096) );
  NAND2_X1 U14002 ( .A1(n11097), .A2(n11123), .ZN(n11104) );
  AND2_X1 U14003 ( .A1(n11099), .A2(n11098), .ZN(n11100) );
  NAND2_X1 U14004 ( .A1(n11101), .A2(n11100), .ZN(n11118) );
  XNOR2_X1 U14005 ( .A(n11118), .B(n11116), .ZN(n11102) );
  NAND2_X1 U14006 ( .A1(n11102), .A2(n11129), .ZN(n11103) );
  NAND2_X1 U14007 ( .A1(n11104), .A2(n11103), .ZN(n11105) );
  INV_X1 U14008 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15679) );
  XNOR2_X1 U14009 ( .A(n11105), .B(n15679), .ZN(n15592) );
  NAND2_X1 U14010 ( .A1(n11105), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11106) );
  NAND2_X1 U14011 ( .A1(n11107), .A2(n11123), .ZN(n11112) );
  INV_X1 U14012 ( .A(n11118), .ZN(n11108) );
  NAND2_X1 U14013 ( .A1(n11108), .A2(n11116), .ZN(n11109) );
  XNOR2_X1 U14014 ( .A(n11109), .B(n11115), .ZN(n11110) );
  NAND2_X1 U14015 ( .A1(n11110), .A2(n11129), .ZN(n11111) );
  NAND2_X1 U14016 ( .A1(n11112), .A2(n11111), .ZN(n15586) );
  OR2_X1 U14017 ( .A1(n15586), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11113) );
  NAND2_X1 U14018 ( .A1(n11114), .A2(n11123), .ZN(n11121) );
  NAND2_X1 U14019 ( .A1(n11116), .A2(n11115), .ZN(n11117) );
  OR2_X1 U14020 ( .A1(n11118), .A2(n11117), .ZN(n11127) );
  XNOR2_X1 U14021 ( .A(n11127), .B(n11128), .ZN(n11119) );
  NAND2_X1 U14022 ( .A1(n11119), .A2(n11129), .ZN(n11120) );
  NAND2_X1 U14023 ( .A1(n11121), .A2(n11120), .ZN(n11122) );
  OR2_X1 U14024 ( .A1(n11122), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15581) );
  NAND2_X1 U14025 ( .A1(n11122), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15580) );
  AND2_X1 U14026 ( .A1(n11124), .A2(n11123), .ZN(n11125) );
  INV_X1 U14027 ( .A(n11127), .ZN(n11130) );
  NAND3_X1 U14028 ( .A1(n11130), .A2(n11129), .A3(n11128), .ZN(n11131) );
  NAND2_X1 U14029 ( .A1(n15572), .A2(n11131), .ZN(n13213) );
  OR2_X1 U14030 ( .A1(n13213), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11132) );
  NAND2_X1 U14031 ( .A1(n13213), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11133) );
  INV_X1 U14032 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11134) );
  INV_X1 U14033 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12330) );
  AND2_X1 U14034 ( .A1(n15572), .A2(n12330), .ZN(n14185) );
  INV_X1 U14035 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15618) );
  NAND2_X1 U14036 ( .A1(n15572), .A2(n15618), .ZN(n11135) );
  NAND2_X1 U14037 ( .A1(n14194), .A2(n11135), .ZN(n14207) );
  INV_X1 U14038 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11136) );
  NAND2_X1 U14039 ( .A1(n15572), .A2(n11136), .ZN(n14204) );
  NAND2_X1 U14040 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11137) );
  NAND2_X1 U14041 ( .A1(n15572), .A2(n11137), .ZN(n13549) );
  NAND2_X1 U14042 ( .A1(n14194), .A2(n11138), .ZN(n14394) );
  INV_X1 U14043 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14380) );
  NOR2_X1 U14044 ( .A1(n15572), .A2(n14380), .ZN(n14393) );
  NOR2_X1 U14045 ( .A1(n14394), .A2(n14393), .ZN(n11141) );
  XNOR2_X1 U14046 ( .A(n15572), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14187) );
  NAND2_X1 U14047 ( .A1(n15572), .A2(n14380), .ZN(n14391) );
  AND2_X1 U14048 ( .A1(n14187), .A2(n14391), .ZN(n11139) );
  INV_X1 U14049 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11140) );
  INV_X1 U14050 ( .A(n11141), .ZN(n14186) );
  NAND2_X1 U14051 ( .A1(n9603), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13550) );
  INV_X1 U14052 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15624) );
  INV_X1 U14053 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15629) );
  NAND2_X1 U14054 ( .A1(n15624), .A2(n15629), .ZN(n11142) );
  NAND2_X1 U14055 ( .A1(n9603), .A2(n11142), .ZN(n13547) );
  NAND2_X1 U14056 ( .A1(n13550), .A2(n13547), .ZN(n14184) );
  INV_X1 U14057 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11143) );
  XNOR2_X1 U14058 ( .A(n15572), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14176) );
  NAND2_X1 U14059 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14329) );
  INV_X1 U14060 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14311) );
  INV_X1 U14061 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n20642) );
  INV_X1 U14062 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14295) );
  NAND3_X1 U14063 ( .A1(n14311), .A2(n20642), .A3(n14295), .ZN(n14099) );
  NAND2_X1 U14064 ( .A1(n11145), .A2(n15572), .ZN(n14129) );
  AND2_X1 U14065 ( .A1(n14129), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11147) );
  AND2_X1 U14066 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14242) );
  NAND2_X1 U14067 ( .A1(n14242), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14231) );
  NAND2_X1 U14068 ( .A1(n14146), .A2(n14231), .ZN(n11146) );
  AND2_X1 U14069 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14245) );
  NOR2_X1 U14070 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11149) );
  MUX2_X1 U14071 ( .A(n14082), .B(n14080), .S(n9603), .Z(n11150) );
  INV_X1 U14072 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14247) );
  MUX2_X1 U14073 ( .A(n19923), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n11166) );
  NAND2_X1 U14074 ( .A1(n20315), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11159) );
  NAND2_X1 U14075 ( .A1(n11166), .A2(n11167), .ZN(n11152) );
  NAND2_X1 U14076 ( .A1(n19923), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11151) );
  NAND2_X1 U14077 ( .A1(n11152), .A2(n11151), .ZN(n11178) );
  XNOR2_X1 U14078 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11177) );
  NAND2_X1 U14079 ( .A1(n11178), .A2(n11177), .ZN(n11154) );
  NAND2_X1 U14080 ( .A1(n20262), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11153) );
  NOR2_X1 U14081 ( .A1(n12926), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11155) );
  INV_X1 U14082 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19833) );
  NAND2_X1 U14083 ( .A1(n19833), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11156) );
  NAND2_X1 U14084 ( .A1(n11191), .A2(n11156), .ZN(n11158) );
  NAND2_X1 U14085 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12637), .ZN(
        n11157) );
  OAI21_X1 U14086 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20315), .A(
        n11159), .ZN(n11162) );
  NOR2_X1 U14087 ( .A1(n11201), .A2(n11162), .ZN(n11165) );
  OAI21_X1 U14088 ( .B1(n11210), .B2(n11162), .A(n11161), .ZN(n11163) );
  INV_X1 U14089 ( .A(n11163), .ZN(n11164) );
  AOI21_X1 U14090 ( .B1(n9865), .B2(n19839), .A(n19853), .ZN(n11180) );
  OAI22_X1 U14091 ( .A1(n11165), .A2(n11203), .B1(n11164), .B2(n11180), .ZN(
        n11172) );
  INV_X1 U14092 ( .A(n11172), .ZN(n11176) );
  XNOR2_X1 U14093 ( .A(n11167), .B(n11166), .ZN(n11249) );
  NOR2_X1 U14094 ( .A1(n19873), .A2(n20446), .ZN(n11169) );
  NOR2_X1 U14095 ( .A1(n11201), .A2(n12597), .ZN(n11168) );
  AOI211_X1 U14096 ( .C1(n11194), .C2(n11249), .A(n11169), .B(n11168), .ZN(
        n11173) );
  INV_X1 U14097 ( .A(n11173), .ZN(n11175) );
  INV_X1 U14098 ( .A(n11169), .ZN(n11170) );
  AND2_X1 U14099 ( .A1(n11170), .A2(n19853), .ZN(n11171) );
  NAND2_X1 U14100 ( .A1(n11201), .A2(n11171), .ZN(n11193) );
  AOI22_X1 U14101 ( .A1(n11173), .A2(n11172), .B1(n11249), .B2(n11193), .ZN(
        n11174) );
  AOI21_X1 U14102 ( .B1(n11176), .B2(n11175), .A(n11174), .ZN(n11184) );
  XNOR2_X1 U14103 ( .A(n11178), .B(n11177), .ZN(n11250) );
  AOI211_X1 U14104 ( .C1(n11194), .C2(n11250), .A(n11180), .B(n11179), .ZN(
        n11183) );
  INV_X1 U14105 ( .A(n11179), .ZN(n11182) );
  INV_X1 U14106 ( .A(n11180), .ZN(n11181) );
  OAI22_X1 U14107 ( .A1(n11184), .A2(n11183), .B1(n11182), .B2(n11181), .ZN(
        n11189) );
  XNOR2_X1 U14108 ( .A(n11186), .B(n11185), .ZN(n11248) );
  NAND2_X1 U14109 ( .A1(n11187), .A2(n11248), .ZN(n11188) );
  AOI22_X1 U14110 ( .A1(n11189), .A2(n11188), .B1(n11203), .B2(n11248), .ZN(
        n11198) );
  NOR2_X1 U14111 ( .A1(n19833), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11190) );
  INV_X1 U14112 ( .A(n11251), .ZN(n11192) );
  INV_X1 U14113 ( .A(n11193), .ZN(n11195) );
  NAND3_X1 U14114 ( .A1(n11195), .A2(n11194), .A3(n11251), .ZN(n11196) );
  INV_X1 U14115 ( .A(n11253), .ZN(n11202) );
  NAND2_X1 U14116 ( .A1(n11203), .A2(n11202), .ZN(n11204) );
  INV_X1 U14117 ( .A(n12899), .ZN(n12486) );
  NAND2_X1 U14118 ( .A1(n12486), .A2(n12701), .ZN(n11208) );
  AND2_X1 U14119 ( .A1(n11208), .A2(n11207), .ZN(n12502) );
  NAND2_X1 U14120 ( .A1(n14422), .A2(n12485), .ZN(n11209) );
  AND2_X1 U14121 ( .A1(n12484), .A2(n11210), .ZN(n15381) );
  NAND2_X1 U14122 ( .A1(n20516), .A2(n11214), .ZN(n20548) );
  AND2_X1 U14123 ( .A1(n20548), .A2(n20446), .ZN(n11211) );
  NAND2_X1 U14124 ( .A1(n20446), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15394) );
  INV_X1 U14125 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20347) );
  NAND2_X1 U14126 ( .A1(n20347), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n11212) );
  AND2_X1 U14127 ( .A1(n15394), .A2(n11212), .ZN(n12677) );
  INV_X1 U14128 ( .A(n12677), .ZN(n11213) );
  NAND2_X1 U14129 ( .A1(n19781), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14261) );
  OAI21_X1 U14130 ( .B1(n14190), .B2(n11215), .A(n14261), .ZN(n11216) );
  AOI22_X1 U14131 ( .A1(n10461), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11218), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11223) );
  AOI22_X1 U14132 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11222) );
  AOI22_X1 U14133 ( .A1(n11038), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11219), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11221) );
  AOI22_X1 U14134 ( .A1(n10544), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11039), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11220) );
  NAND4_X1 U14135 ( .A1(n11223), .A2(n11222), .A3(n11221), .A4(n11220), .ZN(
        n11232) );
  AOI22_X1 U14136 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11230) );
  AOI22_X1 U14137 ( .A1(n10551), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10575), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11229) );
  AOI22_X1 U14138 ( .A1(n10463), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11228) );
  AOI22_X1 U14139 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12914), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11227) );
  NAND4_X1 U14140 ( .A1(n11230), .A2(n11229), .A3(n11228), .A4(n11227), .ZN(
        n11231) );
  NOR2_X1 U14141 ( .A1(n11232), .A2(n11231), .ZN(n11233) );
  XNOR2_X1 U14142 ( .A(n11234), .B(n11233), .ZN(n11240) );
  NAND2_X1 U14143 ( .A1(n20448), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11235) );
  NAND2_X1 U14144 ( .A1(n11028), .A2(n11235), .ZN(n11236) );
  AOI21_X1 U14145 ( .B1(n11237), .B2(P1_EAX_REG_30__SCAN_IN), .A(n11236), .ZN(
        n11238) );
  OAI21_X1 U14146 ( .B1(n11240), .B2(n11239), .A(n11238), .ZN(n11242) );
  XNOR2_X1 U14147 ( .A(n12284), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14093) );
  NAND2_X1 U14148 ( .A1(n14093), .A2(n12280), .ZN(n11241) );
  NAND2_X1 U14149 ( .A1(n11242), .A2(n11241), .ZN(n13906) );
  AOI22_X1 U14150 ( .A1(n10508), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n11243), .ZN(n11244) );
  XNOR2_X1 U14151 ( .A(n11245), .B(n11244), .ZN(n14089) );
  NAND2_X1 U14152 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20546) );
  INV_X1 U14153 ( .A(n20546), .ZN(n20457) );
  AND2_X1 U14154 ( .A1(n12484), .A2(n13056), .ZN(n12515) );
  OR4_X1 U14155 ( .A1(n11251), .A2(n11250), .A3(n11249), .A4(n11248), .ZN(
        n11252) );
  NAND2_X1 U14156 ( .A1(n11253), .A2(n11252), .ZN(n12424) );
  OR2_X1 U14157 ( .A1(n12424), .A2(n20457), .ZN(n12695) );
  OR2_X1 U14158 ( .A1(n11247), .A2(n12695), .ZN(n12491) );
  INV_X1 U14159 ( .A(n13056), .ZN(n12508) );
  NOR2_X1 U14160 ( .A1(n19886), .A2(n19602), .ZN(n11254) );
  NAND4_X1 U14161 ( .A1(n12520), .A2(n11255), .A3(n11254), .A4(n19878), .ZN(
        n12651) );
  OAI22_X1 U14162 ( .A1(n12491), .A2(n19602), .B1(n12508), .B2(n12651), .ZN(
        n11256) );
  AOI21_X1 U14163 ( .B1(n12688), .B2(n12515), .A(n11256), .ZN(n11257) );
  INV_X1 U14164 ( .A(n19886), .ZN(n13724) );
  NAND3_X1 U14165 ( .A1(n14089), .A2(n19713), .A3(n13724), .ZN(n11274) );
  NOR4_X1 U14166 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n11261) );
  NOR4_X1 U14167 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n11260) );
  NOR4_X1 U14168 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n11259) );
  NOR4_X1 U14169 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n11258) );
  AND4_X1 U14170 ( .A1(n11261), .A2(n11260), .A3(n11259), .A4(n11258), .ZN(
        n11266) );
  NOR4_X1 U14171 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n11264) );
  NOR4_X1 U14172 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n11263) );
  NOR4_X1 U14173 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n11262) );
  INV_X1 U14174 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20469) );
  AND4_X1 U14175 ( .A1(n11264), .A2(n11263), .A3(n11262), .A4(n20469), .ZN(
        n11265) );
  NAND2_X1 U14176 ( .A1(n11266), .A2(n11265), .ZN(n11267) );
  NOR3_X1 U14177 ( .A1(n15545), .A2(n19836), .A3(n12684), .ZN(n11268) );
  AOI22_X1 U14178 ( .A1(n14071), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15545), .ZN(n11269) );
  INV_X1 U14179 ( .A(n11269), .ZN(n11272) );
  INV_X1 U14180 ( .A(n19836), .ZN(n19834) );
  NOR2_X1 U14181 ( .A1(n12684), .A2(n19834), .ZN(n11270) );
  NAND2_X1 U14182 ( .A1(n19713), .A2(n11270), .ZN(n14063) );
  INV_X1 U14183 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n15992) );
  NOR2_X1 U14184 ( .A1(n14063), .A2(n15992), .ZN(n11271) );
  NOR2_X1 U14185 ( .A1(n11272), .A2(n11271), .ZN(n11273) );
  NAND2_X1 U14186 ( .A1(n11274), .A2(n11273), .ZN(P1_U2873) );
  AOI22_X1 U14187 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9606), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11279) );
  INV_X2 U14188 ( .A(n11291), .ZN(n11816) );
  AOI22_X1 U14189 ( .A1(n11816), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11804), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11278) );
  AOI22_X1 U14190 ( .A1(n11777), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11654), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11277) );
  AOI22_X1 U14191 ( .A1(n11348), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9627), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11276) );
  NAND4_X1 U14192 ( .A1(n11279), .A2(n11278), .A3(n11277), .A4(n11276), .ZN(
        n11285) );
  AOI22_X1 U14193 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9605), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11283) );
  AOI22_X1 U14194 ( .A1(n11816), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11804), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11282) );
  AOI22_X1 U14195 ( .A1(n11777), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11654), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11281) );
  AOI22_X1 U14196 ( .A1(n11348), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11815), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11280) );
  NAND4_X1 U14197 ( .A1(n11283), .A2(n11282), .A3(n11281), .A4(n11280), .ZN(
        n11284) );
  AOI22_X1 U14198 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(n9607), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11290) );
  AOI22_X1 U14199 ( .A1(n11777), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11804), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11289) );
  AOI22_X1 U14200 ( .A1(n11816), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11654), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11288) );
  AOI22_X1 U14201 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n11815), .B1(
        n11348), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11287) );
  NAND4_X1 U14202 ( .A1(n11290), .A2(n11289), .A3(n11288), .A4(n11287), .ZN(
        n11297) );
  AOI22_X1 U14203 ( .A1(n9624), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9606), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11295) );
  AOI22_X1 U14204 ( .A1(n11816), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11804), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11294) );
  AOI22_X1 U14205 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11654), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11293) );
  AOI22_X1 U14206 ( .A1(n11348), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9627), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11292) );
  NAND4_X1 U14207 ( .A1(n11295), .A2(n11294), .A3(n11293), .A4(n11292), .ZN(
        n11296) );
  AOI22_X1 U14208 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9606), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11302) );
  AOI22_X1 U14209 ( .A1(n9638), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11804), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11301) );
  AOI22_X1 U14210 ( .A1(n11777), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11654), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11300) );
  AOI22_X1 U14211 ( .A1(n11348), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9627), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11299) );
  NAND4_X1 U14212 ( .A1(n11302), .A2(n11301), .A3(n11300), .A4(n11299), .ZN(
        n11308) );
  AOI22_X1 U14213 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9624), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11306) );
  AOI22_X1 U14214 ( .A1(n9638), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11804), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11305) );
  AOI22_X1 U14215 ( .A1(n9605), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11654), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11304) );
  AOI22_X1 U14216 ( .A1(n11348), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11815), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11303) );
  NAND4_X1 U14217 ( .A1(n11306), .A2(n11305), .A3(n11304), .A4(n11303), .ZN(
        n11307) );
  AND3_X2 U14218 ( .A1(n18907), .A2(n12581), .A3(n12630), .ZN(n11375) );
  AOI22_X1 U14219 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11312) );
  AOI22_X1 U14220 ( .A1(n9637), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11804), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11311) );
  AOI22_X1 U14221 ( .A1(n11777), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11654), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11310) );
  AOI22_X1 U14222 ( .A1(n11348), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9627), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11309) );
  AOI22_X1 U14223 ( .A1(n9625), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(n9607), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11317) );
  AOI22_X1 U14224 ( .A1(n9637), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11804), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11316) );
  AOI22_X1 U14225 ( .A1(n9624), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11654), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11315) );
  AOI22_X1 U14226 ( .A1(n11348), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11815), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11314) );
  AOI22_X1 U14227 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9605), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11323) );
  AOI22_X1 U14228 ( .A1(n9638), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11804), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11322) );
  AOI22_X1 U14229 ( .A1(n11777), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11654), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11321) );
  AOI22_X1 U14230 ( .A1(n11348), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9627), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11320) );
  AOI22_X1 U14231 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9606), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11326) );
  AOI22_X1 U14232 ( .A1(n9638), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11804), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11325) );
  AOI22_X1 U14233 ( .A1(n9624), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11654), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11324) );
  AOI22_X1 U14234 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(n9605), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11330) );
  AOI22_X1 U14235 ( .A1(n9638), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11804), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11329) );
  AOI22_X1 U14236 ( .A1(n11777), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11654), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11328) );
  AOI22_X1 U14237 ( .A1(n11348), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11815), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11327) );
  AOI22_X1 U14238 ( .A1(n9624), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11654), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11333) );
  AOI22_X1 U14239 ( .A1(n9638), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11804), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11332) );
  AOI22_X1 U14240 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9606), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11336) );
  AOI22_X1 U14241 ( .A1(n11348), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11815), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11334) );
  NAND3_X1 U14242 ( .A1(n10285), .A2(n11336), .A3(n11335), .ZN(n11337) );
  AOI22_X1 U14243 ( .A1(n9605), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11816), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11343) );
  AOI22_X1 U14244 ( .A1(n9623), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11804), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11342) );
  AOI22_X1 U14245 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11654), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11341) );
  AOI22_X1 U14246 ( .A1(n11348), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11815), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11340) );
  AOI22_X1 U14247 ( .A1(n11348), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11815), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11347) );
  AOI22_X1 U14248 ( .A1(n11816), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11804), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11346) );
  AOI22_X1 U14249 ( .A1(n11777), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11654), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11345) );
  AOI22_X1 U14250 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11344) );
  AOI22_X1 U14251 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9605), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11352) );
  AOI22_X1 U14252 ( .A1(n11816), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11804), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11351) );
  AOI22_X1 U14253 ( .A1(n11777), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11654), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11350) );
  AOI22_X1 U14254 ( .A1(n11348), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9627), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11349) );
  NAND4_X1 U14255 ( .A1(n11352), .A2(n11351), .A3(n11350), .A4(n11349), .ZN(
        n11358) );
  AOI22_X1 U14256 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11356) );
  AOI22_X1 U14257 ( .A1(n11816), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11804), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11355) );
  AOI22_X1 U14258 ( .A1(n11777), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11654), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11354) );
  AOI22_X1 U14259 ( .A1(n11348), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9627), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11353) );
  NAND4_X1 U14260 ( .A1(n11356), .A2(n11355), .A3(n11354), .A4(n11353), .ZN(
        n11357) );
  NAND4_X1 U14261 ( .A1(n18907), .A2(n9808), .A3(n12630), .A4(n12549), .ZN(
        n11359) );
  INV_X2 U14262 ( .A(n18919), .ZN(n12631) );
  NAND2_X2 U14263 ( .A1(n12631), .A2(n9614), .ZN(n11373) );
  AND3_X1 U14264 ( .A1(n9634), .A2(n12003), .A3(n12630), .ZN(n11361) );
  INV_X1 U14265 ( .A(n12065), .ZN(n12045) );
  NAND2_X1 U14266 ( .A1(n12540), .A2(n9634), .ZN(n11840) );
  NAND2_X2 U14267 ( .A1(n11832), .A2(n12005), .ZN(n11382) );
  NAND2_X1 U14268 ( .A1(n12065), .A2(n12541), .ZN(n12534) );
  NAND3_X1 U14269 ( .A1(n11373), .A2(n12536), .A3(n18907), .ZN(n12545) );
  NAND3_X1 U14270 ( .A1(n12534), .A2(n12545), .A3(n12630), .ZN(n12579) );
  NAND2_X1 U14271 ( .A1(n12579), .A2(n12581), .ZN(n11365) );
  NAND2_X1 U14272 ( .A1(n11365), .A2(n11364), .ZN(n11366) );
  NAND2_X1 U14273 ( .A1(n12065), .A2(n12540), .ZN(n12583) );
  MUX2_X1 U14274 ( .A(n12631), .B(n12630), .S(n12541), .Z(n11369) );
  AND2_X1 U14275 ( .A1(n11373), .A2(n18900), .ZN(n11368) );
  NAND2_X1 U14276 ( .A1(n12065), .A2(n12581), .ZN(n11367) );
  NAND3_X1 U14277 ( .A1(n11369), .A2(n11368), .A3(n11367), .ZN(n11372) );
  INV_X1 U14278 ( .A(n11370), .ZN(n11371) );
  NAND3_X1 U14279 ( .A1(n11372), .A2(n9634), .A3(n11371), .ZN(n12588) );
  NAND2_X1 U14280 ( .A1(n11375), .A2(n11374), .ZN(n12443) );
  AND2_X1 U14281 ( .A1(n18900), .A2(n12005), .ZN(n11376) );
  NAND2_X1 U14282 ( .A1(n12443), .A2(n11376), .ZN(n11854) );
  INV_X1 U14283 ( .A(n12859), .ZN(n11377) );
  NAND3_X1 U14284 ( .A1(n11854), .A2(n11832), .A3(n11377), .ZN(n11378) );
  NOR2_X1 U14285 ( .A1(n11382), .A2(n15904), .ZN(n11379) );
  NAND2_X1 U14286 ( .A1(n15904), .A2(n13706), .ZN(n12857) );
  NAND2_X1 U14287 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11380) );
  NAND2_X1 U14288 ( .A1(n12857), .A2(n11380), .ZN(n11381) );
  AOI21_X1 U14289 ( .B1(n11888), .B2(P2_REIP_REG_0__SCAN_IN), .A(n11381), .ZN(
        n11384) );
  NAND2_X1 U14290 ( .A1(n14452), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n11383) );
  NAND4_X1 U14291 ( .A1(n11385), .A2(n11444), .A3(n11384), .A4(n11383), .ZN(
        n11395) );
  NAND2_X1 U14292 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n11386) );
  NAND2_X1 U14293 ( .A1(n11949), .A2(n11386), .ZN(n11387) );
  OAI21_X1 U14294 ( .B1(n11389), .B2(n11388), .A(n11387), .ZN(n11393) );
  NAND2_X1 U14295 ( .A1(n11445), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11390) );
  AND2_X1 U14296 ( .A1(n11391), .A2(n11390), .ZN(n11392) );
  NAND2_X1 U14297 ( .A1(n11393), .A2(n11392), .ZN(n11394) );
  OR2_X1 U14298 ( .A1(n11395), .A2(n11394), .ZN(n11397) );
  NAND2_X1 U14299 ( .A1(n12631), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11398) );
  NOR2_X1 U14300 ( .A1(n19533), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11399) );
  AOI21_X1 U14301 ( .B1(n11459), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n11399), .ZN(n11400) );
  INV_X1 U14302 ( .A(n12664), .ZN(n13709) );
  NAND2_X1 U14303 ( .A1(n11716), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11404) );
  INV_X1 U14304 ( .A(n11404), .ZN(n11403) );
  NAND2_X1 U14305 ( .A1(n13709), .A2(n11403), .ZN(n11405) );
  NAND2_X1 U14306 ( .A1(n12664), .A2(n11404), .ZN(n11415) );
  NAND2_X1 U14307 ( .A1(n12209), .A2(n12846), .ZN(n12832) );
  INV_X1 U14308 ( .A(n11406), .ZN(n11407) );
  OR2_X2 U14309 ( .A1(n12832), .A2(n11407), .ZN(n12811) );
  AOI22_X1 U14310 ( .A1(n12811), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n11445), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11408) );
  INV_X1 U14311 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n11412) );
  NAND2_X1 U14312 ( .A1(n11888), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11411) );
  NAND2_X1 U14313 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11410) );
  OAI211_X1 U14314 ( .C1(n11949), .C2(n11412), .A(n11411), .B(n11410), .ZN(
        n11413) );
  AOI21_X2 U14315 ( .B1(n11448), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n11413), .ZN(n11418) );
  NAND2_X1 U14316 ( .A1(n11459), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11414) );
  XNOR2_X1 U14317 ( .A(n19571), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19021) );
  INV_X1 U14318 ( .A(n19533), .ZN(n19333) );
  NAND2_X1 U14319 ( .A1(n19021), .A2(n19333), .ZN(n19194) );
  NAND2_X1 U14320 ( .A1(n11419), .A2(n11418), .ZN(n11420) );
  NAND2_X2 U14321 ( .A1(n11424), .A2(n11423), .ZN(n11443) );
  AOI21_X1 U14322 ( .B1(n15904), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n11425) );
  INV_X1 U14323 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n11427) );
  NAND2_X1 U14324 ( .A1(n11888), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11426) );
  AOI21_X2 U14325 ( .B1(n11448), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n11428), .ZN(n11431) );
  INV_X1 U14326 ( .A(n11431), .ZN(n11429) );
  NAND2_X1 U14327 ( .A1(n11430), .A2(n11429), .ZN(n11433) );
  INV_X1 U14328 ( .A(n11430), .ZN(n11432) );
  NAND2_X2 U14329 ( .A1(n11432), .A2(n11431), .ZN(n11441) );
  NAND2_X2 U14330 ( .A1(n11433), .A2(n11441), .ZN(n11442) );
  XNOR2_X2 U14331 ( .A(n11443), .B(n11442), .ZN(n13233) );
  NAND2_X1 U14332 ( .A1(n13233), .A2(n12461), .ZN(n11437) );
  NAND2_X1 U14333 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19227) );
  NAND2_X1 U14334 ( .A1(n19227), .A2(n19550), .ZN(n11434) );
  NOR2_X1 U14335 ( .A1(n19550), .A2(n19560), .ZN(n19332) );
  NAND2_X1 U14336 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19332), .ZN(
        n18882) );
  NAND2_X1 U14337 ( .A1(n11434), .A2(n18882), .ZN(n19020) );
  NOR2_X1 U14338 ( .A1(n19020), .A2(n19533), .ZN(n11435) );
  AOI21_X1 U14339 ( .B1(n11459), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11435), .ZN(n11436) );
  NAND2_X1 U14340 ( .A1(n11438), .A2(n9729), .ZN(n11439) );
  NAND2_X1 U14341 ( .A1(n11445), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11446) );
  INV_X1 U14342 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n12222) );
  NAND2_X1 U14343 ( .A1(n11888), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11450) );
  NAND2_X1 U14344 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11449) );
  OAI211_X1 U14345 ( .C1(n11957), .C2(n12222), .A(n11450), .B(n11449), .ZN(
        n11451) );
  NAND2_X1 U14346 ( .A1(n11452), .A2(n11453), .ZN(n11885) );
  INV_X1 U14347 ( .A(n11452), .ZN(n11455) );
  INV_X1 U14348 ( .A(n11453), .ZN(n11454) );
  NAND2_X1 U14349 ( .A1(n11455), .A2(n11454), .ZN(n11456) );
  AND2_X2 U14350 ( .A1(n11885), .A2(n11456), .ZN(n11886) );
  XNOR2_X2 U14351 ( .A(n11887), .B(n11886), .ZN(n13226) );
  NAND2_X1 U14352 ( .A1(n13226), .A2(n12461), .ZN(n11461) );
  NAND2_X1 U14353 ( .A1(n19332), .A2(n12827), .ZN(n19106) );
  INV_X1 U14354 ( .A(n19106), .ZN(n11457) );
  INV_X1 U14355 ( .A(n19135), .ZN(n19132) );
  NAND2_X1 U14356 ( .A1(n18882), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11458) );
  AOI21_X1 U14357 ( .B1(n19132), .B2(n11458), .A(n19533), .ZN(n19258) );
  AOI21_X1 U14358 ( .B1(n11459), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19258), .ZN(n11460) );
  NAND2_X1 U14359 ( .A1(n11716), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n11463) );
  NAND2_X1 U14360 ( .A1(n12658), .A2(n12659), .ZN(n11467) );
  INV_X1 U14361 ( .A(n11463), .ZN(n11465) );
  AND2_X1 U14362 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n12631), .ZN(
        n11464) );
  INV_X1 U14363 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13316) );
  INV_X1 U14364 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11747) );
  INV_X1 U14365 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12765) );
  INV_X1 U14366 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11809) );
  AND2_X2 U14367 ( .A1(n11777), .A2(n9952), .ZN(n12129) );
  AOI22_X1 U14368 ( .A1(n11629), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12129), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11474) );
  AOI22_X1 U14369 ( .A1(n11618), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12032), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11473) );
  AOI22_X1 U14370 ( .A1(n9604), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12034), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11472) );
  AND2_X2 U14371 ( .A1(n11348), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11574) );
  AND2_X2 U14372 ( .A1(n11348), .A2(n9952), .ZN(n12147) );
  AOI22_X1 U14373 ( .A1(n11574), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11471) );
  NAND4_X1 U14374 ( .A1(n11474), .A2(n11473), .A3(n11472), .A4(n11471), .ZN(
        n11481) );
  AOI22_X1 U14375 ( .A1(n11533), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9639), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11479) );
  AND2_X2 U14376 ( .A1(n11815), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12033) );
  AND2_X2 U14377 ( .A1(n9627), .A2(n9952), .ZN(n12148) );
  AOI22_X1 U14378 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12148), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11478) );
  AND2_X2 U14379 ( .A1(n12795), .A2(n11656), .ZN(n12136) );
  AND2_X2 U14380 ( .A1(n11656), .A2(n11475), .ZN(n12135) );
  AOI22_X1 U14381 ( .A1(n12136), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12135), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11477) );
  AND2_X2 U14382 ( .A1(n12796), .A2(n11656), .ZN(n12138) );
  AND2_X2 U14383 ( .A1(n11656), .A2(n12774), .ZN(n12137) );
  AOI22_X1 U14384 ( .A1(n12138), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11476) );
  NAND4_X1 U14385 ( .A1(n11479), .A2(n11478), .A3(n11477), .A4(n11476), .ZN(
        n11480) );
  NOR2_X1 U14386 ( .A1(n11481), .A2(n11480), .ZN(n12947) );
  AOI22_X1 U14387 ( .A1(n11629), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9604), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11485) );
  AOI22_X1 U14388 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n11618), .B1(
        n12034), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11484) );
  AOI22_X1 U14389 ( .A1(n12129), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12032), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11483) );
  AOI22_X1 U14390 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n11574), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11482) );
  NAND4_X1 U14391 ( .A1(n11485), .A2(n11484), .A3(n11483), .A4(n11482), .ZN(
        n11491) );
  AOI22_X1 U14392 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11533), .B1(
        n9639), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11489) );
  AOI22_X1 U14393 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12033), .B1(
        n12148), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11488) );
  AOI22_X1 U14394 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12136), .B1(
        n12135), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11487) );
  AOI22_X1 U14395 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12138), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11486) );
  NAND4_X1 U14396 ( .A1(n11489), .A2(n11488), .A3(n11487), .A4(n11486), .ZN(
        n11490) );
  AOI22_X1 U14397 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n11629), .B1(
        n12129), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11495) );
  AOI22_X1 U14398 ( .A1(n11618), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12032), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11494) );
  AOI22_X1 U14399 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n11573), .B1(
        n12034), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11493) );
  AOI22_X1 U14400 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n11574), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11492) );
  NAND4_X1 U14401 ( .A1(n11495), .A2(n11494), .A3(n11493), .A4(n11492), .ZN(
        n11502) );
  AOI22_X1 U14402 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n11533), .B1(
        n9639), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11500) );
  AOI22_X1 U14403 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n12033), .B1(
        n12148), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11499) );
  AOI22_X1 U14404 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12136), .B1(
        n12135), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11498) );
  AOI22_X1 U14405 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n12138), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11497) );
  NAND4_X1 U14406 ( .A1(n11500), .A2(n11499), .A3(n11498), .A4(n11497), .ZN(
        n11501) );
  NOR2_X1 U14407 ( .A1(n11502), .A2(n11501), .ZN(n12965) );
  AOI22_X1 U14408 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n11629), .B1(
        n12129), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11512) );
  AOI22_X1 U14409 ( .A1(n11618), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12032), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11511) );
  AOI22_X1 U14410 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n12034), .B1(
        n9604), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11510) );
  INV_X1 U14411 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11507) );
  INV_X1 U14412 ( .A(n12147), .ZN(n11506) );
  INV_X1 U14413 ( .A(n11574), .ZN(n11505) );
  INV_X1 U14414 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13230) );
  OAI22_X1 U14415 ( .A1(n11507), .A2(n11506), .B1(n11505), .B2(n13230), .ZN(
        n11508) );
  INV_X1 U14416 ( .A(n11508), .ZN(n11509) );
  NAND4_X1 U14417 ( .A1(n11512), .A2(n11511), .A3(n11510), .A4(n11509), .ZN(
        n11518) );
  AOI22_X1 U14418 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n11533), .B1(
        n9639), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11516) );
  AOI22_X1 U14419 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n12033), .B1(
        n12148), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11515) );
  AOI22_X1 U14420 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n12136), .B1(
        n12135), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11514) );
  AOI22_X1 U14421 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12138), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11513) );
  NAND4_X1 U14422 ( .A1(n11516), .A2(n11515), .A3(n11514), .A4(n11513), .ZN(
        n11517) );
  AOI22_X1 U14423 ( .A1(n11629), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12129), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11522) );
  AOI22_X1 U14424 ( .A1(n11618), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12032), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11521) );
  AOI22_X1 U14425 ( .A1(n9604), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12034), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11520) );
  AOI22_X1 U14426 ( .A1(n11574), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11519) );
  NAND4_X1 U14427 ( .A1(n11522), .A2(n11521), .A3(n11520), .A4(n11519), .ZN(
        n11528) );
  AOI22_X1 U14428 ( .A1(n11533), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9639), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11526) );
  AOI22_X1 U14429 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12148), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11525) );
  AOI22_X1 U14430 ( .A1(n12136), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12135), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11524) );
  AOI22_X1 U14431 ( .A1(n12138), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11523) );
  NAND4_X1 U14432 ( .A1(n11526), .A2(n11525), .A3(n11524), .A4(n11523), .ZN(
        n11527) );
  AOI22_X1 U14433 ( .A1(n12129), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11618), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11532) );
  AOI22_X1 U14434 ( .A1(n11629), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9604), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11531) );
  AOI22_X1 U14435 ( .A1(n12034), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12032), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11530) );
  AOI22_X1 U14436 ( .A1(n11574), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11529) );
  NAND4_X1 U14437 ( .A1(n11532), .A2(n11531), .A3(n11530), .A4(n11529), .ZN(
        n11539) );
  AOI22_X1 U14438 ( .A1(n11533), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9639), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11537) );
  AOI22_X1 U14439 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12148), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11536) );
  AOI22_X1 U14440 ( .A1(n12136), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12135), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11535) );
  AOI22_X1 U14441 ( .A1(n12138), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11534) );
  NAND4_X1 U14442 ( .A1(n11537), .A2(n11536), .A3(n11535), .A4(n11534), .ZN(
        n11538) );
  AOI22_X1 U14443 ( .A1(n11629), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12129), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11543) );
  AOI22_X1 U14444 ( .A1(n11618), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12032), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11542) );
  AOI22_X1 U14445 ( .A1(n11573), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12034), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11541) );
  AOI22_X1 U14446 ( .A1(n11574), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11540) );
  NAND4_X1 U14447 ( .A1(n11543), .A2(n11542), .A3(n11541), .A4(n11540), .ZN(
        n11549) );
  AOI22_X1 U14448 ( .A1(n11533), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9639), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11547) );
  AOI22_X1 U14449 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12148), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11546) );
  AOI22_X1 U14450 ( .A1(n12136), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12135), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11545) );
  AOI22_X1 U14451 ( .A1(n12138), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11544) );
  NAND4_X1 U14452 ( .A1(n11547), .A2(n11546), .A3(n11545), .A4(n11544), .ZN(
        n11548) );
  NOR2_X1 U14453 ( .A1(n11549), .A2(n11548), .ZN(n13118) );
  AOI22_X1 U14454 ( .A1(n11629), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12129), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11555) );
  AOI22_X1 U14455 ( .A1(n11618), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12032), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11554) );
  AOI22_X1 U14456 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n12034), .B1(
        n11573), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11553) );
  AOI22_X1 U14457 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n11574), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11552) );
  NAND4_X1 U14458 ( .A1(n11555), .A2(n11554), .A3(n11553), .A4(n11552), .ZN(
        n11561) );
  AOI22_X1 U14459 ( .A1(n11533), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9639), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11559) );
  AOI22_X1 U14460 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12148), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11558) );
  AOI22_X1 U14461 ( .A1(n12136), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12135), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11557) );
  AOI22_X1 U14462 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n12138), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11556) );
  NAND4_X1 U14463 ( .A1(n11559), .A2(n11558), .A3(n11557), .A4(n11556), .ZN(
        n11560) );
  AOI22_X1 U14464 ( .A1(n11629), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12129), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11566) );
  AOI22_X1 U14465 ( .A1(n11618), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12032), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11565) );
  AOI22_X1 U14466 ( .A1(n11573), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12034), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11564) );
  AOI22_X1 U14467 ( .A1(n11574), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11563) );
  NAND4_X1 U14468 ( .A1(n11566), .A2(n11565), .A3(n11564), .A4(n11563), .ZN(
        n11572) );
  AOI22_X1 U14469 ( .A1(n11533), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9639), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11570) );
  AOI22_X1 U14470 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12148), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11569) );
  AOI22_X1 U14471 ( .A1(n12136), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12135), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11568) );
  AOI22_X1 U14472 ( .A1(n12138), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11567) );
  NAND4_X1 U14473 ( .A1(n11570), .A2(n11569), .A3(n11568), .A4(n11567), .ZN(
        n11571) );
  NOR2_X1 U14474 ( .A1(n11572), .A2(n11571), .ZN(n13196) );
  AOI22_X1 U14475 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n11629), .B1(
        n12129), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11578) );
  AOI22_X1 U14476 ( .A1(n11618), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12032), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11577) );
  AOI22_X1 U14477 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n12034), .B1(
        n9604), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11576) );
  AOI22_X1 U14478 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n11574), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11575) );
  NAND4_X1 U14479 ( .A1(n11578), .A2(n11577), .A3(n11576), .A4(n11575), .ZN(
        n11584) );
  AOI22_X1 U14480 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11533), .B1(
        n9639), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11582) );
  AOI22_X1 U14481 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n12033), .B1(
        n12148), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11581) );
  AOI22_X1 U14482 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12136), .B1(
        n12135), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11580) );
  AOI22_X1 U14483 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12138), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11579) );
  NAND4_X1 U14484 ( .A1(n11582), .A2(n11581), .A3(n11580), .A4(n11579), .ZN(
        n11583) );
  AOI22_X1 U14485 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n11629), .B1(
        n12129), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11591) );
  INV_X1 U14486 ( .A(n11618), .ZN(n11632) );
  INV_X1 U14487 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11586) );
  INV_X1 U14488 ( .A(n12032), .ZN(n11631) );
  INV_X1 U14489 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11585) );
  OAI22_X1 U14490 ( .A1(n11632), .A2(n11586), .B1(n11631), .B2(n11585), .ZN(
        n11587) );
  INV_X1 U14491 ( .A(n11587), .ZN(n11590) );
  AOI22_X1 U14492 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n12034), .B1(
        n11573), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11589) );
  AOI22_X1 U14493 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n11574), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11588) );
  NAND4_X1 U14494 ( .A1(n11591), .A2(n11590), .A3(n11589), .A4(n11588), .ZN(
        n11597) );
  AOI22_X1 U14495 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n11533), .B1(
        n9639), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11595) );
  AOI22_X1 U14496 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n12033), .B1(
        n12148), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11594) );
  AOI22_X1 U14497 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n12136), .B1(
        n12135), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11593) );
  AOI22_X1 U14498 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12138), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11592) );
  NAND4_X1 U14499 ( .A1(n11595), .A2(n11594), .A3(n11593), .A4(n11592), .ZN(
        n11596) );
  NOR2_X1 U14500 ( .A1(n11597), .A2(n11596), .ZN(n13420) );
  AOI22_X1 U14501 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n11629), .B1(
        n12129), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11601) );
  AOI22_X1 U14502 ( .A1(n11618), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12032), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11600) );
  AOI22_X1 U14503 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n12034), .B1(
        n9604), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11599) );
  AOI22_X1 U14504 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n11574), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11598) );
  NAND4_X1 U14505 ( .A1(n11601), .A2(n11600), .A3(n11599), .A4(n11598), .ZN(
        n11607) );
  AOI22_X1 U14506 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n11533), .B1(
        n9639), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11605) );
  AOI22_X1 U14507 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n12033), .B1(
        n12148), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11604) );
  AOI22_X1 U14508 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12136), .B1(
        n12135), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11603) );
  AOI22_X1 U14509 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n12138), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11602) );
  NAND4_X1 U14510 ( .A1(n11605), .A2(n11604), .A3(n11603), .A4(n11602), .ZN(
        n11606) );
  NOR2_X1 U14511 ( .A1(n11607), .A2(n11606), .ZN(n14533) );
  AOI22_X1 U14512 ( .A1(n11629), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12129), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11611) );
  AOI22_X1 U14513 ( .A1(n11618), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12032), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11610) );
  AOI22_X1 U14514 ( .A1(n11573), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12034), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11609) );
  AOI22_X1 U14515 ( .A1(n11574), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11608) );
  NAND4_X1 U14516 ( .A1(n11611), .A2(n11610), .A3(n11609), .A4(n11608), .ZN(
        n11617) );
  AOI22_X1 U14517 ( .A1(n11533), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9639), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11615) );
  AOI22_X1 U14518 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12148), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11614) );
  AOI22_X1 U14519 ( .A1(n12136), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12135), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11613) );
  AOI22_X1 U14520 ( .A1(n12138), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11612) );
  NAND4_X1 U14521 ( .A1(n11615), .A2(n11614), .A3(n11613), .A4(n11612), .ZN(
        n11616) );
  OR2_X1 U14522 ( .A1(n11617), .A2(n11616), .ZN(n14526) );
  AOI22_X1 U14523 ( .A1(n11629), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12129), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11622) );
  AOI22_X1 U14524 ( .A1(n11618), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12032), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11621) );
  AOI22_X1 U14525 ( .A1(n11573), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12034), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11620) );
  AOI22_X1 U14526 ( .A1(n11574), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11619) );
  NAND4_X1 U14527 ( .A1(n11622), .A2(n11621), .A3(n11620), .A4(n11619), .ZN(
        n11628) );
  AOI22_X1 U14528 ( .A1(n11533), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9639), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11626) );
  AOI22_X1 U14529 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12148), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11625) );
  AOI22_X1 U14530 ( .A1(n12136), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12135), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11624) );
  AOI22_X1 U14531 ( .A1(n12138), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11623) );
  NAND4_X1 U14532 ( .A1(n11626), .A2(n11625), .A3(n11624), .A4(n11623), .ZN(
        n11627) );
  OR2_X1 U14533 ( .A1(n11628), .A2(n11627), .ZN(n14520) );
  AOI22_X1 U14534 ( .A1(n11629), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12129), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11637) );
  INV_X1 U14535 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11630) );
  OAI22_X1 U14536 ( .A1(n11632), .A2(n12765), .B1(n11631), .B2(n11630), .ZN(
        n11633) );
  INV_X1 U14537 ( .A(n11633), .ZN(n11636) );
  AOI22_X1 U14538 ( .A1(n9604), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12034), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11635) );
  AOI22_X1 U14539 ( .A1(n11574), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11634) );
  NAND4_X1 U14540 ( .A1(n11637), .A2(n11636), .A3(n11635), .A4(n11634), .ZN(
        n11643) );
  AOI22_X1 U14541 ( .A1(n11533), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9639), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11641) );
  AOI22_X1 U14542 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12148), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11640) );
  AOI22_X1 U14543 ( .A1(n12136), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12135), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11639) );
  AOI22_X1 U14544 ( .A1(n12138), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11638) );
  NAND4_X1 U14545 ( .A1(n11641), .A2(n11640), .A3(n11639), .A4(n11638), .ZN(
        n11642) );
  NOR2_X1 U14546 ( .A1(n11643), .A2(n11642), .ZN(n14516) );
  AOI22_X1 U14547 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n11629), .B1(
        n12129), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11647) );
  AOI22_X1 U14548 ( .A1(n11618), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12032), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11646) );
  AOI22_X1 U14549 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n9604), .B1(
        n12034), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11645) );
  AOI22_X1 U14550 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n11574), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11644) );
  NAND4_X1 U14551 ( .A1(n11647), .A2(n11646), .A3(n11645), .A4(n11644), .ZN(
        n11653) );
  AOI22_X1 U14552 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n11533), .B1(
        n9639), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11651) );
  AOI22_X1 U14553 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n12033), .B1(
        n12148), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11650) );
  AOI22_X1 U14554 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n12136), .B1(
        n12135), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11649) );
  AOI22_X1 U14555 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12138), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11648) );
  NAND4_X1 U14556 ( .A1(n11651), .A2(n11650), .A3(n11649), .A4(n11648), .ZN(
        n11652) );
  NOR2_X1 U14557 ( .A1(n11653), .A2(n11652), .ZN(n11677) );
  INV_X1 U14558 ( .A(n11677), .ZN(n11676) );
  AOI22_X1 U14559 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11816), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11665) );
  AOI22_X1 U14560 ( .A1(n9624), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(n9605), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11664) );
  INV_X1 U14561 ( .A(n11654), .ZN(n11655) );
  AOI22_X1 U14562 ( .A1(n9627), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11801), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11663) );
  INV_X1 U14563 ( .A(n11804), .ZN(n11810) );
  INV_X1 U14564 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11660) );
  NAND2_X1 U14565 ( .A1(n9635), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11659) );
  INV_X1 U14566 ( .A(n11656), .ZN(n11658) );
  NAND2_X1 U14567 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11657) );
  NAND2_X1 U14568 ( .A1(n11658), .A2(n11657), .ZN(n11808) );
  OAI211_X1 U14569 ( .C1(n11810), .C2(n11660), .A(n11659), .B(n11808), .ZN(
        n11661) );
  INV_X1 U14570 ( .A(n11661), .ZN(n11662) );
  NAND4_X1 U14571 ( .A1(n11665), .A2(n11664), .A3(n11663), .A4(n11662), .ZN(
        n11674) );
  AOI22_X1 U14572 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9638), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11672) );
  AOI22_X1 U14573 ( .A1(n9623), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(n9607), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11671) );
  AOI22_X1 U14574 ( .A1(n9627), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11801), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11670) );
  INV_X1 U14575 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11667) );
  NAND2_X1 U14576 ( .A1(n9635), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11666) );
  INV_X1 U14577 ( .A(n11808), .ZN(n11769) );
  OAI211_X1 U14578 ( .C1(n11810), .C2(n11667), .A(n11666), .B(n11769), .ZN(
        n11668) );
  INV_X1 U14579 ( .A(n11668), .ZN(n11669) );
  NAND4_X1 U14580 ( .A1(n11672), .A2(n11671), .A3(n11670), .A4(n11669), .ZN(
        n11673) );
  NAND2_X1 U14581 ( .A1(n11674), .A2(n11673), .ZN(n11680) );
  INV_X1 U14582 ( .A(n11680), .ZN(n11675) );
  NAND2_X1 U14583 ( .A1(n11676), .A2(n11675), .ZN(n11698) );
  OAI21_X1 U14584 ( .B1(n18895), .B2(n11680), .A(n11677), .ZN(n11678) );
  OAI21_X1 U14585 ( .B1(n11698), .B2(n18895), .A(n11678), .ZN(n11700) );
  NOR2_X1 U14586 ( .A1(n9643), .A2(n11680), .ZN(n14507) );
  AOI22_X1 U14587 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11816), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11688) );
  AOI22_X1 U14588 ( .A1(n9623), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(n9606), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11687) );
  AOI22_X1 U14589 ( .A1(n11815), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11801), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11686) );
  INV_X1 U14590 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11683) );
  NAND2_X1 U14591 ( .A1(n9635), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11682) );
  OAI211_X1 U14592 ( .C1(n11810), .C2(n11683), .A(n11682), .B(n11769), .ZN(
        n11684) );
  INV_X1 U14593 ( .A(n11684), .ZN(n11685) );
  NAND4_X1 U14594 ( .A1(n11688), .A2(n11687), .A3(n11686), .A4(n11685), .ZN(
        n11697) );
  AOI22_X1 U14595 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11695) );
  AOI22_X1 U14596 ( .A1(n11816), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11801), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11694) );
  AOI22_X1 U14597 ( .A1(n9624), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(n9635), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11693) );
  INV_X1 U14598 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11690) );
  NAND2_X1 U14599 ( .A1(n11815), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11689) );
  OAI211_X1 U14600 ( .C1(n11810), .C2(n11690), .A(n11689), .B(n11808), .ZN(
        n11691) );
  INV_X1 U14601 ( .A(n11691), .ZN(n11692) );
  NAND4_X1 U14602 ( .A1(n11695), .A2(n11694), .A3(n11693), .A4(n11692), .ZN(
        n11696) );
  NAND2_X1 U14603 ( .A1(n11697), .A2(n11696), .ZN(n14496) );
  NOR2_X1 U14604 ( .A1(n11698), .A2(n14496), .ZN(n11717) );
  AOI211_X1 U14605 ( .C1(n14496), .C2(n11698), .A(n11762), .B(n11717), .ZN(
        n14498) );
  INV_X1 U14606 ( .A(n14507), .ZN(n11699) );
  AOI22_X1 U14607 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11816), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11706) );
  AOI22_X1 U14608 ( .A1(n9624), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(n9606), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11705) );
  AOI22_X1 U14609 ( .A1(n11815), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11801), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11704) );
  NAND2_X1 U14610 ( .A1(n9635), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11701) );
  OAI211_X1 U14611 ( .C1(n11810), .C2(n11586), .A(n11701), .B(n11808), .ZN(
        n11702) );
  INV_X1 U14612 ( .A(n11702), .ZN(n11703) );
  NAND4_X1 U14613 ( .A1(n11706), .A2(n11705), .A3(n11704), .A4(n11703), .ZN(
        n11715) );
  AOI22_X1 U14614 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9638), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11713) );
  AOI22_X1 U14615 ( .A1(n11777), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9605), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11712) );
  AOI22_X1 U14616 ( .A1(n11815), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11801), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11711) );
  INV_X1 U14617 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11708) );
  NAND2_X1 U14618 ( .A1(n9635), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n11707) );
  OAI211_X1 U14619 ( .C1(n11810), .C2(n11708), .A(n11707), .B(n11769), .ZN(
        n11709) );
  INV_X1 U14620 ( .A(n11709), .ZN(n11710) );
  NAND4_X1 U14621 ( .A1(n11713), .A2(n11712), .A3(n11711), .A4(n11710), .ZN(
        n11714) );
  AND2_X1 U14622 ( .A1(n11715), .A2(n11714), .ZN(n11719) );
  NAND2_X1 U14623 ( .A1(n11717), .A2(n11719), .ZN(n11740) );
  OAI211_X1 U14624 ( .C1(n11717), .C2(n11719), .A(n11740), .B(n11716), .ZN(
        n11721) );
  INV_X1 U14625 ( .A(n11721), .ZN(n11718) );
  INV_X1 U14626 ( .A(n11719), .ZN(n11720) );
  NOR2_X1 U14627 ( .A1(n9643), .A2(n11720), .ZN(n14489) );
  AOI22_X1 U14628 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(n9624), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11730) );
  AOI22_X1 U14629 ( .A1(n9605), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11801), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11729) );
  AOI22_X1 U14630 ( .A1(n9638), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(n9635), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11728) );
  INV_X1 U14631 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11725) );
  NAND2_X1 U14632 ( .A1(n11815), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11724) );
  OAI211_X1 U14633 ( .C1(n11810), .C2(n11725), .A(n11724), .B(n11808), .ZN(
        n11726) );
  INV_X1 U14634 ( .A(n11726), .ZN(n11727) );
  NAND4_X1 U14635 ( .A1(n11730), .A2(n11729), .A3(n11728), .A4(n11727), .ZN(
        n11739) );
  AOI22_X1 U14636 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9623), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11737) );
  AOI22_X1 U14637 ( .A1(n9638), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11801), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11736) );
  AOI22_X1 U14638 ( .A1(n9607), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9635), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11735) );
  INV_X1 U14639 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11732) );
  NAND2_X1 U14640 ( .A1(n9627), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11731) );
  OAI211_X1 U14641 ( .C1(n11810), .C2(n11732), .A(n11731), .B(n11769), .ZN(
        n11733) );
  INV_X1 U14642 ( .A(n11733), .ZN(n11734) );
  NAND4_X1 U14643 ( .A1(n11737), .A2(n11736), .A3(n11735), .A4(n11734), .ZN(
        n11738) );
  NAND2_X1 U14644 ( .A1(n11739), .A2(n11738), .ZN(n11742) );
  AOI21_X1 U14645 ( .B1(n11740), .B2(n11742), .A(n11762), .ZN(n11741) );
  NAND2_X1 U14646 ( .A1(n11741), .A2(n11763), .ZN(n11743) );
  NOR2_X1 U14647 ( .A1(n9643), .A2(n11742), .ZN(n14482) );
  INV_X1 U14648 ( .A(n11743), .ZN(n11744) );
  AOI22_X1 U14649 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(n9638), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11752) );
  AOI22_X1 U14650 ( .A1(n9624), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(n9607), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11751) );
  AOI22_X1 U14651 ( .A1(n11815), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11801), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11750) );
  NAND2_X1 U14652 ( .A1(n9635), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11746) );
  OAI211_X1 U14653 ( .C1(n11810), .C2(n11747), .A(n11746), .B(n11808), .ZN(
        n11748) );
  INV_X1 U14654 ( .A(n11748), .ZN(n11749) );
  NAND4_X1 U14655 ( .A1(n11752), .A2(n11751), .A3(n11750), .A4(n11749), .ZN(
        n11761) );
  AOI22_X1 U14656 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11816), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11759) );
  AOI22_X1 U14657 ( .A1(n9624), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n9606), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11758) );
  AOI22_X1 U14658 ( .A1(n9627), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11801), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11757) );
  INV_X1 U14659 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11754) );
  NAND2_X1 U14660 ( .A1(n9635), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11753) );
  OAI211_X1 U14661 ( .C1(n11810), .C2(n11754), .A(n11753), .B(n11769), .ZN(
        n11755) );
  INV_X1 U14662 ( .A(n11755), .ZN(n11756) );
  NAND4_X1 U14663 ( .A1(n11759), .A2(n11758), .A3(n11757), .A4(n11756), .ZN(
        n11760) );
  NAND2_X1 U14664 ( .A1(n11761), .A2(n11760), .ZN(n11765) );
  AOI21_X1 U14665 ( .B1(n11763), .B2(n11765), .A(n11762), .ZN(n11764) );
  NAND2_X1 U14666 ( .A1(n11764), .A2(n11786), .ZN(n11767) );
  INV_X1 U14667 ( .A(n11765), .ZN(n11766) );
  NAND2_X1 U14668 ( .A1(n18895), .A2(n11766), .ZN(n14477) );
  AOI22_X1 U14669 ( .A1(n9625), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9623), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11776) );
  AOI22_X1 U14670 ( .A1(n11816), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11801), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11775) );
  AOI22_X1 U14671 ( .A1(n9606), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9627), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11774) );
  INV_X1 U14672 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11771) );
  NAND2_X1 U14673 ( .A1(n9635), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11770) );
  OAI211_X1 U14674 ( .C1(n11810), .C2(n11771), .A(n11770), .B(n11769), .ZN(
        n11772) );
  INV_X1 U14675 ( .A(n11772), .ZN(n11773) );
  NAND4_X1 U14676 ( .A1(n11776), .A2(n11775), .A3(n11774), .A4(n11773), .ZN(
        n11785) );
  AOI22_X1 U14677 ( .A1(n11777), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11816), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11783) );
  AOI22_X1 U14678 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11801), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11782) );
  AOI22_X1 U14679 ( .A1(n9605), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(n9635), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11781) );
  NAND2_X1 U14680 ( .A1(n9627), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11778) );
  OAI211_X1 U14681 ( .C1(n11810), .C2(n13316), .A(n11778), .B(n11808), .ZN(
        n11779) );
  INV_X1 U14682 ( .A(n11779), .ZN(n11780) );
  NAND4_X1 U14683 ( .A1(n11783), .A2(n11782), .A3(n11781), .A4(n11780), .ZN(
        n11784) );
  AND2_X1 U14684 ( .A1(n11785), .A2(n11784), .ZN(n14469) );
  INV_X1 U14685 ( .A(n11786), .ZN(n14466) );
  NAND3_X1 U14686 ( .A1(n14466), .A2(n14469), .A3(n12005), .ZN(n11800) );
  AOI22_X1 U14687 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9638), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11788) );
  AOI22_X1 U14688 ( .A1(n9624), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(n9607), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11787) );
  NAND2_X1 U14689 ( .A1(n11788), .A2(n11787), .ZN(n11798) );
  INV_X1 U14690 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13452) );
  AOI22_X1 U14691 ( .A1(n9627), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11801), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11790) );
  AOI21_X1 U14692 ( .B1(n11804), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n11808), .ZN(n11789) );
  OAI211_X1 U14693 ( .C1(n9617), .C2(n13452), .A(n11790), .B(n11789), .ZN(
        n11797) );
  OAI21_X1 U14694 ( .B1(n11810), .B2(n12765), .A(n11808), .ZN(n11792) );
  INV_X1 U14695 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13460) );
  INV_X1 U14696 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13444) );
  OAI22_X1 U14697 ( .A1(n9628), .A2(n13460), .B1(n11655), .B2(n13444), .ZN(
        n11791) );
  AOI211_X1 U14698 ( .C1(n9635), .C2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n11792), .B(n11791), .ZN(n11795) );
  AOI22_X1 U14699 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11816), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11794) );
  AOI22_X1 U14700 ( .A1(n9623), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(n9605), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11793) );
  NAND3_X1 U14701 ( .A1(n11795), .A2(n11794), .A3(n11793), .ZN(n11796) );
  OAI21_X1 U14702 ( .B1(n11798), .B2(n11797), .A(n11796), .ZN(n11799) );
  XNOR2_X1 U14703 ( .A(n11800), .B(n11799), .ZN(n14460) );
  AOI22_X1 U14704 ( .A1(n9624), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11816), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11803) );
  AOI22_X1 U14705 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11801), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11802) );
  NAND2_X1 U14706 ( .A1(n11803), .A2(n11802), .ZN(n11822) );
  INV_X1 U14707 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11807) );
  AOI22_X1 U14708 ( .A1(n9606), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9635), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11806) );
  AOI21_X1 U14709 ( .B1(n11804), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n11808), .ZN(n11805) );
  OAI211_X1 U14710 ( .C1(n9628), .C2(n11807), .A(n11806), .B(n11805), .ZN(
        n11821) );
  OAI21_X1 U14711 ( .B1(n11810), .B2(n11809), .A(n11808), .ZN(n11814) );
  INV_X1 U14712 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11812) );
  INV_X1 U14713 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11811) );
  OAI22_X1 U14714 ( .A1(n9617), .A2(n11812), .B1(n11655), .B2(n11811), .ZN(
        n11813) );
  AOI211_X1 U14715 ( .C1(n9627), .C2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n11814), .B(n11813), .ZN(n11819) );
  AOI22_X1 U14716 ( .A1(n9625), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11816), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11818) );
  AOI22_X1 U14717 ( .A1(n9623), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(n9607), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11817) );
  NAND3_X1 U14718 ( .A1(n11819), .A2(n11818), .A3(n11817), .ZN(n11820) );
  OAI21_X1 U14719 ( .B1(n11822), .B2(n11821), .A(n11820), .ZN(n11823) );
  INV_X1 U14720 ( .A(n11837), .ZN(n11824) );
  NAND2_X1 U14721 ( .A1(n12435), .A2(n11824), .ZN(n11826) );
  NAND2_X1 U14722 ( .A1(n19560), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11825) );
  NAND2_X1 U14723 ( .A1(n11826), .A2(n11825), .ZN(n11834) );
  INV_X1 U14724 ( .A(n11833), .ZN(n11828) );
  NAND2_X1 U14725 ( .A1(n11834), .A2(n11828), .ZN(n11830) );
  NAND2_X1 U14726 ( .A1(n19550), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11829) );
  MUX2_X1 U14727 ( .A(n12827), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n11844) );
  NOR2_X1 U14728 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15419), .ZN(
        n11831) );
  INV_X1 U14729 ( .A(n12442), .ZN(n11850) );
  NAND2_X1 U14730 ( .A1(n11852), .A2(n9643), .ZN(n11835) );
  XNOR2_X1 U14731 ( .A(n11834), .B(n11833), .ZN(n12204) );
  MUX2_X1 U14732 ( .A(n11835), .B(n11382), .S(n12204), .Z(n11842) );
  INV_X1 U14733 ( .A(n12204), .ZN(n12216) );
  INV_X1 U14734 ( .A(n12435), .ZN(n11836) );
  OAI21_X1 U14735 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19571), .A(
        n11837), .ZN(n12456) );
  OAI21_X1 U14736 ( .B1(n11836), .B2(n12456), .A(n12455), .ZN(n11839) );
  INV_X1 U14737 ( .A(n12456), .ZN(n12436) );
  XNOR2_X1 U14738 ( .A(n12435), .B(n11837), .ZN(n12206) );
  OAI211_X1 U14739 ( .C1(n9643), .C2(n12436), .A(n9634), .B(n12206), .ZN(
        n11838) );
  OAI211_X1 U14740 ( .C1(n11840), .C2(n12216), .A(n11839), .B(n11838), .ZN(
        n11841) );
  NAND2_X1 U14741 ( .A1(n11842), .A2(n11841), .ZN(n11848) );
  NOR2_X1 U14742 ( .A1(n11845), .A2(n11844), .ZN(n11846) );
  MUX2_X1 U14743 ( .A(n11382), .B(n11848), .S(n12440), .Z(n11849) );
  NAND2_X1 U14744 ( .A1(n11850), .A2(n11849), .ZN(n11851) );
  MUX2_X1 U14745 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n11851), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n12530) );
  NAND2_X1 U14746 ( .A1(n12442), .A2(n18705), .ZN(n11853) );
  NOR2_X1 U14747 ( .A1(n12794), .A2(n11854), .ZN(n12778) );
  NAND2_X1 U14748 ( .A1(n12839), .A2(n12778), .ZN(n12785) );
  INV_X1 U14749 ( .A(n12775), .ZN(n11855) );
  NAND2_X1 U14750 ( .A1(n12785), .A2(n11855), .ZN(n11857) );
  NAND2_X1 U14751 ( .A1(n13706), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19440) );
  INV_X1 U14752 ( .A(n19440), .ZN(n11856) );
  NAND2_X1 U14753 ( .A1(n14552), .A2(n14522), .ZN(n11962) );
  NAND2_X1 U14754 ( .A1(n11933), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11863) );
  INV_X1 U14755 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n11860) );
  NAND2_X1 U14756 ( .A1(n14451), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11859) );
  NAND2_X1 U14757 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11858) );
  OAI211_X1 U14758 ( .C1(n11957), .C2(n11860), .A(n11859), .B(n11858), .ZN(
        n11861) );
  INV_X1 U14759 ( .A(n11861), .ZN(n11862) );
  NAND2_X1 U14760 ( .A1(n11863), .A2(n11862), .ZN(n13120) );
  INV_X4 U14761 ( .A(n11895), .ZN(n11933) );
  INV_X1 U14762 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n11866) );
  NAND2_X1 U14763 ( .A1(n14451), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11865) );
  NAND2_X1 U14764 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11864) );
  OAI211_X1 U14765 ( .C1(n11957), .C2(n11866), .A(n11865), .B(n11864), .ZN(
        n11867) );
  AOI21_X1 U14766 ( .B1(n11933), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n11867), .ZN(n13050) );
  INV_X1 U14767 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n11870) );
  NAND2_X1 U14768 ( .A1(n14451), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n11869) );
  NAND2_X1 U14769 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11868) );
  OAI211_X1 U14770 ( .C1(n11957), .C2(n11870), .A(n11869), .B(n11868), .ZN(
        n11871) );
  AOI21_X1 U14771 ( .B1(n11933), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n11871), .ZN(n13027) );
  INV_X1 U14772 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n11874) );
  NAND2_X1 U14773 ( .A1(n14451), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11873) );
  NAND2_X1 U14774 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11872) );
  OAI211_X1 U14775 ( .C1(n11957), .C2(n11874), .A(n11873), .B(n11872), .ZN(
        n11875) );
  AOI21_X1 U14776 ( .B1(n11933), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n11875), .ZN(n12903) );
  NAND2_X1 U14777 ( .A1(n11933), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11881) );
  INV_X1 U14778 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n11878) );
  NAND2_X1 U14779 ( .A1(n14451), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11877) );
  NAND2_X1 U14780 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11876) );
  OAI211_X1 U14781 ( .C1(n11957), .C2(n11878), .A(n11877), .B(n11876), .ZN(
        n11879) );
  INV_X1 U14782 ( .A(n11879), .ZN(n11880) );
  NAND2_X1 U14783 ( .A1(n11881), .A2(n11880), .ZN(n12734) );
  INV_X1 U14784 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n12732) );
  NAND2_X1 U14785 ( .A1(n14451), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n11883) );
  NAND2_X1 U14786 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11882) );
  OAI211_X1 U14787 ( .C1(n11957), .C2(n12732), .A(n11883), .B(n11882), .ZN(
        n11884) );
  AOI21_X1 U14788 ( .B1(n11933), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n11884), .ZN(n12728) );
  INV_X1 U14789 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n12671) );
  NAND2_X1 U14790 ( .A1(n11933), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11890) );
  AOI22_X1 U14791 ( .A1(n14451), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11889) );
  OAI211_X1 U14792 ( .C1(n11957), .C2(n12671), .A(n11890), .B(n11889), .ZN(
        n12669) );
  INV_X1 U14793 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n12773) );
  NAND2_X1 U14794 ( .A1(n11933), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11892) );
  AOI22_X1 U14795 ( .A1(n14451), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11891) );
  OAI211_X1 U14796 ( .C1(n12773), .C2(n11949), .A(n11892), .B(n11891), .ZN(
        n12768) );
  INV_X1 U14797 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n13752) );
  AOI22_X1 U14798 ( .A1(n14451), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11894) );
  NAND2_X1 U14799 ( .A1(n14452), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11893) );
  OAI211_X1 U14800 ( .C1(n11895), .C2(n13752), .A(n11894), .B(n11893), .ZN(
        n12945) );
  NAND2_X1 U14801 ( .A1(n11933), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11897) );
  AOI22_X1 U14802 ( .A1(n14451), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n11896) );
  OAI211_X1 U14803 ( .C1(n10071), .C2(n11949), .A(n11897), .B(n11896), .ZN(
        n12967) );
  INV_X1 U14804 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n11900) );
  NAND2_X1 U14805 ( .A1(n11933), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11899) );
  AOI22_X1 U14806 ( .A1(n14451), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n11898) );
  OAI211_X1 U14807 ( .C1(n11900), .C2(n11949), .A(n11899), .B(n11898), .ZN(
        n13038) );
  INV_X1 U14808 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n11903) );
  NAND2_X1 U14809 ( .A1(n14451), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11902) );
  NAND2_X1 U14810 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11901) );
  OAI211_X1 U14811 ( .C1(n11957), .C2(n11903), .A(n11902), .B(n11901), .ZN(
        n11904) );
  AOI21_X1 U14812 ( .B1(n11933), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n11904), .ZN(n13175) );
  INV_X1 U14813 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n11907) );
  NAND2_X1 U14814 ( .A1(n14451), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11906) );
  NAND2_X1 U14815 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11905) );
  OAI211_X1 U14816 ( .C1(n11957), .C2(n11907), .A(n11906), .B(n11905), .ZN(
        n11908) );
  AOI21_X1 U14817 ( .B1(n11933), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n11908), .ZN(n13206) );
  INV_X1 U14818 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n11911) );
  NAND2_X1 U14819 ( .A1(n14451), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11910) );
  NAND2_X1 U14820 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11909) );
  OAI211_X1 U14821 ( .C1(n11957), .C2(n11911), .A(n11910), .B(n11909), .ZN(
        n11912) );
  AOI21_X1 U14822 ( .B1(n11933), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n11912), .ZN(n13415) );
  INV_X1 U14823 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n11915) );
  NAND2_X1 U14824 ( .A1(n11933), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11914) );
  AOI22_X1 U14825 ( .A1(n14451), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11913) );
  OAI211_X1 U14826 ( .C1(n11957), .C2(n11915), .A(n11914), .B(n11913), .ZN(
        n14543) );
  INV_X1 U14827 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n11918) );
  NAND2_X1 U14828 ( .A1(n14451), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11917) );
  NAND2_X1 U14829 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11916) );
  OAI211_X1 U14830 ( .C1(n11957), .C2(n11918), .A(n11917), .B(n11916), .ZN(
        n11919) );
  AOI21_X1 U14831 ( .B1(n11933), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n11919), .ZN(n14539) );
  OR2_X2 U14832 ( .A1(n14546), .A2(n14539), .ZN(n14537) );
  INV_X1 U14833 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n11922) );
  NAND2_X1 U14834 ( .A1(n14451), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11921) );
  NAND2_X1 U14835 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11920) );
  OAI211_X1 U14836 ( .C1(n11957), .C2(n11922), .A(n11921), .B(n11920), .ZN(
        n11923) );
  AOI21_X1 U14837 ( .B1(n11933), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n11923), .ZN(n14528) );
  INV_X1 U14838 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n12226) );
  NAND2_X1 U14839 ( .A1(n11933), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11925) );
  AOI22_X1 U14840 ( .A1(n14451), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n11924) );
  OAI211_X1 U14841 ( .C1(n11957), .C2(n12226), .A(n11925), .B(n11924), .ZN(
        n12256) );
  INV_X1 U14842 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n11928) );
  NAND2_X1 U14843 ( .A1(n11933), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11927) );
  AOI22_X1 U14844 ( .A1(n14451), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n11926) );
  OAI211_X1 U14845 ( .C1(n11949), .C2(n11928), .A(n11927), .B(n11926), .ZN(
        n12270) );
  INV_X1 U14846 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n11931) );
  NAND2_X1 U14847 ( .A1(n14451), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11930) );
  NAND2_X1 U14848 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n11929) );
  OAI211_X1 U14849 ( .C1(n11949), .C2(n11931), .A(n11930), .B(n11929), .ZN(
        n11932) );
  AOI21_X1 U14850 ( .B1(n11933), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n11932), .ZN(n14510) );
  NAND2_X1 U14851 ( .A1(n14451), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11935) );
  NAND2_X1 U14852 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11934) );
  OAI211_X1 U14853 ( .C1(n11949), .C2(n10064), .A(n11935), .B(n11934), .ZN(
        n11936) );
  AOI21_X1 U14854 ( .B1(n11933), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n11936), .ZN(n14501) );
  OR2_X2 U14855 ( .A1(n14509), .A2(n14501), .ZN(n14503) );
  INV_X1 U14856 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n14493) );
  NAND2_X1 U14857 ( .A1(n14451), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11938) );
  NAND2_X1 U14858 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11937) );
  OAI211_X1 U14859 ( .C1(n11949), .C2(n14493), .A(n11938), .B(n11937), .ZN(
        n11939) );
  AOI21_X1 U14860 ( .B1(n11933), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n11939), .ZN(n14492) );
  INV_X1 U14861 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n11942) );
  NAND2_X1 U14862 ( .A1(n11933), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11941) );
  AOI22_X1 U14863 ( .A1(n14451), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n11940) );
  OAI211_X1 U14864 ( .C1(n11949), .C2(n11942), .A(n11941), .B(n11940), .ZN(
        n14483) );
  INV_X1 U14865 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n11945) );
  NAND2_X1 U14866 ( .A1(n11933), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11944) );
  AOI22_X1 U14867 ( .A1(n14451), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n11943) );
  OAI211_X1 U14868 ( .C1(n11949), .C2(n11945), .A(n11944), .B(n11943), .ZN(
        n14473) );
  INV_X1 U14869 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n11948) );
  NAND2_X1 U14870 ( .A1(n11933), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11947) );
  AOI22_X1 U14871 ( .A1(n14451), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n11946) );
  OAI211_X1 U14872 ( .C1(n11949), .C2(n11948), .A(n11947), .B(n11946), .ZN(
        n14470) );
  INV_X1 U14873 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n11952) );
  NAND2_X1 U14874 ( .A1(n14451), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11951) );
  NAND2_X1 U14875 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11950) );
  OAI211_X1 U14876 ( .C1(n11957), .C2(n11952), .A(n11951), .B(n11950), .ZN(
        n11953) );
  AOI21_X1 U14877 ( .B1(n11933), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n11953), .ZN(n14463) );
  OR2_X2 U14878 ( .A1(n9681), .A2(n14463), .ZN(n14461) );
  INV_X1 U14879 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n11956) );
  NAND2_X1 U14880 ( .A1(n14451), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n11955) );
  NAND2_X1 U14881 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n11954) );
  OAI211_X1 U14882 ( .C1(n11957), .C2(n11956), .A(n11955), .B(n11954), .ZN(
        n11958) );
  AOI21_X1 U14883 ( .B1(n11933), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n11958), .ZN(n14450) );
  XNOR2_X2 U14884 ( .A(n14461), .B(n14450), .ZN(n14656) );
  NAND2_X1 U14885 ( .A1(n14548), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11959) );
  INV_X1 U14886 ( .A(n11960), .ZN(n11961) );
  NAND2_X1 U14887 ( .A1(n11962), .A2(n11961), .ZN(P2_U2857) );
  INV_X1 U14888 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11967) );
  AND2_X1 U14889 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11963) );
  INV_X1 U14890 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n14818) );
  AND2_X1 U14891 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11964) );
  INV_X1 U14892 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14710) );
  INV_X1 U14893 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14688) );
  INV_X1 U14894 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11968) );
  INV_X1 U14895 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14666) );
  NAND2_X1 U14896 ( .A1(n12000), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11966) );
  INV_X1 U14897 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11965) );
  AOI21_X1 U14898 ( .B1(n14666), .B2(n11970), .A(n12000), .ZN(n15705) );
  NAND2_X1 U14899 ( .A1(n11972), .A2(n11968), .ZN(n11969) );
  NAND2_X1 U14900 ( .A1(n11970), .A2(n11969), .ZN(n14680) );
  INV_X1 U14901 ( .A(n14680), .ZN(n15715) );
  INV_X1 U14902 ( .A(n11972), .ZN(n11973) );
  AOI21_X1 U14903 ( .B1(n14688), .B2(n11971), .A(n11973), .ZN(n15727) );
  OR2_X1 U14904 ( .A1(n11974), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11975) );
  NAND2_X1 U14905 ( .A1(n11971), .A2(n11975), .ZN(n14698) );
  INV_X1 U14906 ( .A(n14698), .ZN(n15736) );
  AOI21_X1 U14907 ( .B1(n14710), .B2(n11976), .A(n11974), .ZN(n15749) );
  OAI21_X1 U14908 ( .B1(n9748), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n11976), .ZN(n14718) );
  INV_X1 U14909 ( .A(n14718), .ZN(n15760) );
  AOI21_X1 U14910 ( .B1(n10114), .B2(n11977), .A(n9748), .ZN(n15768) );
  OAI21_X1 U14911 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n11978), .A(
        n11977), .ZN(n11979) );
  INV_X1 U14912 ( .A(n11979), .ZN(n15784) );
  AOI21_X1 U14913 ( .B1(n14742), .B2(n11981), .A(n11978), .ZN(n14746) );
  OAI21_X1 U14914 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n11980), .A(
        n11981), .ZN(n14755) );
  INV_X1 U14915 ( .A(n14755), .ZN(n18443) );
  AOI21_X1 U14916 ( .B1(n18456), .B2(n11982), .A(n11980), .ZN(n18452) );
  OR2_X1 U14917 ( .A1(n11983), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11984) );
  NAND2_X1 U14918 ( .A1(n11982), .A2(n11984), .ZN(n14778) );
  INV_X1 U14919 ( .A(n14778), .ZN(n18464) );
  INV_X1 U14920 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18479) );
  NAND2_X1 U14921 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n11985), .ZN(
        n11986) );
  AOI21_X1 U14922 ( .B1(n18479), .B2(n11986), .A(n11983), .ZN(n18475) );
  INV_X1 U14923 ( .A(n15696), .ZN(n11999) );
  OAI21_X1 U14924 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n11985), .A(
        n11986), .ZN(n18486) );
  AOI21_X1 U14925 ( .B1(n20697), .B2(n9727), .A(n11985), .ZN(n18501) );
  AOI21_X1 U14926 ( .B1(n18518), .B2(n11987), .A(n11988), .ZN(n18523) );
  AOI21_X1 U14927 ( .B1(n18541), .B2(n11989), .A(n11990), .ZN(n18548) );
  AOI21_X1 U14928 ( .B1(n15824), .B2(n11991), .A(n11992), .ZN(n18571) );
  AOI21_X1 U14929 ( .B1(n14818), .B2(n11993), .A(n11994), .ZN(n18594) );
  INV_X1 U14930 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n15843) );
  NAND2_X1 U14931 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n11995), .ZN(
        n11998) );
  AOI21_X1 U14932 ( .B1(n15843), .B2(n11998), .A(n11996), .ZN(n18621) );
  AOI21_X1 U14933 ( .B1(n15853), .B2(n11997), .A(n11995), .ZN(n15844) );
  OAI22_X1 U14934 ( .A1(n15904), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n13165) );
  INV_X1 U14935 ( .A(n13165), .ZN(n14446) );
  AOI22_X1 U14936 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n15083), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n15904), .ZN(n13110) );
  NOR2_X1 U14937 ( .A1(n14446), .A2(n13110), .ZN(n13109) );
  OAI21_X1 U14938 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n11997), .ZN(n18826) );
  NAND2_X1 U14939 ( .A1(n13109), .A2(n18826), .ZN(n13013) );
  NOR2_X1 U14940 ( .A1(n15844), .A2(n13013), .ZN(n18629) );
  OAI21_X1 U14941 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n11995), .A(
        n11998), .ZN(n18815) );
  NAND2_X1 U14942 ( .A1(n18629), .A2(n18815), .ZN(n18619) );
  NOR2_X1 U14943 ( .A1(n18621), .A2(n18619), .ZN(n18606) );
  OAI21_X1 U14944 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n11996), .A(
        n11993), .ZN(n18607) );
  NAND2_X1 U14945 ( .A1(n18606), .A2(n18607), .ZN(n18592) );
  NOR2_X1 U14946 ( .A1(n18594), .A2(n18592), .ZN(n18581) );
  OAI21_X1 U14947 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n11994), .A(
        n11991), .ZN(n18582) );
  NAND2_X1 U14948 ( .A1(n18581), .A2(n18582), .ZN(n18569) );
  NOR2_X1 U14949 ( .A1(n18571), .A2(n18569), .ZN(n18558) );
  OAI21_X1 U14950 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n11992), .A(
        n11989), .ZN(n18559) );
  NAND2_X1 U14951 ( .A1(n18558), .A2(n18559), .ZN(n18549) );
  NOR2_X1 U14952 ( .A1(n18548), .A2(n18549), .ZN(n18534) );
  OAI21_X1 U14953 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n11990), .A(
        n11987), .ZN(n18535) );
  NAND2_X1 U14954 ( .A1(n18534), .A2(n18535), .ZN(n18521) );
  NOR2_X1 U14955 ( .A1(n18523), .A2(n18521), .ZN(n18510) );
  OAI21_X1 U14956 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n11988), .A(
        n9727), .ZN(n18511) );
  NAND2_X1 U14957 ( .A1(n18510), .A2(n18511), .ZN(n18499) );
  OAI21_X1 U14958 ( .B1(n18501), .B2(n18499), .A(n13164), .ZN(n18485) );
  NOR2_X1 U14959 ( .A1(n18475), .A2(n18474), .ZN(n18473) );
  NOR2_X1 U14960 ( .A1(n18464), .A2(n18463), .ZN(n18462) );
  NOR2_X1 U14961 ( .A1(n18630), .A2(n18462), .ZN(n18451) );
  NOR2_X1 U14962 ( .A1(n18452), .A2(n18451), .ZN(n18450) );
  NOR2_X2 U14963 ( .A1(n18630), .A2(n18450), .ZN(n18442) );
  NOR2_X1 U14964 ( .A1(n15784), .A2(n12264), .ZN(n12263) );
  NOR2_X1 U14965 ( .A1(n18630), .A2(n12263), .ZN(n15767) );
  NOR2_X1 U14966 ( .A1(n15768), .A2(n15767), .ZN(n15766) );
  NOR2_X1 U14967 ( .A1(n15736), .A2(n15735), .ZN(n15734) );
  NOR2_X1 U14968 ( .A1(n18630), .A2(n15734), .ZN(n15726) );
  NOR2_X1 U14969 ( .A1(n15727), .A2(n15726), .ZN(n15725) );
  XNOR2_X1 U14970 ( .A(n12000), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15697) );
  XNOR2_X1 U14971 ( .A(n12001), .B(n15697), .ZN(n12002) );
  NAND4_X1 U14972 ( .A1(n15904), .A2(n19586), .A3(n19263), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19437) );
  NAND2_X1 U14973 ( .A1(n12002), .A2(n18623), .ZN(n12235) );
  AND2_X1 U14974 ( .A1(n12003), .A2(n12630), .ZN(n12629) );
  NOR2_X1 U14975 ( .A1(n12005), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12008) );
  INV_X1 U14976 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19494) );
  AND2_X1 U14977 ( .A1(n12005), .A2(n19535), .ZN(n12006) );
  AOI22_X1 U14978 ( .A1(n12004), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n14826), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12007) );
  OAI21_X1 U14979 ( .B1(n12103), .B2(n19494), .A(n12007), .ZN(n14596) );
  INV_X1 U14980 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n12012) );
  AOI22_X1 U14981 ( .A1(n12163), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n12006), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12011) );
  INV_X1 U14982 ( .A(n13036), .ZN(n12009) );
  OR2_X1 U14983 ( .A1(n12169), .A2(n12009), .ZN(n12010) );
  OAI211_X1 U14984 ( .C1(n12103), .C2(n12012), .A(n12011), .B(n12010), .ZN(
        n12013) );
  INV_X1 U14985 ( .A(n12013), .ZN(n15869) );
  INV_X1 U14986 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n12016) );
  INV_X2 U14987 ( .A(n12187), .ZN(n12163) );
  AOI22_X1 U14988 ( .A1(n12163), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n12006), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12015) );
  OR2_X1 U14989 ( .A1(n12169), .A2(n12947), .ZN(n12014) );
  OAI211_X1 U14990 ( .C1(n12103), .C2(n12016), .A(n12015), .B(n12014), .ZN(
        n12017) );
  INV_X1 U14991 ( .A(n12017), .ZN(n15886) );
  INV_X1 U14992 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15883) );
  INV_X1 U14993 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n18754) );
  INV_X1 U14994 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19470) );
  OAI222_X1 U14995 ( .A1(n15883), .A2(n12186), .B1(n12187), .B2(n18754), .C1(
        n12103), .C2(n19470), .ZN(n12634) );
  INV_X1 U14996 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n12030) );
  AOI22_X1 U14997 ( .A1(n12163), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n14826), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12029) );
  AOI22_X1 U14998 ( .A1(n11629), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12129), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12021) );
  AOI22_X1 U14999 ( .A1(n11618), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12032), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12020) );
  AOI22_X1 U15000 ( .A1(n9604), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12034), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12019) );
  AOI22_X1 U15001 ( .A1(n11574), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12018) );
  NAND4_X1 U15002 ( .A1(n12021), .A2(n12020), .A3(n12019), .A4(n12018), .ZN(
        n12027) );
  AOI22_X1 U15003 ( .A1(n11533), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9639), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12025) );
  AOI22_X1 U15004 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12148), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12024) );
  AOI22_X1 U15005 ( .A1(n12136), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12135), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12023) );
  AOI22_X1 U15006 ( .A1(n12138), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12022) );
  NAND4_X1 U15007 ( .A1(n12025), .A2(n12024), .A3(n12023), .A4(n12022), .ZN(
        n12026) );
  OR2_X1 U15008 ( .A1(n12169), .A2(n13356), .ZN(n12028) );
  OAI211_X1 U15009 ( .C1(n12103), .C2(n12030), .A(n12029), .B(n12028), .ZN(
        n12031) );
  INV_X1 U15010 ( .A(n12031), .ZN(n18633) );
  AOI22_X1 U15011 ( .A1(n11533), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9639), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12038) );
  AOI22_X1 U15012 ( .A1(n9604), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12148), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12037) );
  AOI22_X1 U15013 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12032), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12036) );
  AOI22_X1 U15014 ( .A1(n12034), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11574), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12035) );
  NAND4_X1 U15015 ( .A1(n12038), .A2(n12037), .A3(n12036), .A4(n12035), .ZN(
        n12044) );
  AOI22_X1 U15016 ( .A1(n12138), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12135), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12042) );
  AOI22_X1 U15017 ( .A1(n12136), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12041) );
  AOI22_X1 U15018 ( .A1(n12129), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11618), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12040) );
  AOI22_X1 U15019 ( .A1(n11629), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12039) );
  NAND4_X1 U15020 ( .A1(n12042), .A2(n12041), .A3(n12040), .A4(n12039), .ZN(
        n12043) );
  NOR2_X1 U15021 ( .A1(n12044), .A2(n12043), .ZN(n12468) );
  OR2_X1 U15022 ( .A1(n12468), .A2(n12169), .ZN(n12048) );
  NAND2_X1 U15023 ( .A1(n12045), .A2(n12006), .ZN(n12082) );
  MUX2_X1 U15024 ( .A(n12630), .B(n19571), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12046) );
  AND2_X1 U15025 ( .A1(n12082), .A2(n12046), .ZN(n12047) );
  NAND2_X1 U15026 ( .A1(n12048), .A2(n12047), .ZN(n12564) );
  INV_X1 U15027 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18432) );
  AOI21_X1 U15028 ( .B1(n18926), .B2(P2_EAX_REG_0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12050) );
  NAND2_X1 U15029 ( .A1(n9643), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12049) );
  OAI211_X1 U15030 ( .C1(n12103), .C2(n18432), .A(n12050), .B(n12049), .ZN(
        n12565) );
  INV_X1 U15031 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19462) );
  AOI22_X1 U15032 ( .A1(n12004), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n12006), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12051) );
  OAI21_X1 U15033 ( .B1(n12103), .B2(n19462), .A(n12051), .ZN(n12052) );
  NOR2_X1 U15034 ( .A1(n12563), .A2(n12052), .ZN(n12071) );
  INV_X1 U15035 ( .A(n12052), .ZN(n12053) );
  XNOR2_X1 U15036 ( .A(n12563), .B(n12053), .ZN(n12866) );
  AOI22_X1 U15037 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n11629), .B1(
        n12129), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12058) );
  AOI22_X1 U15038 ( .A1(n11618), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12032), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12057) );
  AOI22_X1 U15039 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n11573), .B1(
        n12034), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12056) );
  AOI22_X1 U15040 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n11574), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12055) );
  NAND4_X1 U15041 ( .A1(n12058), .A2(n12057), .A3(n12056), .A4(n12055), .ZN(
        n12064) );
  AOI22_X1 U15042 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11533), .B1(
        n9639), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12062) );
  AOI22_X1 U15043 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12148), .B1(
        n12033), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12061) );
  AOI22_X1 U15044 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12136), .B1(
        n12135), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12060) );
  AOI22_X1 U15045 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12138), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12059) );
  NAND4_X1 U15046 ( .A1(n12062), .A2(n12061), .A3(n12060), .A4(n12059), .ZN(
        n12063) );
  INV_X1 U15047 ( .A(n13293), .ZN(n12068) );
  NAND2_X1 U15048 ( .A1(n12065), .A2(n12630), .ZN(n12066) );
  MUX2_X1 U15049 ( .A(n12066), .B(n19560), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12067) );
  OAI21_X1 U15050 ( .B1(n12068), .B2(n12169), .A(n12067), .ZN(n12865) );
  INV_X1 U15051 ( .A(n12865), .ZN(n12069) );
  AOI22_X1 U15052 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n11629), .B1(
        n12129), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12075) );
  AOI22_X1 U15053 ( .A1(n11573), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12032), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12074) );
  AOI22_X1 U15054 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n11618), .B1(
        n12034), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12073) );
  AOI22_X1 U15055 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n11574), .B1(
        n12033), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12072) );
  NAND4_X1 U15056 ( .A1(n12075), .A2(n12074), .A3(n12073), .A4(n12072), .ZN(
        n12081) );
  AOI22_X1 U15057 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n11533), .B1(
        n9639), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12079) );
  AOI22_X1 U15058 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n12148), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12078) );
  AOI22_X1 U15059 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n12136), .B1(
        n12135), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12077) );
  AOI22_X1 U15060 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n12138), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12076) );
  NAND4_X1 U15061 ( .A1(n12079), .A2(n12078), .A3(n12077), .A4(n12076), .ZN(
        n12080) );
  NOR2_X1 U15062 ( .A1(n12081), .A2(n12080), .ZN(n13347) );
  NAND2_X1 U15063 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12083) );
  OAI211_X1 U15064 ( .C1(n12169), .C2(n13347), .A(n12083), .B(n12082), .ZN(
        n12084) );
  NOR2_X1 U15065 ( .A1(n12085), .A2(n12084), .ZN(n12087) );
  XNOR2_X1 U15066 ( .A(n12085), .B(n12084), .ZN(n12979) );
  INV_X1 U15067 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19463) );
  INV_X1 U15068 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18878) );
  AOI22_X1 U15069 ( .A1(n12163), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n12006), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12086) );
  OAI21_X1 U15070 ( .B1(n12103), .B2(n19463), .A(n12086), .ZN(n12978) );
  NOR2_X1 U15071 ( .A1(n12979), .A2(n12978), .ZN(n12980) );
  INV_X1 U15072 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n12102) );
  AOI22_X1 U15073 ( .A1(n14826), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12089) );
  NAND2_X1 U15074 ( .A1(n12163), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n12088) );
  AND2_X1 U15075 ( .A1(n12089), .A2(n12088), .ZN(n12101) );
  AOI22_X1 U15076 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n11629), .B1(
        n12129), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12093) );
  AOI22_X1 U15077 ( .A1(n11618), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12032), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12092) );
  AOI22_X1 U15078 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n9604), .B1(
        n12034), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12091) );
  AOI22_X1 U15079 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n11574), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12090) );
  NAND4_X1 U15080 ( .A1(n12093), .A2(n12092), .A3(n12091), .A4(n12090), .ZN(
        n12099) );
  AOI22_X1 U15081 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n11533), .B1(
        n9639), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12097) );
  AOI22_X1 U15082 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n12148), .B1(
        n12033), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12096) );
  AOI22_X1 U15083 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12136), .B1(
        n12135), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12095) );
  AOI22_X1 U15084 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n12138), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12094) );
  NAND4_X1 U15085 ( .A1(n12097), .A2(n12096), .A3(n12095), .A4(n12094), .ZN(
        n12098) );
  INV_X1 U15086 ( .A(n12221), .ZN(n13267) );
  OR2_X1 U15087 ( .A1(n12169), .A2(n13267), .ZN(n12100) );
  OAI211_X1 U15088 ( .C1(n12103), .C2(n12102), .A(n12101), .B(n12100), .ZN(
        n13017) );
  INV_X1 U15089 ( .A(n12103), .ZN(n12198) );
  AOI22_X1 U15090 ( .A1(n12198), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n12006), 
        .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12115) );
  INV_X1 U15091 ( .A(n12169), .ZN(n12174) );
  AOI22_X1 U15092 ( .A1(n11629), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12129), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12107) );
  AOI22_X1 U15093 ( .A1(n11618), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12032), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12106) );
  AOI22_X1 U15094 ( .A1(n9604), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12034), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12105) );
  AOI22_X1 U15095 ( .A1(n11574), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12104) );
  NAND4_X1 U15096 ( .A1(n12107), .A2(n12106), .A3(n12105), .A4(n12104), .ZN(
        n12113) );
  AOI22_X1 U15097 ( .A1(n11533), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9639), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12111) );
  AOI22_X1 U15098 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12148), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12110) );
  AOI22_X1 U15099 ( .A1(n12136), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12135), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12109) );
  AOI22_X1 U15100 ( .A1(n12138), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12108) );
  NAND4_X1 U15101 ( .A1(n12111), .A2(n12110), .A3(n12109), .A4(n12108), .ZN(
        n12112) );
  AOI22_X1 U15102 ( .A1(n12174), .A2(n13323), .B1(n12163), .B2(
        P2_EAX_REG_5__SCAN_IN), .ZN(n12114) );
  NAND2_X1 U15103 ( .A1(n12115), .A2(n12114), .ZN(n13370) );
  AOI22_X1 U15104 ( .A1(n11629), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12129), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12119) );
  AOI22_X1 U15105 ( .A1(n9604), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12032), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12118) );
  AOI22_X1 U15106 ( .A1(n11618), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12034), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12117) );
  AOI22_X1 U15107 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12116) );
  NAND4_X1 U15108 ( .A1(n12119), .A2(n12118), .A3(n12117), .A4(n12116), .ZN(
        n12125) );
  AOI22_X1 U15109 ( .A1(n11533), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9639), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12123) );
  AOI22_X1 U15110 ( .A1(n12148), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11574), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12122) );
  AOI22_X1 U15111 ( .A1(n12136), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12135), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12121) );
  AOI22_X1 U15112 ( .A1(n12138), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12120) );
  NAND4_X1 U15113 ( .A1(n12123), .A2(n12122), .A3(n12121), .A4(n12120), .ZN(
        n12124) );
  OR2_X1 U15114 ( .A1(n12169), .A2(n13467), .ZN(n12126) );
  INV_X1 U15115 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19468) );
  AOI22_X1 U15116 ( .A1(n12163), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n12006), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12127) );
  OAI21_X1 U15117 ( .B1(n12103), .B2(n19468), .A(n12127), .ZN(n12128) );
  INV_X1 U15118 ( .A(n12128), .ZN(n12624) );
  NAND2_X1 U15119 ( .A1(n11629), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n12134) );
  NAND2_X1 U15120 ( .A1(n12129), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n12133) );
  NAND2_X1 U15121 ( .A1(n12032), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n12132) );
  NAND2_X1 U15122 ( .A1(n9604), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n12131) );
  AOI22_X1 U15123 ( .A1(n12136), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12135), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12142) );
  AOI22_X1 U15124 ( .A1(n12138), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12141) );
  NAND2_X1 U15125 ( .A1(n11533), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12140) );
  NAND2_X1 U15126 ( .A1(n9639), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n12139) );
  NAND2_X1 U15127 ( .A1(n11618), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12146) );
  NAND2_X1 U15128 ( .A1(n12034), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12145) );
  NAND2_X1 U15129 ( .A1(n11574), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12144) );
  NAND2_X1 U15130 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12143) );
  AOI22_X1 U15131 ( .A1(n12148), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12149) );
  OAI22_X2 U15132 ( .A1(n12625), .A2(n12624), .B1(n13327), .B2(n12169), .ZN(
        n12635) );
  INV_X1 U15133 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n12156) );
  AOI22_X1 U15134 ( .A1(n12163), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n12006), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12155) );
  INV_X1 U15135 ( .A(n12907), .ZN(n12153) );
  OR2_X1 U15136 ( .A1(n12169), .A2(n12153), .ZN(n12154) );
  OAI211_X1 U15137 ( .C1(n12103), .C2(n12156), .A(n12155), .B(n12154), .ZN(
        n12738) );
  INV_X1 U15138 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n12159) );
  AOI22_X1 U15139 ( .A1(n12163), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n12006), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12158) );
  OR2_X1 U15140 ( .A1(n12169), .A2(n12965), .ZN(n12157) );
  OAI211_X1 U15141 ( .C1(n12103), .C2(n12159), .A(n12158), .B(n12157), .ZN(
        n12160) );
  INV_X1 U15142 ( .A(n12160), .ZN(n12747) );
  INV_X1 U15143 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n12161) );
  OAI22_X1 U15144 ( .A1(n12161), .A2(n12103), .B1(n12169), .B2(n13031), .ZN(
        n12162) );
  INV_X1 U15145 ( .A(n12162), .ZN(n12165) );
  AOI22_X1 U15146 ( .A1(n12163), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n12006), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12164) );
  NAND2_X1 U15147 ( .A1(n12165), .A2(n12164), .ZN(n12910) );
  NAND2_X2 U15148 ( .A1(n12911), .A2(n12910), .ZN(n15870) );
  NOR2_X4 U15149 ( .A1(n15869), .A2(n15870), .ZN(n15868) );
  INV_X1 U15150 ( .A(n13053), .ZN(n12168) );
  NAND2_X1 U15151 ( .A1(n12198), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n12167) );
  AOI22_X1 U15152 ( .A1(n12004), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n12006), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12166) );
  OAI211_X1 U15153 ( .C1(n12168), .C2(n12169), .A(n12167), .B(n12166), .ZN(
        n13004) );
  NAND2_X2 U15154 ( .A1(n15868), .A2(n13004), .ZN(n15855) );
  INV_X1 U15155 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n12172) );
  AOI22_X1 U15156 ( .A1(n12163), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n14826), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12171) );
  OR2_X1 U15157 ( .A1(n12169), .A2(n13118), .ZN(n12170) );
  OAI211_X1 U15158 ( .C1(n12103), .C2(n12172), .A(n12171), .B(n12170), .ZN(
        n12173) );
  INV_X1 U15159 ( .A(n12173), .ZN(n15856) );
  AOI22_X1 U15160 ( .A1(n12198), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n14826), .ZN(n12176) );
  AOI22_X1 U15161 ( .A1(n12174), .A2(n10283), .B1(P2_EAX_REG_15__SCAN_IN), 
        .B2(n12163), .ZN(n12175) );
  NAND2_X1 U15162 ( .A1(n12176), .A2(n12175), .ZN(n13048) );
  INV_X1 U15163 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n12178) );
  AOI22_X1 U15164 ( .A1(n12163), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n14826), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12177) );
  OAI21_X1 U15165 ( .B1(n12103), .B2(n12178), .A(n12177), .ZN(n12179) );
  INV_X1 U15166 ( .A(n12179), .ZN(n13198) );
  INV_X1 U15167 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19483) );
  AOI22_X1 U15168 ( .A1(n12004), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n14826), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12180) );
  OAI21_X1 U15169 ( .B1(n12103), .B2(n19483), .A(n12180), .ZN(n13391) );
  INV_X1 U15170 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19485) );
  AOI22_X1 U15171 ( .A1(n12004), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n14826), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12181) );
  OAI21_X1 U15172 ( .B1(n12103), .B2(n19485), .A(n12181), .ZN(n12182) );
  INV_X1 U15173 ( .A(n12182), .ZN(n13424) );
  OR2_X2 U15174 ( .A1(n9650), .A2(n13424), .ZN(n13423) );
  INV_X1 U15175 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19487) );
  AOI22_X1 U15176 ( .A1(n12004), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n14826), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12183) );
  OAI21_X1 U15177 ( .B1(n12103), .B2(n19487), .A(n12183), .ZN(n14631) );
  INV_X1 U15178 ( .A(n14631), .ZN(n12184) );
  INV_X1 U15179 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n14754) );
  AOI22_X1 U15180 ( .A1(n12004), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n14826), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12185) );
  OAI21_X1 U15181 ( .B1(n12103), .B2(n14754), .A(n12185), .ZN(n14619) );
  INV_X1 U15182 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19490) );
  INV_X1 U15183 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n18725) );
  INV_X1 U15184 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n13877) );
  OAI222_X1 U15185 ( .A1(n12103), .A2(n19490), .B1(n12187), .B2(n18725), .C1(
        n13877), .C2(n12186), .ZN(n12258) );
  NAND2_X1 U15186 ( .A1(n12198), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n12189) );
  AOI22_X1 U15187 ( .A1(n12004), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n14826), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12188) );
  INV_X1 U15188 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19496) );
  AOI22_X1 U15189 ( .A1(n12004), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n14826), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12190) );
  OAI21_X1 U15190 ( .B1(n12103), .B2(n19496), .A(n12190), .ZN(n14894) );
  NAND2_X1 U15191 ( .A1(n12198), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n12192) );
  AOI22_X1 U15192 ( .A1(n12004), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n14826), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12191) );
  AND2_X1 U15193 ( .A1(n12192), .A2(n12191), .ZN(n14586) );
  NAND2_X1 U15194 ( .A1(n12198), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n12194) );
  AOI22_X1 U15195 ( .A1(n12163), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n14826), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12193) );
  AND2_X1 U15196 ( .A1(n12194), .A2(n12193), .ZN(n14579) );
  NOR2_X2 U15197 ( .A1(n9649), .A2(n14579), .ZN(n14581) );
  INV_X1 U15198 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19503) );
  AOI22_X1 U15199 ( .A1(n12163), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n14826), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12195) );
  OAI21_X1 U15200 ( .B1(n12103), .B2(n19503), .A(n12195), .ZN(n14573) );
  NAND2_X1 U15201 ( .A1(n12198), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12197) );
  AOI22_X1 U15202 ( .A1(n12163), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n14826), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12196) );
  AND2_X1 U15203 ( .A1(n12197), .A2(n12196), .ZN(n14565) );
  NAND2_X1 U15204 ( .A1(n12198), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n12200) );
  AOI22_X1 U15205 ( .A1(n12163), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n14826), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12199) );
  AND2_X1 U15206 ( .A1(n12200), .A2(n12199), .ZN(n14558) );
  INV_X1 U15207 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n13872) );
  AOI22_X1 U15208 ( .A1(n12163), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n14826), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12201) );
  OAI21_X1 U15209 ( .B1(n12103), .B2(n13872), .A(n12201), .ZN(n12202) );
  NAND2_X1 U15210 ( .A1(n9713), .A2(n10176), .ZN(n12203) );
  NAND2_X1 U15211 ( .A1(n12204), .A2(n12440), .ZN(n12446) );
  INV_X1 U15212 ( .A(n12446), .ZN(n12205) );
  AND2_X1 U15213 ( .A1(n12206), .A2(n12205), .ZN(n12207) );
  OR2_X1 U15214 ( .A1(n12442), .A2(n12207), .ZN(n12833) );
  INV_X1 U15215 ( .A(n12832), .ZN(n12208) );
  INV_X1 U15216 ( .A(n18414), .ZN(n19590) );
  NOR2_X1 U15217 ( .A1(n9634), .A2(n9643), .ZN(n12538) );
  NAND2_X1 U15218 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19593) );
  INV_X1 U15219 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n18411) );
  NOR2_X1 U15220 ( .A1(n20627), .A2(n18411), .ZN(n19453) );
  NOR2_X1 U15221 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n19454) );
  NOR3_X1 U15222 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19453), .A3(n19454), 
        .ZN(n19582) );
  NAND2_X1 U15223 ( .A1(n19593), .A2(n19582), .ZN(n12840) );
  NOR2_X1 U15224 ( .A1(n12840), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n12210) );
  NAND2_X1 U15225 ( .A1(n12538), .A2(n12210), .ZN(n12856) );
  NOR2_X2 U15226 ( .A1(n19590), .A2(n12856), .ZN(n18647) );
  OR2_X1 U15227 ( .A1(n12833), .A2(n18416), .ZN(n12394) );
  INV_X1 U15228 ( .A(n19593), .ZN(n19587) );
  NOR2_X1 U15229 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19587), .ZN(n12211) );
  OR2_X1 U15230 ( .A1(n18702), .A2(n12210), .ZN(n15690) );
  NOR2_X1 U15231 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n12211), .ZN(n12212) );
  NAND2_X1 U15232 ( .A1(n12397), .A2(n12212), .ZN(n12213) );
  MUX2_X1 U15233 ( .A(n12214), .B(n13356), .S(n12455), .Z(n12215) );
  MUX2_X1 U15234 ( .A(n12215), .B(P2_EBX_REG_4__SCAN_IN), .S(n18911), .Z(
        n13342) );
  MUX2_X1 U15235 ( .A(n12438), .B(P2_EBX_REG_2__SCAN_IN), .S(n18911), .Z(
        n13074) );
  INV_X1 U15236 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n12665) );
  AND2_X1 U15237 ( .A1(n18911), .A2(n12665), .ZN(n12457) );
  NAND2_X1 U15238 ( .A1(n12457), .A2(n11412), .ZN(n12218) );
  NAND2_X1 U15239 ( .A1(n9614), .A2(n13293), .ZN(n12217) );
  INV_X1 U15240 ( .A(n12219), .ZN(n12220) );
  MUX2_X1 U15241 ( .A(n12221), .B(n12220), .S(n11382), .Z(n12223) );
  MUX2_X1 U15242 ( .A(n12223), .B(n12222), .S(n18911), .Z(n13015) );
  NOR2_X2 U15243 ( .A1(n13342), .A2(n13340), .ZN(n13329) );
  MUX2_X1 U15244 ( .A(n13323), .B(n12732), .S(n18911), .Z(n13328) );
  MUX2_X1 U15245 ( .A(n13467), .B(P2_EBX_REG_6__SCAN_IN), .S(n18911), .Z(
        n13473) );
  MUX2_X1 U15246 ( .A(n12224), .B(n12773), .S(n18911), .Z(n13748) );
  NAND2_X1 U15247 ( .A1(n18911), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13745) );
  NOR2_X2 U15248 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n13765), .ZN(n13771) );
  NAND2_X1 U15249 ( .A1(n18911), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13770) );
  NAND2_X1 U15250 ( .A1(n18911), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n13796) );
  NAND2_X1 U15251 ( .A1(n18911), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n13788) );
  NAND2_X1 U15252 ( .A1(n18911), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n13783) );
  AND2_X1 U15253 ( .A1(n18911), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n13785) );
  AND2_X1 U15254 ( .A1(n18911), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n13800) );
  NAND2_X1 U15255 ( .A1(n18911), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n13779) );
  NAND2_X2 U15256 ( .A1(n12265), .A2(n13834), .ZN(n12255) );
  NAND2_X1 U15257 ( .A1(n18911), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12266) );
  NAND2_X2 U15258 ( .A1(n13834), .A2(n9682), .ZN(n14644) );
  NAND2_X1 U15259 ( .A1(n18911), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n13738) );
  AND2_X1 U15260 ( .A1(n18911), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n13840) );
  AND2_X1 U15261 ( .A1(n18911), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n13851) );
  AND2_X1 U15262 ( .A1(n18911), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12227) );
  OAI21_X1 U15263 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n19587), .A(
        P2_EBX_REG_31__SCAN_IN), .ZN(n12228) );
  INV_X1 U15264 ( .A(n12228), .ZN(n12229) );
  NAND2_X1 U15265 ( .A1(n13706), .A2(n19535), .ZN(n19537) );
  NOR2_X1 U15266 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19537), .ZN(n12396) );
  INV_X2 U15267 ( .A(n18496), .ZN(n18850) );
  NOR2_X1 U15268 ( .A1(n19535), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19101) );
  INV_X1 U15269 ( .A(n19101), .ZN(n19433) );
  NOR2_X1 U15270 ( .A1(n19440), .A2(n19433), .ZN(n15907) );
  AOI22_X1 U15271 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n18639), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n9772), .ZN(n12230) );
  OAI21_X1 U15272 ( .B1(n13853), .B2(n18616), .A(n12230), .ZN(n12231) );
  AOI21_X1 U15273 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n18614), .A(n12231), .ZN(
        n12232) );
  OAI21_X1 U15274 ( .B1(n14656), .B2(n18643), .A(n12232), .ZN(n12233) );
  NAND2_X1 U15275 ( .A1(n12235), .A2(n12234), .ZN(P2_U2825) );
  NOR2_X1 U15276 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12237) );
  NOR4_X1 U15277 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12236) );
  NAND4_X1 U15278 ( .A1(P2_W_R_N_REG_SCAN_IN), .A2(P2_M_IO_N_REG_SCAN_IN), 
        .A3(n12237), .A4(n12236), .ZN(n12249) );
  INV_X1 U15279 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20539) );
  NOR3_X1 U15280 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20539), .ZN(n12239) );
  NOR4_X1 U15281 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n12238) );
  NAND4_X1 U15282 ( .A1(n19836), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n12239), .A4(
        n12238), .ZN(U214) );
  NOR4_X1 U15283 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_14__SCAN_IN), .A3(P2_ADDRESS_REG_13__SCAN_IN), .A4(
        P2_ADDRESS_REG_12__SCAN_IN), .ZN(n12243) );
  NOR4_X1 U15284 ( .A1(P2_ADDRESS_REG_19__SCAN_IN), .A2(
        P2_ADDRESS_REG_18__SCAN_IN), .A3(P2_ADDRESS_REG_17__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n12242) );
  NOR4_X1 U15285 ( .A1(P2_ADDRESS_REG_7__SCAN_IN), .A2(
        P2_ADDRESS_REG_6__SCAN_IN), .A3(P2_ADDRESS_REG_5__SCAN_IN), .A4(
        P2_ADDRESS_REG_4__SCAN_IN), .ZN(n12241) );
  NOR4_X1 U15286 ( .A1(P2_ADDRESS_REG_11__SCAN_IN), .A2(
        P2_ADDRESS_REG_10__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n12240) );
  NAND4_X1 U15287 ( .A1(n12243), .A2(n12242), .A3(n12241), .A4(n12240), .ZN(
        n12248) );
  NOR4_X1 U15288 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_3__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n12246) );
  NOR4_X1 U15289 ( .A1(P2_ADDRESS_REG_23__SCAN_IN), .A2(
        P2_ADDRESS_REG_22__SCAN_IN), .A3(P2_ADDRESS_REG_21__SCAN_IN), .A4(
        P2_ADDRESS_REG_20__SCAN_IN), .ZN(n12245) );
  NOR4_X1 U15290 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_26__SCAN_IN), .A3(P2_ADDRESS_REG_25__SCAN_IN), .A4(
        P2_ADDRESS_REG_24__SCAN_IN), .ZN(n12244) );
  INV_X1 U15291 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19465) );
  NAND4_X1 U15292 ( .A1(n12246), .A2(n12245), .A3(n12244), .A4(n19465), .ZN(
        n12247) );
  NOR2_X1 U15293 ( .A1(n14633), .A2(n12249), .ZN(n15991) );
  NAND2_X1 U15294 ( .A1(n15991), .A2(U214), .ZN(U212) );
  AOI211_X1 U15295 ( .C1(n14746), .C2(n12251), .A(n12250), .B(n19437), .ZN(
        n12262) );
  NAND2_X1 U15296 ( .A1(n18911), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12252) );
  NOR2_X1 U15297 ( .A1(n12253), .A2(n12252), .ZN(n12254) );
  OR2_X1 U15298 ( .A1(n12255), .A2(n12254), .ZN(n13806) );
  OAI22_X1 U15299 ( .A1(n14742), .A2(n18540), .B1(n13806), .B2(n18616), .ZN(
        n12261) );
  INV_X1 U15300 ( .A(n18614), .ZN(n18642) );
  OAI22_X1 U15301 ( .A1(n18642), .A2(n12226), .B1(n19490), .B2(n18601), .ZN(
        n12260) );
  NOR2_X1 U15302 ( .A1(n14529), .A2(n12256), .ZN(n12257) );
  OR2_X1 U15303 ( .A1(n12271), .A2(n12257), .ZN(n14743) );
  OAI21_X1 U15304 ( .B1(n14621), .B2(n12258), .A(n12268), .ZN(n14936) );
  INV_X1 U15305 ( .A(n18647), .ZN(n18628) );
  OAI22_X1 U15306 ( .A1(n14743), .A2(n18643), .B1(n14936), .B2(n18628), .ZN(
        n12259) );
  OR4_X1 U15307 ( .A1(n12262), .A2(n12261), .A3(n12260), .A4(n12259), .ZN(
        P2_U2834) );
  AOI211_X1 U15308 ( .C1(n15784), .C2(n12264), .A(n12263), .B(n19437), .ZN(
        n12275) );
  INV_X1 U15309 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n19492) );
  INV_X1 U15310 ( .A(n12265), .ZN(n12267) );
  OAI21_X1 U15311 ( .B1(n12267), .B2(n12266), .A(n13824), .ZN(n13822) );
  OAI22_X1 U15312 ( .A1(n19492), .A2(n18601), .B1(n13822), .B2(n18616), .ZN(
        n12274) );
  OAI22_X1 U15313 ( .A1(n18642), .A2(n11928), .B1(n10113), .B2(n18540), .ZN(
        n12273) );
  XNOR2_X1 U15314 ( .A(n12269), .B(n12268), .ZN(n14920) );
  OAI21_X1 U15315 ( .B1(n12271), .B2(n12270), .A(n9659), .ZN(n14927) );
  OAI22_X1 U15316 ( .A1(n18628), .A2(n14920), .B1(n18643), .B2(n14927), .ZN(
        n12272) );
  OR4_X1 U15317 ( .A1(n12275), .A2(n12274), .A3(n12273), .A4(n12272), .ZN(
        P2_U2833) );
  AOI21_X1 U15318 ( .B1(n12278), .B2(n13930), .A(n12277), .ZN(n14118) );
  AND2_X1 U15319 ( .A1(n12478), .A2(n12485), .ZN(n12483) );
  INV_X1 U15320 ( .A(n12424), .ZN(n12279) );
  NAND2_X1 U15321 ( .A1(n12414), .A2(n12696), .ZN(n12412) );
  NAND2_X1 U15322 ( .A1(n20448), .A2(n20445), .ZN(n15684) );
  INV_X1 U15323 ( .A(n15684), .ZN(n20542) );
  NAND2_X1 U15324 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20542), .ZN(n15397) );
  NOR2_X1 U15325 ( .A1(n15397), .A2(n20446), .ZN(n12283) );
  NAND2_X1 U15326 ( .A1(n20547), .A2(n12280), .ZN(n12281) );
  NAND2_X1 U15327 ( .A1(n19798), .A2(n12281), .ZN(n12282) );
  INV_X1 U15328 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14095) );
  XNOR2_X1 U15329 ( .A(n12285), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14087) );
  NOR2_X1 U15330 ( .A1(n14087), .A2(n20445), .ZN(n12286) );
  NOR2_X1 U15331 ( .A1(n14036), .A2(n15470), .ZN(n12393) );
  AND2_X4 U15332 ( .A1(n19839), .A2(n19853), .ZN(n13715) );
  NAND2_X2 U15333 ( .A1(n9692), .A2(n13715), .ZN(n13718) );
  OR2_X1 U15334 ( .A1(n13718), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n12291) );
  INV_X1 U15335 ( .A(n19863), .ZN(n12287) );
  INV_X1 U15336 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19819) );
  NAND2_X1 U15337 ( .A1(n12302), .A2(n19819), .ZN(n12289) );
  INV_X1 U15338 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n12654) );
  NAND2_X1 U15339 ( .A1(n13715), .A2(n12654), .ZN(n12288) );
  NAND3_X1 U15340 ( .A1(n12289), .A2(n12352), .A3(n12288), .ZN(n12290) );
  NAND2_X1 U15341 ( .A1(n12291), .A2(n12290), .ZN(n12295) );
  NAND2_X1 U15342 ( .A1(n12302), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12294) );
  INV_X1 U15343 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n12292) );
  NAND2_X1 U15344 ( .A1(n12352), .A2(n12292), .ZN(n12293) );
  NAND2_X1 U15345 ( .A1(n12294), .A2(n12293), .ZN(n12718) );
  XNOR2_X1 U15346 ( .A(n12295), .B(n12718), .ZN(n13087) );
  NAND2_X1 U15347 ( .A1(n13087), .A2(n13715), .ZN(n12296) );
  OR2_X1 U15348 ( .A1(n13718), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n12300) );
  NAND2_X1 U15349 ( .A1(n12302), .A2(n19831), .ZN(n12298) );
  INV_X1 U15350 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n12896) );
  NAND2_X1 U15351 ( .A1(n13715), .A2(n12896), .ZN(n12297) );
  NAND3_X1 U15352 ( .A1(n12298), .A2(n12372), .A3(n12297), .ZN(n12299) );
  AND2_X1 U15353 ( .A1(n12300), .A2(n12299), .ZN(n12893) );
  MUX2_X1 U15354 ( .A(n12365), .B(n12372), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n12301) );
  OAI21_X1 U15355 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n13887), .A(
        n12301), .ZN(n12992) );
  MUX2_X1 U15356 ( .A(n13718), .B(n12302), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n12306) );
  INV_X1 U15357 ( .A(n12302), .ZN(n12303) );
  NAND2_X1 U15358 ( .A1(n12303), .A2(n13886), .ZN(n12360) );
  NAND2_X1 U15359 ( .A1(n13886), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12304) );
  AND2_X1 U15360 ( .A1(n12360), .A2(n12304), .ZN(n12305) );
  NAND2_X1 U15361 ( .A1(n12306), .A2(n12305), .ZN(n12974) );
  MUX2_X1 U15362 ( .A(n12365), .B(n12372), .S(P1_EBX_REG_5__SCAN_IN), .Z(
        n12307) );
  OAI21_X1 U15363 ( .B1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n13887), .A(
        n12307), .ZN(n13010) );
  OR2_X1 U15364 ( .A1(n13718), .A2(P1_EBX_REG_6__SCAN_IN), .ZN(n12312) );
  INV_X1 U15365 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12308) );
  NAND2_X1 U15366 ( .A1(n12302), .A2(n12308), .ZN(n12310) );
  INV_X1 U15367 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n19709) );
  NAND2_X1 U15368 ( .A1(n13715), .A2(n19709), .ZN(n12309) );
  NAND3_X1 U15369 ( .A1(n12310), .A2(n12372), .A3(n12309), .ZN(n12311) );
  INV_X1 U15370 ( .A(n12365), .ZN(n12371) );
  INV_X1 U15371 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n19640) );
  NAND2_X1 U15372 ( .A1(n12371), .A2(n19640), .ZN(n12315) );
  NAND2_X1 U15373 ( .A1(n12372), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12313) );
  OAI211_X1 U15374 ( .C1(n13886), .C2(P1_EBX_REG_7__SCAN_IN), .A(n12302), .B(
        n12313), .ZN(n12314) );
  OR2_X1 U15375 ( .A1(n13718), .A2(P1_EBX_REG_8__SCAN_IN), .ZN(n12319) );
  INV_X1 U15376 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n13212) );
  NAND2_X1 U15377 ( .A1(n12302), .A2(n13212), .ZN(n12317) );
  INV_X1 U15378 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13154) );
  NAND2_X1 U15379 ( .A1(n13715), .A2(n13154), .ZN(n12316) );
  NAND3_X1 U15380 ( .A1(n12317), .A2(n12372), .A3(n12316), .ZN(n12318) );
  NAND2_X1 U15381 ( .A1(n12319), .A2(n12318), .ZN(n13148) );
  MUX2_X1 U15382 ( .A(n12365), .B(n12372), .S(P1_EBX_REG_9__SCAN_IN), .Z(
        n12320) );
  OAI21_X1 U15383 ( .B1(n13887), .B2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n12320), .ZN(n13182) );
  OR2_X1 U15384 ( .A1(n13718), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n12324) );
  NAND2_X1 U15385 ( .A1(n12302), .A2(n15629), .ZN(n12322) );
  INV_X1 U15386 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n13401) );
  NAND2_X1 U15387 ( .A1(n13715), .A2(n13401), .ZN(n12321) );
  NAND3_X1 U15388 ( .A1(n12322), .A2(n12372), .A3(n12321), .ZN(n12323) );
  NAND2_X1 U15389 ( .A1(n12324), .A2(n12323), .ZN(n13399) );
  INV_X1 U15390 ( .A(n9692), .ZN(n12372) );
  NAND2_X1 U15391 ( .A1(n12372), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12325) );
  OAI211_X1 U15392 ( .C1(n13886), .C2(P1_EBX_REG_11__SCAN_IN), .A(n12302), .B(
        n12325), .ZN(n12326) );
  OAI21_X1 U15393 ( .B1(n12365), .B2(P1_EBX_REG_11__SCAN_IN), .A(n12326), .ZN(
        n15523) );
  MUX2_X1 U15394 ( .A(n13718), .B(n12302), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n12328) );
  NAND2_X1 U15395 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n13886), .ZN(
        n12327) );
  MUX2_X1 U15396 ( .A(n12365), .B(n12372), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n12329) );
  OAI21_X1 U15397 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n13887), .A(
        n12329), .ZN(n13511) );
  OR3_X2 U15398 ( .A1(n15520), .A2(n13524), .A3(n13511), .ZN(n13534) );
  OR2_X1 U15399 ( .A1(n13718), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n12334) );
  NAND2_X1 U15400 ( .A1(n12302), .A2(n12330), .ZN(n12332) );
  INV_X1 U15401 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n13543) );
  NAND2_X1 U15402 ( .A1(n13715), .A2(n13543), .ZN(n12331) );
  NAND3_X1 U15403 ( .A1(n12332), .A2(n12372), .A3(n12331), .ZN(n12333) );
  INV_X1 U15404 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n15539) );
  NAND2_X1 U15405 ( .A1(n12371), .A2(n15539), .ZN(n12337) );
  NAND2_X1 U15406 ( .A1(n12372), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12335) );
  OAI211_X1 U15407 ( .C1(n13886), .C2(P1_EBX_REG_15__SCAN_IN), .A(n12302), .B(
        n12335), .ZN(n12336) );
  MUX2_X1 U15408 ( .A(n13718), .B(n12302), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n12339) );
  NAND2_X1 U15409 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n13886), .ZN(
        n12338) );
  NAND2_X1 U15410 ( .A1(n12372), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12340) );
  OAI211_X1 U15411 ( .C1(n13886), .C2(P1_EBX_REG_17__SCAN_IN), .A(n12302), .B(
        n12340), .ZN(n12341) );
  OAI21_X1 U15412 ( .B1(n12365), .B2(P1_EBX_REG_17__SCAN_IN), .A(n12341), .ZN(
        n13964) );
  MUX2_X1 U15413 ( .A(n13718), .B(n12302), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n12344) );
  NAND2_X1 U15414 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n13886), .ZN(
        n12342) );
  AND2_X1 U15415 ( .A1(n12360), .A2(n12342), .ZN(n12343) );
  AND2_X1 U15416 ( .A1(n12344), .A2(n12343), .ZN(n14006) );
  MUX2_X1 U15417 ( .A(n12365), .B(n12372), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n12345) );
  OAI21_X1 U15418 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n13887), .A(
        n12345), .ZN(n14007) );
  NOR2_X1 U15419 ( .A1(n14006), .A2(n14007), .ZN(n12346) );
  OR2_X1 U15420 ( .A1(n13718), .A2(P1_EBX_REG_20__SCAN_IN), .ZN(n12351) );
  INV_X1 U15421 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14347) );
  NAND2_X1 U15422 ( .A1(n12302), .A2(n14347), .ZN(n12349) );
  INV_X1 U15423 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n12347) );
  NAND2_X1 U15424 ( .A1(n13715), .A2(n12347), .ZN(n12348) );
  NAND3_X1 U15425 ( .A1(n12349), .A2(n12372), .A3(n12348), .ZN(n12350) );
  NAND2_X1 U15426 ( .A1(n12351), .A2(n12350), .ZN(n14002) );
  NAND2_X1 U15427 ( .A1(n12352), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12353) );
  OAI211_X1 U15428 ( .C1(n13886), .C2(P1_EBX_REG_21__SCAN_IN), .A(n12302), .B(
        n12353), .ZN(n12354) );
  OAI21_X1 U15429 ( .B1(n12365), .B2(P1_EBX_REG_21__SCAN_IN), .A(n12354), .ZN(
        n14335) );
  MUX2_X1 U15430 ( .A(n13718), .B(n12302), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n12356) );
  NAND2_X1 U15431 ( .A1(n13886), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12355) );
  AND3_X1 U15432 ( .A1(n12356), .A2(n12360), .A3(n12355), .ZN(n13992) );
  NAND2_X1 U15433 ( .A1(n12352), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12357) );
  OAI211_X1 U15434 ( .C1(n13886), .C2(P1_EBX_REG_23__SCAN_IN), .A(n12302), .B(
        n12357), .ZN(n12358) );
  OAI21_X1 U15435 ( .B1(n12365), .B2(P1_EBX_REG_23__SCAN_IN), .A(n12358), .ZN(
        n13944) );
  MUX2_X1 U15436 ( .A(n13718), .B(n12302), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n12362) );
  NAND2_X1 U15437 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n13886), .ZN(
        n12359) );
  AND2_X1 U15438 ( .A1(n12360), .A2(n12359), .ZN(n12361) );
  NAND2_X1 U15439 ( .A1(n12362), .A2(n12361), .ZN(n13987) );
  NAND2_X1 U15440 ( .A1(n12372), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12363) );
  OAI211_X1 U15441 ( .C1(n13886), .C2(P1_EBX_REG_25__SCAN_IN), .A(n12302), .B(
        n12363), .ZN(n12364) );
  OAI21_X1 U15442 ( .B1(n12365), .B2(P1_EBX_REG_25__SCAN_IN), .A(n12364), .ZN(
        n13980) );
  OR2_X1 U15443 ( .A1(n13718), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n12370) );
  INV_X1 U15444 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14244) );
  NAND2_X1 U15445 ( .A1(n12302), .A2(n14244), .ZN(n12368) );
  INV_X1 U15446 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n12366) );
  NAND2_X1 U15447 ( .A1(n13715), .A2(n12366), .ZN(n12367) );
  NAND3_X1 U15448 ( .A1(n12368), .A2(n12372), .A3(n12367), .ZN(n12369) );
  INV_X1 U15449 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n13975) );
  NAND2_X1 U15450 ( .A1(n12371), .A2(n13975), .ZN(n12375) );
  NAND2_X1 U15451 ( .A1(n12372), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12373) );
  OAI211_X1 U15452 ( .C1(n13886), .C2(P1_EBX_REG_27__SCAN_IN), .A(n12302), .B(
        n12373), .ZN(n12374) );
  AND2_X1 U15453 ( .A1(n12375), .A2(n12374), .ZN(n12376) );
  NOR2_X1 U15454 ( .A1(n13932), .A2(n12376), .ZN(n12377) );
  OR2_X1 U15455 ( .A1(n13923), .A2(n12377), .ZN(n14282) );
  NAND2_X1 U15456 ( .A1(n13715), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n12381) );
  AND2_X1 U15457 ( .A1(n20546), .A2(n20347), .ZN(n15391) );
  NOR2_X1 U15458 ( .A1(n12381), .A2(n15391), .ZN(n12378) );
  NOR2_X1 U15459 ( .A1(n14282), .A2(n19681), .ZN(n12392) );
  NAND2_X1 U15460 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n12385) );
  INV_X1 U15461 ( .A(n13961), .ZN(n15449) );
  INV_X1 U15462 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20488) );
  INV_X1 U15463 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n13410) );
  INV_X1 U15464 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n19629) );
  NAND4_X1 U15465 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_4__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n13153)
         );
  NAND4_X1 U15466 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .A3(P1_REIP_REG_6__SCAN_IN), .A4(P1_REIP_REG_5__SCAN_IN), .ZN(n19625)
         );
  NOR4_X1 U15467 ( .A1(n13410), .A2(n19629), .A3(n13153), .A4(n19625), .ZN(
        n13406) );
  INV_X1 U15468 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n15610) );
  NAND2_X1 U15469 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n13509) );
  NOR2_X1 U15470 ( .A1(n15610), .A2(n13509), .ZN(n13958) );
  NAND3_X1 U15471 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n13406), .A3(n13958), 
        .ZN(n13531) );
  NAND3_X1 U15472 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .ZN(n15481) );
  NOR2_X1 U15473 ( .A1(n13531), .A2(n15481), .ZN(n13962) );
  NAND4_X1 U15474 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(P1_REIP_REG_19__SCAN_IN), 
        .A3(P1_REIP_REG_18__SCAN_IN), .A4(n13962), .ZN(n15461) );
  NOR2_X1 U15475 ( .A1(n20488), .A2(n15461), .ZN(n13950) );
  NAND3_X1 U15476 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .A3(n13950), .ZN(n12384) );
  NOR2_X1 U15477 ( .A1(n15449), .A2(n12384), .ZN(n13949) );
  NAND2_X1 U15478 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n13949), .ZN(n15427) );
  NOR2_X1 U15479 ( .A1(n12385), .A2(n15427), .ZN(n13727) );
  OR2_X1 U15480 ( .A1(n12379), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n15416) );
  NAND2_X1 U15481 ( .A1(n12597), .A2(n15416), .ZN(n12479) );
  NAND2_X1 U15482 ( .A1(n12479), .A2(n15391), .ZN(n12382) );
  NOR2_X1 U15483 ( .A1(n12382), .A2(n12485), .ZN(n12380) );
  NAND2_X1 U15484 ( .A1(n13963), .A2(n13961), .ZN(n19636) );
  OR2_X1 U15485 ( .A1(n13727), .A2(n19669), .ZN(n13934) );
  INV_X1 U15486 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20496) );
  NOR2_X1 U15487 ( .A1(n13934), .A2(n20496), .ZN(n12391) );
  AND3_X1 U15488 ( .A1(n12382), .A2(n19839), .A3(n12381), .ZN(n12383) );
  NOR2_X1 U15489 ( .A1(n13963), .A2(n12384), .ZN(n15442) );
  NAND2_X1 U15490 ( .A1(n15442), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n15429) );
  NOR2_X1 U15491 ( .A1(n15429), .A2(n12385), .ZN(n13918) );
  NAND2_X1 U15492 ( .A1(n13918), .A2(n20496), .ZN(n12389) );
  AND2_X1 U15493 ( .A1(n14087), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12386) );
  INV_X1 U15494 ( .A(n14116), .ZN(n12387) );
  AOI22_X1 U15495 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n19675), .B1(
        n19644), .B2(n12387), .ZN(n12388) );
  OAI211_X1 U15496 ( .C1(n13975), .C2(n19662), .A(n12389), .B(n12388), .ZN(
        n12390) );
  INV_X1 U15497 ( .A(n12394), .ZN(n12395) );
  INV_X1 U15498 ( .A(n12846), .ZN(n18700) );
  NAND2_X1 U15499 ( .A1(n12395), .A2(n18700), .ZN(n18644) );
  OR2_X1 U15500 ( .A1(n12397), .A2(n12396), .ZN(n12399) );
  AOI21_X1 U15501 ( .B1(P2_MEMORYFETCH_REG_SCAN_IN), .B2(n18644), .A(n12399), 
        .ZN(n12398) );
  INV_X1 U15502 ( .A(n12398), .ZN(P2_U2814) );
  NOR2_X1 U15503 ( .A1(P2_READREQUEST_REG_SCAN_IN), .A2(n12399), .ZN(n12400)
         );
  INV_X1 U15504 ( .A(n12626), .ZN(n19584) );
  AOI22_X1 U15505 ( .A1(n12400), .A2(n18644), .B1(n18414), .B2(n19584), .ZN(
        P2_U3612) );
  INV_X1 U15506 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n18707) );
  NAND2_X2 U15507 ( .A1(n12401), .A2(n19593), .ZN(n18804) );
  INV_X2 U15508 ( .A(n18702), .ZN(n18801) );
  NAND2_X1 U15509 ( .A1(n18773), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n12405) );
  INV_X1 U15510 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n12402) );
  OR2_X1 U15511 ( .A1(n14633), .A2(n12402), .ZN(n12404) );
  NAND2_X1 U15512 ( .A1(n14610), .A2(BUF2_REG_14__SCAN_IN), .ZN(n12403) );
  NAND2_X1 U15513 ( .A1(n12404), .A2(n12403), .ZN(n18656) );
  NAND2_X1 U15514 ( .A1(n12410), .A2(n18656), .ZN(n12622) );
  OAI211_X1 U15515 ( .C1(n18707), .C2(n18702), .A(n12405), .B(n12622), .ZN(
        P2_U2966) );
  INV_X1 U15516 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n18745) );
  NAND2_X1 U15517 ( .A1(n18773), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n12408) );
  INV_X1 U15518 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16023) );
  OR2_X1 U15519 ( .A1(n14610), .A2(n16023), .ZN(n12407) );
  NAND2_X1 U15520 ( .A1(n14610), .A2(BUF2_REG_12__SCAN_IN), .ZN(n12406) );
  NAND2_X1 U15521 ( .A1(n12407), .A2(n12406), .ZN(n18660) );
  NAND2_X1 U15522 ( .A1(n12410), .A2(n18660), .ZN(n12618) );
  OAI211_X1 U15523 ( .C1(n18745), .C2(n18702), .A(n12408), .B(n12618), .ZN(
        P2_U2979) );
  INV_X1 U15524 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n18752) );
  NAND2_X1 U15525 ( .A1(n18773), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n12411) );
  INV_X1 U15526 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n20584) );
  INV_X1 U15527 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n12409) );
  AOI22_X1 U15528 ( .A1(n14634), .A2(n20584), .B1(n12409), .B2(n14610), .ZN(
        n18663) );
  NAND2_X1 U15529 ( .A1(n12410), .A2(n18663), .ZN(n12620) );
  OAI211_X1 U15530 ( .C1(n18752), .C2(n18702), .A(n12411), .B(n12620), .ZN(
        P2_U2975) );
  NOR2_X1 U15531 ( .A1(n20516), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n19600) );
  AOI21_X1 U15532 ( .B1(n12412), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n19600), 
        .ZN(n12413) );
  NAND2_X1 U15533 ( .A1(n12642), .A2(n12413), .ZN(P1_U2801) );
  NOR2_X1 U15534 ( .A1(n12414), .A2(n11246), .ZN(n12415) );
  AOI21_X1 U15535 ( .B1(n12691), .B2(n12508), .A(n12415), .ZN(n19601) );
  NAND3_X1 U15536 ( .A1(n12508), .A2(n15416), .A3(n13886), .ZN(n12416) );
  NAND2_X1 U15537 ( .A1(n12416), .A2(n20546), .ZN(n20544) );
  NAND2_X1 U15538 ( .A1(n19601), .A2(n20544), .ZN(n15386) );
  AND2_X1 U15539 ( .A1(n15386), .A2(n12696), .ZN(n19610) );
  INV_X1 U15540 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n12431) );
  INV_X1 U15541 ( .A(n11063), .ZN(n12417) );
  NAND2_X1 U15542 ( .A1(n12417), .A2(n13887), .ZN(n12419) );
  INV_X1 U15543 ( .A(n12492), .ZN(n13062) );
  NAND2_X1 U15544 ( .A1(n12420), .A2(n13062), .ZN(n12418) );
  AND2_X1 U15545 ( .A1(n12419), .A2(n12418), .ZN(n12504) );
  NOR2_X1 U15546 ( .A1(n14422), .A2(n12597), .ZN(n12690) );
  INV_X1 U15547 ( .A(n12705), .ZN(n12427) );
  NAND2_X1 U15548 ( .A1(n12420), .A2(n12508), .ZN(n12421) );
  NAND2_X1 U15549 ( .A1(n12484), .A2(n12421), .ZN(n12700) );
  INV_X1 U15550 ( .A(n12700), .ZN(n12422) );
  OAI21_X1 U15551 ( .B1(n12423), .B2(n12422), .A(n12691), .ZN(n12426) );
  NAND2_X1 U15552 ( .A1(n12483), .A2(n12424), .ZN(n12425) );
  OAI211_X1 U15553 ( .C1(n12691), .C2(n12427), .A(n12426), .B(n12425), .ZN(
        n12428) );
  NAND2_X1 U15554 ( .A1(n12428), .A2(n19886), .ZN(n15383) );
  INV_X1 U15555 ( .A(n15383), .ZN(n12429) );
  NAND2_X1 U15556 ( .A1(n19610), .A2(n12429), .ZN(n12430) );
  OAI21_X1 U15557 ( .B1(n19610), .B2(n12431), .A(n12430), .ZN(P1_U3484) );
  NOR2_X1 U15558 ( .A1(n19600), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n12433)
         );
  OAI21_X1 U15559 ( .B1(n13056), .B2(n9692), .A(n20550), .ZN(n12432) );
  OAI21_X1 U15560 ( .B1(n12433), .B2(n20550), .A(n12432), .ZN(P1_U3487) );
  NOR2_X1 U15561 ( .A1(n19533), .A2(n19263), .ZN(n19552) );
  NAND2_X1 U15562 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n19563) );
  NAND2_X1 U15563 ( .A1(n13706), .A2(n19586), .ZN(n15905) );
  NAND2_X1 U15564 ( .A1(n15904), .A2(n15905), .ZN(n19585) );
  NAND2_X1 U15565 ( .A1(n12436), .A2(n12435), .ZN(n12437) );
  NAND2_X1 U15566 ( .A1(n12438), .A2(n12437), .ZN(n12439) );
  AND2_X1 U15567 ( .A1(n12440), .A2(n12439), .ZN(n12441) );
  OR2_X1 U15568 ( .A1(n12442), .A2(n12441), .ZN(n19572) );
  INV_X1 U15569 ( .A(n12538), .ZN(n12444) );
  INV_X1 U15570 ( .A(n12833), .ZN(n12445) );
  OAI21_X1 U15571 ( .B1(n12456), .B2(n12446), .A(n12445), .ZN(n12447) );
  INV_X1 U15572 ( .A(n12447), .ZN(n12451) );
  NAND2_X1 U15573 ( .A1(n12815), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12449) );
  NAND2_X1 U15574 ( .A1(n12449), .A2(n15192), .ZN(n12844) );
  INV_X1 U15575 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n12450) );
  OAI21_X1 U15576 ( .B1(n11618), .B2(n12844), .A(n12450), .ZN(n19562) );
  MUX2_X1 U15577 ( .A(n12451), .B(n19562), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n19574) );
  NAND2_X1 U15578 ( .A1(n19574), .A2(n9643), .ZN(n12452) );
  OAI22_X1 U15579 ( .A1(n19572), .A2(n19575), .B1(n12848), .B2(n12452), .ZN(
        n12553) );
  NOR2_X1 U15580 ( .A1(n9634), .A2(n18416), .ZN(n12453) );
  NAND2_X1 U15581 ( .A1(n12553), .A2(n12453), .ZN(n18418) );
  OR2_X1 U15582 ( .A1(n12468), .A2(n9643), .ZN(n12454) );
  INV_X1 U15583 ( .A(n12454), .ZN(n13294) );
  NAND2_X1 U15584 ( .A1(n12454), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13349) );
  INV_X1 U15585 ( .A(n13349), .ZN(n12469) );
  AOI21_X1 U15586 ( .B1(n13294), .B2(n10038), .A(n12469), .ZN(n12573) );
  MUX2_X1 U15587 ( .A(n12456), .B(n12468), .S(n12455), .Z(n12458) );
  AOI21_X1 U15588 ( .B1(n12458), .B2(n9614), .A(n12457), .ZN(n14439) );
  NAND2_X1 U15589 ( .A1(n14439), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13334) );
  OAI21_X1 U15590 ( .B1(n14439), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13334), .ZN(n12570) );
  NAND2_X1 U15591 ( .A1(n18850), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n12560) );
  OAI21_X1 U15592 ( .B1(n18833), .B2(n12570), .A(n12560), .ZN(n12459) );
  AOI21_X1 U15593 ( .B1(n18821), .B2(n12573), .A(n12459), .ZN(n12465) );
  NAND2_X1 U15594 ( .A1(n19533), .A2(n19537), .ZN(n19561) );
  NAND2_X1 U15595 ( .A1(n19561), .A2(n15904), .ZN(n12460) );
  INV_X1 U15596 ( .A(n12461), .ZN(n12463) );
  NAND2_X1 U15597 ( .A1(n19263), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12462) );
  NAND2_X1 U15598 ( .A1(n12463), .A2(n12462), .ZN(n12472) );
  OAI21_X1 U15599 ( .B1(n18820), .B2(n12472), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12464) );
  OAI211_X1 U15600 ( .C1(n18811), .C2(n13221), .A(n12465), .B(n12464), .ZN(
        P2_U3014) );
  NAND3_X1 U15601 ( .A1(n18911), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n12466) );
  NAND2_X1 U15602 ( .A1(n13073), .A2(n12466), .ZN(n13333) );
  NAND2_X1 U15603 ( .A1(n13334), .A2(n13333), .ZN(n13335) );
  OAI21_X1 U15604 ( .B1(n13333), .B2(n13334), .A(n13335), .ZN(n12467) );
  XOR2_X1 U15605 ( .A(n12467), .B(n15083), .Z(n15087) );
  INV_X1 U15606 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12475) );
  XOR2_X1 U15607 ( .A(n12468), .B(n13293), .Z(n13348) );
  XOR2_X1 U15608 ( .A(n12469), .B(n13348), .Z(n12470) );
  NOR2_X1 U15609 ( .A1(n15083), .A2(n12470), .ZN(n13350) );
  AOI21_X1 U15610 ( .B1(n15083), .B2(n12470), .A(n13350), .ZN(n15086) );
  NAND2_X1 U15611 ( .A1(n18850), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n15089) );
  INV_X1 U15612 ( .A(n15089), .ZN(n12471) );
  AOI21_X1 U15613 ( .B1(n18821), .B2(n15086), .A(n12471), .ZN(n12474) );
  NAND2_X1 U15614 ( .A1(n18829), .A2(n12475), .ZN(n12473) );
  OAI211_X1 U15615 ( .C1(n15852), .C2(n12475), .A(n12474), .B(n12473), .ZN(
        n12476) );
  AOI21_X1 U15616 ( .B1(n18808), .B2(n15087), .A(n12476), .ZN(n12477) );
  OAI21_X1 U15617 ( .B1(n15080), .B2(n18811), .A(n12477), .ZN(P2_U3013) );
  INV_X1 U15618 ( .A(n12515), .ZN(n12498) );
  INV_X1 U15619 ( .A(n12691), .ZN(n12495) );
  INV_X1 U15620 ( .A(n12712), .ZN(n14421) );
  INV_X1 U15621 ( .A(n15416), .ZN(n12481) );
  NAND2_X1 U15622 ( .A1(n12479), .A2(n20546), .ZN(n12685) );
  INV_X1 U15623 ( .A(n12685), .ZN(n12480) );
  OAI21_X1 U15624 ( .B1(n11246), .B2(n12481), .A(n12480), .ZN(n12482) );
  AOI21_X1 U15625 ( .B1(n14421), .B2(n12686), .A(n12482), .ZN(n12494) );
  INV_X1 U15626 ( .A(n12483), .ZN(n12490) );
  INV_X1 U15627 ( .A(n12484), .ZN(n12489) );
  AOI21_X1 U15628 ( .B1(n12486), .B2(n19853), .A(n12485), .ZN(n12487) );
  AND2_X1 U15629 ( .A1(n12488), .A2(n12487), .ZN(n12501) );
  AOI21_X1 U15630 ( .B1(n12490), .B2(n12489), .A(n12501), .ZN(n12692) );
  OAI211_X1 U15631 ( .C1(n12492), .C2(n19858), .A(n12692), .B(n12491), .ZN(
        n12493) );
  AOI21_X1 U15632 ( .B1(n12495), .B2(n12494), .A(n12493), .ZN(n12497) );
  INV_X1 U15633 ( .A(n12650), .ZN(n12496) );
  OAI211_X1 U15634 ( .C1(n12691), .C2(n12498), .A(n12497), .B(n12496), .ZN(
        n15374) );
  INV_X1 U15635 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20270) );
  NAND2_X1 U15636 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n15683) );
  INV_X1 U15637 ( .A(n15683), .ZN(n14416) );
  NAND2_X1 U15638 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n14416), .ZN(n15688) );
  INV_X1 U15639 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19609) );
  OAI22_X1 U15640 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20270), .B1(n15688), 
        .B2(n19609), .ZN(n12499) );
  AOI21_X1 U15641 ( .B1(n15374), .B2(n12696), .A(n12499), .ZN(n14437) );
  INV_X1 U15642 ( .A(n12500), .ZN(n12509) );
  INV_X1 U15643 ( .A(n12501), .ZN(n12507) );
  NAND2_X1 U15644 ( .A1(n12502), .A2(n12917), .ZN(n12503) );
  NAND2_X1 U15645 ( .A1(n12503), .A2(n19853), .ZN(n12505) );
  AND2_X1 U15646 ( .A1(n12505), .A2(n12504), .ZN(n12506) );
  OAI211_X1 U15647 ( .C1(n12509), .C2(n12508), .A(n12507), .B(n12506), .ZN(
        n12709) );
  INV_X1 U15648 ( .A(n12510), .ZN(n12512) );
  NAND3_X1 U15649 ( .A1(n12512), .A2(n12686), .A3(n12511), .ZN(n12513) );
  NOR2_X1 U15650 ( .A1(n12709), .A2(n12513), .ZN(n12514) );
  NAND2_X1 U15651 ( .A1(n12514), .A2(n11247), .ZN(n14425) );
  INV_X1 U15652 ( .A(n14425), .ZN(n12523) );
  OR2_X1 U15653 ( .A1(n12515), .A2(n12705), .ZN(n12919) );
  XNOR2_X1 U15654 ( .A(n14427), .B(n12516), .ZN(n12524) );
  INV_X1 U15655 ( .A(n12524), .ZN(n12519) );
  XNOR2_X1 U15656 ( .A(n12517), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12518) );
  AOI22_X1 U15657 ( .A1(n12919), .A2(n12519), .B1(n12712), .B2(n12518), .ZN(
        n12522) );
  NAND3_X1 U15658 ( .A1(n12523), .A2(n12520), .A3(n12524), .ZN(n12521) );
  OAI211_X1 U15659 ( .C1(n20259), .C2(n12523), .A(n12522), .B(n12521), .ZN(
        n12912) );
  INV_X1 U15660 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13554) );
  NOR2_X1 U15661 ( .A1(n20445), .A2(n13554), .ZN(n14430) );
  INV_X1 U15662 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14238) );
  OAI22_X1 U15663 ( .A1(n14238), .A2(n19819), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14431) );
  INV_X1 U15664 ( .A(n14431), .ZN(n12525) );
  AOI222_X1 U15665 ( .A1(n12912), .A2(n12614), .B1(n14430), .B2(n12525), .C1(
        n14426), .C2(n12524), .ZN(n12527) );
  NAND2_X1 U15666 ( .A1(n14437), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12526) );
  OAI21_X1 U15667 ( .B1(n14437), .B2(n12527), .A(n12526), .ZN(P1_U3472) );
  MUX2_X1 U15668 ( .A(n11412), .B(n15080), .S(n14540), .Z(n12529) );
  OAI21_X1 U15669 ( .B1(n19557), .B2(n14550), .A(n12529), .ZN(P2_U2886) );
  NOR2_X1 U15670 ( .A1(n12839), .A2(n18895), .ZN(n18701) );
  INV_X1 U15671 ( .A(n12840), .ZN(n12786) );
  NAND3_X1 U15672 ( .A1(n18701), .A2(n12786), .A3(n12549), .ZN(n12556) );
  INV_X1 U15673 ( .A(n18701), .ZN(n12532) );
  AOI21_X1 U15674 ( .B1(n12530), .B2(n9634), .A(n18907), .ZN(n12531) );
  NAND2_X1 U15675 ( .A1(n12532), .A2(n12531), .ZN(n12555) );
  NAND2_X1 U15676 ( .A1(n12859), .A2(n12786), .ZN(n12533) );
  OR2_X1 U15677 ( .A1(n12833), .A2(n12533), .ZN(n12548) );
  NAND2_X1 U15678 ( .A1(n12534), .A2(n18900), .ZN(n12535) );
  NAND2_X1 U15679 ( .A1(n12846), .A2(n12535), .ZN(n12546) );
  NAND2_X1 U15680 ( .A1(n12536), .A2(n11373), .ZN(n12537) );
  NAND2_X1 U15681 ( .A1(n12537), .A2(n12630), .ZN(n12539) );
  NAND2_X1 U15682 ( .A1(n12539), .A2(n12538), .ZN(n12580) );
  NAND2_X1 U15683 ( .A1(n18895), .A2(n12541), .ZN(n12574) );
  NAND2_X1 U15684 ( .A1(n12574), .A2(n9634), .ZN(n12542) );
  NAND3_X1 U15685 ( .A1(n12542), .A2(n12581), .A3(n12630), .ZN(n12543) );
  NAND2_X1 U15686 ( .A1(n12543), .A2(n18900), .ZN(n12544) );
  NAND4_X1 U15687 ( .A1(n12546), .A2(n12545), .A3(n12580), .A4(n12544), .ZN(
        n12575) );
  INV_X1 U15688 ( .A(n12575), .ZN(n12547) );
  MUX2_X1 U15689 ( .A(n12859), .B(n12549), .S(n18895), .Z(n12550) );
  NAND2_X1 U15690 ( .A1(n12550), .A2(n19593), .ZN(n12551) );
  NOR2_X1 U15691 ( .A1(n12833), .A2(n12551), .ZN(n12552) );
  NOR2_X1 U15692 ( .A1(n12553), .A2(n12552), .ZN(n12554) );
  NAND4_X1 U15693 ( .A1(n12556), .A2(n12555), .A3(n12784), .A4(n12554), .ZN(
        n12557) );
  AOI21_X1 U15694 ( .B1(n18895), .B2(n12811), .A(n12558), .ZN(n12559) );
  OAI21_X1 U15695 ( .B1(n18839), .B2(n13221), .A(n12560), .ZN(n12572) );
  OR2_X1 U15696 ( .A1(n12848), .A2(n11382), .ZN(n19573) );
  AND2_X1 U15697 ( .A1(n12832), .A2(n9643), .ZN(n12561) );
  NOR2_X1 U15698 ( .A1(n12778), .A2(n12561), .ZN(n12562) );
  INV_X1 U15699 ( .A(n12563), .ZN(n12569) );
  INV_X1 U15700 ( .A(n12564), .ZN(n12567) );
  INV_X1 U15701 ( .A(n12565), .ZN(n12566) );
  NAND2_X1 U15702 ( .A1(n12567), .A2(n12566), .ZN(n12568) );
  NAND2_X1 U15703 ( .A1(n12569), .A2(n12568), .ZN(n14443) );
  OAI22_X1 U15704 ( .A1(n18859), .A2(n12570), .B1(n15898), .B2(n14443), .ZN(
        n12571) );
  AOI211_X1 U15705 ( .C1(n18849), .C2(n12573), .A(n12572), .B(n12571), .ZN(
        n12596) );
  INV_X1 U15706 ( .A(n12576), .ZN(n12577) );
  NOR2_X1 U15707 ( .A1(n12578), .A2(n12577), .ZN(n12627) );
  NAND2_X1 U15708 ( .A1(n12579), .A2(n9643), .ZN(n12793) );
  NAND2_X1 U15709 ( .A1(n12793), .A2(n12580), .ZN(n12582) );
  NAND2_X1 U15710 ( .A1(n12582), .A2(n12581), .ZN(n12590) );
  INV_X1 U15711 ( .A(n12583), .ZN(n12585) );
  OAI21_X1 U15712 ( .B1(n12585), .B2(n12584), .A(n12626), .ZN(n12587) );
  OAI22_X1 U15713 ( .A1(n12626), .A2(n18907), .B1(n9634), .B2(n18900), .ZN(
        n12586) );
  AOI21_X1 U15714 ( .B1(n12587), .B2(n9644), .A(n12586), .ZN(n12589) );
  NAND3_X1 U15715 ( .A1(n12590), .A2(n12589), .A3(n12588), .ZN(n12591) );
  OR2_X1 U15716 ( .A1(n12627), .A2(n12591), .ZN(n12806) );
  NOR2_X1 U15717 ( .A1(n12806), .A2(n12775), .ZN(n12592) );
  INV_X1 U15718 ( .A(n14943), .ZN(n15081) );
  AND2_X1 U15719 ( .A1(n12593), .A2(n18496), .ZN(n18855) );
  INV_X1 U15720 ( .A(n18855), .ZN(n12594) );
  MUX2_X1 U15721 ( .A(n15081), .B(n12594), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n12595) );
  NAND2_X1 U15722 ( .A1(n12596), .A2(n12595), .ZN(P2_U3046) );
  INV_X1 U15723 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n12600) );
  NAND2_X1 U15724 ( .A1(n11246), .A2(n12597), .ZN(n12714) );
  AOI21_X1 U15725 ( .B1(n14421), .B2(n12714), .A(n15416), .ZN(n12598) );
  NAND2_X1 U15726 ( .A1(n19716), .A2(n19839), .ZN(n12763) );
  NOR2_X1 U15727 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15683), .ZN(n19736) );
  NOR2_X4 U15728 ( .A1(n19716), .A2(n19746), .ZN(n19745) );
  AOI22_X1 U15729 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n19746), .B1(n19745), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n12599) );
  OAI21_X1 U15730 ( .B1(n12600), .B2(n12763), .A(n12599), .ZN(P1_U2911) );
  INV_X1 U15731 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n12602) );
  AOI22_X1 U15732 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n19746), .B1(n19745), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n12601) );
  OAI21_X1 U15733 ( .B1(n12602), .B2(n12763), .A(n12601), .ZN(P1_U2908) );
  INV_X1 U15734 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n12604) );
  AOI22_X1 U15735 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n19746), .B1(n19745), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12603) );
  OAI21_X1 U15736 ( .B1(n12604), .B2(n12763), .A(n12603), .ZN(P1_U2907) );
  INV_X1 U15737 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n12606) );
  AOI22_X1 U15738 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n19746), .B1(n19745), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12605) );
  OAI21_X1 U15739 ( .B1(n12606), .B2(n12763), .A(n12605), .ZN(P1_U2906) );
  INV_X1 U15740 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n12608) );
  AOI22_X1 U15741 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n19746), .B1(n19745), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n12607) );
  OAI21_X1 U15742 ( .B1(n12608), .B2(n12763), .A(n12607), .ZN(P1_U2910) );
  INV_X1 U15743 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n12610) );
  AOI22_X1 U15744 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n19746), .B1(n19745), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n12609) );
  OAI21_X1 U15745 ( .B1(n12610), .B2(n12763), .A(n12609), .ZN(P1_U2912) );
  AOI22_X1 U15746 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n19746), .B1(n19745), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n12611) );
  OAI21_X1 U15747 ( .B1(n14032), .B2(n12763), .A(n12611), .ZN(P1_U2909) );
  INV_X1 U15748 ( .A(n14437), .ZN(n12640) );
  AOI22_X1 U15749 ( .A1(n19961), .A2(n14425), .B1(n12612), .B2(n12617), .ZN(
        n15369) );
  INV_X1 U15750 ( .A(n12614), .ZN(n14435) );
  AOI22_X1 U15751 ( .A1(n12617), .A2(n14426), .B1(n13554), .B2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n12613) );
  OAI21_X1 U15752 ( .B1(n15369), .B2(n14435), .A(n12613), .ZN(n12615) );
  AND2_X1 U15753 ( .A1(n12712), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15370) );
  AOI22_X1 U15754 ( .A1(n12640), .A2(n12615), .B1(n12614), .B2(n15370), .ZN(
        n12616) );
  OAI21_X1 U15755 ( .B1(n12617), .B2(n12640), .A(n12616), .ZN(P1_U3474) );
  INV_X1 U15756 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n18711) );
  NAND2_X1 U15757 ( .A1(n18802), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n12619) );
  OAI211_X1 U15758 ( .C1(n18711), .C2(n18702), .A(n12619), .B(n12618), .ZN(
        P2_U2964) );
  INV_X1 U15759 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n18719) );
  NAND2_X1 U15760 ( .A1(n18802), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n12621) );
  OAI211_X1 U15761 ( .C1(n18719), .C2(n18702), .A(n12621), .B(n12620), .ZN(
        P2_U2960) );
  INV_X1 U15762 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n18741) );
  NAND2_X1 U15763 ( .A1(n18802), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n12623) );
  OAI211_X1 U15764 ( .C1(n18741), .C2(n18702), .A(n12623), .B(n12622), .ZN(
        P2_U2981) );
  XNOR2_X1 U15765 ( .A(n12625), .B(n12624), .ZN(n18613) );
  NAND2_X1 U15766 ( .A1(n12626), .A2(n19593), .ZN(n12841) );
  OAI22_X1 U15767 ( .A1(n12839), .A2(n12834), .B1(n12841), .B2(n12843), .ZN(
        n12783) );
  INV_X1 U15768 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n18757) );
  AND2_X1 U15769 ( .A1(n18686), .A2(n12629), .ZN(n15778) );
  NAND2_X1 U15770 ( .A1(n12631), .A2(n12630), .ZN(n12632) );
  INV_X1 U15771 ( .A(n13199), .ZN(n12633) );
  AOI22_X1 U15772 ( .A1(n14634), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n14633), .ZN(n18920) );
  OAI222_X1 U15773 ( .A1(n18613), .A2(n18675), .B1(n18686), .B2(n18757), .C1(
        n18698), .C2(n18920), .ZN(P2_U2913) );
  OAI21_X1 U15774 ( .B1(n12635), .B2(n12634), .A(n15885), .ZN(n18599) );
  AOI22_X1 U15775 ( .A1(n14634), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n14633), .ZN(n18928) );
  OAI222_X1 U15776 ( .A1(n18599), .A2(n18675), .B1(n18686), .B2(n18754), .C1(
        n18698), .C2(n18928), .ZN(P2_U2912) );
  INV_X1 U15777 ( .A(n19995), .ZN(n20258) );
  OR2_X1 U15778 ( .A1(n12636), .A2(n20258), .ZN(n12638) );
  XNOR2_X1 U15779 ( .A(n12638), .B(n12637), .ZN(n19680) );
  OR4_X1 U15780 ( .A1(n14437), .A2(n14435), .A3(n11247), .A4(n19680), .ZN(
        n12639) );
  OAI21_X1 U15781 ( .B1(n12640), .B2(n12637), .A(n12639), .ZN(P1_U3468) );
  AND2_X1 U15782 ( .A1(n20541), .A2(n20457), .ZN(n12641) );
  OR2_X2 U15783 ( .A1(n12642), .A2(n12641), .ZN(n19773) );
  INV_X1 U15784 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n12646) );
  INV_X1 U15785 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n12643) );
  NOR2_X1 U15786 ( .A1(n19834), .A2(n12643), .ZN(n12644) );
  AOI21_X1 U15787 ( .B1(DATAI_15_), .B2(n19834), .A(n12644), .ZN(n14078) );
  INV_X1 U15788 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n12645) );
  INV_X1 U15789 ( .A(n19773), .ZN(n12958) );
  OAI222_X1 U15790 ( .A1(n12957), .A2(n12646), .B1(n12959), .B2(n14078), .C1(
        n12645), .C2(n12958), .ZN(P1_U2967) );
  OAI21_X1 U15791 ( .B1(n12649), .B2(n12648), .A(n12647), .ZN(n13090) );
  XNOR2_X1 U15792 ( .A(n13087), .B(n13715), .ZN(n12886) );
  INV_X1 U15793 ( .A(n12886), .ZN(n12655) );
  OAI22_X1 U15794 ( .A1(n14025), .A2(n12655), .B1(n12654), .B2(n19710), .ZN(
        n12656) );
  INV_X1 U15795 ( .A(n12656), .ZN(n12657) );
  OAI21_X1 U15796 ( .B1(n13090), .B2(n14024), .A(n12657), .ZN(P1_U2871) );
  BUF_X4 U15797 ( .A(n13226), .Z(n15895) );
  MUX2_X1 U15798 ( .A(P2_EBX_REG_3__SCAN_IN), .B(n15895), .S(n14540), .Z(
        n12660) );
  INV_X1 U15799 ( .A(n12660), .ZN(n12661) );
  OAI21_X1 U15800 ( .B1(n19540), .B2(n14550), .A(n12661), .ZN(P2_U2884) );
  NAND2_X1 U15801 ( .A1(n9643), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12662) );
  NAND4_X1 U15802 ( .A1(n12662), .A2(n18919), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n19535), .ZN(n12663) );
  INV_X1 U15803 ( .A(n14548), .ZN(n14525) );
  MUX2_X1 U15804 ( .A(n12665), .B(n13221), .S(n14525), .Z(n12666) );
  OAI21_X1 U15805 ( .B1(n14550), .B2(n19566), .A(n12666), .ZN(P2_U2887) );
  NAND2_X1 U15806 ( .A1(n12667), .A2(n12724), .ZN(n12668) );
  OAI21_X1 U15807 ( .B1(n12667), .B2(n12724), .A(n12668), .ZN(n18677) );
  OR2_X1 U15808 ( .A1(n9764), .A2(n12669), .ZN(n12670) );
  NAND2_X1 U15809 ( .A1(n12670), .A2(n12727), .ZN(n18838) );
  MUX2_X1 U15810 ( .A(n12671), .B(n18838), .S(n14540), .Z(n12672) );
  OAI21_X1 U15811 ( .B1(n18677), .B2(n14550), .A(n12672), .ZN(P2_U2883) );
  OR2_X1 U15812 ( .A1(n12674), .A2(n12673), .ZN(n12675) );
  NAND2_X1 U15813 ( .A1(n12676), .A2(n12675), .ZN(n19715) );
  NAND2_X1 U15814 ( .A1(n12677), .A2(n14190), .ZN(n12682) );
  INV_X1 U15815 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13108) );
  NOR2_X1 U15816 ( .A1(n19798), .A2(n13108), .ZN(n12720) );
  OR2_X1 U15817 ( .A1(n12678), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12679) );
  NAND2_X1 U15818 ( .A1(n12680), .A2(n12679), .ZN(n12723) );
  NOR2_X1 U15819 ( .A1(n19608), .A2(n12723), .ZN(n12681) );
  AOI211_X1 U15820 ( .C1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n12682), .A(
        n12720), .B(n12681), .ZN(n12683) );
  OAI21_X1 U15821 ( .B1(n19835), .B2(n19715), .A(n12683), .ZN(P1_U2999) );
  OAI211_X1 U15822 ( .C1(n12686), .C2(n12685), .A(n19839), .B(n12684), .ZN(
        n12687) );
  NAND3_X1 U15823 ( .A1(n12688), .A2(n9615), .A3(n12687), .ZN(n12699) );
  NAND2_X1 U15824 ( .A1(n19853), .A2(n15416), .ZN(n12689) );
  NAND2_X1 U15825 ( .A1(n12689), .A2(n19858), .ZN(n12694) );
  NAND2_X1 U15826 ( .A1(n12691), .A2(n12690), .ZN(n12693) );
  OAI211_X1 U15827 ( .C1(n12695), .C2(n12694), .A(n12693), .B(n12692), .ZN(
        n12697) );
  NAND2_X1 U15828 ( .A1(n12697), .A2(n12696), .ZN(n12698) );
  OAI21_X1 U15829 ( .B1(n12701), .B2(n12715), .A(n12700), .ZN(n12702) );
  OR2_X1 U15830 ( .A1(n12703), .A2(n12702), .ZN(n12704) );
  MUX2_X1 U15831 ( .A(n12706), .B(n9615), .S(n19839), .Z(n12708) );
  NAND2_X1 U15832 ( .A1(n12708), .A2(n12707), .ZN(n12710) );
  OR2_X1 U15833 ( .A1(n12710), .A2(n12709), .ZN(n12711) );
  NAND2_X1 U15834 ( .A1(n12717), .A2(n12711), .ZN(n14326) );
  NAND2_X1 U15835 ( .A1(n19824), .A2(n14326), .ZN(n12883) );
  OR2_X1 U15836 ( .A1(n12717), .A2(n19781), .ZN(n13555) );
  AOI21_X1 U15837 ( .B1(n13555), .B2(n15609), .A(n13554), .ZN(n12713) );
  AOI21_X1 U15838 ( .B1(n13554), .B2(n12883), .A(n12713), .ZN(n12722) );
  OAI21_X1 U15839 ( .B1(n12715), .B2(n10396), .A(n12714), .ZN(n12716) );
  OR2_X1 U15840 ( .A1(n13887), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12719) );
  AND2_X1 U15841 ( .A1(n12719), .A2(n12718), .ZN(n13105) );
  AOI21_X1 U15842 ( .B1(n19807), .B2(n13105), .A(n12720), .ZN(n12721) );
  OAI211_X1 U15843 ( .C1(n19820), .C2(n12723), .A(n12722), .B(n12721), .ZN(
        P1_U3031) );
  AND2_X1 U15844 ( .A1(n12667), .A2(n12724), .ZN(n12726) );
  OAI211_X1 U15845 ( .C1(n12726), .C2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A(
        n14522), .B(n12725), .ZN(n12731) );
  NAND2_X1 U15846 ( .A1(n12728), .A2(n12727), .ZN(n12729) );
  AND2_X1 U15847 ( .A1(n12729), .A2(n10033), .ZN(n18624) );
  NAND2_X1 U15848 ( .A1(n14540), .A2(n18624), .ZN(n12730) );
  OAI211_X1 U15849 ( .C1(n14525), .C2(n12732), .A(n12731), .B(n12730), .ZN(
        P2_U2882) );
  XOR2_X1 U15850 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B(n12725), .Z(n12737)
         );
  NOR2_X1 U15851 ( .A1(n12734), .A2(n12733), .ZN(n12735) );
  OR2_X1 U15852 ( .A1(n12769), .A2(n12735), .ZN(n13492) );
  MUX2_X1 U15853 ( .A(n11878), .B(n13492), .S(n14540), .Z(n12736) );
  OAI21_X1 U15854 ( .B1(n12737), .B2(n14550), .A(n12736), .ZN(P2_U2881) );
  OAI21_X1 U15855 ( .B1(n12738), .B2(n15884), .A(n12746), .ZN(n18576) );
  AOI22_X1 U15856 ( .A1(n14634), .A2(BUF1_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n14633), .ZN(n18794) );
  INV_X1 U15857 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n18750) );
  OAI222_X1 U15858 ( .A1(n18576), .A2(n18675), .B1(n18794), .B2(n18698), .C1(
        n18750), .C2(n18686), .ZN(P2_U2910) );
  INV_X1 U15859 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13082) );
  INV_X1 U15860 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n13060) );
  NOR2_X1 U15861 ( .A1(n19798), .A2(n13060), .ZN(n12885) );
  NOR2_X1 U15862 ( .A1(n14190), .A2(n13082), .ZN(n12739) );
  AOI211_X1 U15863 ( .C1(n15566), .C2(n13082), .A(n12885), .B(n12739), .ZN(
        n12742) );
  OR2_X1 U15864 ( .A1(n12740), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12887) );
  NAND3_X1 U15865 ( .A1(n12887), .A2(n12888), .A3(n19788), .ZN(n12741) );
  OAI211_X1 U15866 ( .C1(n13090), .C2(n19835), .A(n12742), .B(n12741), .ZN(
        P1_U2998) );
  INV_X1 U15867 ( .A(n19546), .ZN(n12743) );
  NAND2_X1 U15868 ( .A1(n12743), .A2(n14522), .ZN(n12745) );
  BUF_X4 U15869 ( .A(n13233), .Z(n13260) );
  NAND2_X1 U15870 ( .A1(n14540), .A2(n13260), .ZN(n12744) );
  OAI211_X1 U15871 ( .C1(n14525), .C2(n11427), .A(n12745), .B(n12744), .ZN(
        P2_U2885) );
  XNOR2_X1 U15872 ( .A(n12747), .B(n12746), .ZN(n18565) );
  AOI22_X1 U15873 ( .A1(n14634), .A2(BUF1_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n14610), .ZN(n18796) );
  INV_X1 U15874 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n20620) );
  OAI222_X1 U15875 ( .A1(n18565), .A2(n18675), .B1(n18796), .B2(n18698), .C1(
        n20620), .C2(n18686), .ZN(P2_U2909) );
  INV_X1 U15876 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n12749) );
  AOI22_X1 U15877 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n19736), .B1(n19745), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n12748) );
  OAI21_X1 U15878 ( .B1(n12749), .B2(n12763), .A(n12748), .ZN(P1_U2920) );
  INV_X1 U15879 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n12751) );
  AOI22_X1 U15880 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n19736), .B1(n19745), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n12750) );
  OAI21_X1 U15881 ( .B1(n12751), .B2(n12763), .A(n12750), .ZN(P1_U2919) );
  INV_X1 U15882 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n12753) );
  AOI22_X1 U15883 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n19736), .B1(n19745), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n12752) );
  OAI21_X1 U15884 ( .B1(n12753), .B2(n12763), .A(n12752), .ZN(P1_U2917) );
  INV_X1 U15885 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n12755) );
  AOI22_X1 U15886 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n19736), .B1(n19745), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n12754) );
  OAI21_X1 U15887 ( .B1(n12755), .B2(n12763), .A(n12754), .ZN(P1_U2918) );
  INV_X1 U15888 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n12757) );
  AOI22_X1 U15889 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n19746), .B1(n19745), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n12756) );
  OAI21_X1 U15890 ( .B1(n12757), .B2(n12763), .A(n12756), .ZN(P1_U2915) );
  INV_X1 U15891 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n12759) );
  AOI22_X1 U15892 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n19746), .B1(n19745), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n12758) );
  OAI21_X1 U15893 ( .B1(n12759), .B2(n12763), .A(n12758), .ZN(P1_U2916) );
  INV_X1 U15894 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n12761) );
  AOI22_X1 U15895 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n19746), .B1(n19745), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n12760) );
  OAI21_X1 U15896 ( .B1(n12761), .B2(n12763), .A(n12760), .ZN(P1_U2913) );
  INV_X1 U15897 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n12764) );
  AOI22_X1 U15898 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n19746), .B1(n19745), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n12762) );
  OAI21_X1 U15899 ( .B1(n12764), .B2(n12763), .A(n12762), .ZN(P1_U2914) );
  NOR2_X1 U15900 ( .A1(n12725), .A2(n12765), .ZN(n12767) );
  OAI211_X1 U15901 ( .C1(n12767), .C2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A(
        n14522), .B(n12766), .ZN(n12772) );
  NOR2_X1 U15902 ( .A1(n12769), .A2(n12768), .ZN(n12770) );
  OR2_X1 U15903 ( .A1(n12946), .A2(n12770), .ZN(n14820) );
  INV_X1 U15904 ( .A(n14820), .ZN(n18596) );
  NAND2_X1 U15905 ( .A1(n14540), .A2(n18596), .ZN(n12771) );
  OAI211_X1 U15906 ( .C1(n14525), .C2(n12773), .A(n12772), .B(n12771), .ZN(
        P2_U2880) );
  NOR2_X1 U15907 ( .A1(n12774), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12812) );
  OR2_X1 U15908 ( .A1(n12558), .A2(n12775), .ZN(n12777) );
  NAND2_X1 U15909 ( .A1(n12777), .A2(n9617), .ZN(n12813) );
  INV_X1 U15910 ( .A(n12778), .ZN(n12838) );
  NAND2_X1 U15911 ( .A1(n12838), .A2(n12834), .ZN(n12808) );
  OAI21_X1 U15912 ( .B1(n9635), .B2(n12812), .A(n12808), .ZN(n12781) );
  NAND2_X1 U15913 ( .A1(n12811), .A2(n12779), .ZN(n12780) );
  OAI211_X1 U15914 ( .C1(n12812), .C2(n12813), .A(n12781), .B(n12780), .ZN(
        n12782) );
  AOI21_X1 U15915 ( .B1(n13233), .B2(n12806), .A(n12782), .ZN(n19524) );
  INV_X1 U15916 ( .A(n12783), .ZN(n12789) );
  AND2_X1 U15917 ( .A1(n12785), .A2(n12784), .ZN(n12788) );
  NAND3_X1 U15918 ( .A1(n18701), .A2(n18700), .A3(n12786), .ZN(n12787) );
  NAND3_X1 U15919 ( .A1(n12789), .A2(n12788), .A3(n12787), .ZN(n13169) );
  NAND2_X1 U15920 ( .A1(n19524), .A2(n13169), .ZN(n12791) );
  OR2_X1 U15921 ( .A1(n13169), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12790) );
  AND2_X1 U15922 ( .A1(n12791), .A2(n12790), .ZN(n12852) );
  INV_X1 U15923 ( .A(n12852), .ZN(n12805) );
  NAND2_X1 U15924 ( .A1(n12811), .A2(n12792), .ZN(n12798) );
  NAND2_X1 U15925 ( .A1(n12794), .A2(n12793), .ZN(n12800) );
  OAI21_X1 U15926 ( .B1(n12796), .B2(n12795), .A(n12800), .ZN(n12797) );
  NAND2_X1 U15927 ( .A1(n12798), .A2(n12797), .ZN(n12799) );
  AOI21_X1 U15928 ( .B1(n13263), .B2(n12806), .A(n12799), .ZN(n13166) );
  MUX2_X1 U15929 ( .A(n12811), .B(n12800), .S(n13713), .Z(n12801) );
  AOI21_X1 U15930 ( .B1(n14440), .B2(n12806), .A(n12801), .ZN(n13708) );
  OAI211_X1 U15931 ( .C1(n13166), .C2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n13708), .ZN(n12803) );
  NAND2_X1 U15932 ( .A1(n13166), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12802) );
  NAND3_X1 U15933 ( .A1(n12803), .A2(n13169), .A3(n12802), .ZN(n12804) );
  AOI21_X1 U15934 ( .B1(n12805), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n12804), .ZN(n12825) );
  NAND2_X1 U15935 ( .A1(n15895), .A2(n12806), .ZN(n12820) );
  INV_X1 U15936 ( .A(n12812), .ZN(n12807) );
  NAND2_X1 U15937 ( .A1(n12808), .A2(n12807), .ZN(n12810) );
  AOI21_X1 U15938 ( .B1(n12811), .B2(n12815), .A(n9635), .ZN(n12809) );
  NAND2_X1 U15939 ( .A1(n12810), .A2(n12809), .ZN(n12817) );
  INV_X1 U15940 ( .A(n12811), .ZN(n12814) );
  OAI211_X1 U15941 ( .C1(n12815), .C2(n12814), .A(n12807), .B(n12813), .ZN(
        n12816) );
  MUX2_X1 U15942 ( .A(n12817), .B(n12816), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n12818) );
  INV_X1 U15943 ( .A(n12818), .ZN(n12819) );
  NAND2_X1 U15944 ( .A1(n12820), .A2(n12819), .ZN(n19519) );
  INV_X1 U15945 ( .A(n13169), .ZN(n12821) );
  OR2_X1 U15946 ( .A1(n19519), .A2(n12821), .ZN(n12823) );
  OR2_X1 U15947 ( .A1(n13169), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12822) );
  NAND2_X1 U15948 ( .A1(n12823), .A2(n12822), .ZN(n12826) );
  NAND2_X1 U15949 ( .A1(n12826), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12824) );
  NAND2_X1 U15950 ( .A1(n12825), .A2(n12824), .ZN(n12830) );
  INV_X1 U15951 ( .A(n12826), .ZN(n12853) );
  NAND2_X1 U15952 ( .A1(n12853), .A2(n12827), .ZN(n12829) );
  NAND3_X1 U15953 ( .A1(n12852), .A2(n12827), .A3(n19550), .ZN(n12828) );
  NAND3_X1 U15954 ( .A1(n12830), .A2(n12829), .A3(n12828), .ZN(n12831) );
  NAND2_X1 U15955 ( .A1(n12831), .A2(n15419), .ZN(n12855) );
  NAND2_X1 U15956 ( .A1(n12833), .A2(n12832), .ZN(n12837) );
  INV_X1 U15957 ( .A(n12834), .ZN(n12835) );
  NAND2_X1 U15958 ( .A1(n12839), .A2(n12835), .ZN(n12836) );
  OAI211_X1 U15959 ( .C1(n12839), .C2(n12838), .A(n12837), .B(n12836), .ZN(
        n19577) );
  NAND2_X1 U15960 ( .A1(n12841), .A2(n12840), .ZN(n12842) );
  NOR2_X1 U15961 ( .A1(n12843), .A2(n12842), .ZN(n18417) );
  OAI21_X1 U15962 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n18417), .ZN(n12847) );
  NAND2_X1 U15963 ( .A1(n18895), .A2(n12844), .ZN(n12845) );
  OR2_X1 U15964 ( .A1(n12846), .A2(n12845), .ZN(n15190) );
  OAI211_X1 U15965 ( .C1(n9634), .C2(n12848), .A(n12847), .B(n15190), .ZN(
        n12849) );
  NOR2_X1 U15966 ( .A1(n19577), .A2(n12849), .ZN(n12850) );
  OAI21_X1 U15967 ( .B1(n13169), .B2(n15192), .A(n12850), .ZN(n12851) );
  AOI21_X1 U15968 ( .B1(n12853), .B2(n12852), .A(n12851), .ZN(n12854) );
  NAND2_X1 U15969 ( .A1(n12855), .A2(n12854), .ZN(n15909) );
  OAI21_X1 U15970 ( .B1(n15909), .B2(P2_STATE2_REG_1__SCAN_IN), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n12862) );
  INV_X1 U15971 ( .A(n12856), .ZN(n12860) );
  AND2_X1 U15972 ( .A1(n12857), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19591) );
  INV_X1 U15973 ( .A(n19591), .ZN(n12858) );
  AOI21_X1 U15974 ( .B1(n12860), .B2(n12859), .A(n12858), .ZN(n12861) );
  AND2_X1 U15975 ( .A1(n12862), .A2(n12861), .ZN(n15910) );
  OAI21_X1 U15976 ( .B1(n15910), .B2(n15904), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12864) );
  NAND2_X1 U15977 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n12863), .ZN(n15906) );
  NAND2_X1 U15978 ( .A1(n12864), .A2(n15906), .ZN(P2_U3593) );
  AOI22_X1 U15979 ( .A1(n14634), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n14633), .ZN(n18896) );
  XNOR2_X1 U15980 ( .A(n12866), .B(n12865), .ZN(n13111) );
  XNOR2_X1 U15981 ( .A(n19538), .B(n13111), .ZN(n12867) );
  INV_X1 U15982 ( .A(n14443), .ZN(n18695) );
  NAND2_X1 U15983 ( .A1(n19128), .A2(n18695), .ZN(n18693) );
  NAND2_X1 U15984 ( .A1(n12867), .A2(n18693), .ZN(n12982) );
  OAI21_X1 U15985 ( .B1(n12867), .B2(n18693), .A(n12982), .ZN(n12868) );
  NAND2_X1 U15986 ( .A1(n12868), .A2(n18694), .ZN(n12870) );
  INV_X1 U15987 ( .A(n13111), .ZN(n19553) );
  AOI22_X1 U15988 ( .A1(n18692), .A2(n19553), .B1(n18691), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n12869) );
  OAI211_X1 U15989 ( .C1(n18896), .C2(n18698), .A(n12870), .B(n12869), .ZN(
        P2_U2918) );
  OAI21_X1 U15990 ( .B1(n12873), .B2(n12872), .A(n12871), .ZN(n13070) );
  NOR2_X1 U15991 ( .A1(n12875), .A2(n12874), .ZN(n19821) );
  INV_X1 U15992 ( .A(n19821), .ZN(n12876) );
  INV_X1 U15993 ( .A(n12877), .ZN(n13064) );
  INV_X1 U15994 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12878) );
  INV_X1 U15995 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n13058) );
  OAI22_X1 U15996 ( .A1(n14190), .A2(n12878), .B1(n19798), .B2(n13058), .ZN(
        n12879) );
  AOI21_X1 U15997 ( .B1(n13064), .B2(n15566), .A(n12879), .ZN(n12880) );
  OAI211_X1 U15998 ( .C1(n19835), .C2(n13070), .A(n12881), .B(n12880), .ZN(
        P1_U2997) );
  INV_X1 U15999 ( .A(n13555), .ZN(n12882) );
  AOI21_X1 U16000 ( .B1(n13554), .B2(n12883), .A(n12882), .ZN(n12891) );
  NAND2_X1 U16001 ( .A1(n19795), .A2(n19824), .ZN(n15652) );
  INV_X1 U16002 ( .A(n15652), .ZN(n14383) );
  NOR3_X1 U16003 ( .A1(n14383), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n13559), .ZN(n12884) );
  AOI211_X1 U16004 ( .C1(n12886), .C2(n19807), .A(n12885), .B(n12884), .ZN(
        n12890) );
  NAND3_X1 U16005 ( .A1(n19810), .A2(n12888), .A3(n12887), .ZN(n12889) );
  OAI211_X1 U16006 ( .C1(n12891), .C2(n19819), .A(n12890), .B(n12889), .ZN(
        P1_U3030) );
  AOI22_X1 U16007 ( .A1(n19705), .A2(n13105), .B1(P1_EBX_REG_0__SCAN_IN), .B2(
        n14004), .ZN(n12892) );
  OAI21_X1 U16008 ( .B1(n14024), .B2(n19715), .A(n12892), .ZN(P1_U2872) );
  NAND2_X1 U16009 ( .A1(n12894), .A2(n12893), .ZN(n12895) );
  NAND2_X1 U16010 ( .A1(n12993), .A2(n12895), .ZN(n19822) );
  OAI22_X1 U16011 ( .A1(n14025), .A2(n19822), .B1(n12896), .B2(n19710), .ZN(
        n12897) );
  INV_X1 U16012 ( .A(n12897), .ZN(n12898) );
  OAI21_X1 U16013 ( .B1(n13070), .B2(n14024), .A(n12898), .ZN(P1_U2870) );
  NAND2_X1 U16014 ( .A1(n12899), .A2(n19886), .ZN(n12900) );
  NAND2_X2 U16015 ( .A1(n19713), .A2(n12900), .ZN(n19714) );
  INV_X1 U16016 ( .A(n12900), .ZN(n12901) );
  MUX2_X1 U16017 ( .A(DATAI_2_), .B(BUF1_REG_2__SCAN_IN), .S(n19836), .Z(
        n19860) );
  INV_X1 U16018 ( .A(n19860), .ZN(n12902) );
  INV_X1 U16019 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n19742) );
  OAI222_X1 U16020 ( .A1(n13070), .A2(n19714), .B1(n19712), .B2(n12902), .C1(
        n19713), .C2(n19742), .ZN(P1_U2902) );
  NAND2_X1 U16021 ( .A1(n12903), .A2(n12944), .ZN(n12905) );
  INV_X1 U16022 ( .A(n12966), .ZN(n12904) );
  AND2_X1 U16023 ( .A1(n12905), .A2(n12904), .ZN(n18573) );
  INV_X1 U16024 ( .A(n18573), .ZN(n15066) );
  OAI211_X1 U16025 ( .C1(n12906), .C2(n12907), .A(n12964), .B(n14522), .ZN(
        n12909) );
  NAND2_X1 U16026 ( .A1(n14548), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12908) );
  OAI211_X1 U16027 ( .C1(n15066), .C2(n14548), .A(n12909), .B(n12908), .ZN(
        P2_U2878) );
  INV_X1 U16028 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n18747) );
  AOI22_X1 U16029 ( .A1(n14634), .A2(BUF1_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n14610), .ZN(n18798) );
  OAI21_X1 U16030 ( .B1(n12911), .B2(n12910), .A(n15870), .ZN(n18539) );
  OAI222_X1 U16031 ( .A1(n18686), .A2(n18747), .B1(n18798), .B2(n18698), .C1(
        n18539), .C2(n18675), .ZN(P2_U2908) );
  NOR2_X1 U16032 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n20445), .ZN(n12932) );
  MUX2_X1 U16033 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n12912), .S(
        n15374), .Z(n15378) );
  AOI22_X1 U16034 ( .A1(n12932), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15378), .B2(n20445), .ZN(n12929) );
  XNOR2_X1 U16035 ( .A(n12913), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12924) );
  INV_X1 U16036 ( .A(n12915), .ZN(n12916) );
  OAI211_X1 U16037 ( .C1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C2(n14427), .A(
        n10553), .B(n12916), .ZN(n14434) );
  OR3_X1 U16038 ( .A1(n14425), .A2(n12917), .A3(n14434), .ZN(n12923) );
  MUX2_X1 U16039 ( .A(n12918), .B(n12926), .S(n14427), .Z(n12920) );
  OAI21_X1 U16040 ( .B1(n12921), .B2(n12920), .A(n12919), .ZN(n12922) );
  OAI211_X1 U16041 ( .C1(n14421), .C2(n12924), .A(n12923), .B(n12922), .ZN(
        n12925) );
  AOI21_X1 U16042 ( .B1(n20517), .B2(n14425), .A(n12925), .ZN(n14436) );
  MUX2_X1 U16043 ( .A(n12926), .B(n14436), .S(n15374), .Z(n15380) );
  INV_X1 U16044 ( .A(n15380), .ZN(n12927) );
  AOI22_X1 U16045 ( .A1(n12932), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n20445), .B2(n12927), .ZN(n12928) );
  NOR2_X1 U16046 ( .A1(n12929), .A2(n12928), .ZN(n15389) );
  INV_X1 U16047 ( .A(n14428), .ZN(n12930) );
  NAND2_X1 U16048 ( .A1(n15389), .A2(n12930), .ZN(n14417) );
  OAI21_X1 U16049 ( .B1(n11247), .B2(n19680), .A(n15374), .ZN(n12931) );
  OAI211_X1 U16050 ( .C1(n15374), .C2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n12931), .B(n20445), .ZN(n12934) );
  NAND2_X1 U16051 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n12932), .ZN(
        n12933) );
  AND2_X1 U16052 ( .A1(n12934), .A2(n12933), .ZN(n15385) );
  NAND3_X1 U16053 ( .A1(n14417), .A2(n15385), .A3(n19609), .ZN(n12936) );
  INV_X1 U16054 ( .A(n15688), .ZN(n12935) );
  NAND2_X1 U16055 ( .A1(n12936), .A2(n12935), .ZN(n12937) );
  NAND2_X1 U16056 ( .A1(n12937), .A2(n19897), .ZN(n20526) );
  NAND2_X1 U16057 ( .A1(n20270), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14418) );
  INV_X1 U16058 ( .A(n14418), .ZN(n20518) );
  NOR2_X1 U16059 ( .A1(n20259), .A2(n20518), .ZN(n12942) );
  AND2_X1 U16060 ( .A1(n9631), .A2(n12939), .ZN(n20387) );
  OR2_X1 U16061 ( .A1(n9631), .A2(n20516), .ZN(n12940) );
  NAND2_X1 U16062 ( .A1(n20316), .A2(n20347), .ZN(n20256) );
  NAND2_X1 U16063 ( .A1(n12940), .A2(n20256), .ZN(n20216) );
  OAI21_X1 U16064 ( .B1(n12942), .B2(n12941), .A(n20526), .ZN(n12943) );
  OAI21_X1 U16065 ( .B1(n20526), .B2(n20262), .A(n12943), .ZN(P1_U3476) );
  OAI21_X1 U16066 ( .B1(n12946), .B2(n12945), .A(n12944), .ZN(n18588) );
  INV_X1 U16067 ( .A(n18588), .ZN(n15890) );
  INV_X1 U16068 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n18578) );
  NOR2_X1 U16069 ( .A1(n14540), .A2(n18578), .ZN(n12949) );
  AOI211_X1 U16070 ( .C1(n12947), .C2(n12766), .A(n14550), .B(n12906), .ZN(
        n12948) );
  AOI211_X1 U16071 ( .C1(n15890), .C2(n14525), .A(n12949), .B(n12948), .ZN(
        n12950) );
  INV_X1 U16072 ( .A(n12950), .ZN(P2_U2879) );
  INV_X1 U16073 ( .A(n20526), .ZN(n20529) );
  INV_X1 U16074 ( .A(n9631), .ZN(n12951) );
  NAND2_X1 U16075 ( .A1(n12951), .A2(n20347), .ZN(n12953) );
  INV_X1 U16076 ( .A(n12952), .ZN(n20349) );
  AOI22_X1 U16077 ( .A1(n20216), .A2(n12953), .B1(n20349), .B2(n14418), .ZN(
        n12955) );
  NAND2_X1 U16078 ( .A1(n20529), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12954) );
  OAI21_X1 U16079 ( .B1(n20529), .B2(n12955), .A(n12954), .ZN(P1_U3477) );
  MUX2_X1 U16080 ( .A(DATAI_1_), .B(BUF1_REG_1__SCAN_IN), .S(n19836), .Z(
        n19855) );
  INV_X1 U16081 ( .A(n19855), .ZN(n12956) );
  INV_X1 U16082 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n19744) );
  OAI222_X1 U16083 ( .A1(n13090), .A2(n19714), .B1(n19712), .B2(n12956), .C1(
        n19713), .C2(n19744), .ZN(P1_U2903) );
  AOI22_X1 U16084 ( .A1(n19774), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n19773), .ZN(n12960) );
  MUX2_X1 U16085 ( .A(DATAI_7_), .B(BUF1_REG_7__SCAN_IN), .S(n19836), .Z(
        n19889) );
  NAND2_X1 U16086 ( .A1(n19763), .A2(n19889), .ZN(n13137) );
  NAND2_X1 U16087 ( .A1(n12960), .A2(n13137), .ZN(P1_U2959) );
  AOI22_X1 U16088 ( .A1(n19774), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n19773), .ZN(n12961) );
  MUX2_X1 U16089 ( .A(DATAI_5_), .B(BUF1_REG_5__SCAN_IN), .S(n19836), .Z(
        n19875) );
  NAND2_X1 U16090 ( .A1(n19763), .A2(n19875), .ZN(n13141) );
  NAND2_X1 U16091 ( .A1(n12961), .A2(n13141), .ZN(P1_U2957) );
  AOI22_X1 U16092 ( .A1(n19774), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n19773), .ZN(n12962) );
  MUX2_X1 U16093 ( .A(DATAI_6_), .B(BUF1_REG_6__SCAN_IN), .S(n19836), .Z(
        n19880) );
  NAND2_X1 U16094 ( .A1(n19763), .A2(n19880), .ZN(n13139) );
  NAND2_X1 U16095 ( .A1(n12962), .A2(n13139), .ZN(P1_U2958) );
  AOI22_X1 U16096 ( .A1(n19774), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n19773), .ZN(n12963) );
  MUX2_X1 U16097 ( .A(DATAI_4_), .B(BUF1_REG_4__SCAN_IN), .S(n19836), .Z(
        n19870) );
  NAND2_X1 U16098 ( .A1(n19763), .A2(n19870), .ZN(n13143) );
  NAND2_X1 U16099 ( .A1(n12963), .A2(n13143), .ZN(P1_U2956) );
  OAI211_X1 U16100 ( .C1(n11504), .C2(n11503), .A(n14522), .B(n13030), .ZN(
        n12970) );
  OR2_X1 U16101 ( .A1(n12967), .A2(n12966), .ZN(n12968) );
  AND2_X1 U16102 ( .A1(n12968), .A2(n13026), .ZN(n18562) );
  NAND2_X1 U16103 ( .A1(n14540), .A2(n18562), .ZN(n12969) );
  OAI211_X1 U16104 ( .C1(n14525), .C2(n10071), .A(n12970), .B(n12969), .ZN(
        P2_U2877) );
  NAND2_X1 U16105 ( .A1(n12972), .A2(n12971), .ZN(n12973) );
  AND2_X1 U16106 ( .A1(n13006), .A2(n12973), .ZN(n19786) );
  INV_X1 U16107 ( .A(n19786), .ZN(n12977) );
  INV_X1 U16108 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n12975) );
  OAI21_X1 U16109 ( .B1(n12991), .B2(n12974), .A(n13009), .ZN(n19799) );
  OAI222_X1 U16110 ( .A1(n12977), .A2(n14024), .B1(n19710), .B2(n12975), .C1(
        n19799), .C2(n14025), .ZN(P1_U2868) );
  INV_X1 U16111 ( .A(n19870), .ZN(n12976) );
  INV_X1 U16112 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n19738) );
  OAI222_X1 U16113 ( .A1(n12977), .A2(n19714), .B1(n19712), .B2(n12976), .C1(
        n19713), .C2(n19738), .ZN(P1_U2900) );
  NAND2_X1 U16114 ( .A1(n12979), .A2(n12978), .ZN(n12981) );
  AND2_X1 U16115 ( .A1(n12981), .A2(n10181), .ZN(n18863) );
  XOR2_X1 U16116 ( .A(n18863), .B(n19546), .Z(n12985) );
  NAND2_X1 U16117 ( .A1(n19557), .A2(n13111), .ZN(n12983) );
  NAND2_X1 U16118 ( .A1(n12983), .A2(n12982), .ZN(n12984) );
  NAND2_X1 U16119 ( .A1(n12985), .A2(n12984), .ZN(n18668) );
  OAI21_X1 U16120 ( .B1(n12985), .B2(n12984), .A(n18668), .ZN(n12986) );
  NAND2_X1 U16121 ( .A1(n12986), .A2(n18694), .ZN(n12988) );
  INV_X1 U16122 ( .A(n18698), .ZN(n18667) );
  AOI22_X1 U16123 ( .A1(n14634), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n14633), .ZN(n18901) );
  INV_X1 U16124 ( .A(n18901), .ZN(n13425) );
  AOI22_X1 U16125 ( .A1(n18667), .A2(n13425), .B1(n18691), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n12987) );
  OAI211_X1 U16126 ( .C1(n18863), .C2(n18687), .A(n12988), .B(n12987), .ZN(
        P2_U2917) );
  XOR2_X1 U16127 ( .A(n12990), .B(n12989), .Z(n19700) );
  INV_X1 U16128 ( .A(n19700), .ZN(n13003) );
  AOI21_X1 U16129 ( .B1(n12993), .B2(n12992), .A(n12991), .ZN(n19806) );
  AOI22_X1 U16130 ( .A1(n19705), .A2(n19806), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n14004), .ZN(n12994) );
  OAI21_X1 U16131 ( .B1(n13003), .B2(n14024), .A(n12994), .ZN(P1_U2869) );
  OAI21_X1 U16132 ( .B1(n12997), .B2(n12996), .A(n12995), .ZN(n19808) );
  INV_X1 U16133 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n12998) );
  NOR2_X1 U16134 ( .A1(n19798), .A2(n12998), .ZN(n19805) );
  AOI21_X1 U16135 ( .B1(n19782), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n19805), .ZN(n12999) );
  OAI21_X1 U16136 ( .B1(n19793), .B2(n19689), .A(n12999), .ZN(n13000) );
  AOI21_X1 U16137 ( .B1(n19700), .B2(n19787), .A(n13000), .ZN(n13001) );
  OAI21_X1 U16138 ( .B1(n19808), .B2(n19608), .A(n13001), .ZN(P1_U2996) );
  MUX2_X1 U16139 ( .A(DATAI_3_), .B(BUF1_REG_3__SCAN_IN), .S(n19836), .Z(
        n19865) );
  INV_X1 U16140 ( .A(n19865), .ZN(n13002) );
  INV_X1 U16141 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n19740) );
  OAI222_X1 U16142 ( .A1(n13003), .A2(n19714), .B1(n19712), .B2(n13002), .C1(
        n19713), .C2(n19740), .ZN(P1_U2901) );
  OAI21_X1 U16143 ( .B1(n13004), .B2(n15868), .A(n15855), .ZN(n18528) );
  AOI22_X1 U16144 ( .A1(n14634), .A2(BUF1_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n14610), .ZN(n18800) );
  INV_X1 U16145 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n18743) );
  OAI222_X1 U16146 ( .A1(n18528), .A2(n18675), .B1(n18800), .B2(n18698), .C1(
        n18743), .C2(n18686), .ZN(P2_U2906) );
  AND2_X1 U16147 ( .A1(n13006), .A2(n13005), .ZN(n13007) );
  OR2_X1 U16148 ( .A1(n13044), .A2(n13007), .ZN(n15595) );
  INV_X1 U16149 ( .A(n15669), .ZN(n13008) );
  AOI21_X1 U16150 ( .B1(n13010), .B2(n13009), .A(n13008), .ZN(n19663) );
  AOI22_X1 U16151 ( .A1(n19705), .A2(n19663), .B1(P1_EBX_REG_5__SCAN_IN), .B2(
        n14004), .ZN(n13011) );
  OAI21_X1 U16152 ( .B1(n15595), .B2(n14024), .A(n13011), .ZN(P1_U2867) );
  INV_X1 U16153 ( .A(n19875), .ZN(n13012) );
  OAI222_X1 U16154 ( .A1(n15595), .A2(n19714), .B1(n19712), .B2(n13012), .C1(
        n19713), .C2(n10616), .ZN(P1_U2899) );
  NAND2_X1 U16155 ( .A1(n15696), .A2(n13013), .ZN(n13014) );
  XNOR2_X1 U16156 ( .A(n15844), .B(n13014), .ZN(n13024) );
  OAI21_X1 U16157 ( .B1(n13016), .B2(n13015), .A(n13340), .ZN(n13332) );
  OAI22_X1 U16158 ( .A1(n12102), .A2(n18601), .B1(n13332), .B2(n18616), .ZN(
        n13020) );
  XNOR2_X1 U16159 ( .A(n13018), .B(n13017), .ZN(n19534) );
  OAI22_X1 U16160 ( .A1(n15853), .A2(n18540), .B1(n18628), .B2(n19534), .ZN(
        n13019) );
  AOI211_X1 U16161 ( .C1(P2_EBX_REG_3__SCAN_IN), .C2(n18614), .A(n13020), .B(
        n13019), .ZN(n13022) );
  NAND2_X1 U16162 ( .A1(n15895), .A2(n18625), .ZN(n13021) );
  OAI211_X1 U16163 ( .C1(n19540), .C2(n18644), .A(n13022), .B(n13021), .ZN(
        n13023) );
  AOI21_X1 U16164 ( .B1(n13024), .B2(n18623), .A(n13023), .ZN(n13025) );
  INV_X1 U16165 ( .A(n13025), .ZN(P2_U2852) );
  NAND2_X1 U16166 ( .A1(n13027), .A2(n13026), .ZN(n13029) );
  INV_X1 U16167 ( .A(n13037), .ZN(n13028) );
  AND2_X1 U16168 ( .A1(n13029), .A2(n13028), .ZN(n18545) );
  INV_X1 U16169 ( .A(n18545), .ZN(n15033) );
  NOR2_X1 U16170 ( .A1(n14548), .A2(n15033), .ZN(n13033) );
  AOI211_X1 U16171 ( .C1(n13031), .C2(n13030), .A(n14550), .B(n9647), .ZN(
        n13032) );
  AOI211_X1 U16172 ( .C1(P2_EBX_REG_11__SCAN_IN), .C2(n14548), .A(n13033), .B(
        n13032), .ZN(n13034) );
  INV_X1 U16173 ( .A(n13034), .ZN(P2_U2876) );
  OAI211_X1 U16174 ( .C1(n9647), .C2(n13036), .A(n10154), .B(n14522), .ZN(
        n13041) );
  OR2_X1 U16175 ( .A1(n13038), .A2(n13037), .ZN(n13039) );
  NAND2_X1 U16176 ( .A1(n13039), .A2(n13049), .ZN(n18538) );
  INV_X1 U16177 ( .A(n18538), .ZN(n15805) );
  NAND2_X1 U16178 ( .A1(n14540), .A2(n15805), .ZN(n13040) );
  OAI211_X1 U16179 ( .C1(n14525), .C2(n11900), .A(n13041), .B(n13040), .ZN(
        P2_U2875) );
  OR2_X1 U16180 ( .A1(n13044), .A2(n13043), .ZN(n13045) );
  AND2_X1 U16181 ( .A1(n13042), .A2(n13045), .ZN(n19707) );
  INV_X1 U16182 ( .A(n19707), .ZN(n13047) );
  INV_X1 U16183 ( .A(n19880), .ZN(n13046) );
  INV_X1 U16184 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n19734) );
  OAI222_X1 U16185 ( .A1(n13047), .A2(n19714), .B1(n19712), .B2(n13046), .C1(
        n19713), .C2(n19734), .ZN(P1_U2898) );
  INV_X1 U16186 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n18739) );
  OAI21_X1 U16187 ( .B1(n15854), .B2(n13048), .A(n9728), .ZN(n18506) );
  AOI22_X1 U16188 ( .A1(n14634), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n14610), .ZN(n18805) );
  OAI222_X1 U16189 ( .A1(n18686), .A2(n18739), .B1(n18506), .B2(n18675), .C1(
        n18698), .C2(n18805), .ZN(P2_U2904) );
  NAND2_X1 U16190 ( .A1(n13050), .A2(n13049), .ZN(n13052) );
  INV_X1 U16191 ( .A(n13119), .ZN(n13051) );
  AND2_X1 U16192 ( .A1(n13052), .A2(n13051), .ZN(n18525) );
  INV_X1 U16193 ( .A(n18525), .ZN(n15016) );
  OAI211_X1 U16194 ( .C1(n13035), .C2(n13053), .A(n13117), .B(n14522), .ZN(
        n13055) );
  NAND2_X1 U16195 ( .A1(n14548), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n13054) );
  OAI211_X1 U16196 ( .C1(n15016), .C2(n14548), .A(n13055), .B(n13054), .ZN(
        P2_U2874) );
  NAND2_X1 U16197 ( .A1(n13063), .A2(n13056), .ZN(n13057) );
  NAND2_X1 U16198 ( .A1(n15470), .A2(n13057), .ZN(n19699) );
  INV_X1 U16199 ( .A(n19699), .ZN(n13091) );
  INV_X1 U16200 ( .A(n13963), .ZN(n15450) );
  NAND2_X1 U16201 ( .A1(n15450), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n19696) );
  INV_X1 U16202 ( .A(n19696), .ZN(n13059) );
  NAND2_X1 U16203 ( .A1(n13059), .A2(n13058), .ZN(n13068) );
  OAI21_X1 U16204 ( .B1(n15449), .B2(n13060), .A(n19636), .ZN(n19703) );
  OAI22_X1 U16205 ( .A1(n19703), .A2(n13058), .B1(n19681), .B2(n19822), .ZN(
        n13061) );
  AOI21_X1 U16206 ( .B1(n19675), .B2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n13061), .ZN(n13067) );
  INV_X1 U16207 ( .A(n20259), .ZN(n19842) );
  NAND2_X1 U16208 ( .A1(n13063), .A2(n13062), .ZN(n19679) );
  INV_X1 U16209 ( .A(n19679), .ZN(n19694) );
  AOI22_X1 U16210 ( .A1(n19842), .A2(n19694), .B1(n19687), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n13066) );
  NAND2_X1 U16211 ( .A1(n19644), .A2(n13064), .ZN(n13065) );
  AND4_X1 U16212 ( .A1(n13068), .A2(n13067), .A3(n13066), .A4(n13065), .ZN(
        n13069) );
  OAI21_X1 U16213 ( .B1(n13091), .B2(n13070), .A(n13069), .ZN(P1_U2838) );
  NOR2_X1 U16214 ( .A1(n18630), .A2(n13109), .ZN(n13071) );
  XNOR2_X1 U16215 ( .A(n13071), .B(n18826), .ZN(n13072) );
  NAND2_X1 U16216 ( .A1(n13072), .A2(n18623), .ZN(n13081) );
  XNOR2_X1 U16217 ( .A(n13074), .B(n13073), .ZN(n13337) );
  INV_X1 U16218 ( .A(n13337), .ZN(n13338) );
  OAI22_X1 U16219 ( .A1(n18642), .A2(n11427), .B1(n18863), .B2(n18628), .ZN(
        n13075) );
  AOI21_X1 U16220 ( .B1(n18637), .B2(n13338), .A(n13075), .ZN(n13076) );
  INV_X1 U16221 ( .A(n13076), .ZN(n13079) );
  AOI22_X1 U16222 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n18639), .B1(
        P2_REIP_REG_2__SCAN_IN), .B2(n9772), .ZN(n13077) );
  INV_X1 U16223 ( .A(n13077), .ZN(n13078) );
  AOI211_X1 U16224 ( .C1(n18625), .C2(n13260), .A(n13079), .B(n13078), .ZN(
        n13080) );
  OAI211_X1 U16225 ( .C1(n19546), .C2(n18644), .A(n13081), .B(n13080), .ZN(
        P2_U2853) );
  AOI22_X1 U16226 ( .A1(P1_EBX_REG_1__SCAN_IN), .A2(n19687), .B1(n15449), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n13089) );
  NOR2_X1 U16227 ( .A1(n19679), .A2(n12952), .ZN(n13086) );
  NAND2_X1 U16228 ( .A1(n19675), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13084) );
  NAND2_X1 U16229 ( .A1(n19644), .A2(n13082), .ZN(n13083) );
  OAI211_X1 U16230 ( .C1(n13963), .C2(P1_REIP_REG_1__SCAN_IN), .A(n13084), .B(
        n13083), .ZN(n13085) );
  AOI211_X1 U16231 ( .C1(n19686), .C2(n13087), .A(n13086), .B(n13085), .ZN(
        n13088) );
  OAI211_X1 U16232 ( .C1(n13091), .C2(n13090), .A(n13089), .B(n13088), .ZN(
        P1_U2839) );
  NAND2_X1 U16233 ( .A1(n13042), .A2(n13092), .ZN(n13093) );
  AND2_X1 U16234 ( .A1(n13146), .A2(n13093), .ZN(n19638) );
  INV_X1 U16235 ( .A(n19638), .ZN(n13095) );
  INV_X1 U16236 ( .A(n19889), .ZN(n13094) );
  OAI222_X1 U16237 ( .A1(n13095), .A2(n19714), .B1(n19712), .B2(n13094), .C1(
        n19713), .C2(n10647), .ZN(P1_U2897) );
  NOR2_X1 U16238 ( .A1(n13097), .A2(n13096), .ZN(n13098) );
  OR2_X1 U16239 ( .A1(n13149), .A2(n13098), .ZN(n19639) );
  OAI22_X1 U16240 ( .A1(n14025), .A2(n19639), .B1(n19640), .B2(n19710), .ZN(
        n13099) );
  AOI21_X1 U16241 ( .B1(n19638), .B2(n19706), .A(n13099), .ZN(n13100) );
  INV_X1 U16242 ( .A(n13100), .ZN(P1_U2865) );
  INV_X1 U16243 ( .A(n19715), .ZN(n13104) );
  INV_X1 U16244 ( .A(n19961), .ZN(n13102) );
  OAI21_X1 U16245 ( .B1(n19675), .B2(n19644), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13101) );
  OAI21_X1 U16246 ( .B1(n19679), .B2(n13102), .A(n13101), .ZN(n13103) );
  AOI21_X1 U16247 ( .B1(n13104), .B2(n19699), .A(n13103), .ZN(n13107) );
  AOI22_X1 U16248 ( .A1(P1_EBX_REG_0__SCAN_IN), .A2(n19687), .B1(n19686), .B2(
        n13105), .ZN(n13106) );
  OAI211_X1 U16249 ( .C1(n19669), .C2(n13108), .A(n13107), .B(n13106), .ZN(
        P1_U2840) );
  AOI211_X1 U16250 ( .C1(n14446), .C2(n13110), .A(n18630), .B(n13109), .ZN(
        n13163) );
  NOR2_X1 U16251 ( .A1(n19437), .A2(n15696), .ZN(n18544) );
  AOI22_X1 U16252 ( .A1(n13163), .A2(n18623), .B1(n18544), .B2(n12475), .ZN(
        n13116) );
  OAI22_X1 U16253 ( .A1(n18628), .A2(n13111), .B1(n18616), .B2(n13333), .ZN(
        n13114) );
  AOI22_X1 U16254 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18639), .B1(
        P2_REIP_REG_1__SCAN_IN), .B2(n9772), .ZN(n13112) );
  OAI21_X1 U16255 ( .B1(n18642), .B2(n11412), .A(n13112), .ZN(n13113) );
  AOI211_X1 U16256 ( .C1(n13263), .C2(n18625), .A(n13114), .B(n13113), .ZN(
        n13115) );
  OAI211_X1 U16257 ( .C1(n19557), .C2(n18644), .A(n13116), .B(n13115), .ZN(
        P2_U2854) );
  OAI211_X1 U16258 ( .C1(n11551), .C2(n11550), .A(n14522), .B(n13178), .ZN(
        n13122) );
  OAI21_X1 U16259 ( .B1(n13120), .B2(n13119), .A(n13176), .ZN(n18516) );
  INV_X1 U16260 ( .A(n18516), .ZN(n15858) );
  NAND2_X1 U16261 ( .A1(n14540), .A2(n15858), .ZN(n13121) );
  OAI211_X1 U16262 ( .C1(n14525), .C2(n11860), .A(n13122), .B(n13121), .ZN(
        P2_U2873) );
  AOI22_X1 U16263 ( .A1(n19774), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n19773), .ZN(n13123) );
  NAND2_X1 U16264 ( .A1(n19763), .A2(n19860), .ZN(n13124) );
  NAND2_X1 U16265 ( .A1(n13123), .A2(n13124), .ZN(P1_U2954) );
  AOI22_X1 U16266 ( .A1(n19774), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n19773), .ZN(n13125) );
  NAND2_X1 U16267 ( .A1(n13125), .A2(n13124), .ZN(P1_U2939) );
  AOI22_X1 U16268 ( .A1(n19774), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n19773), .ZN(n13126) );
  NAND2_X1 U16269 ( .A1(n19763), .A2(n19865), .ZN(n13127) );
  NAND2_X1 U16270 ( .A1(n13126), .A2(n13127), .ZN(P1_U2955) );
  AOI22_X1 U16271 ( .A1(n19774), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n19773), .ZN(n13128) );
  NAND2_X1 U16272 ( .A1(n13128), .A2(n13127), .ZN(P1_U2940) );
  AOI22_X1 U16273 ( .A1(n19774), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n19773), .ZN(n13131) );
  INV_X1 U16274 ( .A(DATAI_0_), .ZN(n13130) );
  NAND2_X1 U16275 ( .A1(n19836), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13129) );
  OAI21_X1 U16276 ( .B1(n19836), .B2(n13130), .A(n13129), .ZN(n19846) );
  NAND2_X1 U16277 ( .A1(n19763), .A2(n19846), .ZN(n13135) );
  NAND2_X1 U16278 ( .A1(n13131), .A2(n13135), .ZN(P1_U2952) );
  AOI22_X1 U16279 ( .A1(n19774), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n19773), .ZN(n13132) );
  NAND2_X1 U16280 ( .A1(n19763), .A2(n19855), .ZN(n13133) );
  NAND2_X1 U16281 ( .A1(n13132), .A2(n13133), .ZN(P1_U2953) );
  AOI22_X1 U16282 ( .A1(n19774), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n19773), .ZN(n13134) );
  NAND2_X1 U16283 ( .A1(n13134), .A2(n13133), .ZN(P1_U2938) );
  AOI22_X1 U16284 ( .A1(n19774), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n19773), .ZN(n13136) );
  NAND2_X1 U16285 ( .A1(n13136), .A2(n13135), .ZN(P1_U2937) );
  AOI22_X1 U16286 ( .A1(n19774), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n19773), .ZN(n13138) );
  NAND2_X1 U16287 ( .A1(n13138), .A2(n13137), .ZN(P1_U2944) );
  AOI22_X1 U16288 ( .A1(n19774), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n19773), .ZN(n13140) );
  NAND2_X1 U16289 ( .A1(n13140), .A2(n13139), .ZN(P1_U2943) );
  AOI22_X1 U16290 ( .A1(n19774), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n19773), .ZN(n13142) );
  NAND2_X1 U16291 ( .A1(n13142), .A2(n13141), .ZN(P1_U2942) );
  AOI22_X1 U16292 ( .A1(n19774), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n19773), .ZN(n13144) );
  NAND2_X1 U16293 ( .A1(n13144), .A2(n13143), .ZN(P1_U2941) );
  AOI21_X1 U16294 ( .B1(n13147), .B2(n13146), .A(n13145), .ZN(n13219) );
  OR2_X1 U16295 ( .A1(n13149), .A2(n13148), .ZN(n13150) );
  NAND2_X1 U16296 ( .A1(n13183), .A2(n13150), .ZN(n15656) );
  OAI22_X1 U16297 ( .A1(n14025), .A2(n15656), .B1(n13154), .B2(n19710), .ZN(
        n13151) );
  AOI21_X1 U16298 ( .B1(n13219), .B2(n19706), .A(n13151), .ZN(n13152) );
  INV_X1 U16299 ( .A(n13152), .ZN(P1_U2864) );
  INV_X1 U16300 ( .A(n13219), .ZN(n13162) );
  INV_X1 U16301 ( .A(n13217), .ZN(n13159) );
  NOR2_X1 U16302 ( .A1(n13963), .A2(n13153), .ZN(n19651) );
  NAND4_X1 U16303 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .A4(n19651), .ZN(n13157) );
  INV_X1 U16304 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n15655) );
  OR2_X1 U16305 ( .A1(n13153), .A2(n15449), .ZN(n19667) );
  OAI21_X1 U16306 ( .B1(n19625), .B2(n19667), .A(n19636), .ZN(n19628) );
  NAND2_X1 U16307 ( .A1(n13961), .A2(n19600), .ZN(n19653) );
  OAI22_X1 U16308 ( .A1(n13154), .A2(n19662), .B1(n19681), .B2(n15656), .ZN(
        n13155) );
  AOI211_X1 U16309 ( .C1(n19675), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n19678), .B(n13155), .ZN(n13156) );
  OAI221_X1 U16310 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(n13157), .C1(n15655), 
        .C2(n19628), .A(n13156), .ZN(n13158) );
  AOI21_X1 U16311 ( .B1(n19644), .B2(n13159), .A(n13158), .ZN(n13160) );
  OAI21_X1 U16312 ( .B1(n13162), .B2(n15470), .A(n13160), .ZN(P1_U2832) );
  MUX2_X1 U16313 ( .A(DATAI_8_), .B(BUF1_REG_8__SCAN_IN), .S(n19836), .Z(
        n19750) );
  AOI22_X1 U16314 ( .A1(n15544), .A2(n19750), .B1(n15545), .B2(
        P1_EAX_REG_8__SCAN_IN), .ZN(n13161) );
  OAI21_X1 U16315 ( .B1(n13162), .B2(n19714), .A(n13161), .ZN(P1_U2896) );
  AOI21_X1 U16316 ( .B1(n18630), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n13163), .ZN(n19529) );
  AOI22_X1 U16317 ( .A1(n18630), .A2(n10038), .B1(n13165), .B2(n15696), .ZN(
        n13707) );
  NAND2_X1 U16318 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n13707), .ZN(n19528) );
  INV_X1 U16319 ( .A(n19528), .ZN(n13168) );
  OAI22_X1 U16320 ( .A1(n19557), .A2(n19525), .B1(n19537), .B2(n13166), .ZN(
        n13167) );
  AOI21_X1 U16321 ( .B1(n19529), .B2(n13168), .A(n13167), .ZN(n13174) );
  NAND2_X1 U16322 ( .A1(n13169), .A2(n18699), .ZN(n13172) );
  OAI22_X1 U16323 ( .A1(n15906), .A2(n12450), .B1(P2_STATE2_REG_0__SCAN_IN), 
        .B2(n19535), .ZN(n13170) );
  INV_X1 U16324 ( .A(n13170), .ZN(n13171) );
  NAND2_X1 U16325 ( .A1(n13172), .A2(n13171), .ZN(n19530) );
  INV_X1 U16326 ( .A(n19530), .ZN(n19521) );
  NAND2_X1 U16327 ( .A1(n19521), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13173) );
  OAI21_X1 U16328 ( .B1(n13174), .B2(n19521), .A(n13173), .ZN(P2_U3600) );
  NAND2_X1 U16329 ( .A1(n13176), .A2(n13175), .ZN(n13177) );
  AND2_X1 U16330 ( .A1(n13207), .A2(n13177), .ZN(n18503) );
  OAI211_X1 U16331 ( .C1(n11562), .C2(n10283), .A(n14522), .B(n13195), .ZN(
        n13180) );
  NAND2_X1 U16332 ( .A1(n14548), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n13179) );
  OAI211_X1 U16333 ( .C1(n15002), .C2(n14548), .A(n13180), .B(n13179), .ZN(
        P2_U2872) );
  AOI21_X1 U16334 ( .B1(n13181), .B2(n9850), .A(n13398), .ZN(n19632) );
  INV_X1 U16335 ( .A(n19632), .ZN(n13437) );
  AOI21_X1 U16336 ( .B1(n13183), .B2(n13182), .A(n9750), .ZN(n19626) );
  AOI22_X1 U16337 ( .A1(n19705), .A2(n19626), .B1(P1_EBX_REG_9__SCAN_IN), .B2(
        n14004), .ZN(n13184) );
  OAI21_X1 U16338 ( .B1(n13437), .B2(n14024), .A(n13184), .ZN(P1_U2863) );
  MUX2_X1 U16339 ( .A(DATAI_9_), .B(BUF1_REG_9__SCAN_IN), .S(n19836), .Z(
        n19752) );
  AOI22_X1 U16340 ( .A1(n15544), .A2(n19752), .B1(n15545), .B2(
        P1_EAX_REG_9__SCAN_IN), .ZN(n13185) );
  OAI21_X1 U16341 ( .B1(n13437), .B2(n19714), .A(n13185), .ZN(P1_U2895) );
  NAND3_X1 U16342 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n12827), .A3(
        n19560), .ZN(n19056) );
  NOR2_X1 U16343 ( .A1(n19571), .A2(n19056), .ZN(n19073) );
  AOI21_X1 U16344 ( .B1(n19092), .B2(n19127), .A(n19263), .ZN(n13186) );
  NOR2_X1 U16345 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19106), .ZN(
        n19093) );
  AOI221_X1 U16346 ( .B1(n19073), .B2(n19535), .C1(n13186), .C2(n19535), .A(
        n19093), .ZN(n13188) );
  NAND2_X1 U16347 ( .A1(n13260), .A2(n13187), .ZN(n13222) );
  NOR3_X1 U16348 ( .A1(n13442), .A2(n19093), .A3(n19586), .ZN(n13189) );
  INV_X1 U16349 ( .A(n19096), .ZN(n13194) );
  INV_X1 U16350 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13193) );
  AOI22_X1 U16351 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n18924), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n18923), .ZN(n19383) );
  AOI22_X1 U16352 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n18924), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n18923), .ZN(n19306) );
  INV_X1 U16353 ( .A(n19306), .ZN(n19380) );
  AOI22_X1 U16354 ( .A1(n19095), .A2(n19303), .B1(n19089), .B2(n19380), .ZN(
        n13192) );
  NOR2_X1 U16355 ( .A1(n19073), .A2(n19093), .ZN(n13190) );
  AOI211_X2 U16356 ( .C1(n13190), .C2(n19586), .A(n19101), .B(n13189), .ZN(
        n19094) );
  AOI22_X1 U16357 ( .A1(n14634), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n14633), .ZN(n18785) );
  NOR2_X2 U16358 ( .A1(n18785), .A2(n19104), .ZN(n19371) );
  NOR2_X2 U16359 ( .A1(n9634), .A2(n18925), .ZN(n19370) );
  AOI22_X1 U16360 ( .A1(n19094), .A2(n19371), .B1(n19370), .B2(n19093), .ZN(
        n13191) );
  OAI211_X1 U16361 ( .C1(n13194), .C2(n13193), .A(n13192), .B(n13191), .ZN(
        P2_U3096) );
  AOI21_X1 U16362 ( .B1(n13196), .B2(n13195), .A(n13386), .ZN(n13197) );
  INV_X1 U16363 ( .A(n13197), .ZN(n13211) );
  AOI21_X1 U16364 ( .B1(n13198), .B2(n9728), .A(n13392), .ZN(n18491) );
  NAND2_X1 U16365 ( .A1(n18651), .A2(BUF2_REG_16__SCAN_IN), .ZN(n13203) );
  NAND2_X1 U16366 ( .A1(n18652), .A2(BUF1_REG_16__SCAN_IN), .ZN(n13202) );
  INV_X1 U16367 ( .A(n18785), .ZN(n13200) );
  AOI22_X1 U16368 ( .A1(n15778), .A2(n13200), .B1(n18691), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n13201) );
  NAND3_X1 U16369 ( .A1(n13203), .A2(n13202), .A3(n13201), .ZN(n13204) );
  AOI21_X1 U16370 ( .B1(n18491), .B2(n18692), .A(n13204), .ZN(n13205) );
  OAI21_X1 U16371 ( .B1(n18671), .B2(n13211), .A(n13205), .ZN(P2_U2903) );
  NAND2_X1 U16372 ( .A1(n14548), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n13210) );
  NAND2_X1 U16373 ( .A1(n13207), .A2(n13206), .ZN(n13208) );
  AND2_X1 U16374 ( .A1(n13416), .A2(n13208), .ZN(n18490) );
  NAND2_X1 U16375 ( .A1(n14540), .A2(n18490), .ZN(n13209) );
  OAI211_X1 U16376 ( .C1(n13211), .C2(n14550), .A(n13210), .B(n13209), .ZN(
        P2_U2871) );
  XNOR2_X1 U16377 ( .A(n13213), .B(n13212), .ZN(n13214) );
  XNOR2_X1 U16378 ( .A(n13215), .B(n13214), .ZN(n15653) );
  AOI22_X1 U16379 ( .A1(n19782), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n19781), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n13216) );
  OAI21_X1 U16380 ( .B1(n19793), .B2(n13217), .A(n13216), .ZN(n13218) );
  AOI21_X1 U16381 ( .B1(n13219), .B2(n19787), .A(n13218), .ZN(n13220) );
  OAI21_X1 U16382 ( .B1(n15653), .B2(n19608), .A(n13220), .ZN(P1_U2991) );
  INV_X1 U16383 ( .A(n13222), .ZN(n13223) );
  AOI22_X1 U16384 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n13442), .B1(
        n19340), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13256) );
  NAND2_X1 U16385 ( .A1(n15080), .A2(n13260), .ZN(n13224) );
  NOR2_X2 U16386 ( .A1(n13257), .A2(n13224), .ZN(n19023) );
  INV_X1 U16387 ( .A(n13224), .ZN(n13225) );
  AOI22_X1 U16388 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19023), .B1(
        n19259), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13255) );
  NAND2_X1 U16389 ( .A1(n14440), .A2(n13231), .ZN(n13227) );
  INV_X1 U16390 ( .A(n13227), .ZN(n13228) );
  NAND2_X1 U16391 ( .A1(n13260), .A2(n13228), .ZN(n13248) );
  OR2_X2 U16392 ( .A1(n15895), .A2(n13248), .ZN(n19053) );
  INV_X1 U16393 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13229) );
  OAI22_X1 U16394 ( .A1(n13230), .A2(n18933), .B1(n19053), .B2(n13229), .ZN(
        n13239) );
  INV_X1 U16395 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13237) );
  INV_X1 U16396 ( .A(n13231), .ZN(n13232) );
  NAND2_X1 U16397 ( .A1(n13232), .A2(n14440), .ZN(n13240) );
  OR2_X2 U16398 ( .A1(n13234), .A2(n15895), .ZN(n18992) );
  INV_X1 U16399 ( .A(n13234), .ZN(n13235) );
  INV_X1 U16400 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13236) );
  OAI22_X1 U16401 ( .A1(n13237), .A2(n18992), .B1(n19225), .B2(n13236), .ZN(
        n13238) );
  NOR2_X1 U16402 ( .A1(n13239), .A2(n13238), .ZN(n13254) );
  INV_X1 U16403 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13245) );
  INV_X1 U16404 ( .A(n13240), .ZN(n13241) );
  NAND2_X1 U16405 ( .A1(n13260), .A2(n13241), .ZN(n13242) );
  OR2_X2 U16406 ( .A1(n15895), .A2(n13242), .ZN(n19099) );
  INV_X1 U16407 ( .A(n13242), .ZN(n13243) );
  NAND2_X1 U16408 ( .A1(n15895), .A2(n13243), .ZN(n19368) );
  INV_X1 U16409 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13244) );
  OAI22_X1 U16410 ( .A1(n13245), .A2(n19099), .B1(n19368), .B2(n13244), .ZN(
        n13252) );
  INV_X1 U16411 ( .A(n13246), .ZN(n13247) );
  NAND2_X2 U16412 ( .A1(n15895), .A2(n13247), .ZN(n19165) );
  INV_X1 U16413 ( .A(n13248), .ZN(n13249) );
  NAND2_X1 U16414 ( .A1(n15895), .A2(n13249), .ZN(n19293) );
  INV_X1 U16415 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13250) );
  OAI22_X1 U16416 ( .A1(n11507), .A2(n19165), .B1(n19293), .B2(n13250), .ZN(
        n13251) );
  NOR2_X1 U16417 ( .A1(n13252), .A2(n13251), .ZN(n13253) );
  NAND2_X1 U16418 ( .A1(n18887), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13259) );
  NAND2_X1 U16419 ( .A1(n13459), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n13258) );
  NAND2_X1 U16420 ( .A1(n13259), .A2(n13258), .ZN(n13265) );
  INV_X1 U16421 ( .A(n13260), .ZN(n13261) );
  NOR2_X2 U16422 ( .A1(n13264), .A2(n15080), .ZN(n19195) );
  NOR3_X1 U16423 ( .A1(n13265), .A2(n10286), .A3(n10284), .ZN(n13266) );
  NAND2_X1 U16424 ( .A1(n10289), .A2(n13266), .ZN(n13269) );
  NAND2_X1 U16425 ( .A1(n13267), .A2(n18895), .ZN(n13268) );
  INV_X1 U16426 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13272) );
  INV_X1 U16427 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13270) );
  OAI211_X1 U16428 ( .C1(n19099), .C2(n13272), .A(n13271), .B(n9643), .ZN(
        n13273) );
  AOI21_X1 U16429 ( .B1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n19340), .A(
        n13273), .ZN(n13277) );
  NAND2_X1 U16430 ( .A1(n18887), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13276) );
  NAND2_X1 U16431 ( .A1(n13459), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n13275) );
  NAND2_X1 U16432 ( .A1(n19195), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n13274) );
  NAND4_X1 U16433 ( .A1(n13277), .A2(n13276), .A3(n13275), .A4(n13274), .ZN(
        n13297) );
  NAND2_X1 U16434 ( .A1(n19136), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n13291) );
  INV_X1 U16435 ( .A(n19259), .ZN(n19265) );
  INV_X1 U16436 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13278) );
  NOR2_X1 U16437 ( .A1(n19265), .A2(n13278), .ZN(n13282) );
  INV_X1 U16438 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13280) );
  INV_X1 U16439 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13279) );
  OAI22_X1 U16440 ( .A1(n13280), .A2(n18992), .B1(n19368), .B2(n13279), .ZN(
        n13281) );
  NOR2_X1 U16441 ( .A1(n13282), .A2(n13281), .ZN(n13290) );
  INV_X1 U16442 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13284) );
  INV_X1 U16443 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13283) );
  OAI22_X1 U16444 ( .A1(n13284), .A2(n18933), .B1(n19053), .B2(n13283), .ZN(
        n13288) );
  INV_X1 U16445 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13286) );
  INV_X1 U16446 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13285) );
  OAI22_X1 U16447 ( .A1(n13286), .A2(n19293), .B1(n19165), .B2(n13285), .ZN(
        n13287) );
  NOR2_X1 U16448 ( .A1(n13288), .A2(n13287), .ZN(n13289) );
  NAND4_X1 U16449 ( .A1(n13292), .A2(n13291), .A3(n13290), .A4(n13289), .ZN(
        n13296) );
  NAND2_X1 U16450 ( .A1(n13294), .A2(n13293), .ZN(n13346) );
  NAND2_X1 U16451 ( .A1(n13346), .A2(n13347), .ZN(n13295) );
  AOI22_X1 U16452 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n13442), .B1(
        n19340), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13315) );
  AOI22_X1 U16453 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19023), .B1(
        n19259), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13314) );
  INV_X1 U16454 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13301) );
  INV_X1 U16455 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13300) );
  OAI22_X1 U16456 ( .A1(n13301), .A2(n19099), .B1(n19293), .B2(n13300), .ZN(
        n13305) );
  INV_X1 U16457 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13303) );
  INV_X1 U16458 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13302) );
  OAI22_X1 U16459 ( .A1(n13303), .A2(n19368), .B1(n19225), .B2(n13302), .ZN(
        n13304) );
  NOR2_X1 U16460 ( .A1(n13305), .A2(n13304), .ZN(n13313) );
  INV_X1 U16461 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13307) );
  INV_X1 U16462 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13306) );
  OAI22_X1 U16463 ( .A1(n13307), .A2(n18992), .B1(n19053), .B2(n13306), .ZN(
        n13311) );
  INV_X1 U16464 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13309) );
  INV_X1 U16465 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13308) );
  OAI22_X1 U16466 ( .A1(n13309), .A2(n18933), .B1(n19165), .B2(n13308), .ZN(
        n13310) );
  NOR2_X1 U16467 ( .A1(n13311), .A2(n13310), .ZN(n13312) );
  NAND4_X1 U16468 ( .A1(n13315), .A2(n13314), .A3(n13313), .A4(n13312), .ZN(
        n13322) );
  NAND2_X1 U16469 ( .A1(n19195), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n13320) );
  NAND2_X1 U16470 ( .A1(n13459), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n13319) );
  NAND2_X1 U16471 ( .A1(n19136), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n13318) );
  INV_X1 U16472 ( .A(n18887), .ZN(n18884) );
  NAND4_X1 U16473 ( .A1(n13320), .A2(n13319), .A3(n13318), .A4(n13317), .ZN(
        n13321) );
  INV_X1 U16474 ( .A(n13323), .ZN(n13324) );
  NAND2_X1 U16475 ( .A1(n13324), .A2(n18895), .ZN(n13325) );
  OAI21_X1 U16476 ( .B1(n13329), .B2(n13328), .A(n13475), .ZN(n18617) );
  INV_X1 U16477 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13373) );
  XNOR2_X1 U16478 ( .A(n13479), .B(n13373), .ZN(n13478) );
  NOR2_X1 U16479 ( .A1(n13334), .A2(n13333), .ZN(n13336) );
  OAI21_X1 U16480 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13336), .A(
        n13335), .ZN(n18823) );
  XNOR2_X1 U16481 ( .A(n13337), .B(n18878), .ZN(n18822) );
  OR2_X1 U16482 ( .A1(n18823), .A2(n18822), .ZN(n18825) );
  NAND2_X1 U16483 ( .A1(n13338), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13339) );
  NAND2_X1 U16484 ( .A1(n18825), .A2(n13339), .ZN(n15845) );
  INV_X1 U16485 ( .A(n13340), .ZN(n13341) );
  XNOR2_X1 U16486 ( .A(n13342), .B(n13341), .ZN(n18638) );
  INV_X1 U16487 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18844) );
  NAND2_X1 U16488 ( .A1(n18638), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13343) );
  NAND2_X1 U16489 ( .A1(n13344), .A2(n13343), .ZN(n13477) );
  XNOR2_X1 U16490 ( .A(n13478), .B(n13477), .ZN(n15837) );
  XOR2_X1 U16491 ( .A(n13347), .B(n13346), .Z(n18819) );
  NOR2_X1 U16492 ( .A1(n13349), .A2(n13348), .ZN(n13351) );
  NOR2_X1 U16493 ( .A1(n13351), .A2(n13350), .ZN(n13352) );
  XOR2_X1 U16494 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n13352), .Z(
        n18818) );
  NOR2_X1 U16495 ( .A1(n18819), .A2(n18818), .ZN(n18817) );
  NOR2_X1 U16496 ( .A1(n13352), .A2(n18878), .ZN(n13353) );
  OR2_X1 U16497 ( .A1(n18817), .A2(n13353), .ZN(n13354) );
  INV_X1 U16498 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n15903) );
  XNOR2_X1 U16499 ( .A(n13354), .B(n15903), .ZN(n15849) );
  NAND2_X1 U16500 ( .A1(n13354), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13355) );
  NAND2_X1 U16501 ( .A1(n13357), .A2(n13356), .ZN(n13358) );
  NAND2_X1 U16502 ( .A1(n13439), .A2(n13358), .ZN(n13360) );
  INV_X1 U16503 ( .A(n13359), .ZN(n13361) );
  NAND2_X1 U16504 ( .A1(n13361), .A2(n13360), .ZN(n13362) );
  OAI21_X1 U16505 ( .B1(n9966), .B2(n13366), .A(n13365), .ZN(n13367) );
  OAI21_X1 U16506 ( .B1(n13471), .B2(n9966), .A(n13367), .ZN(n15839) );
  INV_X1 U16507 ( .A(n15839), .ZN(n13382) );
  NAND2_X1 U16508 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18869) );
  NAND2_X1 U16509 ( .A1(n18878), .A2(n18869), .ZN(n18865) );
  INV_X1 U16510 ( .A(n18870), .ZN(n18856) );
  NOR2_X1 U16511 ( .A1(n18878), .A2(n18869), .ZN(n13371) );
  INV_X1 U16512 ( .A(n13371), .ZN(n18866) );
  AOI21_X1 U16513 ( .B1(n18856), .B2(n18866), .A(n18855), .ZN(n13368) );
  OAI21_X1 U16514 ( .B1(n18864), .B2(n18865), .A(n13368), .ZN(n13488) );
  NOR2_X1 U16515 ( .A1(n15903), .A2(n13488), .ZN(n18841) );
  NAND2_X1 U16516 ( .A1(n18837), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13380) );
  OAI21_X1 U16517 ( .B1(n18634), .B2(n13370), .A(n13369), .ZN(n18674) );
  INV_X1 U16518 ( .A(n18674), .ZN(n13378) );
  INV_X1 U16519 ( .A(n18624), .ZN(n13376) );
  INV_X1 U16520 ( .A(n18864), .ZN(n13372) );
  OAI211_X1 U16521 ( .C1(n13372), .C2(n13371), .A(n18865), .B(n14943), .ZN(
        n15902) );
  NOR2_X1 U16522 ( .A1(n15903), .A2(n15902), .ZN(n18845) );
  OAI221_X1 U16523 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(n13373), .C2(n18844), .A(
        n18845), .ZN(n13375) );
  NAND2_X1 U16524 ( .A1(n18850), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n13374) );
  OAI211_X1 U16525 ( .C1(n18839), .C2(n13376), .A(n13375), .B(n13374), .ZN(
        n13377) );
  AOI21_X1 U16526 ( .B1(n13378), .B2(n18875), .A(n13377), .ZN(n13379) );
  OAI21_X1 U16527 ( .B1(n18841), .B2(n13380), .A(n13379), .ZN(n13381) );
  AOI21_X1 U16528 ( .B1(n13382), .B2(n18849), .A(n13381), .ZN(n13383) );
  OAI21_X1 U16529 ( .B1(n18859), .B2(n15837), .A(n13383), .ZN(P2_U3041) );
  OR2_X1 U16530 ( .A1(n13386), .A2(n13385), .ZN(n13387) );
  NAND2_X1 U16531 ( .A1(n13384), .A2(n13387), .ZN(n13419) );
  NAND2_X1 U16532 ( .A1(n18652), .A2(BUF1_REG_17__SCAN_IN), .ZN(n13390) );
  INV_X1 U16533 ( .A(n18896), .ZN(n13388) );
  AOI22_X1 U16534 ( .A1(n15778), .A2(n13388), .B1(n18691), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n13389) );
  NAND2_X1 U16535 ( .A1(n13390), .A2(n13389), .ZN(n13394) );
  OAI21_X1 U16536 ( .B1(n13392), .B2(n13391), .A(n9650), .ZN(n18484) );
  NOR2_X1 U16537 ( .A1(n18484), .A2(n18687), .ZN(n13393) );
  AOI211_X1 U16538 ( .C1(n18651), .C2(BUF2_REG_17__SCAN_IN), .A(n13394), .B(
        n13393), .ZN(n13395) );
  OAI21_X1 U16539 ( .B1(n18671), .B2(n13419), .A(n13395), .ZN(P2_U2902) );
  INV_X1 U16540 ( .A(n13501), .ZN(n13396) );
  OAI21_X1 U16541 ( .B1(n13398), .B2(n13397), .A(n13396), .ZN(n14219) );
  OR2_X1 U16542 ( .A1(n9750), .A2(n13399), .ZN(n13400) );
  AND2_X1 U16543 ( .A1(n15522), .A2(n13400), .ZN(n15631) );
  INV_X1 U16544 ( .A(n15631), .ZN(n13402) );
  OAI22_X1 U16545 ( .A1(n14025), .A2(n13402), .B1(n13401), .B2(n19710), .ZN(
        n13403) );
  INV_X1 U16546 ( .A(n13403), .ZN(n13404) );
  OAI21_X1 U16547 ( .B1(n14219), .B2(n14024), .A(n13404), .ZN(P1_U2862) );
  MUX2_X1 U16548 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n19836), .Z(
        n19754) );
  AOI22_X1 U16549 ( .A1(n15544), .A2(n19754), .B1(n15545), .B2(
        P1_EAX_REG_10__SCAN_IN), .ZN(n13405) );
  OAI21_X1 U16550 ( .B1(n14219), .B2(n19714), .A(n13405), .ZN(P1_U2894) );
  INV_X1 U16551 ( .A(n14215), .ZN(n13413) );
  INV_X1 U16552 ( .A(n13406), .ZN(n13508) );
  NAND2_X1 U16553 ( .A1(n15450), .A2(n13508), .ZN(n13407) );
  AND2_X1 U16554 ( .A1(n13407), .A2(n13961), .ZN(n13507) );
  AOI21_X1 U16555 ( .B1(n19675), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n19678), .ZN(n13409) );
  AOI22_X1 U16556 ( .A1(P1_EBX_REG_10__SCAN_IN), .A2(n19687), .B1(n19686), 
        .B2(n15631), .ZN(n13408) );
  OAI211_X1 U16557 ( .C1(n13410), .C2(n13507), .A(n13409), .B(n13408), .ZN(
        n13412) );
  INV_X1 U16558 ( .A(n19651), .ZN(n19665) );
  NOR4_X1 U16559 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n19629), .A3(n19625), 
        .A4(n19665), .ZN(n13411) );
  AOI211_X1 U16560 ( .C1(n19644), .C2(n13413), .A(n13412), .B(n13411), .ZN(
        n13414) );
  OAI21_X1 U16561 ( .B1(n14219), .B2(n15470), .A(n13414), .ZN(P1_U2830) );
  AND2_X1 U16562 ( .A1(n13416), .A2(n13415), .ZN(n13417) );
  NOR2_X1 U16563 ( .A1(n14544), .A2(n13417), .ZN(n18482) );
  INV_X1 U16564 ( .A(n18482), .ZN(n14982) );
  MUX2_X1 U16565 ( .A(n11911), .B(n14982), .S(n14525), .Z(n13418) );
  OAI21_X1 U16566 ( .B1(n13419), .B2(n14550), .A(n13418), .ZN(P2_U2870) );
  INV_X1 U16567 ( .A(n13384), .ZN(n13422) );
  INV_X1 U16568 ( .A(n13420), .ZN(n13421) );
  OAI21_X1 U16569 ( .B1(n13422), .B2(n13421), .A(n14534), .ZN(n14551) );
  INV_X1 U16570 ( .A(n13423), .ZN(n14632) );
  AOI21_X1 U16571 ( .B1(n13424), .B2(n9650), .A(n14632), .ZN(n18470) );
  NAND2_X1 U16572 ( .A1(n18651), .A2(BUF2_REG_18__SCAN_IN), .ZN(n13428) );
  NAND2_X1 U16573 ( .A1(n18652), .A2(BUF1_REG_18__SCAN_IN), .ZN(n13427) );
  AOI22_X1 U16574 ( .A1(n15778), .A2(n13425), .B1(n18691), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n13426) );
  NAND3_X1 U16575 ( .A1(n13428), .A2(n13427), .A3(n13426), .ZN(n13429) );
  AOI21_X1 U16576 ( .B1(n18470), .B2(n18692), .A(n13429), .ZN(n13430) );
  OAI21_X1 U16577 ( .B1(n18671), .B2(n14551), .A(n13430), .ZN(P2_U2901) );
  MUX2_X1 U16578 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n11134), .S(
        n15572), .Z(n13431) );
  XNOR2_X1 U16579 ( .A(n13432), .B(n13431), .ZN(n15644) );
  NAND2_X1 U16580 ( .A1(n15644), .A2(n19788), .ZN(n13436) );
  INV_X1 U16581 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n13433) );
  NAND2_X1 U16582 ( .A1(n19781), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n15641) );
  OAI21_X1 U16583 ( .B1(n14190), .B2(n13433), .A(n15641), .ZN(n13434) );
  AOI21_X1 U16584 ( .B1(n15566), .B2(n19631), .A(n13434), .ZN(n13435) );
  OAI211_X1 U16585 ( .C1(n19835), .C2(n13437), .A(n13436), .B(n13435), .ZN(
        P1_U2990) );
  INV_X1 U16586 ( .A(n13439), .ZN(n13441) );
  AOI22_X1 U16587 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19023), .B1(
        n19259), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13458) );
  AOI22_X1 U16588 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n13442), .B1(
        n19340), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13457) );
  INV_X1 U16589 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13443) );
  OAI22_X1 U16590 ( .A1(n13444), .A2(n19099), .B1(n19165), .B2(n13443), .ZN(
        n13448) );
  INV_X1 U16591 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13446) );
  INV_X1 U16592 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13445) );
  OAI22_X1 U16593 ( .A1(n13446), .A2(n18933), .B1(n19293), .B2(n13445), .ZN(
        n13447) );
  NOR2_X1 U16594 ( .A1(n13448), .A2(n13447), .ZN(n13456) );
  INV_X1 U16595 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13450) );
  INV_X1 U16596 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13449) );
  OAI22_X1 U16597 ( .A1(n13450), .A2(n18992), .B1(n19053), .B2(n13449), .ZN(
        n13454) );
  INV_X1 U16598 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13451) );
  OAI22_X1 U16599 ( .A1(n13452), .A2(n19225), .B1(n19368), .B2(n13451), .ZN(
        n13453) );
  NOR2_X1 U16600 ( .A1(n13454), .A2(n13453), .ZN(n13455) );
  NAND4_X1 U16601 ( .A1(n13458), .A2(n13457), .A3(n13456), .A4(n13455), .ZN(
        n13466) );
  NAND2_X1 U16602 ( .A1(n19136), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n13464) );
  NAND2_X1 U16603 ( .A1(n18887), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n13463) );
  NAND2_X1 U16604 ( .A1(n19195), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n13462) );
  INV_X1 U16605 ( .A(n13459), .ZN(n18962) );
  NAND4_X1 U16606 ( .A1(n13464), .A2(n13463), .A3(n13462), .A4(n13461), .ZN(
        n13465) );
  NAND2_X1 U16607 ( .A1(n13467), .A2(n18895), .ZN(n13468) );
  INV_X1 U16608 ( .A(n13856), .ZN(n13470) );
  INV_X1 U16609 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13491) );
  XNOR2_X1 U16610 ( .A(n13855), .B(n13491), .ZN(n13498) );
  INV_X1 U16611 ( .A(n13473), .ZN(n13474) );
  XNOR2_X1 U16612 ( .A(n13475), .B(n13474), .ZN(n18602) );
  INV_X1 U16613 ( .A(n18602), .ZN(n13476) );
  NAND2_X1 U16614 ( .A1(n13478), .A2(n13477), .ZN(n13481) );
  NAND2_X1 U16615 ( .A1(n13479), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13480) );
  XNOR2_X1 U16616 ( .A(n13741), .B(n13742), .ZN(n13496) );
  INV_X1 U16617 ( .A(n13492), .ZN(n18610) );
  AOI22_X1 U16618 ( .A1(n18830), .A2(n18610), .B1(n18820), .B2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n13485) );
  OAI22_X1 U16619 ( .A1(n19468), .A2(n18600), .B1(n18816), .B2(n18607), .ZN(
        n13483) );
  INV_X1 U16620 ( .A(n13483), .ZN(n13484) );
  OAI211_X1 U16621 ( .C1(n13496), .C2(n18833), .A(n13485), .B(n13484), .ZN(
        n13486) );
  AOI21_X1 U16622 ( .B1(n13498), .B2(n18821), .A(n13486), .ZN(n13487) );
  INV_X1 U16623 ( .A(n13487), .ZN(P2_U3008) );
  NAND3_X1 U16624 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13489) );
  NOR2_X1 U16625 ( .A1(n13489), .A2(n15902), .ZN(n13873) );
  AOI221_X1 U16626 ( .B1(n13491), .B2(n14943), .C1(n13489), .C2(n14943), .A(
        n13488), .ZN(n15894) );
  INV_X1 U16627 ( .A(n15894), .ZN(n15071) );
  NOR2_X1 U16628 ( .A1(n19468), .A2(n18600), .ZN(n13490) );
  AOI221_X1 U16629 ( .B1(n13873), .B2(n13491), .C1(n15071), .C2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(n13490), .ZN(n13495) );
  OAI22_X1 U16630 ( .A1(n18613), .A2(n15898), .B1(n18839), .B2(n13492), .ZN(
        n13493) );
  INV_X1 U16631 ( .A(n13493), .ZN(n13494) );
  OAI211_X1 U16632 ( .C1(n13496), .C2(n18859), .A(n13495), .B(n13494), .ZN(
        n13497) );
  AOI21_X1 U16633 ( .B1(n13498), .B2(n18849), .A(n13497), .ZN(n13499) );
  INV_X1 U16634 ( .A(n13499), .ZN(P2_U3040) );
  OR2_X1 U16635 ( .A1(n13501), .A2(n13500), .ZN(n13502) );
  NAND2_X1 U16636 ( .A1(n13503), .A2(n13502), .ZN(n15529) );
  INV_X1 U16637 ( .A(n15528), .ZN(n13504) );
  OAI21_X1 U16638 ( .B1(n15529), .B2(n13504), .A(n13503), .ZN(n13521) );
  AND2_X1 U16639 ( .A1(n13521), .A2(n13520), .ZN(n13523) );
  OAI21_X1 U16640 ( .B1(n13523), .B2(n13505), .A(n13527), .ZN(n14211) );
  MUX2_X1 U16641 ( .A(DATAI_13_), .B(BUF1_REG_13__SCAN_IN), .S(n19836), .Z(
        n19760) );
  AOI22_X1 U16642 ( .A1(n15544), .A2(n19760), .B1(n15545), .B2(
        P1_EAX_REG_13__SCAN_IN), .ZN(n13506) );
  OAI21_X1 U16643 ( .B1(n14211), .B2(n19714), .A(n13506), .ZN(P1_U2891) );
  INV_X1 U16644 ( .A(n13507), .ZN(n15530) );
  AOI21_X1 U16645 ( .B1(n13509), .B2(n19636), .A(n15530), .ZN(n15514) );
  NOR2_X1 U16646 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n13509), .ZN(n13510) );
  AOI22_X1 U16647 ( .A1(n15525), .A2(n13510), .B1(n19644), .B2(n14208), .ZN(
        n13516) );
  OAI21_X1 U16648 ( .B1(n15520), .B2(n13524), .A(n13511), .ZN(n13512) );
  AND2_X1 U16649 ( .A1(n13512), .A2(n13534), .ZN(n15614) );
  AOI22_X1 U16650 ( .A1(P1_EBX_REG_13__SCAN_IN), .A2(n19687), .B1(n19686), 
        .B2(n15614), .ZN(n13513) );
  OAI211_X1 U16651 ( .C1(n19691), .C2(n20629), .A(n13513), .B(n19653), .ZN(
        n13514) );
  INV_X1 U16652 ( .A(n13514), .ZN(n13515) );
  OAI211_X1 U16653 ( .C1(n15514), .C2(n15610), .A(n13516), .B(n13515), .ZN(
        n13517) );
  INV_X1 U16654 ( .A(n13517), .ZN(n13518) );
  OAI21_X1 U16655 ( .B1(n14211), .B2(n15470), .A(n13518), .ZN(P1_U2827) );
  AOI22_X1 U16656 ( .A1(n19705), .A2(n15614), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n14004), .ZN(n13519) );
  OAI21_X1 U16657 ( .B1(n14211), .B2(n14024), .A(n13519), .ZN(P1_U2859) );
  NOR2_X1 U16658 ( .A1(n13521), .A2(n13520), .ZN(n13522) );
  XOR2_X1 U16659 ( .A(n13524), .B(n15520), .Z(n15513) );
  AOI22_X1 U16660 ( .A1(n15513), .A2(n19705), .B1(P1_EBX_REG_12__SCAN_IN), 
        .B2(n14004), .ZN(n13525) );
  OAI21_X1 U16661 ( .B1(n15543), .B2(n14024), .A(n13525), .ZN(P1_U2860) );
  AOI21_X1 U16662 ( .B1(n13528), .B2(n13527), .A(n13526), .ZN(n14201) );
  INV_X1 U16663 ( .A(n14201), .ZN(n13542) );
  MUX2_X1 U16664 ( .A(DATAI_14_), .B(BUF1_REG_14__SCAN_IN), .S(n19836), .Z(
        n19762) );
  AOI22_X1 U16665 ( .A1(n15544), .A2(n19762), .B1(n15545), .B2(
        P1_EAX_REG_14__SCAN_IN), .ZN(n13529) );
  OAI21_X1 U16666 ( .B1(n13542), .B2(n19714), .A(n13529), .ZN(P1_U2890) );
  INV_X1 U16667 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n14408) );
  NAND2_X1 U16668 ( .A1(n13958), .A2(n15525), .ZN(n13530) );
  NAND2_X1 U16669 ( .A1(n14408), .A2(n13530), .ZN(n13540) );
  INV_X1 U16670 ( .A(n13531), .ZN(n13532) );
  OAI21_X1 U16671 ( .B1(n13963), .B2(n13532), .A(n13961), .ZN(n15506) );
  INV_X1 U16672 ( .A(n14399), .ZN(n13536) );
  NAND2_X1 U16673 ( .A1(n13534), .A2(n13533), .ZN(n13535) );
  NAND2_X1 U16674 ( .A1(n13536), .A2(n13535), .ZN(n14409) );
  OAI22_X1 U16675 ( .A1(n13543), .A2(n19662), .B1(n19681), .B2(n14409), .ZN(
        n13537) );
  AOI211_X1 U16676 ( .C1(n19675), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n13537), .B(n19678), .ZN(n13538) );
  OAI21_X1 U16677 ( .B1(n14199), .B2(n19690), .A(n13538), .ZN(n13539) );
  AOI21_X1 U16678 ( .B1(n13540), .B2(n15506), .A(n13539), .ZN(n13541) );
  OAI21_X1 U16679 ( .B1(n13542), .B2(n15470), .A(n13541), .ZN(P1_U2826) );
  OAI22_X1 U16680 ( .A1(n14409), .A2(n14025), .B1(n13543), .B2(n19710), .ZN(
        n13544) );
  AOI21_X1 U16681 ( .B1(n14201), .B2(n19706), .A(n13544), .ZN(n13545) );
  INV_X1 U16682 ( .A(n13545), .ZN(P1_U2858) );
  INV_X1 U16683 ( .A(n13547), .ZN(n13548) );
  AOI21_X1 U16684 ( .B1(n9915), .B2(n13549), .A(n13548), .ZN(n13552) );
  AND2_X1 U16685 ( .A1(n13550), .A2(n14204), .ZN(n13551) );
  NAND2_X1 U16686 ( .A1(n13552), .A2(n13551), .ZN(n14205) );
  OAI21_X1 U16687 ( .B1(n13552), .B2(n13551), .A(n14205), .ZN(n13553) );
  INV_X1 U16688 ( .A(n13553), .ZN(n15569) );
  INV_X1 U16689 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n13561) );
  NAND2_X1 U16690 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15649) );
  INV_X1 U16691 ( .A(n15649), .ZN(n19794) );
  NAND2_X1 U16692 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n19801) );
  NOR2_X1 U16693 ( .A1(n15679), .A2(n19801), .ZN(n13562) );
  NAND2_X1 U16694 ( .A1(n19794), .A2(n13562), .ZN(n15633) );
  INV_X1 U16695 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15665) );
  NOR3_X1 U16696 ( .A1(n13212), .A2(n15665), .A3(n12308), .ZN(n15636) );
  NAND3_X1 U16697 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n15636), .ZN(n14222) );
  NOR2_X1 U16698 ( .A1(n15633), .A2(n14222), .ZN(n14223) );
  INV_X1 U16699 ( .A(n19824), .ZN(n13557) );
  OAI21_X1 U16700 ( .B1(n13554), .B2(n19819), .A(n19831), .ZN(n19826) );
  NAND2_X1 U16701 ( .A1(n13562), .A2(n19826), .ZN(n14221) );
  OR2_X1 U16702 ( .A1(n14326), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13556) );
  NAND2_X1 U16703 ( .A1(n13556), .A2(n13555), .ZN(n19817) );
  AOI21_X1 U16704 ( .B1(n13557), .B2(n14221), .A(n19817), .ZN(n15632) );
  OAI21_X1 U16705 ( .B1(n15624), .B2(n14222), .A(n13557), .ZN(n13558) );
  OAI211_X1 U16706 ( .C1(n19795), .C2(n14223), .A(n15632), .B(n13558), .ZN(
        n15621) );
  OAI221_X1 U16707 ( .B1(n15621), .B2(n19816), .C1(n15621), .C2(n15624), .A(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n13560) );
  OAI21_X1 U16708 ( .B1(n19798), .B2(n13561), .A(n13560), .ZN(n13564) );
  NAND3_X1 U16709 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n19816), .ZN(n15651) );
  NAND2_X1 U16710 ( .A1(n19824), .A2(n15651), .ZN(n15623) );
  NAND2_X1 U16711 ( .A1(n13562), .A2(n19809), .ZN(n15674) );
  NOR4_X1 U16712 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15624), .A3(
        n14222), .A4(n15674), .ZN(n13563) );
  AOI211_X1 U16713 ( .C1(n19807), .C2(n15513), .A(n13564), .B(n13563), .ZN(
        n13565) );
  OAI21_X1 U16714 ( .B1(n15569), .B2(n19820), .A(n13565), .ZN(P1_U3019) );
  NAND2_X1 U16715 ( .A1(n18348), .A2(n18339), .ZN(n18343) );
  AOI22_X1 U16716 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13569) );
  INV_X2 U16717 ( .A(n9680), .ZN(n16682) );
  NOR2_X2 U16718 ( .A1(n13573), .A2(n18205), .ZN(n15269) );
  AOI22_X1 U16719 ( .A1(n16682), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9620), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13568) );
  AOI22_X1 U16720 ( .A1(n15219), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9622), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13567) );
  AOI22_X1 U16721 ( .A1(n16733), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9642), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13566) );
  NAND4_X1 U16722 ( .A1(n13569), .A2(n13568), .A3(n13567), .A4(n13566), .ZN(
        n13581) );
  INV_X2 U16723 ( .A(n15251), .ZN(n16435) );
  AOI22_X1 U16724 ( .A1(n15248), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n16610), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13579) );
  AOI22_X1 U16725 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9629), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13578) );
  AOI22_X1 U16726 ( .A1(n9616), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(n9613), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13577) );
  INV_X2 U16727 ( .A(n9683), .ZN(n16723) );
  AOI22_X1 U16728 ( .A1(n16738), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n16723), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13576) );
  NAND4_X1 U16729 ( .A1(n13579), .A2(n13578), .A3(n13577), .A4(n13576), .ZN(
        n13580) );
  AOI22_X1 U16730 ( .A1(n16682), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n16668), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13585) );
  AOI22_X1 U16731 ( .A1(n15219), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13584) );
  AOI22_X1 U16732 ( .A1(n9616), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(n9622), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13583) );
  AOI22_X1 U16733 ( .A1(n16508), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9640), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13582) );
  NAND4_X1 U16734 ( .A1(n13585), .A2(n13584), .A3(n13583), .A4(n13582), .ZN(
        n13591) );
  AOI22_X1 U16735 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n16723), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13589) );
  AOI22_X1 U16736 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9629), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13588) );
  AOI22_X1 U16737 ( .A1(n9612), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16738), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13587) );
  AOI22_X1 U16738 ( .A1(n16634), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9620), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13586) );
  NAND4_X1 U16739 ( .A1(n13589), .A2(n13588), .A3(n13587), .A4(n13586), .ZN(
        n13590) );
  INV_X4 U16740 ( .A(n16435), .ZN(n16634) );
  AOI22_X1 U16741 ( .A1(n15248), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n16634), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13595) );
  AOI22_X1 U16742 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(n9620), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13594) );
  AOI22_X1 U16743 ( .A1(n16682), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n16738), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13593) );
  AOI22_X1 U16744 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9642), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13592) );
  NAND4_X1 U16745 ( .A1(n13595), .A2(n13594), .A3(n13593), .A4(n13592), .ZN(
        n13601) );
  INV_X2 U16746 ( .A(n9683), .ZN(n16741) );
  AOI22_X1 U16747 ( .A1(n16508), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n16741), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13599) );
  AOI22_X1 U16748 ( .A1(n15219), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9629), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13598) );
  AOI22_X1 U16749 ( .A1(n9612), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13597) );
  AOI22_X1 U16750 ( .A1(n9616), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n15241), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13596) );
  NAND4_X1 U16751 ( .A1(n13599), .A2(n13598), .A3(n13597), .A4(n13596), .ZN(
        n13600) );
  AOI22_X1 U16752 ( .A1(n9629), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n16721), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13605) );
  AOI22_X1 U16753 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13604) );
  AOI22_X1 U16754 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n16716), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13603) );
  AOI22_X1 U16755 ( .A1(n9622), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(n9641), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13602) );
  NAND4_X1 U16756 ( .A1(n13605), .A2(n13604), .A3(n13603), .A4(n13602), .ZN(
        n13612) );
  AOI22_X1 U16757 ( .A1(n9630), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(n9616), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13610) );
  AOI22_X1 U16758 ( .A1(n16733), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9613), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13609) );
  AOI22_X1 U16759 ( .A1(n16723), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n16634), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13608) );
  AOI22_X1 U16761 ( .A1(n15219), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n16739), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13607) );
  NAND4_X1 U16762 ( .A1(n13610), .A2(n13609), .A3(n13608), .A4(n13607), .ZN(
        n13611) );
  NAND2_X1 U16763 ( .A1(n16111), .A2(n16890), .ZN(n13662) );
  AOI22_X1 U16764 ( .A1(n16682), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9620), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13616) );
  AOI22_X1 U16765 ( .A1(n9616), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n15241), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13615) );
  AOI22_X1 U16766 ( .A1(n16634), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13614) );
  AOI22_X1 U16767 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(n9642), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13613) );
  NAND4_X1 U16768 ( .A1(n13616), .A2(n13615), .A3(n13614), .A4(n13613), .ZN(
        n13622) );
  AOI22_X1 U16769 ( .A1(n15219), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n16739), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13620) );
  AOI22_X1 U16770 ( .A1(n9611), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n16723), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13619) );
  AOI22_X1 U16771 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9629), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13618) );
  AOI22_X1 U16772 ( .A1(n16508), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n16738), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13617) );
  NAND4_X1 U16773 ( .A1(n13620), .A2(n13619), .A3(n13618), .A4(n13617), .ZN(
        n13621) );
  AOI22_X1 U16774 ( .A1(n15219), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9621), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13632) );
  AOI22_X1 U16775 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n16634), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13631) );
  AOI22_X1 U16776 ( .A1(n16716), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13623) );
  OAI21_X1 U16777 ( .B1(n9679), .B2(n20623), .A(n13623), .ZN(n13629) );
  AOI22_X1 U16778 ( .A1(n16508), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n16663), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13627) );
  AOI22_X1 U16779 ( .A1(n16623), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n16668), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13626) );
  AOI22_X1 U16780 ( .A1(n16723), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9640), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13625) );
  AOI22_X1 U16781 ( .A1(n16738), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n15241), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13624) );
  NAND4_X1 U16782 ( .A1(n13627), .A2(n13626), .A3(n13625), .A4(n13624), .ZN(
        n13628) );
  AOI211_X1 U16783 ( .C1(n9613), .C2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A(
        n13629), .B(n13628), .ZN(n13630) );
  NAND3_X1 U16784 ( .A1(n13632), .A2(n13631), .A3(n13630), .ZN(n15206) );
  NAND2_X1 U16785 ( .A1(n16784), .A2(n15206), .ZN(n13656) );
  AOI22_X1 U16786 ( .A1(n16508), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n15241), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13642) );
  AOI22_X1 U16787 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n16723), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13641) );
  AOI22_X1 U16788 ( .A1(n16663), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n16610), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13633) );
  OAI21_X1 U16789 ( .B1(n9680), .B2(n20650), .A(n13633), .ZN(n13639) );
  AOI22_X1 U16790 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13637) );
  AOI22_X1 U16791 ( .A1(n15219), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n16668), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13636) );
  AOI22_X1 U16792 ( .A1(n16738), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9620), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13635) );
  AOI22_X1 U16793 ( .A1(n9611), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9640), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13634) );
  NAND4_X1 U16794 ( .A1(n13637), .A2(n13636), .A3(n13635), .A4(n13634), .ZN(
        n13638) );
  AOI211_X2 U16795 ( .C1(n9616), .C2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n13639), .B(n13638), .ZN(n13640) );
  NAND2_X1 U16796 ( .A1(n17772), .A2(n17760), .ZN(n13654) );
  AOI22_X1 U16797 ( .A1(n16723), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9622), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13646) );
  AOI22_X1 U16798 ( .A1(n9629), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n16738), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13645) );
  AOI22_X1 U16799 ( .A1(n16716), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13644) );
  AOI22_X1 U16800 ( .A1(n9642), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n16634), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13643) );
  NAND4_X1 U16801 ( .A1(n13646), .A2(n13645), .A3(n13644), .A4(n13643), .ZN(
        n13652) );
  AOI22_X1 U16802 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n16508), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13650) );
  AOI22_X1 U16803 ( .A1(n15219), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n16722), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13649) );
  AOI22_X1 U16804 ( .A1(n9616), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(n9613), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13648) );
  AOI22_X1 U16805 ( .A1(n16682), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n16668), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13647) );
  NAND4_X1 U16806 ( .A1(n13650), .A2(n13649), .A3(n13648), .A4(n13647), .ZN(
        n13651) );
  OAI211_X1 U16807 ( .C1(n17778), .C2(n15423), .A(n17741), .B(n17736), .ZN(
        n13689) );
  OAI21_X1 U16808 ( .B1(n15205), .B2(n13664), .A(n13689), .ZN(n13661) );
  INV_X1 U16809 ( .A(n13662), .ZN(n13660) );
  NOR2_X1 U16810 ( .A1(n17741), .A2(n17736), .ZN(n13666) );
  OR2_X1 U16811 ( .A1(n15200), .A2(n13666), .ZN(n13684) );
  INV_X1 U16812 ( .A(n15200), .ZN(n17748) );
  AOI21_X1 U16813 ( .B1(n13654), .B2(n13656), .A(n13653), .ZN(n13655) );
  AOI21_X1 U16814 ( .B1(n13656), .B2(n13684), .A(n13655), .ZN(n13659) );
  INV_X1 U16815 ( .A(n13656), .ZN(n13657) );
  OAI21_X1 U16816 ( .B1(n17778), .B2(n13657), .A(n15093), .ZN(n13658) );
  OAI211_X1 U16817 ( .C1(n13660), .C2(n13663), .A(n13659), .B(n13658), .ZN(
        n13688) );
  AOI21_X1 U16818 ( .B1(n13663), .B2(n13661), .A(n13688), .ZN(n15195) );
  NAND2_X1 U16819 ( .A1(n13665), .A2(n15195), .ZN(n15194) );
  NOR2_X1 U16820 ( .A1(n17772), .A2(n16784), .ZN(n13685) );
  NAND2_X1 U16821 ( .A1(n18180), .A2(n13685), .ZN(n15092) );
  NOR2_X1 U16822 ( .A1(n13662), .A2(n15092), .ZN(n13667) );
  NAND4_X2 U16823 ( .A1(n15197), .A2(n17766), .A3(n13664), .A4(n17736), .ZN(
        n16976) );
  NAND2_X1 U16824 ( .A1(n13665), .A2(n15200), .ZN(n13687) );
  NAND2_X1 U16825 ( .A1(n16976), .A2(n13687), .ZN(n16094) );
  NAND2_X1 U16826 ( .A1(n13666), .A2(n16094), .ZN(n13691) );
  OAI21_X1 U16827 ( .B1(n13700), .B2(n18362), .A(n18228), .ZN(n13668) );
  NAND2_X1 U16828 ( .A1(n18216), .A2(n13668), .ZN(n18227) );
  NOR2_X1 U16829 ( .A1(n18343), .A2(n18227), .ZN(n13699) );
  INV_X1 U16830 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18403) );
  INV_X1 U16831 ( .A(n18235), .ZN(n18243) );
  AOI22_X1 U16832 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n17987), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18362), .ZN(n13695) );
  XOR2_X1 U16833 ( .A(n13693), .B(n13695), .Z(n13681) );
  AOI22_X1 U16834 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(n18209), .B2(n18355), .ZN(
        n13676) );
  NOR2_X1 U16835 ( .A1(n13677), .A2(n13676), .ZN(n13670) );
  NOR2_X1 U16836 ( .A1(n13671), .A2(n18345), .ZN(n13674) );
  AOI22_X1 U16837 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18228), .B1(
        n13671), .B2(n18345), .ZN(n13675) );
  OAI21_X1 U16838 ( .B1(n18196), .B2(n13674), .A(n13675), .ZN(n13672) );
  NAND2_X1 U16839 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18228), .ZN(
        n13673) );
  OAI22_X1 U16840 ( .A1(n13675), .A2(n18196), .B1(n13674), .B2(n13673), .ZN(
        n13692) );
  XOR2_X1 U16841 ( .A(n13677), .B(n13676), .Z(n15198) );
  INV_X1 U16842 ( .A(n15198), .ZN(n13679) );
  INV_X1 U16843 ( .A(n13680), .ZN(n13678) );
  NAND2_X1 U16844 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18385) );
  NAND2_X1 U16845 ( .A1(n18222), .A2(n18385), .ZN(n13696) );
  NOR3_X1 U16846 ( .A1(n13685), .A2(n13684), .A3(n13683), .ZN(n13686) );
  OAI21_X1 U16847 ( .B1(n17760), .B2(n15423), .A(n13686), .ZN(n15211) );
  OAI21_X1 U16848 ( .B1(n15211), .B2(n13688), .A(n13687), .ZN(n13690) );
  NAND2_X1 U16849 ( .A1(n13690), .A2(n13689), .ZN(n15203) );
  OAI211_X1 U16850 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n20637), .B(n18328), .ZN(n18262) );
  INV_X1 U16851 ( .A(n18262), .ZN(n18390) );
  NAND2_X1 U16852 ( .A1(n18391), .A2(n13691), .ZN(n15196) );
  NAND3_X1 U16853 ( .A1(n18390), .A2(n18215), .A3(n15196), .ZN(n16936) );
  AOI211_X1 U16854 ( .C1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .C2(n18369), .A(
        n13693), .B(n13692), .ZN(n15199) );
  AOI21_X1 U16855 ( .B1(n13695), .B2(n15199), .A(n13694), .ZN(n18219) );
  INV_X1 U16856 ( .A(n18219), .ZN(n15917) );
  NOR2_X1 U16857 ( .A1(n17760), .A2(n15206), .ZN(n18181) );
  NAND3_X1 U16858 ( .A1(n15197), .A2(n15205), .A3(n18181), .ZN(n15193) );
  OAI21_X1 U16859 ( .B1(n13696), .B2(n16936), .A(n15095), .ZN(n13697) );
  NOR3_X1 U16860 ( .A1(n15422), .A2(n15203), .A3(n13697), .ZN(n18186) );
  NAND2_X1 U16861 ( .A1(n18394), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n17735) );
  INV_X1 U16862 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n17725) );
  NAND3_X1 U16863 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATE2_REG_0__SCAN_IN), .ZN(n18337)
         );
  OR2_X1 U16864 ( .A1(n17725), .A2(n18337), .ZN(n13698) );
  OAI211_X1 U16865 ( .C1(n18243), .C2(n18186), .A(n17735), .B(n13698), .ZN(
        n18367) );
  INV_X1 U16866 ( .A(n18367), .ZN(n18370) );
  MUX2_X1 U16867 ( .A(n13699), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n18370), .Z(P3_U3284) );
  OAI211_X1 U16868 ( .C1(n13700), .C2(n18362), .A(n15218), .B(n18228), .ZN(
        n17724) );
  NOR2_X1 U16869 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n17724), .ZN(n13701) );
  NOR2_X1 U16870 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18397) );
  AOI21_X1 U16871 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(n18397), .ZN(n18253) );
  OAI21_X1 U16872 ( .B1(n13701), .B2(n18337), .A(n17896), .ZN(n17730) );
  INV_X1 U16873 ( .A(n17730), .ZN(n13703) );
  INV_X1 U16874 ( .A(n18343), .ZN(n18404) );
  NOR2_X1 U16875 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n16088) );
  NOR2_X1 U16876 ( .A1(n18404), .A2(n16088), .ZN(n18388) );
  INV_X1 U16877 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n16113) );
  NOR2_X1 U16878 ( .A1(n18348), .A2(n16113), .ZN(n17044) );
  OAI22_X1 U16879 ( .A1(n17988), .A2(n18339), .B1(n18388), .B2(n17044), .ZN(
        n13702) );
  INV_X1 U16880 ( .A(n13702), .ZN(n15187) );
  NOR2_X1 U16881 ( .A1(n13703), .A2(n15187), .ZN(n13705) );
  NAND3_X1 U16882 ( .A1(n18403), .A2(n18339), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18035) );
  INV_X1 U16883 ( .A(n18035), .ZN(n15188) );
  NOR2_X1 U16884 ( .A1(n18339), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n17785) );
  OR2_X1 U16885 ( .A1(n17785), .A2(n13703), .ZN(n15185) );
  OR2_X1 U16886 ( .A1(n15188), .A2(n15185), .ZN(n13704) );
  MUX2_X1 U16887 ( .A(n13705), .B(n13704), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  NOR2_X1 U16888 ( .A1(n13707), .A2(n13706), .ZN(n13711) );
  OAI22_X1 U16889 ( .A1(n13709), .A2(n19525), .B1(n19537), .B2(n13708), .ZN(
        n13710) );
  OAI21_X1 U16890 ( .B1(n13711), .B2(n13710), .A(n19530), .ZN(n13712) );
  OAI21_X1 U16891 ( .B1(n19530), .B2(n13713), .A(n13712), .ZN(P2_U3601) );
  INV_X1 U16892 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n13714) );
  NAND2_X1 U16893 ( .A1(n13715), .A2(n13714), .ZN(n13717) );
  OR2_X1 U16894 ( .A1(n13887), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13716) );
  NAND2_X1 U16895 ( .A1(n13716), .A2(n13717), .ZN(n13899) );
  MUX2_X1 U16896 ( .A(n13717), .B(n13899), .S(n12372), .Z(n13722) );
  OR2_X1 U16897 ( .A1(n13718), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n13721) );
  INV_X1 U16898 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14103) );
  NAND2_X1 U16899 ( .A1(n12302), .A2(n14103), .ZN(n13719) );
  OAI211_X1 U16900 ( .C1(P1_EBX_REG_28__SCAN_IN), .C2(n13886), .A(n13719), .B(
        n12352), .ZN(n13720) );
  NAND2_X1 U16901 ( .A1(n13721), .A2(n13720), .ZN(n13922) );
  AOI21_X1 U16902 ( .B1(n13722), .B2(n9653), .A(n9978), .ZN(n14260) );
  AOI22_X1 U16903 ( .A1(n14260), .A2(n19705), .B1(n14004), .B2(
        P1_EBX_REG_29__SCAN_IN), .ZN(n13723) );
  OAI21_X1 U16904 ( .B1(n13737), .B2(n14024), .A(n13723), .ZN(P1_U2843) );
  AOI22_X1 U16905 ( .A1(n14069), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n15545), .ZN(n13726) );
  NOR3_X4 U16906 ( .A1(n15545), .A2(n13724), .A3(n19873), .ZN(n14070) );
  AOI22_X1 U16907 ( .A1(n14071), .A2(DATAI_29_), .B1(n14070), .B2(n19760), 
        .ZN(n13725) );
  OAI211_X1 U16908 ( .C1(n13737), .C2(n19714), .A(n13726), .B(n13725), .ZN(
        P1_U2875) );
  INV_X1 U16909 ( .A(n13727), .ZN(n13728) );
  NAND2_X1 U16910 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n13729) );
  NOR2_X1 U16911 ( .A1(n13728), .A2(n13729), .ZN(n13890) );
  NOR2_X1 U16912 ( .A1(n13890), .A2(n19669), .ZN(n13928) );
  INV_X1 U16913 ( .A(n13729), .ZN(n13730) );
  NAND2_X1 U16914 ( .A1(n13918), .A2(n13730), .ZN(n13908) );
  AOI22_X1 U16915 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19675), .B1(
        n19644), .B2(n13731), .ZN(n13733) );
  NAND2_X1 U16916 ( .A1(n19687), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n13732) );
  OAI211_X1 U16917 ( .C1(n13908), .C2(P1_REIP_REG_29__SCAN_IN), .A(n13733), 
        .B(n13732), .ZN(n13734) );
  AOI21_X1 U16918 ( .B1(n13928), .B2(P1_REIP_REG_29__SCAN_IN), .A(n13734), 
        .ZN(n13736) );
  NAND2_X1 U16919 ( .A1(n14260), .A2(n19686), .ZN(n13735) );
  OAI211_X1 U16920 ( .C1(n13737), .C2(n15470), .A(n13736), .B(n13735), .ZN(
        P1_U2811) );
  INV_X1 U16921 ( .A(n13738), .ZN(n13739) );
  NAND2_X1 U16922 ( .A1(n13739), .A2(n9682), .ZN(n13740) );
  NAND2_X1 U16923 ( .A1(n13839), .A2(n13740), .ZN(n15729) );
  NAND2_X1 U16924 ( .A1(n13743), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13744) );
  OR2_X1 U16925 ( .A1(n13746), .A2(n13745), .ZN(n13747) );
  NAND2_X1 U16926 ( .A1(n13757), .A2(n13747), .ZN(n18577) );
  NOR2_X1 U16927 ( .A1(n18577), .A2(n13327), .ZN(n13751) );
  AND2_X1 U16928 ( .A1(n13751), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15829) );
  INV_X1 U16929 ( .A(n13748), .ZN(n13749) );
  XNOR2_X1 U16930 ( .A(n13750), .B(n13749), .ZN(n18589) );
  AND2_X1 U16931 ( .A1(n18589), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15825) );
  INV_X1 U16932 ( .A(n13751), .ZN(n13753) );
  NAND2_X1 U16933 ( .A1(n13753), .A2(n13752), .ZN(n15828) );
  OR2_X1 U16934 ( .A1(n18589), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15826) );
  AND2_X1 U16935 ( .A1(n15828), .A2(n15826), .ZN(n13754) );
  NAND2_X1 U16936 ( .A1(n18911), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n13756) );
  XNOR2_X1 U16937 ( .A(n13757), .B(n13756), .ZN(n18566) );
  NAND2_X1 U16938 ( .A1(n18566), .A2(n12224), .ZN(n13763) );
  INV_X1 U16939 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15061) );
  AND2_X1 U16940 ( .A1(n13763), .A2(n15061), .ZN(n15056) );
  NAND3_X1 U16941 ( .A1(n13759), .A2(n18911), .A3(P2_EBX_REG_10__SCAN_IN), 
        .ZN(n13758) );
  OAI211_X1 U16942 ( .C1(n13759), .C2(P2_EBX_REG_10__SCAN_IN), .A(n13834), .B(
        n13758), .ZN(n18555) );
  OR2_X1 U16943 ( .A1(n18555), .A2(n13327), .ZN(n13761) );
  INV_X1 U16944 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n13760) );
  NAND2_X1 U16945 ( .A1(n13761), .A2(n13760), .ZN(n15040) );
  NAND2_X1 U16946 ( .A1(n12224), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13762) );
  OR2_X1 U16947 ( .A1(n18555), .A2(n13762), .ZN(n15039) );
  OR2_X1 U16948 ( .A1(n13763), .A2(n15061), .ZN(n15052) );
  NAND2_X1 U16949 ( .A1(n15039), .A2(n15052), .ZN(n13764) );
  AND3_X1 U16950 ( .A1(n18911), .A2(P2_EBX_REG_11__SCAN_IN), .A3(n13765), .ZN(
        n13766) );
  OR2_X1 U16951 ( .A1(n13767), .A2(n13766), .ZN(n13768) );
  NAND2_X1 U16952 ( .A1(n10282), .A2(n12224), .ZN(n15025) );
  INV_X1 U16953 ( .A(n15025), .ZN(n13769) );
  INV_X1 U16954 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15030) );
  OR2_X1 U16955 ( .A1(n13771), .A2(n13770), .ZN(n13772) );
  NAND2_X1 U16956 ( .A1(n13793), .A2(n13772), .ZN(n18531) );
  NOR2_X1 U16957 ( .A1(n18531), .A2(n13327), .ZN(n13773) );
  AND2_X1 U16958 ( .A1(n13773), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15802) );
  INV_X1 U16959 ( .A(n13773), .ZN(n13775) );
  INV_X1 U16960 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n13774) );
  INV_X1 U16961 ( .A(n13806), .ZN(n13776) );
  AOI21_X1 U16962 ( .B1(n13776), .B2(n12224), .A(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14740) );
  NAND2_X1 U16963 ( .A1(n18911), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n13777) );
  XNOR2_X1 U16964 ( .A(n13781), .B(n13777), .ZN(n18445) );
  INV_X1 U16965 ( .A(n18445), .ZN(n13778) );
  AOI21_X1 U16966 ( .B1(n13778), .B2(n12224), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14749) );
  NOR2_X1 U16967 ( .A1(n13802), .A2(n13779), .ZN(n13780) );
  OR2_X1 U16968 ( .A1(n13781), .A2(n13780), .ZN(n18453) );
  INV_X1 U16969 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14956) );
  OAI21_X1 U16970 ( .B1(n18453), .B2(n13327), .A(n14956), .ZN(n14762) );
  MUX2_X1 U16971 ( .A(n13783), .B(P2_EBX_REG_16__SCAN_IN), .S(n13782), .Z(
        n13784) );
  AND2_X1 U16972 ( .A1(n13784), .A2(n13834), .ZN(n18487) );
  NAND2_X1 U16973 ( .A1(n18487), .A2(n12224), .ZN(n13811) );
  XNOR2_X1 U16974 ( .A(n13811), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14790) );
  NAND2_X1 U16975 ( .A1(n13786), .A2(n13785), .ZN(n13787) );
  NAND2_X1 U16976 ( .A1(n13801), .A2(n13787), .ZN(n18476) );
  INV_X1 U16977 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14985) );
  OAI21_X1 U16978 ( .B1(n18476), .B2(n13327), .A(n14985), .ZN(n14736) );
  INV_X1 U16979 ( .A(n13788), .ZN(n13789) );
  XNOR2_X1 U16980 ( .A(n13790), .B(n13789), .ZN(n18495) );
  NAND2_X1 U16981 ( .A1(n18495), .A2(n12224), .ZN(n13791) );
  INV_X1 U16982 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15004) );
  NAND2_X1 U16983 ( .A1(n13791), .A2(n15004), .ZN(n14801) );
  AND2_X1 U16984 ( .A1(n13793), .A2(n13792), .ZN(n13794) );
  OR2_X1 U16985 ( .A1(n13794), .A2(n13798), .ZN(n18517) );
  INV_X1 U16986 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n13795) );
  OAI21_X1 U16987 ( .B1(n18517), .B2(n13327), .A(n13795), .ZN(n14809) );
  INV_X1 U16988 ( .A(n13796), .ZN(n13797) );
  XNOR2_X1 U16989 ( .A(n13798), .B(n13797), .ZN(n18507) );
  NAND2_X1 U16990 ( .A1(n18507), .A2(n12224), .ZN(n13799) );
  INV_X1 U16991 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15861) );
  NAND2_X1 U16992 ( .A1(n13799), .A2(n15861), .ZN(n15794) );
  AND4_X1 U16993 ( .A1(n14736), .A2(n14801), .A3(n14809), .A4(n15794), .ZN(
        n13804) );
  AND2_X1 U16994 ( .A1(n13801), .A2(n13800), .ZN(n13803) );
  OR2_X1 U16995 ( .A1(n13803), .A2(n13802), .ZN(n18467) );
  INV_X1 U16996 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14971) );
  OAI21_X1 U16997 ( .B1(n18467), .B2(n13327), .A(n14971), .ZN(n14771) );
  NAND2_X1 U16998 ( .A1(n12224), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13805) );
  OR2_X1 U16999 ( .A1(n13806), .A2(n13805), .ZN(n14741) );
  INV_X1 U17000 ( .A(n18453), .ZN(n13808) );
  AND2_X1 U17001 ( .A1(n12224), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13807) );
  NAND2_X1 U17002 ( .A1(n13808), .A2(n13807), .ZN(n14761) );
  INV_X1 U17003 ( .A(n18467), .ZN(n13810) );
  AND2_X1 U17004 ( .A1(n12224), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13809) );
  NAND2_X1 U17005 ( .A1(n13810), .A2(n13809), .ZN(n14770) );
  AND2_X1 U17006 ( .A1(n14761), .A2(n14770), .ZN(n14738) );
  INV_X1 U17007 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n20666) );
  NOR2_X1 U17008 ( .A1(n13811), .A2(n20666), .ZN(n14734) );
  INV_X1 U17009 ( .A(n18476), .ZN(n13813) );
  AND2_X1 U17010 ( .A1(n12224), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n13812) );
  NAND2_X1 U17011 ( .A1(n13813), .A2(n13812), .ZN(n14735) );
  AND2_X1 U17012 ( .A1(n12224), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13814) );
  NAND2_X1 U17013 ( .A1(n18495), .A2(n13814), .ZN(n14800) );
  AND2_X1 U17014 ( .A1(n12224), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13815) );
  NAND2_X1 U17015 ( .A1(n18507), .A2(n13815), .ZN(n15793) );
  INV_X1 U17016 ( .A(n18517), .ZN(n13817) );
  AND2_X1 U17017 ( .A1(n12224), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13816) );
  NAND2_X1 U17018 ( .A1(n13817), .A2(n13816), .ZN(n14808) );
  NAND4_X1 U17019 ( .A1(n14735), .A2(n14800), .A3(n15793), .A4(n14808), .ZN(
        n13818) );
  NOR2_X1 U17020 ( .A1(n14734), .A2(n13818), .ZN(n13820) );
  NAND2_X1 U17021 ( .A1(n12224), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13819) );
  NAND4_X1 U17022 ( .A1(n14741), .A2(n14738), .A3(n13820), .A4(n14750), .ZN(
        n13821) );
  NOR2_X1 U17023 ( .A1(n13822), .A2(n13327), .ZN(n13823) );
  NOR2_X1 U17024 ( .A1(n13823), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14915) );
  NAND2_X1 U17025 ( .A1(n13823), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14914) );
  INV_X1 U17026 ( .A(n13824), .ZN(n13825) );
  OAI21_X1 U17027 ( .B1(n13825), .B2(n9758), .A(n13828), .ZN(n15770) );
  NOR2_X1 U17028 ( .A1(n15770), .A2(n13327), .ZN(n13826) );
  XOR2_X1 U17029 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n13826), .Z(
        n14724) );
  INV_X1 U17030 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n13827) );
  INV_X1 U17031 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14721) );
  NOR2_X1 U17032 ( .A1(n9614), .A2(n10064), .ZN(n13829) );
  MUX2_X1 U17033 ( .A(n10064), .B(n13829), .S(n13828), .Z(n13830) );
  NOR2_X1 U17034 ( .A1(n13830), .A2(n13767), .ZN(n15755) );
  NAND2_X1 U17035 ( .A1(n15755), .A2(n12224), .ZN(n14714) );
  NOR2_X1 U17036 ( .A1(n9684), .A2(n14493), .ZN(n13832) );
  NAND2_X1 U17037 ( .A1(n18911), .A2(n13832), .ZN(n13833) );
  NAND2_X1 U17038 ( .A1(n13834), .A2(n13833), .ZN(n13835) );
  AOI21_X1 U17039 ( .B1(n9684), .B2(n14493), .A(n13835), .ZN(n15745) );
  AND2_X1 U17040 ( .A1(n15745), .A2(n12224), .ZN(n13846) );
  OR2_X1 U17041 ( .A1(n13846), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14705) );
  AND2_X1 U17042 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n13836), .ZN(n13837) );
  AOI21_X1 U17043 ( .B1(n18911), .B2(n13837), .A(n14644), .ZN(n15737) );
  NAND2_X1 U17044 ( .A1(n13838), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13848) );
  OAI21_X1 U17045 ( .B1(n13838), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n13848), .ZN(n14694) );
  INV_X1 U17046 ( .A(n13839), .ZN(n13842) );
  INV_X1 U17047 ( .A(n13840), .ZN(n13841) );
  OAI21_X1 U17048 ( .B1(n13842), .B2(n13841), .A(n13850), .ZN(n15712) );
  NOR2_X1 U17049 ( .A1(n15712), .A2(n13327), .ZN(n14676) );
  OAI21_X1 U17050 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n14676), .ZN(n13844) );
  INV_X1 U17051 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14850) );
  INV_X1 U17052 ( .A(n14676), .ZN(n13843) );
  AOI22_X1 U17053 ( .A1(n13845), .A2(n13844), .B1(n14850), .B2(n13843), .ZN(
        n13849) );
  INV_X1 U17054 ( .A(n13846), .ZN(n13847) );
  INV_X1 U17055 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14886) );
  NAND2_X1 U17056 ( .A1(n14707), .A2(n13848), .ZN(n14672) );
  XOR2_X1 U17057 ( .A(n13851), .B(n13850), .Z(n15701) );
  AOI21_X1 U17058 ( .B1(n15701), .B2(n12224), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14662) );
  NAND2_X1 U17059 ( .A1(n12224), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13852) );
  NOR2_X1 U17060 ( .A1(n13853), .A2(n13852), .ZN(n14642) );
  INV_X1 U17061 ( .A(n14642), .ZN(n13854) );
  INV_X1 U17062 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14832) );
  NAND2_X1 U17063 ( .A1(n13857), .A2(n13856), .ZN(n13858) );
  XNOR2_X1 U17064 ( .A(n13865), .B(n13327), .ZN(n13861) );
  INV_X1 U17065 ( .A(n13861), .ZN(n13862) );
  NAND2_X1 U17066 ( .A1(n13863), .A2(n13862), .ZN(n13864) );
  INV_X1 U17067 ( .A(n13865), .ZN(n13867) );
  NAND2_X1 U17068 ( .A1(n13867), .A2(n12224), .ZN(n13866) );
  XNOR2_X1 U17069 ( .A(n13866), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15834) );
  NAND3_X1 U17070 ( .A1(n13867), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n12224), .ZN(n13868) );
  NOR2_X1 U17071 ( .A1(n13774), .A2(n13795), .ZN(n15015) );
  NOR3_X1 U17072 ( .A1(n15061), .A2(n13760), .A3(n15030), .ZN(n15013) );
  AND2_X1 U17073 ( .A1(n15015), .A2(n15013), .ZN(n15863) );
  NAND2_X1 U17074 ( .A1(n15863), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13874) );
  AND2_X1 U17075 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14774) );
  AND2_X1 U17076 ( .A1(n14774), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14972) );
  NAND2_X1 U17077 ( .A1(n14972), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14732) );
  OR2_X1 U17078 ( .A1(n13874), .A2(n14732), .ZN(n14944) );
  AND2_X1 U17079 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n13875) );
  NAND2_X1 U17080 ( .A1(n13875), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13869) );
  NOR2_X1 U17081 ( .A1(n14944), .A2(n13869), .ZN(n14905) );
  AND2_X1 U17082 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14893) );
  INV_X1 U17083 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14877) );
  INV_X1 U17084 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14851) );
  INV_X1 U17085 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14669) );
  XNOR2_X1 U17086 ( .A(n14668), .B(n14832), .ZN(n14658) );
  NAND3_X1 U17087 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14833) );
  AND2_X1 U17088 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n13879) );
  AOI21_X1 U17089 ( .B1(n14893), .B2(n14905), .A(n15081), .ZN(n13871) );
  NAND2_X1 U17090 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15880) );
  NAND2_X1 U17091 ( .A1(n14943), .A2(n15880), .ZN(n13870) );
  NOR3_X1 U17092 ( .A1(n13871), .A2(n15068), .A3(n14721), .ZN(n14900) );
  OR2_X1 U17093 ( .A1(n14900), .A2(n15028), .ZN(n14887) );
  OAI21_X1 U17094 ( .B1(n15028), .B2(n13879), .A(n14887), .ZN(n14861) );
  AOI21_X1 U17095 ( .B1(n14833), .B2(n18837), .A(n14861), .ZN(n14824) );
  NOR2_X1 U17096 ( .A1(n14824), .A2(n14832), .ZN(n13883) );
  NOR2_X1 U17097 ( .A1(n18600), .A2(n13872), .ZN(n14654) );
  NAND2_X1 U17098 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13873), .ZN(
        n15881) );
  INV_X1 U17099 ( .A(n13874), .ZN(n14968) );
  NAND2_X1 U17100 ( .A1(n15862), .A2(n14968), .ZN(n14992) );
  INV_X1 U17101 ( .A(n13875), .ZN(n13876) );
  NOR2_X1 U17102 ( .A1(n13877), .A2(n14935), .ZN(n14924) );
  AND2_X1 U17103 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n14924), .ZN(
        n13878) );
  NAND2_X1 U17104 ( .A1(n14871), .A2(n13879), .ZN(n14863) );
  NOR3_X1 U17105 ( .A1(n14863), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n14833), .ZN(n13880) );
  OAI21_X1 U17106 ( .B1(n14656), .B2(n18839), .A(n13881), .ZN(n13882) );
  AOI211_X1 U17107 ( .C1(n14658), .C2(n18849), .A(n13883), .B(n13882), .ZN(
        n13884) );
  OAI21_X1 U17108 ( .B1(n14660), .B2(n18859), .A(n13884), .ZN(P2_U3016) );
  AND2_X1 U17109 ( .A1(n13886), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13885) );
  AOI21_X1 U17110 ( .B1(n13887), .B2(P1_EBX_REG_30__SCAN_IN), .A(n13885), .ZN(
        n13902) );
  MUX2_X1 U17111 ( .A(n13902), .B(n12372), .S(n13898), .Z(n13889) );
  AOI22_X1 U17112 ( .A1(n13887), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n13886), .ZN(n13888) );
  NAND2_X1 U17113 ( .A1(n14089), .A2(n19659), .ZN(n13897) );
  AND2_X1 U17114 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n13892) );
  AOI21_X1 U17115 ( .B1(n13890), .B2(n13892), .A(n19669), .ZN(n13912) );
  INV_X1 U17116 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n13972) );
  INV_X1 U17117 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13891) );
  OAI22_X1 U17118 ( .A1(n19662), .A2(n13972), .B1(n13891), .B2(n19691), .ZN(
        n13895) );
  INV_X1 U17119 ( .A(n13892), .ZN(n13893) );
  NOR3_X1 U17120 ( .A1(n13908), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n13893), 
        .ZN(n13894) );
  AOI211_X1 U17121 ( .C1(n13912), .C2(P1_REIP_REG_31__SCAN_IN), .A(n13895), 
        .B(n13894), .ZN(n13896) );
  OAI211_X1 U17122 ( .C1(n14220), .C2(n19681), .A(n13897), .B(n13896), .ZN(
        P1_U2809) );
  NAND2_X1 U17123 ( .A1(n13898), .A2(n9692), .ZN(n13901) );
  OR2_X1 U17124 ( .A1(n9653), .A2(n13899), .ZN(n13900) );
  NAND2_X1 U17125 ( .A1(n13901), .A2(n13900), .ZN(n13904) );
  INV_X1 U17126 ( .A(n13902), .ZN(n13903) );
  XNOR2_X1 U17127 ( .A(n13904), .B(n13903), .ZN(n14251) );
  NAND2_X1 U17128 ( .A1(n14097), .A2(n19659), .ZN(n13914) );
  INV_X1 U17129 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20502) );
  INV_X1 U17130 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n13907) );
  OAI21_X1 U17131 ( .B1(n13908), .B2(n20502), .A(n13907), .ZN(n13911) );
  INV_X1 U17132 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n13973) );
  AOI22_X1 U17133 ( .A1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19675), .B1(
        n19644), .B2(n14093), .ZN(n13909) );
  OAI21_X1 U17134 ( .B1(n19662), .B2(n13973), .A(n13909), .ZN(n13910) );
  AOI21_X1 U17135 ( .B1(n13912), .B2(n13911), .A(n13910), .ZN(n13913) );
  OAI211_X1 U17136 ( .C1(n19681), .C2(n14251), .A(n13914), .B(n13913), .ZN(
        P1_U2810) );
  AOI21_X1 U17137 ( .B1(n13917), .B2(n13916), .A(n13915), .ZN(n14109) );
  INV_X1 U17138 ( .A(n14109), .ZN(n14031) );
  INV_X1 U17139 ( .A(n13918), .ZN(n13920) );
  INV_X1 U17140 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n13919) );
  OAI21_X1 U17141 ( .B1(n13920), .B2(n20496), .A(n13919), .ZN(n13927) );
  INV_X1 U17142 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n13974) );
  AOI22_X1 U17143 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19675), .B1(
        n19644), .B2(n14105), .ZN(n13921) );
  OAI21_X1 U17144 ( .B1(n19662), .B2(n13974), .A(n13921), .ZN(n13926) );
  OR2_X1 U17145 ( .A1(n13923), .A2(n13922), .ZN(n13924) );
  NAND2_X1 U17146 ( .A1(n9653), .A2(n13924), .ZN(n14273) );
  NOR2_X1 U17147 ( .A1(n14273), .A2(n19681), .ZN(n13925) );
  AOI211_X1 U17148 ( .C1(n13928), .C2(n13927), .A(n13926), .B(n13925), .ZN(
        n13929) );
  OAI21_X1 U17149 ( .B1(n14031), .B2(n15470), .A(n13929), .ZN(P1_U2812) );
  AOI21_X1 U17150 ( .B1(n13931), .B2(n13978), .A(n12276), .ZN(n14127) );
  INV_X1 U17151 ( .A(n14127), .ZN(n14039) );
  AOI21_X1 U17152 ( .B1(n13933), .B2(n13982), .A(n13932), .ZN(n14286) );
  INV_X1 U17153 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n13935) );
  NOR2_X1 U17154 ( .A1(n13934), .A2(n13935), .ZN(n13940) );
  NAND2_X1 U17155 ( .A1(n13935), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n13938) );
  AOI22_X1 U17156 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19675), .B1(
        n19644), .B2(n14123), .ZN(n13937) );
  NAND2_X1 U17157 ( .A1(n19687), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n13936) );
  OAI211_X1 U17158 ( .C1(n15429), .C2(n13938), .A(n13937), .B(n13936), .ZN(
        n13939) );
  AOI211_X1 U17159 ( .C1(n14286), .C2(n19686), .A(n13940), .B(n13939), .ZN(
        n13941) );
  OAI21_X1 U17160 ( .B1(n14039), .B2(n15470), .A(n13941), .ZN(P1_U2814) );
  AOI21_X1 U17161 ( .B1(n13943), .B2(n13995), .A(n13942), .ZN(n14151) );
  INV_X1 U17162 ( .A(n13988), .ZN(n13946) );
  NAND2_X1 U17163 ( .A1(n13994), .A2(n13944), .ZN(n13945) );
  NAND2_X1 U17164 ( .A1(n13946), .A2(n13945), .ZN(n14315) );
  OAI22_X1 U17165 ( .A1(n13947), .A2(n19691), .B1(n14149), .B2(n19690), .ZN(
        n13948) );
  AOI21_X1 U17166 ( .B1(n19687), .B2(P1_EBX_REG_23__SCAN_IN), .A(n13948), .ZN(
        n13953) );
  NOR2_X1 U17167 ( .A1(n19669), .A2(n13949), .ZN(n15443) );
  INV_X1 U17168 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n15459) );
  NAND2_X1 U17169 ( .A1(n15450), .A2(n13950), .ZN(n15453) );
  INV_X1 U17170 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n14147) );
  OAI21_X1 U17171 ( .B1(n15459), .B2(n15453), .A(n14147), .ZN(n13951) );
  NAND2_X1 U17172 ( .A1(n15443), .A2(n13951), .ZN(n13952) );
  OAI211_X1 U17173 ( .C1(n14315), .C2(n19681), .A(n13953), .B(n13952), .ZN(
        n13954) );
  AOI21_X1 U17174 ( .B1(n14151), .B2(n19659), .A(n13954), .ZN(n13955) );
  INV_X1 U17175 ( .A(n13955), .ZN(P1_U2817) );
  OAI21_X1 U17176 ( .B1(n13956), .B2(n13957), .A(n9699), .ZN(n15553) );
  NAND2_X1 U17177 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n13960) );
  NAND3_X1 U17178 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n13958), .A3(n15525), 
        .ZN(n15502) );
  INV_X1 U17179 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n13959) );
  OAI21_X1 U17180 ( .B1(n13960), .B2(n15502), .A(n13959), .ZN(n13970) );
  OAI21_X1 U17181 ( .B1(n13963), .B2(n13962), .A(n13961), .ZN(n15485) );
  AND2_X1 U17182 ( .A1(n14021), .A2(n13964), .ZN(n13965) );
  OR2_X1 U17183 ( .A1(n13965), .A2(n14016), .ZN(n14376) );
  NOR2_X1 U17184 ( .A1(n19681), .A2(n14376), .ZN(n13969) );
  INV_X1 U17185 ( .A(n15554), .ZN(n13967) );
  AOI22_X1 U17186 ( .A1(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19675), .B1(
        P1_EBX_REG_17__SCAN_IN), .B2(n19687), .ZN(n13966) );
  OAI211_X1 U17187 ( .C1(n19690), .C2(n13967), .A(n19653), .B(n13966), .ZN(
        n13968) );
  AOI211_X1 U17188 ( .C1(n13970), .C2(n15485), .A(n13969), .B(n13968), .ZN(
        n13971) );
  OAI21_X1 U17189 ( .B1(n15553), .B2(n15470), .A(n13971), .ZN(P1_U2823) );
  OAI22_X1 U17190 ( .A1(n14220), .A2(n14025), .B1(n13972), .B2(n19710), .ZN(
        P1_U2841) );
  OAI222_X1 U17191 ( .A1(n14024), .A2(n14028), .B1(n19710), .B2(n13973), .C1(
        n14251), .C2(n14025), .ZN(P1_U2842) );
  OAI222_X1 U17192 ( .A1(n13974), .A2(n19710), .B1(n14025), .B2(n14273), .C1(
        n14031), .C2(n14024), .ZN(P1_U2844) );
  OAI222_X1 U17193 ( .A1(n13975), .A2(n19710), .B1(n14025), .B2(n14282), .C1(
        n14036), .C2(n14024), .ZN(P1_U2845) );
  AOI22_X1 U17194 ( .A1(n14286), .A2(n19705), .B1(n14004), .B2(
        P1_EBX_REG_26__SCAN_IN), .ZN(n13976) );
  OAI21_X1 U17195 ( .B1(n14039), .B2(n14024), .A(n13976), .ZN(P1_U2846) );
  OAI21_X1 U17196 ( .B1(n13977), .B2(n13979), .A(n13978), .ZN(n14133) );
  NAND2_X1 U17197 ( .A1(n13990), .A2(n13980), .ZN(n13981) );
  NAND2_X1 U17198 ( .A1(n13982), .A2(n13981), .ZN(n15437) );
  INV_X1 U17199 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n15428) );
  OAI22_X1 U17200 ( .A1(n15437), .A2(n14025), .B1(n15428), .B2(n19710), .ZN(
        n13983) );
  INV_X1 U17201 ( .A(n13983), .ZN(n13984) );
  OAI21_X1 U17202 ( .B1(n14133), .B2(n14024), .A(n13984), .ZN(P1_U2847) );
  NOR2_X1 U17203 ( .A1(n13942), .A2(n13985), .ZN(n13986) );
  OR2_X1 U17204 ( .A1(n13977), .A2(n13986), .ZN(n14141) );
  INV_X1 U17205 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n15438) );
  OR2_X1 U17206 ( .A1(n13988), .A2(n13987), .ZN(n13989) );
  NAND2_X1 U17207 ( .A1(n13990), .A2(n13989), .ZN(n15448) );
  OAI222_X1 U17208 ( .A1(n14024), .A2(n14141), .B1(n19710), .B2(n15438), .C1(
        n15448), .C2(n14025), .ZN(P1_U2848) );
  INV_X1 U17209 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n13991) );
  INV_X1 U17210 ( .A(n14151), .ZN(n14048) );
  OAI222_X1 U17211 ( .A1(n14315), .A2(n14025), .B1(n13991), .B2(n19710), .C1(
        n14048), .C2(n14024), .ZN(P1_U2849) );
  NAND2_X1 U17212 ( .A1(n14334), .A2(n13992), .ZN(n13993) );
  NAND2_X1 U17213 ( .A1(n13994), .A2(n13993), .ZN(n15454) );
  INV_X1 U17214 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n13998) );
  INV_X1 U17215 ( .A(n13995), .ZN(n13996) );
  AOI21_X1 U17216 ( .B1(n13997), .B2(n14051), .A(n13996), .ZN(n14157) );
  INV_X1 U17217 ( .A(n14157), .ZN(n15455) );
  OAI222_X1 U17218 ( .A1(n15454), .A2(n14025), .B1(n19710), .B2(n13998), .C1(
        n14024), .C2(n15455), .ZN(P1_U2850) );
  NOR2_X1 U17219 ( .A1(n13999), .A2(n14000), .ZN(n14001) );
  OR2_X1 U17220 ( .A1(n14053), .A2(n14001), .ZN(n15471) );
  OR2_X1 U17221 ( .A1(n14010), .A2(n14002), .ZN(n14003) );
  AND2_X1 U17222 ( .A1(n9671), .A2(n14003), .ZN(n15473) );
  AOI22_X1 U17223 ( .A1(n15473), .A2(n19705), .B1(n14004), .B2(
        P1_EBX_REG_20__SCAN_IN), .ZN(n14005) );
  OAI21_X1 U17224 ( .B1(n15471), .B2(n14024), .A(n14005), .ZN(P1_U2852) );
  INV_X1 U17225 ( .A(n14006), .ZN(n14015) );
  INV_X1 U17226 ( .A(n14007), .ZN(n14008) );
  AOI21_X1 U17227 ( .B1(n14016), .B2(n14015), .A(n14008), .ZN(n14009) );
  OR2_X1 U17228 ( .A1(n14010), .A2(n14009), .ZN(n15484) );
  INV_X1 U17229 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14013) );
  AOI21_X1 U17230 ( .B1(n14012), .B2(n14011), .A(n13999), .ZN(n15548) );
  INV_X1 U17231 ( .A(n15548), .ZN(n14062) );
  OAI222_X1 U17232 ( .A1(n14025), .A2(n15484), .B1(n19710), .B2(n14013), .C1(
        n14024), .C2(n14062), .ZN(P1_U2853) );
  XNOR2_X1 U17233 ( .A(n9699), .B(n14014), .ZN(n15491) );
  XNOR2_X1 U17234 ( .A(n14016), .B(n14015), .ZN(n15599) );
  INV_X1 U17235 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14017) );
  OAI222_X1 U17236 ( .A1(n15491), .A2(n14024), .B1(n14025), .B2(n15599), .C1(
        n14017), .C2(n19710), .ZN(P1_U2854) );
  INV_X1 U17237 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14018) );
  OAI222_X1 U17238 ( .A1(n15553), .A2(n14024), .B1(n19710), .B2(n14018), .C1(
        n14376), .C2(n14025), .ZN(P1_U2855) );
  NAND2_X1 U17239 ( .A1(n14401), .A2(n14019), .ZN(n14020) );
  NAND2_X1 U17240 ( .A1(n14021), .A2(n14020), .ZN(n15505) );
  INV_X1 U17241 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n20600) );
  AND2_X1 U17242 ( .A1(n14074), .A2(n14022), .ZN(n14023) );
  OR2_X1 U17243 ( .A1(n14023), .A2(n13956), .ZN(n15495) );
  OAI222_X1 U17244 ( .A1(n15505), .A2(n14025), .B1(n19710), .B2(n20600), .C1(
        n14024), .C2(n15495), .ZN(P1_U2856) );
  AOI22_X1 U17245 ( .A1(n14069), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n15545), .ZN(n14027) );
  AOI22_X1 U17246 ( .A1(n14071), .A2(DATAI_30_), .B1(n14070), .B2(n19762), 
        .ZN(n14026) );
  OAI211_X1 U17247 ( .C1(n14028), .C2(n19714), .A(n14027), .B(n14026), .ZN(
        P1_U2874) );
  AOI22_X1 U17248 ( .A1(n14069), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n15545), .ZN(n14030) );
  MUX2_X1 U17249 ( .A(DATAI_12_), .B(BUF1_REG_12__SCAN_IN), .S(n19836), .Z(
        n19758) );
  AOI22_X1 U17250 ( .A1(n14071), .A2(DATAI_28_), .B1(n14070), .B2(n19758), 
        .ZN(n14029) );
  OAI211_X1 U17251 ( .C1(n14031), .C2(n19714), .A(n14030), .B(n14029), .ZN(
        P1_U2876) );
  INV_X1 U17252 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n15999) );
  OAI22_X1 U17253 ( .A1(n14063), .A2(n15999), .B1(n14032), .B2(n19713), .ZN(
        n14033) );
  INV_X1 U17254 ( .A(n14033), .ZN(n14035) );
  MUX2_X1 U17255 ( .A(DATAI_11_), .B(BUF1_REG_11__SCAN_IN), .S(n19836), .Z(
        n19756) );
  AOI22_X1 U17256 ( .A1(n14071), .A2(DATAI_27_), .B1(n14070), .B2(n19756), 
        .ZN(n14034) );
  OAI211_X1 U17257 ( .C1(n14036), .C2(n19714), .A(n14035), .B(n14034), .ZN(
        P1_U2877) );
  AOI22_X1 U17258 ( .A1(n14069), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n15545), .ZN(n14038) );
  AOI22_X1 U17259 ( .A1(n14071), .A2(DATAI_26_), .B1(n14070), .B2(n19754), 
        .ZN(n14037) );
  OAI211_X1 U17260 ( .C1(n14039), .C2(n19714), .A(n14038), .B(n14037), .ZN(
        P1_U2878) );
  AOI22_X1 U17261 ( .A1(n14069), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n15545), .ZN(n14041) );
  AOI22_X1 U17262 ( .A1(n14071), .A2(DATAI_25_), .B1(n14070), .B2(n19752), 
        .ZN(n14040) );
  OAI211_X1 U17263 ( .C1(n14133), .C2(n19714), .A(n14041), .B(n14040), .ZN(
        P1_U2879) );
  INV_X1 U17264 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n14042) );
  OAI22_X1 U17265 ( .A1(n14063), .A2(n14042), .B1(n12610), .B2(n19713), .ZN(
        n14043) );
  INV_X1 U17266 ( .A(n14043), .ZN(n14045) );
  AOI22_X1 U17267 ( .A1(n14071), .A2(DATAI_24_), .B1(n14070), .B2(n19750), 
        .ZN(n14044) );
  OAI211_X1 U17268 ( .C1(n14141), .C2(n19714), .A(n14045), .B(n14044), .ZN(
        P1_U2880) );
  AOI22_X1 U17269 ( .A1(n14069), .A2(BUF1_REG_23__SCAN_IN), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(n15545), .ZN(n14047) );
  AOI22_X1 U17270 ( .A1(n14071), .A2(DATAI_23_), .B1(n14070), .B2(n19889), 
        .ZN(n14046) );
  OAI211_X1 U17271 ( .C1(n14048), .C2(n19714), .A(n14047), .B(n14046), .ZN(
        P1_U2881) );
  AOI22_X1 U17272 ( .A1(n14069), .A2(BUF1_REG_22__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n15545), .ZN(n14050) );
  AOI22_X1 U17273 ( .A1(n14071), .A2(DATAI_22_), .B1(n14070), .B2(n19880), 
        .ZN(n14049) );
  OAI211_X1 U17274 ( .C1(n15455), .C2(n19714), .A(n14050), .B(n14049), .ZN(
        P1_U2882) );
  OAI21_X1 U17275 ( .B1(n14053), .B2(n14052), .A(n14051), .ZN(n14165) );
  INV_X1 U17276 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n16009) );
  OAI22_X1 U17277 ( .A1(n14063), .A2(n16009), .B1(n12757), .B2(n19713), .ZN(
        n14054) );
  INV_X1 U17278 ( .A(n14054), .ZN(n14056) );
  AOI22_X1 U17279 ( .A1(n14071), .A2(DATAI_21_), .B1(n14070), .B2(n19875), 
        .ZN(n14055) );
  OAI211_X1 U17280 ( .C1(n14165), .C2(n19714), .A(n14056), .B(n14055), .ZN(
        P1_U2883) );
  AOI22_X1 U17281 ( .A1(n14069), .A2(BUF1_REG_20__SCAN_IN), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(n15545), .ZN(n14058) );
  AOI22_X1 U17282 ( .A1(n14071), .A2(DATAI_20_), .B1(n14070), .B2(n19870), 
        .ZN(n14057) );
  OAI211_X1 U17283 ( .C1(n15471), .C2(n19714), .A(n14058), .B(n14057), .ZN(
        P1_U2884) );
  INV_X1 U17284 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16013) );
  OAI22_X1 U17285 ( .A1(n14063), .A2(n16013), .B1(n12753), .B2(n19713), .ZN(
        n14059) );
  INV_X1 U17286 ( .A(n14059), .ZN(n14061) );
  AOI22_X1 U17287 ( .A1(n14071), .A2(DATAI_19_), .B1(n14070), .B2(n19865), 
        .ZN(n14060) );
  OAI211_X1 U17288 ( .C1(n14062), .C2(n19714), .A(n14061), .B(n14060), .ZN(
        P1_U2885) );
  INV_X1 U17289 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n18899) );
  OAI22_X1 U17290 ( .A1(n14063), .A2(n18899), .B1(n12755), .B2(n19713), .ZN(
        n14064) );
  INV_X1 U17291 ( .A(n14064), .ZN(n14066) );
  AOI22_X1 U17292 ( .A1(n14071), .A2(DATAI_18_), .B1(n14070), .B2(n19860), 
        .ZN(n14065) );
  OAI211_X1 U17293 ( .C1(n15491), .C2(n19714), .A(n14066), .B(n14065), .ZN(
        P1_U2886) );
  AOI22_X1 U17294 ( .A1(n14069), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n15545), .ZN(n14068) );
  AOI22_X1 U17295 ( .A1(n14071), .A2(DATAI_17_), .B1(n14070), .B2(n19855), 
        .ZN(n14067) );
  OAI211_X1 U17296 ( .C1(n15553), .C2(n19714), .A(n14068), .B(n14067), .ZN(
        P1_U2887) );
  AOI22_X1 U17297 ( .A1(n14069), .A2(BUF1_REG_16__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n15545), .ZN(n14073) );
  AOI22_X1 U17298 ( .A1(n14071), .A2(DATAI_16_), .B1(n14070), .B2(n19846), 
        .ZN(n14072) );
  OAI211_X1 U17299 ( .C1(n15495), .C2(n19714), .A(n14073), .B(n14072), .ZN(
        P1_U2888) );
  INV_X1 U17300 ( .A(n14074), .ZN(n14075) );
  AOI21_X1 U17301 ( .B1(n14077), .B2(n14076), .A(n14075), .ZN(n15560) );
  INV_X1 U17302 ( .A(n15560), .ZN(n14079) );
  OAI222_X1 U17303 ( .A1(n14079), .A2(n19714), .B1(n19712), .B2(n14078), .C1(
        n19713), .C2(n12646), .ZN(P1_U2889) );
  NOR3_X1 U17304 ( .A1(n14080), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n15572), .ZN(n14083) );
  NAND2_X1 U17305 ( .A1(n15572), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14081) );
  INV_X1 U17306 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20507) );
  NOR2_X1 U17307 ( .A1(n19798), .A2(n20507), .ZN(n14249) );
  AOI21_X1 U17308 ( .B1(n19782), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14249), .ZN(n14086) );
  OAI21_X1 U17309 ( .B1(n19793), .B2(n14087), .A(n14086), .ZN(n14088) );
  AOI21_X1 U17310 ( .B1(n14089), .B2(n19787), .A(n14088), .ZN(n14090) );
  AOI21_X1 U17311 ( .B1(n14092), .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n14091), .ZN(n14259) );
  NAND2_X1 U17312 ( .A1(n15566), .A2(n14093), .ZN(n14094) );
  NAND2_X1 U17313 ( .A1(n19781), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14253) );
  OAI211_X1 U17314 ( .C1(n14190), .C2(n14095), .A(n14094), .B(n14253), .ZN(
        n14096) );
  AOI21_X1 U17315 ( .B1(n14097), .B2(n19787), .A(n14096), .ZN(n14098) );
  OAI21_X1 U17316 ( .B1(n14259), .B2(n19608), .A(n14098), .ZN(P1_U2969) );
  NAND2_X1 U17317 ( .A1(n15572), .A2(n14231), .ZN(n14120) );
  NAND2_X1 U17318 ( .A1(n14146), .A2(n14120), .ZN(n14102) );
  OAI21_X1 U17319 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n14099), .A(
        n14102), .ZN(n14101) );
  INV_X1 U17320 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14279) );
  MUX2_X1 U17321 ( .A(n14279), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n15572), .Z(n14100) );
  OAI211_X1 U17322 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n14102), .A(
        n14101), .B(n14100), .ZN(n14104) );
  XNOR2_X1 U17323 ( .A(n14104), .B(n14103), .ZN(n14274) );
  NAND2_X1 U17324 ( .A1(n15566), .A2(n14105), .ZN(n14106) );
  NAND2_X1 U17325 ( .A1(n19781), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14269) );
  OAI211_X1 U17326 ( .C1(n14190), .C2(n14107), .A(n14106), .B(n14269), .ZN(
        n14108) );
  AOI21_X1 U17327 ( .B1(n14109), .B2(n19787), .A(n14108), .ZN(n14110) );
  OAI21_X1 U17328 ( .B1(n19608), .B2(n14274), .A(n14110), .ZN(P1_U2971) );
  INV_X1 U17329 ( .A(n14111), .ZN(n14113) );
  MUX2_X1 U17330 ( .A(n14113), .B(n14112), .S(n9603), .Z(n14114) );
  NOR2_X1 U17331 ( .A1(n19798), .A2(n20496), .ZN(n14278) );
  AOI21_X1 U17332 ( .B1(n19782), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n14278), .ZN(n14115) );
  OAI21_X1 U17333 ( .B1(n19793), .B2(n14116), .A(n14115), .ZN(n14117) );
  AOI21_X1 U17334 ( .B1(n14118), .B2(n19787), .A(n14117), .ZN(n14119) );
  OAI21_X1 U17335 ( .B1(n19608), .B2(n14283), .A(n14119), .ZN(P1_U2972) );
  OAI211_X1 U17336 ( .C1(n9603), .C2(n14146), .A(n14121), .B(n14120), .ZN(
        n14122) );
  XNOR2_X1 U17337 ( .A(n14122), .B(n14244), .ZN(n14292) );
  INV_X1 U17338 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14125) );
  NAND2_X1 U17339 ( .A1(n15566), .A2(n14123), .ZN(n14124) );
  NAND2_X1 U17340 ( .A1(n19781), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14287) );
  OAI211_X1 U17341 ( .C1(n14190), .C2(n14125), .A(n14124), .B(n14287), .ZN(
        n14126) );
  AOI21_X1 U17342 ( .B1(n14127), .B2(n19787), .A(n14126), .ZN(n14128) );
  OAI21_X1 U17343 ( .B1(n19608), .B2(n14292), .A(n14128), .ZN(P1_U2973) );
  NOR3_X1 U17344 ( .A1(n14146), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14131) );
  NAND2_X1 U17345 ( .A1(n14129), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14139) );
  NOR2_X1 U17346 ( .A1(n14139), .A2(n20642), .ZN(n14130) );
  MUX2_X1 U17347 ( .A(n14131), .B(n14130), .S(n15572), .Z(n14132) );
  XNOR2_X1 U17348 ( .A(n14132), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14300) );
  INV_X1 U17349 ( .A(n14133), .ZN(n15434) );
  INV_X1 U17350 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20494) );
  NOR2_X1 U17351 ( .A1(n19798), .A2(n20494), .ZN(n14293) );
  AOI21_X1 U17352 ( .B1(n19782), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n14293), .ZN(n14134) );
  OAI21_X1 U17353 ( .B1(n19793), .B2(n15432), .A(n14134), .ZN(n14135) );
  AOI21_X1 U17354 ( .B1(n15434), .B2(n19787), .A(n14135), .ZN(n14136) );
  OAI21_X1 U17355 ( .B1(n19608), .B2(n14300), .A(n14136), .ZN(P1_U2974) );
  INV_X1 U17356 ( .A(n14146), .ZN(n14137) );
  NAND2_X1 U17357 ( .A1(n14137), .A2(n14139), .ZN(n14138) );
  MUX2_X1 U17358 ( .A(n14139), .B(n14138), .S(n9603), .Z(n14140) );
  XNOR2_X1 U17359 ( .A(n14140), .B(n20642), .ZN(n14309) );
  INV_X1 U17360 ( .A(n14141), .ZN(n15445) );
  NAND2_X1 U17361 ( .A1(n15566), .A2(n15444), .ZN(n14142) );
  NAND2_X1 U17362 ( .A1(n19781), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14304) );
  OAI211_X1 U17363 ( .C1(n14190), .C2(n15439), .A(n14142), .B(n14304), .ZN(
        n14143) );
  AOI21_X1 U17364 ( .B1(n15445), .B2(n19787), .A(n14143), .ZN(n14144) );
  OAI21_X1 U17365 ( .B1(n19608), .B2(n14309), .A(n14144), .ZN(P1_U2975) );
  XNOR2_X1 U17366 ( .A(n15572), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14145) );
  XNOR2_X1 U17367 ( .A(n14146), .B(n14145), .ZN(n14319) );
  NOR2_X1 U17368 ( .A1(n19798), .A2(n14147), .ZN(n14310) );
  AOI21_X1 U17369 ( .B1(n19782), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n14310), .ZN(n14148) );
  OAI21_X1 U17370 ( .B1(n19793), .B2(n14149), .A(n14148), .ZN(n14150) );
  AOI21_X1 U17371 ( .B1(n14151), .B2(n19787), .A(n14150), .ZN(n14152) );
  OAI21_X1 U17372 ( .B1(n14319), .B2(n19608), .A(n14152), .ZN(P1_U2976) );
  NAND2_X1 U17373 ( .A1(n14154), .A2(n14153), .ZN(n14156) );
  INV_X1 U17374 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14155) );
  XNOR2_X1 U17375 ( .A(n14156), .B(n14155), .ZN(n14333) );
  NAND2_X1 U17376 ( .A1(n14157), .A2(n19787), .ZN(n14161) );
  NOR2_X1 U17377 ( .A1(n19798), .A2(n15459), .ZN(n14321) );
  NOR2_X1 U17378 ( .A1(n14190), .A2(n14158), .ZN(n14159) );
  AOI211_X1 U17379 ( .C1(n15566), .C2(n15451), .A(n14321), .B(n14159), .ZN(
        n14160) );
  OAI211_X1 U17380 ( .C1(n14333), .C2(n19608), .A(n14161), .B(n14160), .ZN(
        P1_U2977) );
  INV_X1 U17381 ( .A(n14353), .ZN(n14162) );
  NAND3_X1 U17382 ( .A1(n14162), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n15572), .ZN(n14169) );
  AOI22_X1 U17383 ( .A1(n14169), .A2(n14163), .B1(n15572), .B2(n14347), .ZN(
        n14164) );
  XNOR2_X1 U17384 ( .A(n14164), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14342) );
  INV_X1 U17385 ( .A(n14165), .ZN(n15534) );
  NAND2_X1 U17386 ( .A1(n19781), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n14336) );
  NAND2_X1 U17387 ( .A1(n19782), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14166) );
  OAI211_X1 U17388 ( .C1(n19793), .C2(n15466), .A(n14336), .B(n14166), .ZN(
        n14167) );
  AOI21_X1 U17389 ( .B1(n15534), .B2(n19787), .A(n14167), .ZN(n14168) );
  OAI21_X1 U17390 ( .B1(n14342), .B2(n19608), .A(n14168), .ZN(P1_U2978) );
  OAI21_X1 U17391 ( .B1(n14170), .B2(n15572), .A(n14169), .ZN(n14171) );
  XNOR2_X1 U17392 ( .A(n14171), .B(n14347), .ZN(n14350) );
  NAND2_X1 U17393 ( .A1(n14350), .A2(n19788), .ZN(n14175) );
  INV_X1 U17394 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n14172) );
  NOR2_X1 U17395 ( .A1(n19798), .A2(n14172), .ZN(n14343) );
  NOR2_X1 U17396 ( .A1(n14190), .A2(n15476), .ZN(n14173) );
  AOI211_X1 U17397 ( .C1(n15566), .C2(n15467), .A(n14343), .B(n14173), .ZN(
        n14174) );
  OAI211_X1 U17398 ( .C1(n19835), .C2(n15471), .A(n14175), .B(n14174), .ZN(
        P1_U2979) );
  OAI21_X1 U17399 ( .B1(n14177), .B2(n14176), .A(n14353), .ZN(n15600) );
  INV_X1 U17400 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n14178) );
  OAI22_X1 U17401 ( .A1(n14190), .A2(n15487), .B1(n19798), .B2(n14178), .ZN(
        n14180) );
  NOR2_X1 U17402 ( .A1(n15491), .A2(n19835), .ZN(n14179) );
  AOI211_X1 U17403 ( .C1(n15566), .C2(n15490), .A(n14180), .B(n14179), .ZN(
        n14181) );
  OAI21_X1 U17404 ( .B1(n19608), .B2(n15600), .A(n14181), .ZN(P1_U2981) );
  INV_X1 U17405 ( .A(n14182), .ZN(n14183) );
  OAI21_X1 U17406 ( .B1(n9915), .B2(n14184), .A(n14183), .ZN(n14195) );
  NOR2_X1 U17407 ( .A1(n14195), .A2(n14185), .ZN(n14395) );
  OAI21_X1 U17408 ( .B1(n14395), .B2(n14186), .A(n14391), .ZN(n14188) );
  XNOR2_X1 U17409 ( .A(n14188), .B(n14187), .ZN(n14389) );
  NAND2_X1 U17410 ( .A1(n14389), .A2(n19788), .ZN(n14193) );
  INV_X1 U17411 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n14189) );
  NOR2_X1 U17412 ( .A1(n19798), .A2(n14189), .ZN(n14384) );
  NOR2_X1 U17413 ( .A1(n14190), .A2(n15498), .ZN(n14191) );
  AOI211_X1 U17414 ( .C1(n15566), .C2(n15496), .A(n14384), .B(n14191), .ZN(
        n14192) );
  OAI211_X1 U17415 ( .C1(n19835), .C2(n15495), .A(n14193), .B(n14192), .ZN(
        P1_U2983) );
  NAND2_X1 U17416 ( .A1(n14195), .A2(n14194), .ZN(n14197) );
  MUX2_X1 U17417 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n12330), .S(
        n15572), .Z(n14196) );
  XNOR2_X1 U17418 ( .A(n14197), .B(n14196), .ZN(n14414) );
  INV_X1 U17419 ( .A(n14414), .ZN(n14203) );
  AOI22_X1 U17420 ( .A1(n19782), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n19781), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n14198) );
  OAI21_X1 U17421 ( .B1(n19793), .B2(n14199), .A(n14198), .ZN(n14200) );
  AOI21_X1 U17422 ( .B1(n14201), .B2(n19787), .A(n14200), .ZN(n14202) );
  OAI21_X1 U17423 ( .B1(n14203), .B2(n19608), .A(n14202), .ZN(P1_U2985) );
  NAND2_X1 U17424 ( .A1(n14205), .A2(n14204), .ZN(n14206) );
  XOR2_X1 U17425 ( .A(n14207), .B(n14206), .Z(n15615) );
  AOI22_X1 U17426 ( .A1(n19782), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n19781), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n14210) );
  NAND2_X1 U17427 ( .A1(n15566), .A2(n14208), .ZN(n14209) );
  OAI211_X1 U17428 ( .C1(n14211), .C2(n19835), .A(n14210), .B(n14209), .ZN(
        n14212) );
  AOI21_X1 U17429 ( .B1(n15615), .B2(n19788), .A(n14212), .ZN(n14213) );
  INV_X1 U17430 ( .A(n14213), .ZN(P1_U2986) );
  MUX2_X1 U17431 ( .A(n15570), .B(n15571), .S(n15572), .Z(n14214) );
  XOR2_X1 U17432 ( .A(n15629), .B(n14214), .Z(n15637) );
  NAND2_X1 U17433 ( .A1(n15637), .A2(n19788), .ZN(n14218) );
  NOR2_X1 U17434 ( .A1(n19798), .A2(n13410), .ZN(n15630) );
  NOR2_X1 U17435 ( .A1(n19793), .A2(n14215), .ZN(n14216) );
  AOI211_X1 U17436 ( .C1(n19782), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n15630), .B(n14216), .ZN(n14217) );
  OAI211_X1 U17437 ( .C1(n19835), .C2(n14219), .A(n14218), .B(n14217), .ZN(
        P1_U2989) );
  INV_X1 U17438 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14246) );
  INV_X1 U17439 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15606) );
  NAND4_X1 U17440 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15598) );
  NOR2_X1 U17441 ( .A1(n15606), .A2(n15598), .ZN(n14327) );
  NOR2_X1 U17442 ( .A1(n14222), .A2(n14221), .ZN(n15625) );
  NAND3_X1 U17443 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n15625), .ZN(n14240) );
  NOR2_X1 U17444 ( .A1(n15618), .A2(n14240), .ZN(n14407) );
  AOI21_X1 U17445 ( .B1(n14327), .B2(n14407), .A(n19824), .ZN(n14227) );
  NAND3_X1 U17446 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n14223), .ZN(n15608) );
  NOR2_X1 U17447 ( .A1(n15618), .A2(n15608), .ZN(n14372) );
  NAND2_X1 U17448 ( .A1(n14372), .A2(n14327), .ZN(n14359) );
  INV_X1 U17449 ( .A(n14359), .ZN(n14225) );
  INV_X1 U17450 ( .A(n19817), .ZN(n14224) );
  OAI21_X1 U17451 ( .B1(n19795), .B2(n14225), .A(n14224), .ZN(n14226) );
  OR2_X1 U17452 ( .A1(n14227), .A2(n14226), .ZN(n14357) );
  NOR2_X1 U17453 ( .A1(n15652), .A2(n19817), .ZN(n15634) );
  INV_X1 U17454 ( .A(n15634), .ZN(n14228) );
  OAI21_X1 U17455 ( .B1(n14357), .B2(n14329), .A(n14228), .ZN(n14338) );
  NAND2_X1 U17456 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14330) );
  NAND2_X1 U17457 ( .A1(n15652), .A2(n14330), .ZN(n14229) );
  AND2_X1 U17458 ( .A1(n14338), .A2(n14229), .ZN(n14233) );
  OR2_X1 U17459 ( .A1(n19824), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14230) );
  AND2_X1 U17460 ( .A1(n14233), .A2(n14230), .ZN(n14301) );
  NAND2_X1 U17461 ( .A1(n15652), .A2(n14231), .ZN(n14232) );
  NAND2_X1 U17462 ( .A1(n14301), .A2(n14232), .ZN(n14297) );
  OR2_X1 U17463 ( .A1(n14297), .A2(n14244), .ZN(n14234) );
  INV_X1 U17464 ( .A(n14233), .ZN(n14317) );
  OR2_X1 U17465 ( .A1(n14317), .A2(n15652), .ZN(n14237) );
  NAND2_X1 U17466 ( .A1(n14234), .A2(n14237), .ZN(n14268) );
  INV_X1 U17467 ( .A(n14245), .ZN(n14235) );
  NAND2_X1 U17468 ( .A1(n14237), .A2(n14235), .ZN(n14236) );
  NAND2_X1 U17469 ( .A1(n14268), .A2(n14236), .ZN(n14265) );
  AOI211_X1 U17470 ( .C1(n14247), .C2(n15652), .A(n14246), .B(n14265), .ZN(
        n14255) );
  INV_X1 U17471 ( .A(n14237), .ZN(n14239) );
  NOR3_X1 U17472 ( .A1(n14255), .A2(n14239), .A3(n14238), .ZN(n14250) );
  NAND2_X1 U17473 ( .A1(n19816), .A2(n14372), .ZN(n14302) );
  OAI21_X1 U17474 ( .B1(n14324), .B2(n15618), .A(n14302), .ZN(n15603) );
  NOR2_X1 U17475 ( .A1(n14329), .A2(n14330), .ZN(n14312) );
  AND3_X1 U17476 ( .A1(n14327), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n14312), .ZN(n14241) );
  NAND2_X1 U17477 ( .A1(n15603), .A2(n14241), .ZN(n14303) );
  INV_X1 U17478 ( .A(n14242), .ZN(n14243) );
  NOR2_X1 U17479 ( .A1(n14289), .A2(n14244), .ZN(n14280) );
  NAND2_X1 U17480 ( .A1(n14280), .A2(n14245), .ZN(n14263) );
  NOR4_X1 U17481 ( .A1(n14263), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14247), .A4(n14246), .ZN(n14248) );
  INV_X1 U17482 ( .A(n14251), .ZN(n14257) );
  INV_X1 U17483 ( .A(n14263), .ZN(n14252) );
  AOI21_X1 U17484 ( .B1(n14252), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14254) );
  OAI21_X1 U17485 ( .B1(n14255), .B2(n14254), .A(n14253), .ZN(n14256) );
  AOI21_X1 U17486 ( .B1(n14257), .B2(n19807), .A(n14256), .ZN(n14258) );
  OAI21_X1 U17487 ( .B1(n14259), .B2(n19820), .A(n14258), .ZN(P1_U3001) );
  NAND2_X1 U17488 ( .A1(n14260), .A2(n19807), .ZN(n14262) );
  OAI211_X1 U17489 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n14263), .A(
        n14262), .B(n14261), .ZN(n14264) );
  AOI21_X1 U17490 ( .B1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n14265), .A(
        n14264), .ZN(n14266) );
  OAI21_X1 U17491 ( .B1(n14267), .B2(n19820), .A(n14266), .ZN(P1_U3002) );
  INV_X1 U17492 ( .A(n14268), .ZN(n14285) );
  XNOR2_X1 U17493 ( .A(n14279), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14271) );
  INV_X1 U17494 ( .A(n14269), .ZN(n14270) );
  AOI21_X1 U17495 ( .B1(n14280), .B2(n14271), .A(n14270), .ZN(n14272) );
  OAI21_X1 U17496 ( .B1(n14273), .B2(n19823), .A(n14272), .ZN(n14276) );
  NOR2_X1 U17497 ( .A1(n14274), .A2(n19820), .ZN(n14275) );
  AOI211_X1 U17498 ( .C1(n14285), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14276), .B(n14275), .ZN(n14277) );
  INV_X1 U17499 ( .A(n14277), .ZN(P1_U3003) );
  AOI21_X1 U17500 ( .B1(n14280), .B2(n14279), .A(n14278), .ZN(n14281) );
  OAI21_X1 U17501 ( .B1(n14282), .B2(n19823), .A(n14281), .ZN(n14284) );
  NAND2_X1 U17502 ( .A1(n14286), .A2(n19807), .ZN(n14288) );
  OAI211_X1 U17503 ( .C1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n14289), .A(
        n14288), .B(n14287), .ZN(n14290) );
  AOI21_X1 U17504 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n14297), .A(
        n14290), .ZN(n14291) );
  OAI21_X1 U17505 ( .B1(n14292), .B2(n19820), .A(n14291), .ZN(P1_U3005) );
  INV_X1 U17506 ( .A(n15437), .ZN(n14294) );
  AOI21_X1 U17507 ( .B1(n14294), .B2(n19807), .A(n14293), .ZN(n14299) );
  OAI21_X1 U17508 ( .B1(n14303), .B2(n20642), .A(n14295), .ZN(n14296) );
  NAND2_X1 U17509 ( .A1(n14297), .A2(n14296), .ZN(n14298) );
  OAI211_X1 U17510 ( .C1(n14300), .C2(n19820), .A(n14299), .B(n14298), .ZN(
        P1_U3006) );
  OAI21_X1 U17511 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n14302), .A(
        n14301), .ZN(n14307) );
  NOR2_X1 U17512 ( .A1(n14303), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14306) );
  OAI21_X1 U17513 ( .B1(n15448), .B2(n19823), .A(n14304), .ZN(n14305) );
  AOI211_X1 U17514 ( .C1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n14307), .A(
        n14306), .B(n14305), .ZN(n14308) );
  OAI21_X1 U17515 ( .B1(n14309), .B2(n19820), .A(n14308), .ZN(P1_U3007) );
  INV_X1 U17516 ( .A(n14310), .ZN(n14314) );
  NAND4_X1 U17517 ( .A1(n15603), .A2(n14327), .A3(n14312), .A4(n14311), .ZN(
        n14313) );
  OAI211_X1 U17518 ( .C1(n14315), .C2(n19823), .A(n14314), .B(n14313), .ZN(
        n14316) );
  AOI21_X1 U17519 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n14317), .A(
        n14316), .ZN(n14318) );
  OAI21_X1 U17520 ( .B1(n14319), .B2(n19820), .A(n14318), .ZN(P1_U3008) );
  INV_X1 U17521 ( .A(n14338), .ZN(n14322) );
  NOR2_X1 U17522 ( .A1(n15454), .A2(n19823), .ZN(n14320) );
  AOI211_X1 U17523 ( .C1(n14322), .C2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n14321), .B(n14320), .ZN(n14332) );
  INV_X1 U17524 ( .A(n15608), .ZN(n14323) );
  NAND2_X1 U17525 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n14323), .ZN(
        n14325) );
  OAI21_X1 U17526 ( .B1(n14326), .B2(n14325), .A(n14324), .ZN(n15612) );
  AND2_X1 U17527 ( .A1(n14327), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14328) );
  NAND2_X1 U17528 ( .A1(n15612), .A2(n14328), .ZN(n14358) );
  OAI21_X1 U17529 ( .B1(n14359), .B2(n15609), .A(n14358), .ZN(n14344) );
  AND2_X1 U17530 ( .A1(n14344), .A2(n10280), .ZN(n14340) );
  OAI211_X1 U17531 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n14340), .B(n14330), .ZN(
        n14331) );
  OAI211_X1 U17532 ( .C1(n14333), .C2(n19820), .A(n14332), .B(n14331), .ZN(
        P1_U3009) );
  AOI21_X1 U17533 ( .B1(n14335), .B2(n9671), .A(n9984), .ZN(n15533) );
  NAND2_X1 U17534 ( .A1(n15533), .A2(n19807), .ZN(n14337) );
  OAI211_X1 U17535 ( .C1(n14338), .C2(n11143), .A(n14337), .B(n14336), .ZN(
        n14339) );
  AOI21_X1 U17536 ( .B1(n14340), .B2(n11143), .A(n14339), .ZN(n14341) );
  OAI21_X1 U17537 ( .B1(n14342), .B2(n19820), .A(n14341), .ZN(P1_U3010) );
  NAND2_X1 U17538 ( .A1(n14358), .A2(n15609), .ZN(n14362) );
  INV_X1 U17539 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14360) );
  AOI21_X1 U17540 ( .B1(n14362), .B2(n14360), .A(n14357), .ZN(n14348) );
  AOI21_X1 U17541 ( .B1(n15473), .B2(n19807), .A(n14343), .ZN(n14346) );
  NAND3_X1 U17542 ( .A1(n14344), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n14347), .ZN(n14345) );
  OAI211_X1 U17543 ( .C1(n14348), .C2(n14347), .A(n14346), .B(n14345), .ZN(
        n14349) );
  AOI21_X1 U17544 ( .B1(n14350), .B2(n19810), .A(n14349), .ZN(n14351) );
  INV_X1 U17545 ( .A(n14351), .ZN(P1_U3011) );
  NAND2_X1 U17546 ( .A1(n14353), .A2(n15606), .ZN(n14352) );
  MUX2_X1 U17547 ( .A(n14353), .B(n14352), .S(n9603), .Z(n14354) );
  XNOR2_X1 U17548 ( .A(n14354), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15549) );
  INV_X1 U17549 ( .A(n15549), .ZN(n14365) );
  INV_X1 U17550 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n14355) );
  OAI22_X1 U17551 ( .A1(n15484), .A2(n19823), .B1(n19798), .B2(n14355), .ZN(
        n14356) );
  AOI21_X1 U17552 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n14357), .A(
        n14356), .ZN(n14364) );
  NAND2_X1 U17553 ( .A1(n14359), .A2(n14358), .ZN(n14361) );
  NAND3_X1 U17554 ( .A1(n14362), .A2(n14361), .A3(n14360), .ZN(n14363) );
  OAI211_X1 U17555 ( .C1(n14365), .C2(n19820), .A(n14364), .B(n14363), .ZN(
        P1_U3012) );
  AOI21_X1 U17556 ( .B1(n15571), .B2(n14367), .A(n14366), .ZN(n14370) );
  NOR2_X1 U17557 ( .A1(n14370), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14369) );
  MUX2_X1 U17558 ( .A(n14370), .B(n14369), .S(n9603), .Z(n14371) );
  XNOR2_X1 U17559 ( .A(n14371), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15558) );
  NOR2_X1 U17560 ( .A1(n15558), .A2(n19820), .ZN(n14379) );
  NAND2_X1 U17561 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14375) );
  NAND2_X1 U17562 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15603), .ZN(
        n14381) );
  INV_X1 U17563 ( .A(n14372), .ZN(n14373) );
  AOI21_X1 U17564 ( .B1(n19818), .B2(n14373), .A(n19817), .ZN(n14374) );
  OAI21_X1 U17565 ( .B1(n14407), .B2(n19824), .A(n14374), .ZN(n14382) );
  AOI21_X1 U17566 ( .B1(n15652), .B2(n15598), .A(n14382), .ZN(n15607) );
  AOI221_X1 U17567 ( .B1(n14375), .B2(n9996), .C1(n14381), .C2(n9996), .A(
        n15607), .ZN(n14378) );
  OAI22_X1 U17568 ( .A1(n14376), .A2(n19823), .B1(n19798), .B2(n13959), .ZN(
        n14377) );
  OR3_X1 U17569 ( .A1(n14379), .A2(n14378), .A3(n14377), .ZN(P1_U3014) );
  NOR3_X1 U17570 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n14380), .A3(
        n14381), .ZN(n14388) );
  NOR2_X1 U17571 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n14381), .ZN(
        n14403) );
  INV_X1 U17572 ( .A(n14382), .ZN(n15619) );
  OAI21_X1 U17573 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n14383), .A(
        n15619), .ZN(n14405) );
  OAI21_X1 U17574 ( .B1(n14403), .B2(n14405), .A(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14386) );
  INV_X1 U17575 ( .A(n14384), .ZN(n14385) );
  OAI211_X1 U17576 ( .C1(n15505), .C2(n19823), .A(n14386), .B(n14385), .ZN(
        n14387) );
  AOI211_X1 U17577 ( .C1(n14389), .C2(n19810), .A(n14388), .B(n14387), .ZN(
        n14390) );
  INV_X1 U17578 ( .A(n14390), .ZN(P1_U3015) );
  INV_X1 U17579 ( .A(n14391), .ZN(n14392) );
  NOR2_X1 U17580 ( .A1(n14393), .A2(n14392), .ZN(n14397) );
  NOR2_X1 U17581 ( .A1(n14395), .A2(n14394), .ZN(n14396) );
  XOR2_X1 U17582 ( .A(n14397), .B(n14396), .Z(n15563) );
  OR2_X1 U17583 ( .A1(n14399), .A2(n14398), .ZN(n14400) );
  NAND2_X1 U17584 ( .A1(n14401), .A2(n14400), .ZN(n15510) );
  INV_X1 U17585 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n14402) );
  OAI22_X1 U17586 ( .A1(n15510), .A2(n19823), .B1(n19798), .B2(n14402), .ZN(
        n14404) );
  AOI211_X1 U17587 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n14405), .A(
        n14404), .B(n14403), .ZN(n14406) );
  OAI21_X1 U17588 ( .B1(n15563), .B2(n19820), .A(n14406), .ZN(P1_U3016) );
  NAND3_X1 U17589 ( .A1(n14407), .A2(n12330), .A3(n15623), .ZN(n14412) );
  OAI22_X1 U17590 ( .A1(n14409), .A2(n19823), .B1(n14408), .B2(n19798), .ZN(
        n14410) );
  INV_X1 U17591 ( .A(n14410), .ZN(n14411) );
  OAI211_X1 U17592 ( .C1(n15619), .C2(n12330), .A(n14412), .B(n14411), .ZN(
        n14413) );
  AOI21_X1 U17593 ( .B1(n14414), .B2(n19810), .A(n14413), .ZN(n14415) );
  INV_X1 U17594 ( .A(n14415), .ZN(P1_U3017) );
  NAND3_X1 U17595 ( .A1(n14417), .A2(n15385), .A3(n14416), .ZN(n15398) );
  NAND2_X1 U17596 ( .A1(n19961), .A2(n14418), .ZN(n14419) );
  OAI211_X1 U17597 ( .C1(n20516), .C2(n19922), .A(n15398), .B(n14419), .ZN(
        n14420) );
  MUX2_X1 U17598 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n14420), .S(
        n20526), .Z(P1_U3478) );
  NOR2_X1 U17599 ( .A1(n14421), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14424) );
  NOR3_X1 U17600 ( .A1(n14422), .A2(n14427), .A3(n14428), .ZN(n14423) );
  AOI211_X1 U17601 ( .C1(n20349), .C2(n14425), .A(n14424), .B(n14423), .ZN(
        n15372) );
  INV_X1 U17602 ( .A(n14426), .ZN(n15399) );
  NOR3_X1 U17603 ( .A1(n14428), .A2(n14427), .A3(n15399), .ZN(n14429) );
  AOI21_X1 U17604 ( .B1(n14431), .B2(n14430), .A(n14429), .ZN(n14432) );
  OAI21_X1 U17605 ( .B1(n15372), .B2(n14435), .A(n14432), .ZN(n14433) );
  MUX2_X1 U17606 ( .A(n14433), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n14437), .Z(P1_U3473) );
  OAI22_X1 U17607 ( .A1(n14436), .A2(n14435), .B1(n14434), .B2(n15399), .ZN(
        n14438) );
  MUX2_X1 U17608 ( .A(n14438), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n14437), .Z(P1_U3469) );
  NAND2_X1 U17609 ( .A1(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18639), .ZN(
        n14449) );
  NOR2_X1 U17610 ( .A1(n19566), .A2(n18644), .ZN(n14445) );
  AOI22_X1 U17611 ( .A1(n14440), .A2(n18625), .B1(n18637), .B2(n14439), .ZN(
        n14442) );
  NAND2_X1 U17612 ( .A1(n18614), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n14441) );
  OAI211_X1 U17613 ( .C1(n18628), .C2(n14443), .A(n14442), .B(n14441), .ZN(
        n14444) );
  NAND2_X1 U17614 ( .A1(n18623), .A2(n14446), .ZN(n14447) );
  NAND3_X1 U17615 ( .A1(n14449), .A2(n14448), .A3(n14447), .ZN(P2_U2855) );
  INV_X1 U17616 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n15691) );
  NOR2_X1 U17617 ( .A1(n14461), .A2(n14450), .ZN(n14457) );
  NAND2_X1 U17618 ( .A1(n11933), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14455) );
  AOI22_X1 U17619 ( .A1(n14451), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n14454) );
  NAND2_X1 U17620 ( .A1(n14452), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n14453) );
  NAND3_X1 U17621 ( .A1(n14455), .A2(n14454), .A3(n14453), .ZN(n14456) );
  INV_X1 U17622 ( .A(n15700), .ZN(n14458) );
  NAND2_X1 U17623 ( .A1(n14458), .A2(n14540), .ZN(n14459) );
  OAI21_X1 U17624 ( .B1(n14540), .B2(n15691), .A(n14459), .ZN(P2_U2856) );
  NAND2_X1 U17625 ( .A1(n14548), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14465) );
  INV_X1 U17626 ( .A(n14461), .ZN(n14462) );
  NAND2_X1 U17627 ( .A1(n15703), .A2(n14540), .ZN(n14464) );
  OAI211_X1 U17628 ( .C1(n14562), .C2(n14550), .A(n14465), .B(n14464), .ZN(
        P2_U2858) );
  NOR2_X1 U17629 ( .A1(n14467), .A2(n14466), .ZN(n14468) );
  XOR2_X1 U17630 ( .A(n14469), .B(n14468), .Z(n14570) );
  OAI21_X1 U17631 ( .B1(n14475), .B2(n14470), .A(n9681), .ZN(n15721) );
  NOR2_X1 U17632 ( .A1(n15721), .A2(n14548), .ZN(n14471) );
  AOI21_X1 U17633 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n14548), .A(n14471), .ZN(
        n14472) );
  OAI21_X1 U17634 ( .B1(n14570), .B2(n14550), .A(n14472), .ZN(P2_U2859) );
  NOR2_X1 U17635 ( .A1(n14485), .A2(n14473), .ZN(n14474) );
  OR2_X1 U17636 ( .A1(n14475), .A2(n14474), .ZN(n15722) );
  AOI21_X1 U17637 ( .B1(n14478), .B2(n14477), .A(n14476), .ZN(n14571) );
  NAND2_X1 U17638 ( .A1(n14571), .A2(n14522), .ZN(n14480) );
  NAND2_X1 U17639 ( .A1(n14548), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n14479) );
  OAI211_X1 U17640 ( .C1(n14548), .C2(n15722), .A(n14480), .B(n14479), .ZN(
        P2_U2860) );
  XNOR2_X1 U17641 ( .A(n14481), .B(n14482), .ZN(n14585) );
  NOR2_X1 U17642 ( .A1(n14491), .A2(n14483), .ZN(n14484) );
  OR2_X1 U17643 ( .A1(n14485), .A2(n14484), .ZN(n15740) );
  NOR2_X1 U17644 ( .A1(n15740), .A2(n14548), .ZN(n14486) );
  AOI21_X1 U17645 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n14548), .A(n14486), .ZN(
        n14487) );
  OAI21_X1 U17646 ( .B1(n14585), .B2(n14550), .A(n14487), .ZN(P2_U2861) );
  OAI21_X1 U17647 ( .B1(n14490), .B2(n14489), .A(n14488), .ZN(n14594) );
  AOI21_X1 U17648 ( .B1(n14492), .B2(n14503), .A(n14491), .ZN(n15747) );
  NOR2_X1 U17649 ( .A1(n14525), .A2(n14493), .ZN(n14494) );
  AOI21_X1 U17650 ( .B1(n15747), .B2(n14540), .A(n14494), .ZN(n14495) );
  OAI21_X1 U17651 ( .B1(n14594), .B2(n14550), .A(n14495), .ZN(P2_U2862) );
  NOR2_X1 U17652 ( .A1(n12005), .A2(n14496), .ZN(n14497) );
  XNOR2_X1 U17653 ( .A(n14498), .B(n14497), .ZN(n14499) );
  XNOR2_X1 U17654 ( .A(n14500), .B(n14499), .ZN(n15780) );
  NAND2_X1 U17655 ( .A1(n15780), .A2(n14522), .ZN(n14505) );
  NAND2_X1 U17656 ( .A1(n14509), .A2(n14501), .ZN(n14502) );
  AND2_X1 U17657 ( .A1(n14503), .A2(n14502), .ZN(n15757) );
  NAND2_X1 U17658 ( .A1(n15757), .A2(n14540), .ZN(n14504) );
  OAI211_X1 U17659 ( .C1(n14525), .C2(n10064), .A(n14505), .B(n14504), .ZN(
        P2_U2863) );
  OAI21_X1 U17660 ( .B1(n14508), .B2(n14507), .A(n14506), .ZN(n14603) );
  AOI21_X1 U17661 ( .B1(n14510), .B2(n9659), .A(n10047), .ZN(n15775) );
  INV_X1 U17662 ( .A(n15775), .ZN(n14726) );
  NOR2_X1 U17663 ( .A1(n14726), .A2(n14548), .ZN(n14511) );
  AOI21_X1 U17664 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n14548), .A(n14511), .ZN(
        n14512) );
  OAI21_X1 U17665 ( .B1(n14603), .B2(n14550), .A(n14512), .ZN(P2_U2864) );
  INV_X1 U17666 ( .A(n14514), .ZN(n14515) );
  AOI21_X1 U17667 ( .B1(n14516), .B2(n14513), .A(n14515), .ZN(n14608) );
  NAND2_X1 U17668 ( .A1(n14608), .A2(n14522), .ZN(n14518) );
  INV_X1 U17669 ( .A(n14927), .ZN(n15786) );
  NAND2_X1 U17670 ( .A1(n15786), .A2(n14540), .ZN(n14517) );
  OAI211_X1 U17671 ( .C1(n14525), .C2(n11928), .A(n14518), .B(n14517), .ZN(
        P2_U2865) );
  OR2_X1 U17672 ( .A1(n14519), .A2(n14520), .ZN(n14521) );
  AND2_X1 U17673 ( .A1(n14513), .A2(n14521), .ZN(n14616) );
  NAND2_X1 U17674 ( .A1(n14616), .A2(n14522), .ZN(n14524) );
  INV_X1 U17675 ( .A(n14743), .ZN(n14932) );
  NAND2_X1 U17676 ( .A1(n14932), .A2(n14540), .ZN(n14523) );
  OAI211_X1 U17677 ( .C1(n14525), .C2(n12226), .A(n14524), .B(n14523), .ZN(
        P2_U2866) );
  NOR2_X1 U17678 ( .A1(n14535), .A2(n14526), .ZN(n14527) );
  OR2_X1 U17679 ( .A1(n14519), .A2(n14527), .ZN(n14628) );
  AND2_X1 U17680 ( .A1(n14537), .A2(n14528), .ZN(n14530) );
  OR2_X1 U17681 ( .A1(n14530), .A2(n14529), .ZN(n14945) );
  NOR2_X1 U17682 ( .A1(n14945), .A2(n14548), .ZN(n14531) );
  AOI21_X1 U17683 ( .B1(P2_EBX_REG_20__SCAN_IN), .B2(n14548), .A(n14531), .ZN(
        n14532) );
  OAI21_X1 U17684 ( .B1(n14628), .B2(n14550), .A(n14532), .ZN(P2_U2867) );
  AND2_X1 U17685 ( .A1(n14534), .A2(n14533), .ZN(n14536) );
  OR2_X1 U17686 ( .A1(n14536), .A2(n14535), .ZN(n14641) );
  INV_X1 U17687 ( .A(n14537), .ZN(n14538) );
  AOI21_X1 U17688 ( .B1(n14539), .B2(n14546), .A(n14538), .ZN(n18459) );
  NOR2_X1 U17689 ( .A1(n14540), .A2(n11918), .ZN(n14541) );
  AOI21_X1 U17690 ( .B1(n18459), .B2(n14540), .A(n14541), .ZN(n14542) );
  OAI21_X1 U17691 ( .B1(n14641), .B2(n14550), .A(n14542), .ZN(P2_U2868) );
  OR2_X1 U17692 ( .A1(n14544), .A2(n14543), .ZN(n14545) );
  NAND2_X1 U17693 ( .A1(n14546), .A2(n14545), .ZN(n18472) );
  NOR2_X1 U17694 ( .A1(n14548), .A2(n18472), .ZN(n14547) );
  AOI21_X1 U17695 ( .B1(P2_EBX_REG_18__SCAN_IN), .B2(n14548), .A(n14547), .ZN(
        n14549) );
  OAI21_X1 U17696 ( .B1(n14551), .B2(n14550), .A(n14549), .ZN(P2_U2869) );
  AOI22_X1 U17697 ( .A1(n15778), .A2(n18656), .B1(P2_EAX_REG_30__SCAN_IN), 
        .B2(n18691), .ZN(n14556) );
  AOI22_X1 U17698 ( .A1(n18651), .A2(BUF2_REG_30__SCAN_IN), .B1(n18652), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n14555) );
  NAND2_X1 U17699 ( .A1(n18692), .A2(n14553), .ZN(n14554) );
  NAND4_X1 U17700 ( .A1(n14557), .A2(n14556), .A3(n14555), .A4(n14554), .ZN(
        P2_U2889) );
  XOR2_X1 U17701 ( .A(n14558), .B(n14563), .Z(n15702) );
  INV_X1 U17702 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n18709) );
  OAI22_X1 U17703 ( .A1(n14611), .A2(n18800), .B1(n18686), .B2(n18709), .ZN(
        n14559) );
  AOI21_X1 U17704 ( .B1(n18692), .B2(n15702), .A(n14559), .ZN(n14561) );
  AOI22_X1 U17705 ( .A1(n18651), .A2(BUF2_REG_29__SCAN_IN), .B1(n18652), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n14560) );
  OAI211_X1 U17706 ( .C1(n14562), .C2(n18671), .A(n14561), .B(n14560), .ZN(
        P2_U2890) );
  INV_X1 U17707 ( .A(n14563), .ZN(n14564) );
  AOI21_X1 U17708 ( .B1(n14565), .B2(n14572), .A(n14564), .ZN(n15718) );
  INV_X1 U17709 ( .A(n15718), .ZN(n14566) );
  OAI22_X1 U17710 ( .A1(n18687), .A2(n14566), .B1(n18686), .B2(n18711), .ZN(
        n14567) );
  AOI21_X1 U17711 ( .B1(n15778), .B2(n18660), .A(n14567), .ZN(n14569) );
  AOI22_X1 U17712 ( .A1(n18651), .A2(BUF2_REG_28__SCAN_IN), .B1(n18652), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n14568) );
  OAI211_X1 U17713 ( .C1(n14570), .C2(n18671), .A(n14569), .B(n14568), .ZN(
        P2_U2891) );
  INV_X1 U17714 ( .A(n14571), .ZN(n14578) );
  OAI21_X1 U17715 ( .B1(n14581), .B2(n14573), .A(n14572), .ZN(n14574) );
  INV_X1 U17716 ( .A(n14574), .ZN(n15723) );
  INV_X1 U17717 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n18713) );
  OAI22_X1 U17718 ( .A1(n14611), .A2(n18798), .B1(n18686), .B2(n18713), .ZN(
        n14575) );
  AOI21_X1 U17719 ( .B1(n18692), .B2(n15723), .A(n14575), .ZN(n14577) );
  AOI22_X1 U17720 ( .A1(n18651), .A2(BUF2_REG_27__SCAN_IN), .B1(n18652), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n14576) );
  OAI211_X1 U17721 ( .C1(n14578), .C2(n18671), .A(n14577), .B(n14576), .ZN(
        P2_U2892) );
  AND2_X1 U17722 ( .A1(n9649), .A2(n14579), .ZN(n14580) );
  NOR2_X1 U17723 ( .A1(n14581), .A2(n14580), .ZN(n15743) );
  INV_X1 U17724 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n18715) );
  OAI22_X1 U17725 ( .A1(n14611), .A2(n18796), .B1(n18686), .B2(n18715), .ZN(
        n14582) );
  AOI21_X1 U17726 ( .B1(n18692), .B2(n15743), .A(n14582), .ZN(n14584) );
  AOI22_X1 U17727 ( .A1(n18651), .A2(BUF2_REG_26__SCAN_IN), .B1(n18652), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n14583) );
  OAI211_X1 U17728 ( .C1(n14585), .C2(n18671), .A(n14584), .B(n14583), .ZN(
        P2_U2893) );
  NAND2_X1 U17729 ( .A1(n9689), .A2(n14586), .ZN(n14587) );
  AND2_X1 U17730 ( .A1(n9649), .A2(n14587), .ZN(n15746) );
  INV_X1 U17731 ( .A(n15746), .ZN(n14591) );
  AOI22_X1 U17732 ( .A1(n18651), .A2(BUF2_REG_25__SCAN_IN), .B1(n18652), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n14590) );
  INV_X1 U17733 ( .A(n18794), .ZN(n14588) );
  AOI22_X1 U17734 ( .A1(n15778), .A2(n14588), .B1(n18691), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n14589) );
  OAI211_X1 U17735 ( .C1(n18687), .C2(n14591), .A(n14590), .B(n14589), .ZN(
        n14592) );
  INV_X1 U17736 ( .A(n14592), .ZN(n14593) );
  OAI21_X1 U17737 ( .B1(n14594), .B2(n18671), .A(n14593), .ZN(P2_U2894) );
  NOR2_X1 U17738 ( .A1(n14596), .A2(n14595), .ZN(n14597) );
  OR2_X1 U17739 ( .A1(n14895), .A2(n14597), .ZN(n15773) );
  AOI22_X1 U17740 ( .A1(n18651), .A2(BUF2_REG_23__SCAN_IN), .B1(n18652), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n14600) );
  INV_X1 U17741 ( .A(n18928), .ZN(n14598) );
  AOI22_X1 U17742 ( .A1(n15778), .A2(n14598), .B1(n18691), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n14599) );
  OAI211_X1 U17743 ( .C1(n18687), .C2(n15773), .A(n14600), .B(n14599), .ZN(
        n14601) );
  INV_X1 U17744 ( .A(n14601), .ZN(n14602) );
  OAI21_X1 U17745 ( .B1(n14603), .B2(n18671), .A(n14602), .ZN(P2_U2896) );
  AOI22_X1 U17746 ( .A1(n18651), .A2(BUF2_REG_22__SCAN_IN), .B1(n18652), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n14606) );
  INV_X1 U17747 ( .A(n18920), .ZN(n14604) );
  AOI22_X1 U17748 ( .A1(n15778), .A2(n14604), .B1(n18691), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n14605) );
  OAI211_X1 U17749 ( .C1(n18687), .C2(n14920), .A(n14606), .B(n14605), .ZN(
        n14607) );
  AOI21_X1 U17750 ( .B1(n14608), .B2(n18694), .A(n14607), .ZN(n14609) );
  INV_X1 U17751 ( .A(n14609), .ZN(P2_U2897) );
  INV_X1 U17752 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16036) );
  INV_X1 U17753 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n17764) );
  OAI22_X1 U17754 ( .A1(n14610), .A2(n16036), .B1(n17764), .B2(n14634), .ZN(
        n18666) );
  INV_X1 U17755 ( .A(n18666), .ZN(n18912) );
  OAI22_X1 U17756 ( .A1(n14611), .A2(n18912), .B1(n18686), .B2(n18725), .ZN(
        n14615) );
  INV_X1 U17757 ( .A(n18651), .ZN(n14613) );
  INV_X1 U17758 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n14612) );
  NOR2_X1 U17759 ( .A1(n14613), .A2(n14612), .ZN(n14614) );
  AOI211_X1 U17760 ( .C1(n18652), .C2(BUF1_REG_21__SCAN_IN), .A(n14615), .B(
        n14614), .ZN(n14618) );
  NAND2_X1 U17761 ( .A1(n14616), .A2(n18694), .ZN(n14617) );
  OAI211_X1 U17762 ( .C1(n14936), .C2(n18687), .A(n14618), .B(n14617), .ZN(
        P2_U2898) );
  NOR2_X1 U17763 ( .A1(n14629), .A2(n14619), .ZN(n14620) );
  NAND2_X1 U17764 ( .A1(n18651), .A2(BUF2_REG_20__SCAN_IN), .ZN(n14625) );
  NAND2_X1 U17765 ( .A1(n18652), .A2(BUF1_REG_20__SCAN_IN), .ZN(n14624) );
  AOI22_X1 U17766 ( .A1(n14634), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n14633), .ZN(n18908) );
  INV_X1 U17767 ( .A(n18908), .ZN(n14622) );
  AOI22_X1 U17768 ( .A1(n15778), .A2(n14622), .B1(n18691), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n14623) );
  NAND3_X1 U17769 ( .A1(n14625), .A2(n14624), .A3(n14623), .ZN(n14626) );
  AOI21_X1 U17770 ( .B1(n9725), .B2(n18692), .A(n14626), .ZN(n14627) );
  OAI21_X1 U17771 ( .B1(n18671), .B2(n14628), .A(n14627), .ZN(P2_U2899) );
  INV_X1 U17772 ( .A(n14629), .ZN(n14630) );
  OAI21_X1 U17773 ( .B1(n14632), .B2(n14631), .A(n14630), .ZN(n18461) );
  INV_X1 U17774 ( .A(n18461), .ZN(n14963) );
  NAND2_X1 U17775 ( .A1(n18651), .A2(BUF2_REG_19__SCAN_IN), .ZN(n14638) );
  NAND2_X1 U17776 ( .A1(n18652), .A2(BUF1_REG_19__SCAN_IN), .ZN(n14637) );
  AOI22_X1 U17777 ( .A1(n14634), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n14633), .ZN(n18904) );
  INV_X1 U17778 ( .A(n18904), .ZN(n14635) );
  AOI22_X1 U17779 ( .A1(n15778), .A2(n14635), .B1(n18691), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n14636) );
  NAND3_X1 U17780 ( .A1(n14638), .A2(n14637), .A3(n14636), .ZN(n14639) );
  AOI21_X1 U17781 ( .B1(n14963), .B2(n18692), .A(n14639), .ZN(n14640) );
  OAI21_X1 U17782 ( .B1(n18671), .B2(n14641), .A(n14640), .ZN(P2_U2900) );
  INV_X1 U17783 ( .A(n14644), .ZN(n14647) );
  NOR2_X1 U17784 ( .A1(n14645), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14646) );
  MUX2_X1 U17785 ( .A(n14647), .B(n14646), .S(n18911), .Z(n15692) );
  NAND2_X1 U17786 ( .A1(n15692), .A2(n12224), .ZN(n14648) );
  NOR2_X1 U17787 ( .A1(n15700), .A2(n18811), .ZN(n14652) );
  NAND2_X1 U17788 ( .A1(n18850), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14831) );
  NAND2_X1 U17789 ( .A1(n18820), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14649) );
  OAI211_X1 U17790 ( .C1(n18816), .C2(n14650), .A(n14831), .B(n14649), .ZN(
        n14651) );
  NOR2_X1 U17791 ( .A1(n18816), .A2(n15697), .ZN(n14653) );
  AOI211_X1 U17792 ( .C1(n18820), .C2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n14654), .B(n14653), .ZN(n14655) );
  OAI21_X1 U17793 ( .B1(n14656), .B2(n18811), .A(n14655), .ZN(n14657) );
  AOI21_X1 U17794 ( .B1(n14658), .B2(n18821), .A(n14657), .ZN(n14659) );
  OAI21_X1 U17795 ( .B1(n14660), .B2(n18833), .A(n14659), .ZN(P2_U2984) );
  NOR2_X1 U17796 ( .A1(n14662), .A2(n14661), .ZN(n14664) );
  XOR2_X1 U17797 ( .A(n14664), .B(n14663), .Z(n14849) );
  NAND2_X1 U17798 ( .A1(n18829), .A2(n15705), .ZN(n14665) );
  NAND2_X1 U17799 ( .A1(n13482), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n14840) );
  OAI211_X1 U17800 ( .C1(n15852), .C2(n14666), .A(n14665), .B(n14840), .ZN(
        n14667) );
  AOI21_X1 U17801 ( .B1(n15703), .B2(n18830), .A(n14667), .ZN(n14671) );
  AOI21_X1 U17802 ( .B1(n14669), .B2(n14681), .A(n14668), .ZN(n14847) );
  NAND2_X1 U17803 ( .A1(n14847), .A2(n18821), .ZN(n14670) );
  OAI211_X1 U17804 ( .C1(n14849), .C2(n18833), .A(n14671), .B(n14670), .ZN(
        P2_U2985) );
  INV_X1 U17805 ( .A(n14673), .ZN(n14674) );
  AOI22_X1 U17806 ( .A1(n14686), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n14675), .B2(n14674), .ZN(n14678) );
  XNOR2_X1 U17807 ( .A(n14676), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14677) );
  XNOR2_X1 U17808 ( .A(n14678), .B(n14677), .ZN(n14860) );
  INV_X1 U17809 ( .A(n15721), .ZN(n14684) );
  NAND2_X1 U17810 ( .A1(n13482), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n14853) );
  NAND2_X1 U17811 ( .A1(n18820), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14679) );
  OAI211_X1 U17812 ( .C1(n18816), .C2(n14680), .A(n14853), .B(n14679), .ZN(
        n14683) );
  OAI21_X1 U17813 ( .B1(n14687), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14681), .ZN(n14854) );
  NOR2_X1 U17814 ( .A1(n14854), .A2(n15838), .ZN(n14682) );
  AOI211_X1 U17815 ( .C1(n14684), .C2(n18830), .A(n14683), .B(n14682), .ZN(
        n14685) );
  OAI21_X1 U17816 ( .B1(n14860), .B2(n18833), .A(n14685), .ZN(P2_U2986) );
  XNOR2_X1 U17817 ( .A(n14686), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14870) );
  AOI21_X1 U17818 ( .B1(n14851), .B2(n14695), .A(n14687), .ZN(n14868) );
  NAND2_X1 U17819 ( .A1(n13482), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n14862) );
  OAI21_X1 U17820 ( .B1(n15852), .B2(n14688), .A(n14862), .ZN(n14689) );
  AOI21_X1 U17821 ( .B1(n18829), .B2(n15727), .A(n14689), .ZN(n14690) );
  OAI21_X1 U17822 ( .B1(n15722), .B2(n18811), .A(n14690), .ZN(n14691) );
  AOI21_X1 U17823 ( .B1(n14868), .B2(n18821), .A(n14691), .ZN(n14692) );
  OAI21_X1 U17824 ( .B1(n14870), .B2(n18833), .A(n14692), .ZN(P2_U2987) );
  NAND2_X1 U17825 ( .A1(n14703), .A2(n14707), .ZN(n14693) );
  XOR2_X1 U17826 ( .A(n14694), .B(n14693), .Z(n14881) );
  INV_X1 U17827 ( .A(n14695), .ZN(n14696) );
  AOI21_X1 U17828 ( .B1(n14877), .B2(n14702), .A(n14696), .ZN(n14879) );
  NOR2_X1 U17829 ( .A1(n15740), .A2(n18811), .ZN(n14700) );
  NAND2_X1 U17830 ( .A1(n13482), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n14872) );
  NAND2_X1 U17831 ( .A1(n18820), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14697) );
  OAI211_X1 U17832 ( .C1(n18816), .C2(n14698), .A(n14872), .B(n14697), .ZN(
        n14699) );
  AOI211_X1 U17833 ( .C1(n14879), .C2(n18821), .A(n14700), .B(n14699), .ZN(
        n14701) );
  OAI21_X1 U17834 ( .B1(n14881), .B2(n18833), .A(n14701), .ZN(P2_U2988) );
  OAI21_X1 U17835 ( .B1(n14720), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n14702), .ZN(n14892) );
  INV_X1 U17836 ( .A(n14703), .ZN(n14708) );
  AOI21_X1 U17837 ( .B1(n14705), .B2(n14707), .A(n14704), .ZN(n14706) );
  AOI21_X1 U17838 ( .B1(n14708), .B2(n14707), .A(n14706), .ZN(n14882) );
  NAND2_X1 U17839 ( .A1(n14882), .A2(n18808), .ZN(n14713) );
  NAND2_X1 U17840 ( .A1(n18829), .A2(n15749), .ZN(n14709) );
  NAND2_X1 U17841 ( .A1(n13482), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n14883) );
  OAI211_X1 U17842 ( .C1(n15852), .C2(n14710), .A(n14709), .B(n14883), .ZN(
        n14711) );
  AOI21_X1 U17843 ( .B1(n15747), .B2(n18830), .A(n14711), .ZN(n14712) );
  OAI211_X1 U17844 ( .C1(n15838), .C2(n14892), .A(n14713), .B(n14712), .ZN(
        P2_U2989) );
  XNOR2_X1 U17845 ( .A(n14714), .B(n14721), .ZN(n14715) );
  XNOR2_X1 U17846 ( .A(n14716), .B(n14715), .ZN(n14904) );
  NAND2_X1 U17847 ( .A1(n13482), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n14896) );
  NAND2_X1 U17848 ( .A1(n18820), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14717) );
  OAI211_X1 U17849 ( .C1(n18816), .C2(n14718), .A(n14896), .B(n14717), .ZN(
        n14719) );
  AOI21_X1 U17850 ( .B1(n15757), .B2(n18830), .A(n14719), .ZN(n14723) );
  AOI21_X1 U17851 ( .B1(n14721), .B2(n14729), .A(n14720), .ZN(n14902) );
  NAND2_X1 U17852 ( .A1(n14902), .A2(n18821), .ZN(n14722) );
  OAI211_X1 U17853 ( .C1(n14904), .C2(n18833), .A(n14723), .B(n14722), .ZN(
        P2_U2990) );
  XNOR2_X1 U17854 ( .A(n14725), .B(n14724), .ZN(n14913) );
  OAI22_X1 U17855 ( .A1(n15852), .A2(n10114), .B1(n19494), .B2(n18600), .ZN(
        n14728) );
  NOR2_X1 U17856 ( .A1(n14726), .A2(n18811), .ZN(n14727) );
  AOI211_X1 U17857 ( .C1(n18829), .C2(n15768), .A(n14728), .B(n14727), .ZN(
        n14731) );
  INV_X1 U17858 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14923) );
  NOR2_X1 U17859 ( .A1(n14919), .A2(n14923), .ZN(n14918) );
  OAI21_X1 U17860 ( .B1(n14918), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n14729), .ZN(n14909) );
  OR2_X1 U17861 ( .A1(n14909), .A2(n15838), .ZN(n14730) );
  OAI211_X1 U17862 ( .C1(n14913), .C2(n18833), .A(n14731), .B(n14730), .ZN(
        P2_U2991) );
  NAND2_X2 U17863 ( .A1(n15060), .A2(n14968), .ZN(n14993) );
  NOR2_X2 U17864 ( .A1(n14993), .A2(n14732), .ZN(n14775) );
  NAND2_X1 U17865 ( .A1(n14775), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14766) );
  INV_X1 U17866 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14951) );
  NOR2_X1 U17867 ( .A1(n14766), .A2(n14951), .ZN(n14753) );
  OAI21_X1 U17868 ( .B1(n14753), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n14919), .ZN(n14942) );
  INV_X1 U17869 ( .A(n15793), .ZN(n14733) );
  AOI21_X1 U17870 ( .B1(n14791), .B2(n14790), .A(n14734), .ZN(n14782) );
  AND2_X1 U17871 ( .A1(n14736), .A2(n14735), .ZN(n14783) );
  INV_X1 U17872 ( .A(n14736), .ZN(n14737) );
  INV_X1 U17873 ( .A(n14738), .ZN(n14739) );
  NAND2_X1 U17874 ( .A1(n14931), .A2(n18808), .ZN(n14748) );
  NAND2_X1 U17875 ( .A1(n18850), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n14933) );
  OAI21_X1 U17876 ( .B1(n15852), .B2(n14742), .A(n14933), .ZN(n14745) );
  NOR2_X1 U17877 ( .A1(n14743), .A2(n18811), .ZN(n14744) );
  AOI211_X1 U17878 ( .C1(n18829), .C2(n14746), .A(n14745), .B(n14744), .ZN(
        n14747) );
  OAI211_X1 U17879 ( .C1(n15838), .C2(n14942), .A(n14748), .B(n14747), .ZN(
        P2_U2993) );
  NAND2_X1 U17880 ( .A1(n9929), .A2(n14750), .ZN(n14751) );
  XNOR2_X1 U17881 ( .A(n14752), .B(n14751), .ZN(n14955) );
  AOI21_X1 U17882 ( .B1(n14951), .B2(n14766), .A(n14753), .ZN(n14953) );
  NOR2_X1 U17883 ( .A1(n18600), .A2(n14754), .ZN(n14948) );
  NOR2_X1 U17884 ( .A1(n18816), .A2(n14755), .ZN(n14756) );
  AOI211_X1 U17885 ( .C1(n18820), .C2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n14948), .B(n14756), .ZN(n14757) );
  OAI21_X1 U17886 ( .B1(n14945), .B2(n18811), .A(n14757), .ZN(n14758) );
  AOI21_X1 U17887 ( .B1(n14953), .B2(n18821), .A(n14758), .ZN(n14759) );
  OAI21_X1 U17888 ( .B1(n14955), .B2(n18833), .A(n14759), .ZN(P2_U2994) );
  INV_X1 U17889 ( .A(n14770), .ZN(n14760) );
  OAI21_X1 U17890 ( .B1(n14772), .B2(n14760), .A(n14771), .ZN(n14764) );
  NAND2_X1 U17891 ( .A1(n14762), .A2(n14761), .ZN(n14763) );
  XNOR2_X1 U17892 ( .A(n14764), .B(n14763), .ZN(n14967) );
  NAND2_X1 U17893 ( .A1(n18452), .A2(n18829), .ZN(n14765) );
  NAND2_X1 U17894 ( .A1(n18850), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n14958) );
  OAI211_X1 U17895 ( .C1(n15852), .C2(n18456), .A(n14765), .B(n14958), .ZN(
        n14768) );
  OAI21_X1 U17896 ( .B1(n14775), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n14766), .ZN(n14964) );
  NOR2_X1 U17897 ( .A1(n14964), .A2(n15838), .ZN(n14767) );
  OAI21_X1 U17898 ( .B1(n14967), .B2(n18833), .A(n14769), .ZN(P2_U2995) );
  NAND2_X1 U17899 ( .A1(n14771), .A2(n14770), .ZN(n14773) );
  XOR2_X1 U17900 ( .A(n14773), .B(n14772), .Z(n14980) );
  INV_X1 U17901 ( .A(n14774), .ZN(n14981) );
  AOI21_X1 U17902 ( .B1(n14987), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14776) );
  NOR2_X1 U17903 ( .A1(n14776), .A2(n14775), .ZN(n14977) );
  NOR2_X1 U17904 ( .A1(n18472), .A2(n18811), .ZN(n14780) );
  NAND2_X1 U17905 ( .A1(n18850), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n14973) );
  NAND2_X1 U17906 ( .A1(n18820), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14777) );
  OAI211_X1 U17907 ( .C1(n14778), .C2(n18816), .A(n14973), .B(n14777), .ZN(
        n14779) );
  AOI211_X1 U17908 ( .C1(n14977), .C2(n18821), .A(n14780), .B(n14779), .ZN(
        n14781) );
  OAI21_X1 U17909 ( .B1(n14980), .B2(n18833), .A(n14781), .ZN(P2_U2996) );
  XOR2_X1 U17910 ( .A(n14783), .B(n14782), .Z(n14991) );
  XNOR2_X1 U17911 ( .A(n14987), .B(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14787) );
  AOI22_X1 U17912 ( .A1(n18820), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n18829), .B2(n18475), .ZN(n14786) );
  NOR2_X1 U17913 ( .A1(n19483), .A2(n18600), .ZN(n14784) );
  AOI21_X1 U17914 ( .B1(n18482), .B2(n18830), .A(n14784), .ZN(n14785) );
  OAI211_X1 U17915 ( .C1(n14787), .C2(n15838), .A(n14786), .B(n14785), .ZN(
        n14788) );
  INV_X1 U17916 ( .A(n14788), .ZN(n14789) );
  OAI21_X1 U17917 ( .B1(n14991), .B2(n18833), .A(n14789), .ZN(P2_U2997) );
  XNOR2_X1 U17918 ( .A(n14791), .B(n14790), .ZN(n15001) );
  OR2_X1 U17919 ( .A1(n15001), .A2(n18833), .ZN(n14799) );
  NOR2_X1 U17920 ( .A1(n12178), .A2(n18496), .ZN(n14792) );
  AOI21_X1 U17921 ( .B1(n18490), .B2(n18830), .A(n14792), .ZN(n14798) );
  INV_X1 U17922 ( .A(n14993), .ZN(n15791) );
  AOI21_X1 U17923 ( .B1(n15791), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14793) );
  OR3_X1 U17924 ( .A1(n14793), .A2(n14987), .A3(n15838), .ZN(n14797) );
  INV_X1 U17925 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n14794) );
  OAI22_X1 U17926 ( .A1(n15852), .A2(n14794), .B1(n18816), .B2(n18486), .ZN(
        n14795) );
  INV_X1 U17927 ( .A(n14795), .ZN(n14796) );
  NAND4_X1 U17928 ( .A1(n14799), .A2(n14798), .A3(n14797), .A4(n14796), .ZN(
        P2_U2998) );
  NAND2_X1 U17929 ( .A1(n14801), .A2(n14800), .ZN(n14802) );
  XNOR2_X1 U17930 ( .A(n14803), .B(n14802), .ZN(n15012) );
  XNOR2_X1 U17931 ( .A(n14993), .B(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15010) );
  INV_X1 U17932 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19480) );
  OAI22_X1 U17933 ( .A1(n15852), .A2(n20697), .B1(n19480), .B2(n18600), .ZN(
        n14806) );
  INV_X1 U17934 ( .A(n18501), .ZN(n14804) );
  OAI22_X1 U17935 ( .A1(n18816), .A2(n14804), .B1(n18811), .B2(n15002), .ZN(
        n14805) );
  AOI211_X1 U17936 ( .C1(n15010), .C2(n18821), .A(n14806), .B(n14805), .ZN(
        n14807) );
  OAI21_X1 U17937 ( .B1(n15012), .B2(n18833), .A(n14807), .ZN(P2_U2999) );
  NAND2_X1 U17938 ( .A1(n14809), .A2(n14808), .ZN(n14810) );
  XNOR2_X1 U17939 ( .A(n14811), .B(n14810), .ZN(n15022) );
  INV_X1 U17940 ( .A(n18523), .ZN(n14813) );
  NAND2_X1 U17941 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15799), .ZN(
        n15800) );
  AND2_X1 U17942 ( .A1(n15799), .A2(n15015), .ZN(n15790) );
  AOI21_X1 U17943 ( .B1(n13795), .B2(n15800), .A(n15790), .ZN(n14812) );
  INV_X1 U17944 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n19477) );
  OAI22_X1 U17945 ( .A1(n15852), .A2(n18518), .B1(n19477), .B2(n18496), .ZN(
        n14814) );
  XNOR2_X1 U17946 ( .A(n14815), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15079) );
  INV_X1 U17947 ( .A(n15825), .ZN(n14816) );
  NAND2_X1 U17948 ( .A1(n14816), .A2(n15826), .ZN(n14817) );
  XNOR2_X1 U17949 ( .A(n15827), .B(n14817), .ZN(n15077) );
  OAI22_X1 U17950 ( .A1(n15852), .A2(n14818), .B1(n19470), .B2(n18600), .ZN(
        n14822) );
  INV_X1 U17951 ( .A(n18594), .ZN(n14819) );
  OAI22_X1 U17952 ( .A1(n18811), .A2(n14820), .B1(n18816), .B2(n14819), .ZN(
        n14821) );
  AOI211_X1 U17953 ( .C1(n15077), .C2(n18808), .A(n14822), .B(n14821), .ZN(
        n14823) );
  OAI21_X1 U17954 ( .B1(n15079), .B2(n15838), .A(n14823), .ZN(P2_U3007) );
  OAI21_X1 U17955 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15081), .A(
        n14824), .ZN(n14825) );
  INV_X1 U17956 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n14828) );
  AOI22_X1 U17957 ( .A1(n12163), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n14826), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14827) );
  OAI21_X1 U17958 ( .B1(n12103), .B2(n14828), .A(n14827), .ZN(n14829) );
  XNOR2_X1 U17959 ( .A(n14830), .B(n14829), .ZN(n18650) );
  INV_X1 U17960 ( .A(n14831), .ZN(n14835) );
  NOR4_X1 U17961 ( .A1(n14863), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14833), .A4(n14832), .ZN(n14834) );
  AOI211_X1 U17962 ( .C1(n18875), .C2(n18650), .A(n14835), .B(n14834), .ZN(
        n14836) );
  INV_X1 U17963 ( .A(n15703), .ZN(n14845) );
  AOI21_X1 U17964 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n14863), .ZN(n14838) );
  OR2_X1 U17965 ( .A1(n14861), .A2(n14838), .ZN(n14858) );
  NAND2_X1 U17966 ( .A1(n14858), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14844) );
  NAND2_X1 U17967 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14839) );
  NOR3_X1 U17968 ( .A1(n14863), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14839), .ZN(n14842) );
  INV_X1 U17969 ( .A(n14840), .ZN(n14841) );
  OAI211_X1 U17970 ( .C1(n18839), .C2(n14845), .A(n14844), .B(n14843), .ZN(
        n14846) );
  AOI21_X1 U17971 ( .B1(n14847), .B2(n18849), .A(n14846), .ZN(n14848) );
  OAI21_X1 U17972 ( .B1(n14849), .B2(n18859), .A(n14848), .ZN(P2_U3017) );
  OAI21_X1 U17973 ( .B1(n14863), .B2(n14851), .A(n14850), .ZN(n14857) );
  NAND2_X1 U17974 ( .A1(n18875), .A2(n15718), .ZN(n14852) );
  OAI211_X1 U17975 ( .C1(n15721), .C2(n18839), .A(n14853), .B(n14852), .ZN(
        n14856) );
  NOR2_X1 U17976 ( .A1(n14854), .A2(n18861), .ZN(n14855) );
  AOI211_X1 U17977 ( .C1(n14858), .C2(n14857), .A(n14856), .B(n14855), .ZN(
        n14859) );
  OAI21_X1 U17978 ( .B1(n14860), .B2(n18859), .A(n14859), .ZN(P2_U3018) );
  NAND2_X1 U17979 ( .A1(n14861), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14866) );
  OAI21_X1 U17980 ( .B1(n14863), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n14862), .ZN(n14864) );
  AOI21_X1 U17981 ( .B1(n18875), .B2(n15723), .A(n14864), .ZN(n14865) );
  OAI211_X1 U17982 ( .C1(n18839), .C2(n15722), .A(n14866), .B(n14865), .ZN(
        n14867) );
  AOI21_X1 U17983 ( .B1(n14868), .B2(n18849), .A(n14867), .ZN(n14869) );
  OAI21_X1 U17984 ( .B1(n14870), .B2(n18859), .A(n14869), .ZN(P2_U3019) );
  INV_X1 U17985 ( .A(n14871), .ZN(n14885) );
  XNOR2_X1 U17986 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14873) );
  OAI21_X1 U17987 ( .B1(n14885), .B2(n14873), .A(n14872), .ZN(n14875) );
  NOR2_X1 U17988 ( .A1(n15740), .A2(n18839), .ZN(n14874) );
  AOI211_X1 U17989 ( .C1(n15743), .C2(n18875), .A(n14875), .B(n14874), .ZN(
        n14876) );
  OAI21_X1 U17990 ( .B1(n14887), .B2(n14877), .A(n14876), .ZN(n14878) );
  AOI21_X1 U17991 ( .B1(n14879), .B2(n18849), .A(n14878), .ZN(n14880) );
  OAI21_X1 U17992 ( .B1(n14881), .B2(n18859), .A(n14880), .ZN(P2_U3020) );
  NAND2_X1 U17993 ( .A1(n14882), .A2(n18846), .ZN(n14891) );
  NAND2_X1 U17994 ( .A1(n18875), .A2(n15746), .ZN(n14884) );
  OAI211_X1 U17995 ( .C1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n14885), .A(
        n14884), .B(n14883), .ZN(n14889) );
  NOR2_X1 U17996 ( .A1(n14887), .A2(n14886), .ZN(n14888) );
  AOI211_X1 U17997 ( .C1(n15747), .C2(n18868), .A(n14889), .B(n14888), .ZN(
        n14890) );
  OAI211_X1 U17998 ( .C1(n14892), .C2(n18861), .A(n14891), .B(n14890), .ZN(
        P2_U3021) );
  AOI21_X1 U17999 ( .B1(n14893), .B2(n14924), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14899) );
  OAI21_X1 U18000 ( .B1(n14895), .B2(n14894), .A(n9689), .ZN(n15756) );
  OAI21_X1 U18001 ( .B1(n15898), .B2(n15756), .A(n14896), .ZN(n14897) );
  AOI21_X1 U18002 ( .B1(n15757), .B2(n18868), .A(n14897), .ZN(n14898) );
  OAI21_X1 U18003 ( .B1(n14900), .B2(n14899), .A(n14898), .ZN(n14901) );
  AOI21_X1 U18004 ( .B1(n14902), .B2(n18849), .A(n14901), .ZN(n14903) );
  OAI21_X1 U18005 ( .B1(n14904), .B2(n18859), .A(n14903), .ZN(P2_U3022) );
  OAI21_X1 U18006 ( .B1(n14905), .B2(n15081), .A(n15029), .ZN(n14939) );
  NAND2_X1 U18007 ( .A1(n15775), .A2(n18868), .ZN(n14908) );
  XOR2_X1 U18008 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(n14906) );
  AOI22_X1 U18009 ( .A1(n14924), .A2(n14906), .B1(n18850), .B2(
        P2_REIP_REG_23__SCAN_IN), .ZN(n14907) );
  OAI211_X1 U18010 ( .C1(n15898), .C2(n15773), .A(n14908), .B(n14907), .ZN(
        n14911) );
  NOR2_X1 U18011 ( .A1(n14909), .A2(n18861), .ZN(n14910) );
  AOI211_X1 U18012 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n14939), .A(
        n14911), .B(n14910), .ZN(n14912) );
  OAI21_X1 U18013 ( .B1(n14913), .B2(n18859), .A(n14912), .ZN(P2_U3023) );
  NOR2_X1 U18014 ( .A1(n14915), .A2(n9938), .ZN(n14916) );
  XNOR2_X1 U18015 ( .A(n14917), .B(n14916), .ZN(n15787) );
  INV_X1 U18016 ( .A(n15787), .ZN(n14930) );
  AOI21_X1 U18017 ( .B1(n14923), .B2(n14919), .A(n14918), .ZN(n15785) );
  NAND2_X1 U18018 ( .A1(n14939), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14926) );
  NOR2_X1 U18019 ( .A1(n19492), .A2(n18600), .ZN(n14922) );
  NOR2_X1 U18020 ( .A1(n15898), .A2(n14920), .ZN(n14921) );
  AOI211_X1 U18021 ( .C1(n14924), .C2(n14923), .A(n14922), .B(n14921), .ZN(
        n14925) );
  OAI211_X1 U18022 ( .C1(n14927), .C2(n18839), .A(n14926), .B(n14925), .ZN(
        n14928) );
  AOI21_X1 U18023 ( .B1(n15785), .B2(n18849), .A(n14928), .ZN(n14929) );
  OAI21_X1 U18024 ( .B1(n14930), .B2(n18859), .A(n14929), .ZN(P2_U3024) );
  NAND2_X1 U18025 ( .A1(n14931), .A2(n18846), .ZN(n14941) );
  NAND2_X1 U18026 ( .A1(n14932), .A2(n18868), .ZN(n14934) );
  OAI211_X1 U18027 ( .C1(n14935), .C2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n14934), .B(n14933), .ZN(n14938) );
  NOR2_X1 U18028 ( .A1(n14936), .A2(n15898), .ZN(n14937) );
  AOI211_X1 U18029 ( .C1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n14939), .A(
        n14938), .B(n14937), .ZN(n14940) );
  OAI211_X1 U18030 ( .C1(n14942), .C2(n18861), .A(n14941), .B(n14940), .ZN(
        P2_U3025) );
  AOI21_X1 U18031 ( .B1(n14944), .B2(n14943), .A(n15068), .ZN(n14957) );
  NAND2_X1 U18032 ( .A1(n9725), .A2(n18875), .ZN(n14950) );
  INV_X1 U18033 ( .A(n14945), .ZN(n18440) );
  XNOR2_X1 U18034 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14946) );
  NOR2_X1 U18035 ( .A1(n14960), .A2(n14946), .ZN(n14947) );
  AOI211_X1 U18036 ( .C1(n18440), .C2(n18868), .A(n14948), .B(n14947), .ZN(
        n14949) );
  OAI211_X1 U18037 ( .C1(n14957), .C2(n14951), .A(n14950), .B(n14949), .ZN(
        n14952) );
  AOI21_X1 U18038 ( .B1(n14953), .B2(n18849), .A(n14952), .ZN(n14954) );
  OAI21_X1 U18039 ( .B1(n14955), .B2(n18859), .A(n14954), .ZN(P2_U3026) );
  NOR2_X1 U18040 ( .A1(n14957), .A2(n14956), .ZN(n14962) );
  NAND2_X1 U18041 ( .A1(n18459), .A2(n18868), .ZN(n14959) );
  OAI211_X1 U18042 ( .C1(n14960), .C2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n14959), .B(n14958), .ZN(n14961) );
  AOI211_X1 U18043 ( .C1(n14963), .C2(n18875), .A(n14962), .B(n14961), .ZN(
        n14966) );
  OR2_X1 U18044 ( .A1(n14964), .A2(n18861), .ZN(n14965) );
  OAI211_X1 U18045 ( .C1(n14967), .C2(n18859), .A(n14966), .B(n14965), .ZN(
        P2_U3027) );
  INV_X1 U18046 ( .A(n14972), .ZN(n14969) );
  AOI21_X1 U18047 ( .B1(n15029), .B2(n14968), .A(n15028), .ZN(n15006) );
  AOI21_X1 U18048 ( .B1(n14969), .B2(n18837), .A(n15006), .ZN(n14970) );
  NOR2_X1 U18049 ( .A1(n14970), .A2(n14971), .ZN(n14976) );
  INV_X1 U18050 ( .A(n14992), .ZN(n15005) );
  NAND3_X1 U18051 ( .A1(n15005), .A2(n14972), .A3(n14971), .ZN(n14974) );
  OAI211_X1 U18052 ( .C1(n18472), .C2(n18839), .A(n14974), .B(n14973), .ZN(
        n14975) );
  AOI211_X1 U18053 ( .C1(n18470), .C2(n18875), .A(n14976), .B(n14975), .ZN(
        n14979) );
  NAND2_X1 U18054 ( .A1(n14977), .A2(n18849), .ZN(n14978) );
  OAI211_X1 U18055 ( .C1(n14980), .C2(n18859), .A(n14979), .B(n14978), .ZN(
        P2_U3028) );
  OAI22_X1 U18056 ( .A1(n9884), .A2(n18861), .B1(n14981), .B2(n14992), .ZN(
        n14986) );
  NOR2_X1 U18057 ( .A1(n18484), .A2(n15898), .ZN(n14984) );
  OAI22_X1 U18058 ( .A1(n18839), .A2(n14982), .B1(n19483), .B2(n18600), .ZN(
        n14983) );
  AOI211_X1 U18059 ( .C1(n14986), .C2(n14985), .A(n14984), .B(n14983), .ZN(
        n14990) );
  OAI21_X1 U18060 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15081), .A(
        n14996), .ZN(n14988) );
  NAND2_X1 U18061 ( .A1(n14988), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14989) );
  OAI211_X1 U18062 ( .C1(n14991), .C2(n18859), .A(n14990), .B(n14989), .ZN(
        P2_U3029) );
  NOR2_X1 U18063 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n15004), .ZN(
        n14999) );
  OAI21_X1 U18064 ( .B1(n14993), .B2(n18861), .A(n14992), .ZN(n14998) );
  INV_X1 U18065 ( .A(n18491), .ZN(n14995) );
  AOI22_X1 U18066 ( .A1(n18868), .A2(n18490), .B1(P2_REIP_REG_16__SCAN_IN), 
        .B2(n13482), .ZN(n14994) );
  OAI21_X1 U18067 ( .B1(n14995), .B2(n15898), .A(n14994), .ZN(n14997) );
  OAI21_X1 U18068 ( .B1(n18859), .B2(n15001), .A(n15000), .ZN(P2_U3030) );
  OAI22_X1 U18069 ( .A1(n18839), .A2(n15002), .B1(n19480), .B2(n18600), .ZN(
        n15003) );
  AOI21_X1 U18070 ( .B1(n15005), .B2(n15004), .A(n15003), .ZN(n15008) );
  NAND2_X1 U18071 ( .A1(n15006), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15007) );
  OAI211_X1 U18072 ( .C1(n18506), .C2(n15898), .A(n15008), .B(n15007), .ZN(
        n15009) );
  AOI21_X1 U18073 ( .B1(n15010), .B2(n18849), .A(n15009), .ZN(n15011) );
  OAI21_X1 U18074 ( .B1(n15012), .B2(n18859), .A(n15011), .ZN(P2_U3031) );
  NAND2_X1 U18075 ( .A1(n15013), .A2(n15862), .ZN(n15873) );
  INV_X1 U18076 ( .A(n15013), .ZN(n15014) );
  OAI21_X1 U18077 ( .B1(n15014), .B2(n15068), .A(n18837), .ZN(n15872) );
  OAI21_X1 U18078 ( .B1(n15015), .B2(n15873), .A(n15872), .ZN(n15857) );
  OAI21_X1 U18079 ( .B1(n13774), .B2(n15873), .A(n13795), .ZN(n15020) );
  OAI22_X1 U18080 ( .A1(n15898), .A2(n18528), .B1(n19477), .B2(n18600), .ZN(
        n15019) );
  OAI22_X1 U18081 ( .A1(n18861), .A2(n15017), .B1(n18839), .B2(n15016), .ZN(
        n15018) );
  AOI211_X1 U18082 ( .C1(n15857), .C2(n15020), .A(n15019), .B(n15018), .ZN(
        n15021) );
  OAI21_X1 U18083 ( .B1(n15022), .B2(n18859), .A(n15021), .ZN(P2_U3033) );
  INV_X1 U18084 ( .A(n15023), .ZN(n15043) );
  INV_X1 U18085 ( .A(n15799), .ZN(n15024) );
  OAI21_X1 U18086 ( .B1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n15043), .A(
        n15024), .ZN(n15810) );
  XNOR2_X1 U18087 ( .A(n15025), .B(n15030), .ZN(n15026) );
  XNOR2_X1 U18088 ( .A(n15027), .B(n15026), .ZN(n15809) );
  AOI21_X1 U18089 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15029), .A(
        n15028), .ZN(n15045) );
  NOR2_X1 U18090 ( .A1(n12161), .A2(n18600), .ZN(n15032) );
  NAND2_X1 U18091 ( .A1(n15862), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15047) );
  AOI221_X1 U18092 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C1(n13760), .C2(n15030), .A(
        n15047), .ZN(n15031) );
  AOI211_X1 U18093 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n15045), .A(
        n15032), .B(n15031), .ZN(n15036) );
  OAI22_X1 U18094 ( .A1(n18539), .A2(n15898), .B1(n18839), .B2(n15033), .ZN(
        n15034) );
  INV_X1 U18095 ( .A(n15034), .ZN(n15035) );
  OAI211_X1 U18096 ( .C1(n15809), .C2(n18859), .A(n15036), .B(n15035), .ZN(
        n15037) );
  INV_X1 U18097 ( .A(n15037), .ZN(n15038) );
  OAI21_X1 U18098 ( .B1(n15810), .B2(n18861), .A(n15038), .ZN(P2_U3035) );
  INV_X1 U18099 ( .A(n15052), .ZN(n15055) );
  NOR2_X1 U18100 ( .A1(n15053), .A2(n15055), .ZN(n15042) );
  NAND2_X1 U18101 ( .A1(n15040), .A2(n15039), .ZN(n15041) );
  XNOR2_X1 U18102 ( .A(n15042), .B(n15041), .ZN(n15814) );
  AOI21_X1 U18103 ( .B1(n13760), .B2(n15059), .A(n15043), .ZN(n15815) );
  NAND2_X1 U18104 ( .A1(n15815), .A2(n18849), .ZN(n15051) );
  NOR2_X1 U18105 ( .A1(n12159), .A2(n18600), .ZN(n15044) );
  AOI21_X1 U18106 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n15045), .A(
        n15044), .ZN(n15046) );
  OAI21_X1 U18107 ( .B1(n15898), .B2(n18565), .A(n15046), .ZN(n15049) );
  NOR2_X1 U18108 ( .A1(n15047), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15048) );
  AOI211_X1 U18109 ( .C1(n18562), .C2(n18868), .A(n15049), .B(n15048), .ZN(
        n15050) );
  OAI211_X1 U18110 ( .C1(n15814), .C2(n18859), .A(n15051), .B(n15050), .ZN(
        P2_U3036) );
  NAND2_X1 U18111 ( .A1(n15053), .A2(n15052), .ZN(n15058) );
  OAI21_X1 U18112 ( .B1(n15056), .B2(n15055), .A(n15054), .ZN(n15057) );
  NAND2_X1 U18113 ( .A1(n15058), .A2(n15057), .ZN(n15819) );
  OAI21_X1 U18114 ( .B1(n15060), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15059), .ZN(n15820) );
  OR2_X1 U18115 ( .A1(n15820), .A2(n18861), .ZN(n15070) );
  NAND2_X1 U18116 ( .A1(n15862), .A2(n15061), .ZN(n15065) );
  INV_X1 U18117 ( .A(n18576), .ZN(n15063) );
  NOR2_X1 U18118 ( .A1(n12156), .A2(n18600), .ZN(n15062) );
  AOI21_X1 U18119 ( .B1(n18875), .B2(n15063), .A(n15062), .ZN(n15064) );
  OAI211_X1 U18120 ( .C1(n18839), .C2(n15066), .A(n15065), .B(n15064), .ZN(
        n15067) );
  AOI21_X1 U18121 ( .B1(n15068), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15067), .ZN(n15069) );
  OAI211_X1 U18122 ( .C1(n15819), .C2(n18859), .A(n15070), .B(n15069), .ZN(
        P2_U3037) );
  NAND2_X1 U18123 ( .A1(n15071), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15075) );
  NOR2_X1 U18124 ( .A1(n19470), .A2(n18600), .ZN(n15073) );
  NOR2_X1 U18125 ( .A1(n18599), .A2(n15898), .ZN(n15072) );
  AOI211_X1 U18126 ( .C1(n18868), .C2(n18596), .A(n15073), .B(n15072), .ZN(
        n15074) );
  OAI211_X1 U18127 ( .C1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n15881), .A(
        n15075), .B(n15074), .ZN(n15076) );
  AOI21_X1 U18128 ( .B1(n15077), .B2(n18846), .A(n15076), .ZN(n15078) );
  OAI21_X1 U18129 ( .B1(n15079), .B2(n18861), .A(n15078), .ZN(P2_U3039) );
  NOR2_X1 U18130 ( .A1(n18839), .A2(n15080), .ZN(n15085) );
  INV_X1 U18131 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15083) );
  INV_X1 U18132 ( .A(n18869), .ZN(n15082) );
  AOI211_X1 U18133 ( .C1(n15083), .C2(n10038), .A(n15082), .B(n15081), .ZN(
        n15084) );
  AOI211_X1 U18134 ( .C1(n18849), .C2(n15086), .A(n15085), .B(n15084), .ZN(
        n15091) );
  AOI22_X1 U18135 ( .A1(n18875), .A2(n19553), .B1(n18855), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15090) );
  NAND2_X1 U18136 ( .A1(n18846), .A2(n15087), .ZN(n15088) );
  NAND4_X1 U18137 ( .A1(n15091), .A2(n15090), .A3(n15089), .A4(n15088), .ZN(
        P2_U3045) );
  INV_X1 U18138 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16577) );
  INV_X1 U18139 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n16604) );
  INV_X1 U18140 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n16647) );
  INV_X1 U18141 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n16308) );
  INV_X1 U18142 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n15096) );
  INV_X1 U18143 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n16759) );
  INV_X1 U18144 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n16767) );
  INV_X1 U18145 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n16480) );
  AOI21_X2 U18146 ( .B1(n15095), .B2(n15094), .A(n18243), .ZN(n15420) );
  NAND2_X1 U18147 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16752), .ZN(n16748) );
  AND4_X1 U18148 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(P3_EBX_REG_12__SCAN_IN), 
        .A3(P3_EBX_REG_11__SCAN_IN), .A4(P3_EBX_REG_10__SCAN_IN), .ZN(n16645)
         );
  NAND2_X1 U18149 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16589), .ZN(n16578) );
  NAND4_X1 U18150 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(P3_EBX_REG_24__SCAN_IN), .A4(P3_EBX_REG_23__SCAN_IN), .ZN(n16523)
         );
  NOR2_X2 U18151 ( .A1(n16546), .A2(n16523), .ZN(n16537) );
  NAND2_X1 U18152 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n16537), .ZN(n15172) );
  INV_X1 U18153 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n16172) );
  NOR2_X1 U18154 ( .A1(n16890), .A2(n16772), .ZN(n16775) );
  NAND2_X1 U18155 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n16522) );
  NOR2_X1 U18156 ( .A1(n16765), .A2(n16537), .ZN(n16535) );
  AOI22_X1 U18157 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15101) );
  AOI22_X1 U18158 ( .A1(n9616), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16721), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15100) );
  AOI22_X1 U18159 ( .A1(n9630), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n15241), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15099) );
  AOI22_X1 U18160 ( .A1(n9612), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9641), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15098) );
  NAND4_X1 U18161 ( .A1(n15101), .A2(n15100), .A3(n15099), .A4(n15098), .ZN(
        n15107) );
  AOI22_X1 U18162 ( .A1(n15248), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n16634), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15105) );
  AOI22_X1 U18163 ( .A1(n15219), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n16741), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15104) );
  AOI22_X1 U18164 ( .A1(n16508), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9620), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15103) );
  AOI22_X1 U18165 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9629), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15102) );
  NAND4_X1 U18166 ( .A1(n15105), .A2(n15104), .A3(n15103), .A4(n15102), .ZN(
        n15106) );
  NOR2_X1 U18167 ( .A1(n15107), .A2(n15106), .ZN(n16519) );
  AOI22_X1 U18168 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9629), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15111) );
  AOI22_X1 U18169 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9620), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15110) );
  AOI22_X1 U18170 ( .A1(n16741), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15109) );
  AOI22_X1 U18171 ( .A1(n9613), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9642), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15108) );
  NAND4_X1 U18172 ( .A1(n15111), .A2(n15110), .A3(n15109), .A4(n15108), .ZN(
        n15117) );
  AOI22_X1 U18173 ( .A1(n9630), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n16634), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15115) );
  AOI22_X1 U18174 ( .A1(n9616), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(n9622), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15114) );
  AOI22_X1 U18175 ( .A1(n16733), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n16668), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15113) );
  AOI22_X1 U18176 ( .A1(n15219), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n16721), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15112) );
  NAND4_X1 U18177 ( .A1(n15115), .A2(n15114), .A3(n15113), .A4(n15112), .ZN(
        n15116) );
  NOR2_X1 U18178 ( .A1(n15117), .A2(n15116), .ZN(n16534) );
  AOI22_X1 U18179 ( .A1(n15219), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9621), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n15121) );
  AOI22_X1 U18180 ( .A1(n16733), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n16723), .ZN(n15120) );
  AOI22_X1 U18181 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n9616), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n16716), .ZN(n15119) );
  AOI22_X1 U18182 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n9640), .B1(n9611), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15118) );
  NAND4_X1 U18183 ( .A1(n15121), .A2(n15120), .A3(n15119), .A4(n15118), .ZN(
        n15127) );
  AOI22_X1 U18184 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n9622), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n15217), .ZN(n15125) );
  AOI22_X1 U18185 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n15248), .B1(
        n16721), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n15124) );
  AOI22_X1 U18186 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n9630), .B1(
        n16634), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n15123) );
  AOI22_X1 U18187 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n9629), .ZN(n15122) );
  NAND4_X1 U18188 ( .A1(n15125), .A2(n15124), .A3(n15123), .A4(n15122), .ZN(
        n15126) );
  NOR2_X1 U18189 ( .A1(n15127), .A2(n15126), .ZN(n16543) );
  AOI22_X1 U18190 ( .A1(n9613), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9620), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15138) );
  AOI22_X1 U18191 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15137) );
  INV_X1 U18192 ( .A(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n20695) );
  AOI22_X1 U18193 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n15241), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15129) );
  OAI21_X1 U18194 ( .B1(n16435), .B2(n20695), .A(n15129), .ZN(n15135) );
  AOI22_X1 U18195 ( .A1(n9616), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(n9629), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15133) );
  AOI22_X1 U18196 ( .A1(n9630), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n16668), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15132) );
  AOI22_X1 U18197 ( .A1(n16733), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n16721), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15131) );
  AOI22_X1 U18198 ( .A1(n16741), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9641), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15130) );
  NAND4_X1 U18199 ( .A1(n15133), .A2(n15132), .A3(n15131), .A4(n15130), .ZN(
        n15134) );
  AOI211_X1 U18200 ( .C1(n15219), .C2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A(
        n15135), .B(n15134), .ZN(n15136) );
  NAND3_X1 U18201 ( .A1(n15138), .A2(n15137), .A3(n15136), .ZN(n16548) );
  AOI22_X1 U18202 ( .A1(n15248), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9612), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15149) );
  AOI22_X1 U18203 ( .A1(n16733), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9620), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15148) );
  INV_X1 U18204 ( .A(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n20577) );
  AOI22_X1 U18205 ( .A1(n16738), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n16741), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15139) );
  OAI21_X1 U18206 ( .B1(n16435), .B2(n20577), .A(n15139), .ZN(n15146) );
  AOI22_X1 U18207 ( .A1(n15219), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9629), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15144) );
  AOI22_X1 U18208 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n15241), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15143) );
  AOI22_X1 U18209 ( .A1(n9642), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15142) );
  AOI22_X1 U18210 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9616), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15141) );
  NAND4_X1 U18211 ( .A1(n15144), .A2(n15143), .A3(n15142), .A4(n15141), .ZN(
        n15145) );
  AOI211_X1 U18212 ( .C1(n16682), .C2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n15146), .B(n15145), .ZN(n15147) );
  NAND3_X1 U18213 ( .A1(n15149), .A2(n15148), .A3(n15147), .ZN(n16549) );
  NAND2_X1 U18214 ( .A1(n16548), .A2(n16549), .ZN(n16547) );
  NOR2_X1 U18215 ( .A1(n16543), .A2(n16547), .ZN(n16540) );
  AOI22_X1 U18216 ( .A1(n15219), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15160) );
  AOI22_X1 U18217 ( .A1(n16733), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9630), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n15159) );
  AOI22_X1 U18218 ( .A1(n9612), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n16721), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15150) );
  OAI21_X1 U18219 ( .B1(n15151), .B2(n20650), .A(n15150), .ZN(n15157) );
  AOI22_X1 U18220 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9620), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15155) );
  AOI22_X1 U18221 ( .A1(n16723), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n16634), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n15154) );
  AOI22_X1 U18222 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n15248), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15153) );
  AOI22_X1 U18223 ( .A1(n15241), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9642), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15152) );
  NAND4_X1 U18224 ( .A1(n15155), .A2(n15154), .A3(n15153), .A4(n15152), .ZN(
        n15156) );
  AOI211_X1 U18225 ( .C1(n9616), .C2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A(
        n15157), .B(n15156), .ZN(n15158) );
  NAND3_X1 U18226 ( .A1(n15160), .A2(n15159), .A3(n15158), .ZN(n16539) );
  NAND2_X1 U18227 ( .A1(n16540), .A2(n16539), .ZN(n16538) );
  NOR2_X1 U18228 ( .A1(n16534), .A2(n16538), .ZN(n16533) );
  AOI22_X1 U18229 ( .A1(n16682), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9616), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15170) );
  AOI22_X1 U18230 ( .A1(n9611), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9629), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n15169) );
  AOI22_X1 U18231 ( .A1(n9641), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n16634), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15161) );
  OAI21_X1 U18232 ( .B1(n9683), .B2(n20658), .A(n15161), .ZN(n15167) );
  AOI22_X1 U18233 ( .A1(n16733), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9622), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15165) );
  AOI22_X1 U18234 ( .A1(n15219), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9621), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15164) );
  AOI22_X1 U18235 ( .A1(n15248), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9620), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15163) );
  AOI22_X1 U18236 ( .A1(n16738), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15162) );
  NAND4_X1 U18237 ( .A1(n15165), .A2(n15164), .A3(n15163), .A4(n15162), .ZN(
        n15166) );
  AOI211_X1 U18238 ( .C1(n16722), .C2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A(
        n15167), .B(n15166), .ZN(n15168) );
  NAND3_X1 U18239 ( .A1(n15170), .A2(n15169), .A3(n15168), .ZN(n16529) );
  NAND2_X1 U18240 ( .A1(n16533), .A2(n16529), .ZN(n16528) );
  XOR2_X1 U18241 ( .A(n16519), .B(n16528), .Z(n16794) );
  NAND2_X1 U18242 ( .A1(n16765), .A2(n16794), .ZN(n15171) );
  OAI221_X1 U18243 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n15172), .C1(n16172), 
        .C2(n16527), .A(n15171), .ZN(P3_U2675) );
  AOI22_X1 U18244 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n16634), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15176) );
  AOI22_X1 U18245 ( .A1(n15248), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n16738), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15175) );
  AOI22_X1 U18246 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9616), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15174) );
  AOI22_X1 U18247 ( .A1(n9641), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(n9620), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15173) );
  NAND4_X1 U18248 ( .A1(n15176), .A2(n15175), .A3(n15174), .A4(n15173), .ZN(
        n15182) );
  AOI22_X1 U18249 ( .A1(n16733), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9622), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15180) );
  AOI22_X1 U18250 ( .A1(n15219), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16741), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15179) );
  AOI22_X1 U18251 ( .A1(n9630), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9611), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15178) );
  AOI22_X1 U18252 ( .A1(n9629), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15177) );
  NAND4_X1 U18253 ( .A1(n15180), .A2(n15179), .A3(n15178), .A4(n15177), .ZN(
        n15181) );
  NOR2_X1 U18254 ( .A1(n15182), .A2(n15181), .ZN(n16873) );
  INV_X1 U18255 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n16337) );
  INV_X1 U18256 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16348) );
  INV_X1 U18257 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n16701) );
  NOR4_X1 U18258 ( .A1(n16890), .A2(n16348), .A3(n16701), .A4(n16730), .ZN(
        n16677) );
  INV_X1 U18259 ( .A(n16677), .ZN(n16702) );
  NOR2_X1 U18260 ( .A1(n16337), .A2(n16702), .ZN(n16690) );
  OAI211_X1 U18261 ( .C1(n16690), .C2(P3_EBX_REG_13__SCAN_IN), .A(n16774), .B(
        n15183), .ZN(n15184) );
  OAI21_X1 U18262 ( .B1(n16873), .B2(n16774), .A(n15184), .ZN(P3_U2690) );
  NAND2_X1 U18263 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n17895) );
  NOR2_X1 U18264 ( .A1(n18388), .A2(n17044), .ZN(n15186) );
  AOI221_X1 U18265 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n17895), .C1(n15186), 
        .C2(n17895), .A(n15185), .ZN(n17729) );
  NOR2_X1 U18266 ( .A1(n15187), .A2(n17987), .ZN(n15189) );
  OAI21_X1 U18267 ( .B1(n15189), .B2(n15188), .A(n17730), .ZN(n17727) );
  AOI22_X1 U18268 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n17729), .B1(
        n17727), .B2(n18209), .ZN(P3_U2865) );
  OR3_X1 U18269 ( .A1(n19521), .A2(n19537), .A3(n15190), .ZN(n15191) );
  OAI21_X1 U18270 ( .B1(n19530), .B2(n15192), .A(n15191), .ZN(P2_U3595) );
  XNOR2_X1 U18271 ( .A(n18391), .B(n16111), .ZN(n18407) );
  NOR2_X2 U18272 ( .A1(n18407), .A2(n15193), .ZN(n18218) );
  NAND2_X1 U18273 ( .A1(n18176), .A2(n15194), .ZN(n18190) );
  OAI21_X1 U18274 ( .B1(n15197), .B2(n15196), .A(n15195), .ZN(n18179) );
  INV_X1 U18275 ( .A(n17630), .ZN(n17534) );
  INV_X1 U18276 ( .A(n18222), .ZN(n15202) );
  AOI21_X1 U18277 ( .B1(n15199), .B2(n15198), .A(n15202), .ZN(n18223) );
  INV_X1 U18278 ( .A(n18223), .ZN(n15916) );
  NOR2_X1 U18279 ( .A1(n17741), .A2(n15200), .ZN(n15207) );
  OAI21_X1 U18280 ( .B1(n17748), .B2(n18391), .A(n18262), .ZN(n15201) );
  OAI21_X1 U18281 ( .B1(n15207), .B2(n15201), .A(n18385), .ZN(n16093) );
  NOR3_X1 U18282 ( .A1(n15205), .A2(n15202), .A3(n16093), .ZN(n15204) );
  AOI211_X1 U18283 ( .C1(n15205), .C2(n18219), .A(n15204), .B(n15203), .ZN(
        n15208) );
  NAND2_X1 U18284 ( .A1(n15207), .A2(n15206), .ZN(n15212) );
  AOI221_X4 U18285 ( .B1(n15916), .B2(n15208), .C1(n15212), .C2(n15208), .A(
        n18243), .ZN(n17716) );
  NAND2_X1 U18286 ( .A1(n17534), .A2(n17716), .ZN(n17706) );
  INV_X1 U18287 ( .A(n17706), .ZN(n17631) );
  INV_X1 U18288 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15984) );
  INV_X1 U18289 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15361) );
  INV_X1 U18290 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18366) );
  INV_X1 U18291 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17435) );
  INV_X1 U18292 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17418) );
  NAND2_X1 U18293 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17431) );
  NOR3_X1 U18294 ( .A1(n17435), .A2(n17418), .A3(n17431), .ZN(n15939) );
  NAND2_X1 U18295 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n15939), .ZN(
        n15972) );
  INV_X1 U18296 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17539) );
  INV_X1 U18297 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17522) );
  NOR2_X1 U18298 ( .A1(n17539), .A2(n17522), .ZN(n17513) );
  NAND2_X1 U18299 ( .A1(n17513), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17484) );
  INV_X1 U18300 ( .A(n17484), .ZN(n17467) );
  INV_X1 U18301 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17491) );
  NAND2_X1 U18302 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17482) );
  NOR2_X1 U18303 ( .A1(n17491), .A2(n17482), .ZN(n17475) );
  NAND2_X1 U18304 ( .A1(n17467), .A2(n17475), .ZN(n17473) );
  INV_X1 U18305 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17480) );
  NOR2_X1 U18306 ( .A1(n17473), .A2(n17480), .ZN(n15971) );
  INV_X1 U18307 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17609) );
  NOR2_X1 U18308 ( .A1(n17609), .A2(n17616), .ZN(n17604) );
  NAND2_X1 U18309 ( .A1(n17604), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17586) );
  NAND2_X1 U18310 ( .A1(n17597), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17580) );
  INV_X1 U18311 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17562) );
  INV_X1 U18312 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15341) );
  INV_X1 U18313 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17660) );
  INV_X1 U18314 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17634) );
  NOR3_X1 U18315 ( .A1(n15341), .A2(n17660), .A3(n17634), .ZN(n17509) );
  NAND3_X1 U18316 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n17508) );
  NAND2_X1 U18317 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17670) );
  NOR2_X1 U18318 ( .A1(n17508), .A2(n17670), .ZN(n17626) );
  NAND2_X1 U18319 ( .A1(n17509), .A2(n17626), .ZN(n17557) );
  NOR2_X1 U18320 ( .A1(n17507), .A2(n17557), .ZN(n17511) );
  NAND2_X1 U18321 ( .A1(n15971), .A2(n17511), .ZN(n17446) );
  NOR3_X1 U18322 ( .A1(n18366), .A2(n15972), .A3(n17446), .ZN(n15210) );
  INV_X1 U18323 ( .A(n15939), .ZN(n17413) );
  OAI21_X1 U18324 ( .B1(n17413), .B2(n17446), .A(n18190), .ZN(n15209) );
  AOI21_X1 U18325 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n17692) );
  NOR2_X1 U18326 ( .A1(n17692), .A2(n17508), .ZN(n17628) );
  NAND2_X1 U18327 ( .A1(n17628), .A2(n17509), .ZN(n17529) );
  NOR2_X1 U18328 ( .A1(n17507), .A2(n17529), .ZN(n17512) );
  NAND2_X1 U18329 ( .A1(n15971), .A2(n17512), .ZN(n17452) );
  OAI21_X1 U18330 ( .B1(n17413), .B2(n17452), .A(n18218), .ZN(n17416) );
  OAI211_X1 U18331 ( .C1(n18188), .C2(n15210), .A(n15209), .B(n17416), .ZN(
        n15409) );
  AOI21_X1 U18332 ( .B1(n17610), .B2(n15361), .A(n15409), .ZN(n15973) );
  AOI22_X1 U18333 ( .A1(n9616), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(n9620), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15216) );
  AOI22_X1 U18334 ( .A1(n9611), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n16721), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15215) );
  AOI22_X1 U18335 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n16741), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n15214) );
  AOI22_X1 U18336 ( .A1(n15241), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9642), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15213) );
  NAND4_X1 U18337 ( .A1(n15216), .A2(n15215), .A3(n15214), .A4(n15213), .ZN(
        n15225) );
  AOI22_X1 U18338 ( .A1(n9629), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15223) );
  AOI22_X1 U18339 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n15248), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15222) );
  AOI22_X1 U18340 ( .A1(n15219), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9630), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n15221) );
  AOI22_X1 U18341 ( .A1(n16733), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n16634), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15220) );
  NAND4_X1 U18342 ( .A1(n15223), .A2(n15222), .A3(n15221), .A4(n15220), .ZN(
        n15224) );
  NAND2_X1 U18343 ( .A1(n15980), .A2(n16902), .ZN(n17573) );
  NAND2_X1 U18344 ( .A1(n17716), .A2(n17472), .ZN(n17566) );
  INV_X1 U18345 ( .A(n17566), .ZN(n17639) );
  INV_X1 U18346 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n20668) );
  NOR3_X1 U18347 ( .A1(n15361), .A2(n15984), .A3(n20668), .ZN(n15940) );
  INV_X1 U18348 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17103) );
  NAND2_X1 U18349 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n15971), .ZN(
        n15348) );
  INV_X1 U18350 ( .A(n15348), .ZN(n15319) );
  AOI22_X1 U18351 ( .A1(n9612), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15230) );
  AOI22_X1 U18352 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9621), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15229) );
  AOI22_X1 U18353 ( .A1(n16740), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n16721), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15228) );
  AOI22_X1 U18354 ( .A1(n16682), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9642), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15227) );
  NAND4_X1 U18355 ( .A1(n15230), .A2(n15229), .A3(n15228), .A4(n15227), .ZN(
        n15236) );
  AOI22_X1 U18356 ( .A1(n9616), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(n9629), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15234) );
  AOI22_X1 U18357 ( .A1(n15248), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n16634), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15233) );
  AOI22_X1 U18358 ( .A1(n16723), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9620), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15232) );
  AOI22_X1 U18359 ( .A1(n16733), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n15241), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15231) );
  NAND4_X1 U18360 ( .A1(n15234), .A2(n15233), .A3(n15232), .A4(n15231), .ZN(
        n15235) );
  AOI22_X1 U18361 ( .A1(n9630), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9611), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15240) );
  AOI22_X1 U18362 ( .A1(n15248), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9620), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15239) );
  AOI22_X1 U18363 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9629), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15238) );
  AOI22_X1 U18364 ( .A1(n16733), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9640), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15237) );
  NAND4_X1 U18365 ( .A1(n15240), .A2(n15239), .A3(n15238), .A4(n15237), .ZN(
        n15247) );
  AOI22_X1 U18366 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n16741), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15245) );
  AOI22_X1 U18367 ( .A1(n9616), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(n9622), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15244) );
  AOI22_X1 U18368 ( .A1(n16740), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15243) );
  AOI22_X1 U18369 ( .A1(n16738), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16634), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15242) );
  NAND4_X1 U18370 ( .A1(n15245), .A2(n15244), .A3(n15243), .A4(n15242), .ZN(
        n15246) );
  AOI22_X1 U18371 ( .A1(n9616), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n16741), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15258) );
  AOI22_X1 U18372 ( .A1(n15248), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n16721), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15257) );
  AOI22_X1 U18373 ( .A1(n16682), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9620), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15249) );
  OAI21_X1 U18374 ( .B1(n9633), .B2(n20650), .A(n15249), .ZN(n15256) );
  AOI22_X1 U18375 ( .A1(n16740), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15255) );
  AOI22_X1 U18376 ( .A1(n13570), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9629), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15254) );
  AOI22_X1 U18377 ( .A1(n16508), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15251), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15253) );
  AOI22_X1 U18378 ( .A1(n9612), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9640), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15252) );
  AOI22_X1 U18379 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n9629), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n16723), .ZN(n15262) );
  AOI22_X1 U18380 ( .A1(n16682), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9612), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n15261) );
  AOI22_X1 U18381 ( .A1(n16740), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9616), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n15260) );
  AOI22_X1 U18382 ( .A1(n13570), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n9641), .ZN(n15259) );
  NAND4_X1 U18383 ( .A1(n15262), .A2(n15261), .A3(n15260), .A4(n15259), .ZN(
        n15268) );
  AOI22_X1 U18384 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n15241), .ZN(n15266) );
  AOI22_X1 U18385 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n16508), .B1(
        n16668), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15265) );
  AOI22_X1 U18386 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n16721), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n16716), .ZN(n15264) );
  AOI22_X1 U18387 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n15217), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n15251), .ZN(n15263) );
  NAND4_X1 U18388 ( .A1(n15266), .A2(n15265), .A3(n15264), .A4(n15263), .ZN(
        n15267) );
  NAND2_X1 U18389 ( .A1(n15321), .A2(n16930), .ZN(n15311) );
  AOI22_X1 U18390 ( .A1(n9622), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n9620), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15279) );
  AOI22_X1 U18391 ( .A1(n16738), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n16741), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15278) );
  AOI22_X1 U18392 ( .A1(n16634), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15270) );
  OAI21_X1 U18393 ( .B1(n9679), .B2(n20658), .A(n15270), .ZN(n15276) );
  AOI22_X1 U18394 ( .A1(n16740), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n16508), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15274) );
  AOI22_X1 U18395 ( .A1(n16739), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9629), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15273) );
  AOI22_X1 U18396 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(n9630), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15272) );
  AOI22_X1 U18397 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9641), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15271) );
  NAND4_X1 U18398 ( .A1(n15274), .A2(n15273), .A3(n15272), .A4(n15271), .ZN(
        n15275) );
  AOI211_X1 U18399 ( .C1(n9613), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n15276), .B(n15275), .ZN(n15277) );
  NAND3_X1 U18400 ( .A1(n15279), .A2(n15278), .A3(n15277), .ZN(n16914) );
  NAND2_X1 U18401 ( .A1(n15294), .A2(n16914), .ZN(n15293) );
  AOI22_X1 U18402 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(n9611), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n15290) );
  AOI22_X1 U18403 ( .A1(n16740), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n16722), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n15289) );
  AOI22_X1 U18404 ( .A1(n9642), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n16610), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n15280) );
  OAI21_X1 U18405 ( .B1(n15281), .B2(n20623), .A(n15280), .ZN(n15287) );
  AOI22_X1 U18406 ( .A1(n16723), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n16716), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n15285) );
  AOI22_X1 U18407 ( .A1(n16739), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n16721), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n15284) );
  AOI22_X1 U18408 ( .A1(n9616), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(n9629), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n15283) );
  AOI22_X1 U18409 ( .A1(n16733), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n16682), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n15282) );
  NAND4_X1 U18410 ( .A1(n15285), .A2(n15284), .A3(n15283), .A4(n15282), .ZN(
        n15286) );
  AOI211_X1 U18411 ( .C1(n15241), .C2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n15287), .B(n15286), .ZN(n15288) );
  NAND3_X1 U18412 ( .A1(n15290), .A2(n15289), .A3(n15288), .ZN(n16906) );
  NAND2_X1 U18413 ( .A1(n15292), .A2(n16906), .ZN(n15291) );
  AOI21_X1 U18414 ( .B1(n16902), .B2(n15291), .A(n17318), .ZN(n15317) );
  XOR2_X1 U18415 ( .A(n16906), .B(n15292), .Z(n15314) );
  NAND2_X1 U18416 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15314), .ZN(
        n15315) );
  INV_X1 U18417 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17667) );
  XOR2_X1 U18418 ( .A(n16910), .B(n15293), .Z(n17356) );
  XOR2_X1 U18419 ( .A(n16914), .B(n15294), .Z(n15295) );
  NAND2_X1 U18420 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n15295), .ZN(
        n15313) );
  XOR2_X1 U18421 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n15295), .Z(
        n17370) );
  NAND2_X1 U18422 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n15297), .ZN(
        n15309) );
  NAND2_X1 U18423 ( .A1(n15320), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15308) );
  AOI22_X1 U18424 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n16610), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15301) );
  AOI22_X1 U18425 ( .A1(n16738), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15300) );
  AOI22_X1 U18426 ( .A1(n9616), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(n9620), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15299) );
  AOI22_X1 U18427 ( .A1(n16682), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9641), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15298) );
  NAND4_X1 U18428 ( .A1(n15301), .A2(n15300), .A3(n15299), .A4(n15298), .ZN(
        n15307) );
  AOI22_X1 U18429 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n16741), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15305) );
  AOI22_X1 U18430 ( .A1(n9629), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(n9622), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15304) );
  AOI22_X1 U18431 ( .A1(n16740), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n16508), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n15303) );
  AOI22_X1 U18432 ( .A1(n16739), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9611), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15302) );
  NAND4_X1 U18433 ( .A1(n15305), .A2(n15304), .A3(n15303), .A4(n15302), .ZN(
        n15306) );
  NOR2_X1 U18434 ( .A1(n17407), .A2(n18366), .ZN(n17406) );
  NAND2_X1 U18435 ( .A1(n15308), .A2(n17398), .ZN(n17390) );
  NAND2_X1 U18436 ( .A1(n15309), .A2(n17389), .ZN(n15310) );
  NAND2_X1 U18437 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15310), .ZN(
        n15312) );
  INV_X1 U18438 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n17682) );
  XNOR2_X1 U18439 ( .A(n15310), .B(n17682), .ZN(n17380) );
  XOR2_X1 U18440 ( .A(n16918), .B(n15311), .Z(n17379) );
  NAND2_X1 U18441 ( .A1(n17380), .A2(n17379), .ZN(n17378) );
  NAND2_X1 U18442 ( .A1(n15312), .A2(n17378), .ZN(n17369) );
  NAND2_X1 U18443 ( .A1(n17370), .A2(n17369), .ZN(n17368) );
  NAND2_X1 U18444 ( .A1(n17356), .A2(n17357), .ZN(n17355) );
  XOR2_X1 U18445 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n15314), .Z(
        n17340) );
  NAND2_X1 U18446 ( .A1(n15317), .A2(n15316), .ZN(n15318) );
  NAND2_X1 U18447 ( .A1(n15319), .A2(n17541), .ZN(n17447) );
  NOR2_X1 U18448 ( .A1(n17103), .A2(n17447), .ZN(n17082) );
  NAND2_X1 U18449 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17082), .ZN(
        n17081) );
  NAND2_X1 U18450 ( .A1(n15940), .A2(n17042), .ZN(n15931) );
  NOR2_X1 U18451 ( .A1(n17468), .A2(n17680), .ZN(n17719) );
  NOR2_X1 U18452 ( .A1(n17407), .A2(n15320), .ZN(n15329) );
  NOR2_X1 U18453 ( .A1(n15329), .A2(n15321), .ZN(n15327) );
  NOR2_X1 U18454 ( .A1(n15327), .A2(n16918), .ZN(n15326) );
  NAND2_X1 U18455 ( .A1(n15326), .A2(n16914), .ZN(n15324) );
  NOR2_X1 U18456 ( .A1(n16910), .A2(n15324), .ZN(n15323) );
  NAND2_X1 U18457 ( .A1(n15323), .A2(n16906), .ZN(n15322) );
  NOR2_X1 U18458 ( .A1(n16902), .A2(n15322), .ZN(n15346) );
  XOR2_X1 U18459 ( .A(n15322), .B(n16902), .Z(n17334) );
  XOR2_X1 U18460 ( .A(n15323), .B(n16906), .Z(n15338) );
  XOR2_X1 U18461 ( .A(n15324), .B(n16910), .Z(n15325) );
  NAND2_X1 U18462 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n15325), .ZN(
        n15337) );
  XOR2_X1 U18463 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n15325), .Z(
        n17351) );
  XOR2_X1 U18464 ( .A(n15326), .B(n16914), .Z(n15335) );
  XOR2_X1 U18465 ( .A(n16918), .B(n15327), .Z(n15328) );
  NAND2_X1 U18466 ( .A1(n15328), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n15333) );
  XOR2_X1 U18467 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n15328), .Z(
        n17377) );
  INV_X1 U18468 ( .A(n17407), .ZN(n15424) );
  AOI21_X1 U18469 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n16930), .A(
        n15424), .ZN(n15331) );
  NOR2_X1 U18470 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n16930), .ZN(
        n15330) );
  AOI221_X1 U18471 ( .B1(n15424), .B2(n16930), .C1(n15331), .C2(n18366), .A(
        n15330), .ZN(n17387) );
  NAND2_X1 U18472 ( .A1(n17388), .A2(n17387), .ZN(n17386) );
  NAND2_X1 U18473 ( .A1(n15332), .A2(n17386), .ZN(n17376) );
  NAND2_X1 U18474 ( .A1(n17377), .A2(n17376), .ZN(n17375) );
  NAND2_X1 U18475 ( .A1(n15333), .A2(n17375), .ZN(n15334) );
  NAND2_X1 U18476 ( .A1(n15335), .A2(n15334), .ZN(n15336) );
  XOR2_X1 U18477 ( .A(n15335), .B(n15334), .Z(n17365) );
  NAND2_X1 U18478 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n17365), .ZN(
        n17364) );
  NAND2_X1 U18479 ( .A1(n15338), .A2(n15339), .ZN(n15340) );
  NAND2_X1 U18480 ( .A1(n17343), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17342) );
  NAND2_X1 U18481 ( .A1(n15346), .A2(n15342), .ZN(n15347) );
  NAND2_X1 U18482 ( .A1(n17334), .A2(n17333), .ZN(n15344) );
  NAND2_X1 U18483 ( .A1(n15346), .A2(n15345), .ZN(n15343) );
  OAI211_X1 U18484 ( .C1(n15346), .C2(n15345), .A(n15344), .B(n15343), .ZN(
        n17321) );
  NAND2_X1 U18485 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17321), .ZN(
        n17320) );
  NAND2_X1 U18486 ( .A1(n17450), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17091) );
  INV_X1 U18487 ( .A(n15940), .ZN(n15349) );
  NOR2_X1 U18488 ( .A1(n17415), .A2(n15349), .ZN(n15914) );
  INV_X1 U18489 ( .A(n15914), .ZN(n15932) );
  AOI22_X1 U18490 ( .A1(n17639), .A2(n15931), .B1(n17719), .B2(n15932), .ZN(
        n15410) );
  OAI211_X1 U18491 ( .C1(n15973), .C2(n17680), .A(n15410), .B(n17705), .ZN(
        n15350) );
  AOI21_X1 U18492 ( .B1(n17631), .B2(n15984), .A(n15350), .ZN(n15368) );
  NOR2_X1 U18493 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15352) );
  INV_X1 U18494 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17591) );
  INV_X1 U18495 ( .A(n17513), .ZN(n15355) );
  OR2_X1 U18496 ( .A1(n15355), .A2(n17200), .ZN(n17144) );
  INV_X1 U18497 ( .A(n17447), .ZN(n15358) );
  INV_X1 U18498 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17180) );
  NAND2_X1 U18499 ( .A1(n17180), .A2(n17235), .ZN(n17179) );
  NOR2_X1 U18500 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17179), .ZN(
        n15357) );
  INV_X1 U18501 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17474) );
  NAND2_X1 U18502 ( .A1(n15357), .A2(n17474), .ZN(n17145) );
  NOR2_X1 U18503 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17145), .ZN(
        n17127) );
  INV_X1 U18504 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17451) );
  NAND3_X1 U18505 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17109), .A3(
        n17102), .ZN(n17093) );
  NAND3_X1 U18506 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17318), .A3(
        n17060), .ZN(n15405) );
  NOR2_X1 U18507 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17318), .ZN(
        n15969) );
  XOR2_X1 U18508 ( .A(n15362), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .Z(
        n15951) );
  NAND2_X1 U18509 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15363) );
  NOR2_X1 U18510 ( .A1(n17415), .A2(n15363), .ZN(n15974) );
  INV_X1 U18511 ( .A(n17468), .ZN(n18217) );
  AOI21_X1 U18512 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n17602), .A(
        n18190), .ZN(n17690) );
  INV_X1 U18513 ( .A(n17690), .ZN(n15364) );
  AOI22_X1 U18514 ( .A1(n18218), .A2(n17512), .B1(n15364), .B2(n17511), .ZN(
        n15970) );
  INV_X1 U18515 ( .A(n15970), .ZN(n15365) );
  NAND2_X1 U18516 ( .A1(n15971), .A2(n15365), .ZN(n17428) );
  NOR3_X1 U18517 ( .A1(n15984), .A2(n17428), .A3(n15972), .ZN(n15960) );
  AOI21_X1 U18518 ( .B1(n15974), .B2(n18217), .A(n15960), .ZN(n15366) );
  NAND3_X1 U18519 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(n17042), .ZN(n15976) );
  OAI22_X1 U18520 ( .A1(n15366), .A2(n17680), .B1(n15976), .B2(n17566), .ZN(
        n15412) );
  AOI22_X1 U18521 ( .A1(n17613), .A2(n15951), .B1(n20668), .B2(n15412), .ZN(
        n15367) );
  NAND2_X1 U18522 ( .A1(n17715), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n15948) );
  OAI211_X1 U18523 ( .C1(n15368), .C2(n20668), .A(n15367), .B(n15948), .ZN(
        P3_U2833) );
  INV_X1 U18524 ( .A(n15369), .ZN(n15371) );
  NOR3_X1 U18525 ( .A1(n15371), .A2(n15370), .A3(n20315), .ZN(n15376) );
  AOI21_X1 U18526 ( .B1(n15376), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n15372), .ZN(n15373) );
  NAND2_X1 U18527 ( .A1(n15374), .A2(n15373), .ZN(n15375) );
  OAI21_X1 U18528 ( .B1(n15376), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n15375), .ZN(n15377) );
  AOI222_X1 U18529 ( .A1(n15378), .A2(n20262), .B1(n15378), .B2(n15377), .C1(
        n20262), .C2(n15377), .ZN(n15379) );
  AOI222_X1 U18530 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n15380), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15379), .C1(n15380), 
        .C2(n15379), .ZN(n15390) );
  NOR2_X1 U18531 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(P1_MORE_REG_SCAN_IN), .ZN(
        n15387) );
  INV_X1 U18532 ( .A(n15381), .ZN(n15382) );
  AND2_X1 U18533 ( .A1(n15383), .A2(n15382), .ZN(n15384) );
  OAI211_X1 U18534 ( .C1(n15387), .C2(n15386), .A(n15385), .B(n15384), .ZN(
        n15388) );
  AOI211_X1 U18535 ( .C1(n15390), .C2(n19833), .A(n15389), .B(n15388), .ZN(
        n15404) );
  INV_X1 U18536 ( .A(n11246), .ZN(n15393) );
  INV_X1 U18537 ( .A(n15391), .ZN(n15392) );
  NOR4_X1 U18538 ( .A1(n15393), .A2(n19853), .A3(n15416), .A4(n15392), .ZN(
        n15396) );
  OAI22_X1 U18539 ( .A1(n15396), .A2(n15395), .B1(n15394), .B2(n20546), .ZN(
        n15682) );
  AOI21_X1 U18540 ( .B1(n15404), .B2(n15682), .A(n20446), .ZN(n15689) );
  INV_X1 U18541 ( .A(n15689), .ZN(n15687) );
  OAI211_X1 U18542 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20546), .A(n15398), 
        .B(n15397), .ZN(n15402) );
  NOR2_X1 U18543 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15399), .ZN(n15400) );
  AOI22_X1 U18544 ( .A1(n20547), .A2(n15682), .B1(n20542), .B2(n15400), .ZN(
        n15401) );
  OAI21_X1 U18545 ( .B1(n15687), .B2(n15402), .A(n15401), .ZN(n15403) );
  OAI21_X1 U18546 ( .B1(n15404), .B2(n19602), .A(n15403), .ZN(P1_U3161) );
  NOR2_X1 U18547 ( .A1(n15927), .A2(n15926), .ZN(n15407) );
  XOR2_X1 U18548 ( .A(n15407), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .Z(
        n15943) );
  OAI21_X1 U18549 ( .B1(n17630), .B2(n15940), .A(n17716), .ZN(n15408) );
  OAI21_X1 U18550 ( .B1(n15409), .B2(n15408), .A(n9746), .ZN(n15968) );
  INV_X1 U18551 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15938) );
  AOI21_X1 U18552 ( .B1(n15410), .B2(n15968), .A(n15938), .ZN(n15411) );
  AOI21_X1 U18553 ( .B1(P3_REIP_REG_30__SCAN_IN), .B2(n17715), .A(n15411), 
        .ZN(n15414) );
  NAND3_X1 U18554 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15938), .A3(
        n15412), .ZN(n15413) );
  OAI211_X1 U18555 ( .C1(n15943), .C2(n17636), .A(n15414), .B(n15413), .ZN(
        P3_U2832) );
  INV_X1 U18556 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n19598) );
  INV_X1 U18557 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20462) );
  NOR2_X1 U18558 ( .A1(n20451), .A2(n20462), .ZN(n20456) );
  INV_X1 U18559 ( .A(HOLD), .ZN(n19451) );
  NOR2_X1 U18560 ( .A1(n19598), .A2(n19451), .ZN(n20454) );
  NAND2_X1 U18561 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n20452) );
  OAI21_X1 U18562 ( .B1(n20456), .B2(n20454), .A(n20452), .ZN(n15415) );
  OAI211_X1 U18563 ( .C1(n20546), .C2(n19598), .A(n15416), .B(n15415), .ZN(
        P1_U3195) );
  AND2_X1 U18564 ( .A1(n19745), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR2_X1 U18565 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15418) );
  NOR3_X1 U18566 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n15904), .A3(n19593), 
        .ZN(n19435) );
  NAND2_X1 U18567 ( .A1(n15905), .A2(n15906), .ZN(n15417) );
  AOI211_X1 U18568 ( .C1(n15418), .C2(n19263), .A(n19435), .B(n15417), .ZN(
        P2_U3178) );
  OAI221_X1 U18569 ( .B1(n15906), .B2(n19574), .C1(n15906), .C2(n12450), .A(
        n19104), .ZN(n19570) );
  NOR2_X1 U18570 ( .A1(n15419), .A2(n19570), .ZN(P2_U3047) );
  AND3_X1 U18571 ( .A1(n17741), .A2(n16111), .A3(n15420), .ZN(n15421) );
  NAND2_X1 U18572 ( .A1(n17778), .A2(n15426), .ZN(n16928) );
  INV_X1 U18573 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17009) );
  NOR2_X1 U18574 ( .A1(n16922), .A2(n15423), .ZN(n16932) );
  AOI22_X1 U18575 ( .A1(n16932), .A2(BUF2_REG_0__SCAN_IN), .B1(n16931), .B2(
        n15424), .ZN(n15425) );
  OAI221_X1 U18576 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n16928), .C1(n17009), 
        .C2(n15426), .A(n15425), .ZN(P3_U2735) );
  AND3_X1 U18577 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n19636), .A3(n15427), 
        .ZN(n15431) );
  OAI22_X1 U18578 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n15429), .B1(n15428), 
        .B2(n19662), .ZN(n15430) );
  AOI211_X1 U18579 ( .C1(n19675), .C2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n15431), .B(n15430), .ZN(n15436) );
  INV_X1 U18580 ( .A(n15432), .ZN(n15433) );
  AOI22_X1 U18581 ( .A1(n15434), .A2(n19659), .B1(n15433), .B2(n19644), .ZN(
        n15435) );
  OAI211_X1 U18582 ( .C1(n15437), .C2(n19681), .A(n15436), .B(n15435), .ZN(
        P1_U2815) );
  INV_X1 U18583 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n15441) );
  OAI22_X1 U18584 ( .A1(n15439), .A2(n19691), .B1(n15438), .B2(n19662), .ZN(
        n15440) );
  AOI221_X1 U18585 ( .B1(n15443), .B2(P1_REIP_REG_24__SCAN_IN), .C1(n15442), 
        .C2(n15441), .A(n15440), .ZN(n15447) );
  AOI22_X1 U18586 ( .A1(n15445), .A2(n19659), .B1(n15444), .B2(n19644), .ZN(
        n15446) );
  OAI211_X1 U18587 ( .C1(n15448), .C2(n19681), .A(n15447), .B(n15446), .ZN(
        P1_U2816) );
  OAI21_X1 U18588 ( .B1(n15449), .B2(n15461), .A(n19636), .ZN(n15468) );
  NAND2_X1 U18589 ( .A1(n15450), .A2(n20488), .ZN(n15460) );
  AOI22_X1 U18590 ( .A1(n15451), .A2(n19644), .B1(P1_EBX_REG_22__SCAN_IN), 
        .B2(n19687), .ZN(n15452) );
  OAI21_X1 U18591 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(n15453), .A(n15452), 
        .ZN(n15457) );
  OAI22_X1 U18592 ( .A1(n15455), .A2(n15470), .B1(n19681), .B2(n15454), .ZN(
        n15456) );
  AOI211_X1 U18593 ( .C1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(n19675), .A(
        n15457), .B(n15456), .ZN(n15458) );
  OAI221_X1 U18594 ( .B1(n15459), .B2(n15468), .C1(n15459), .C2(n15460), .A(
        n15458), .ZN(P1_U2818) );
  NOR2_X1 U18595 ( .A1(n15468), .A2(n20488), .ZN(n15463) );
  INV_X1 U18596 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n15536) );
  OAI22_X1 U18597 ( .A1(n15536), .A2(n19662), .B1(n15461), .B2(n15460), .ZN(
        n15462) );
  AOI211_X1 U18598 ( .C1(n19675), .C2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15463), .B(n15462), .ZN(n15465) );
  AOI22_X1 U18599 ( .A1(n15534), .A2(n19659), .B1(n19686), .B2(n15533), .ZN(
        n15464) );
  OAI211_X1 U18600 ( .C1(n15466), .C2(n19690), .A(n15465), .B(n15464), .ZN(
        P1_U2819) );
  AOI22_X1 U18601 ( .A1(n15467), .A2(n19644), .B1(P1_EBX_REG_20__SCAN_IN), 
        .B2(n19687), .ZN(n15475) );
  NOR3_X1 U18602 ( .A1(n14178), .A2(n15481), .A3(n15502), .ZN(n15477) );
  AOI21_X1 U18603 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(n15477), .A(
        P1_REIP_REG_20__SCAN_IN), .ZN(n15469) );
  OAI22_X1 U18604 ( .A1(n15471), .A2(n15470), .B1(n15469), .B2(n15468), .ZN(
        n15472) );
  AOI21_X1 U18605 ( .B1(n19686), .B2(n15473), .A(n15472), .ZN(n15474) );
  OAI211_X1 U18606 ( .C1(n15476), .C2(n19691), .A(n15475), .B(n15474), .ZN(
        P1_U2820) );
  AOI22_X1 U18607 ( .A1(P1_EBX_REG_19__SCAN_IN), .A2(n19687), .B1(n15477), 
        .B2(n14355), .ZN(n15479) );
  AOI21_X1 U18608 ( .B1(n19675), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n19678), .ZN(n15478) );
  OAI211_X1 U18609 ( .C1(n15552), .C2(n19690), .A(n15479), .B(n15478), .ZN(
        n15480) );
  AOI21_X1 U18610 ( .B1(n15548), .B2(n19659), .A(n15480), .ZN(n15483) );
  NOR3_X1 U18611 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n15481), .A3(n15502), 
        .ZN(n15489) );
  OAI21_X1 U18612 ( .B1(n15489), .B2(n15485), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n15482) );
  OAI211_X1 U18613 ( .C1(n15484), .C2(n19681), .A(n15483), .B(n15482), .ZN(
        P1_U2821) );
  AOI22_X1 U18614 ( .A1(P1_EBX_REG_18__SCAN_IN), .A2(n19687), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n15485), .ZN(n15486) );
  OAI211_X1 U18615 ( .C1(n19691), .C2(n15487), .A(n15486), .B(n19653), .ZN(
        n15488) );
  AOI211_X1 U18616 ( .C1(n19644), .C2(n15490), .A(n15489), .B(n15488), .ZN(
        n15494) );
  INV_X1 U18617 ( .A(n15491), .ZN(n15492) );
  NAND2_X1 U18618 ( .A1(n15492), .A2(n19659), .ZN(n15493) );
  OAI211_X1 U18619 ( .C1(n15599), .C2(n19681), .A(n15494), .B(n15493), .ZN(
        P1_U2822) );
  INV_X1 U18620 ( .A(n15495), .ZN(n15501) );
  NOR3_X1 U18621 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n14402), .A3(n15502), 
        .ZN(n15500) );
  AOI22_X1 U18622 ( .A1(n15496), .A2(n19644), .B1(P1_EBX_REG_16__SCAN_IN), 
        .B2(n19687), .ZN(n15497) );
  OAI211_X1 U18623 ( .C1(n19691), .C2(n15498), .A(n19653), .B(n15497), .ZN(
        n15499) );
  AOI211_X1 U18624 ( .C1(n15501), .C2(n19659), .A(n15500), .B(n15499), .ZN(
        n15504) );
  NOR2_X1 U18625 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n15502), .ZN(n15509) );
  OAI21_X1 U18626 ( .B1(n15509), .B2(n15506), .A(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n15503) );
  OAI211_X1 U18627 ( .C1(n15505), .C2(n19681), .A(n15504), .B(n15503), .ZN(
        P1_U2824) );
  AOI22_X1 U18628 ( .A1(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n19675), .B1(
        P1_REIP_REG_15__SCAN_IN), .B2(n15506), .ZN(n15507) );
  OAI211_X1 U18629 ( .C1(n19662), .C2(n15539), .A(n15507), .B(n19653), .ZN(
        n15508) );
  AOI211_X1 U18630 ( .C1(n19644), .C2(n15559), .A(n15509), .B(n15508), .ZN(
        n15512) );
  INV_X1 U18631 ( .A(n15510), .ZN(n15537) );
  AOI22_X1 U18632 ( .A1(n15560), .A2(n19659), .B1(n19686), .B2(n15537), .ZN(
        n15511) );
  NAND2_X1 U18633 ( .A1(n15512), .A2(n15511), .ZN(P1_U2825) );
  AOI22_X1 U18634 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19675), .B1(
        P1_EBX_REG_12__SCAN_IN), .B2(n19687), .ZN(n15519) );
  AOI21_X1 U18635 ( .B1(n15513), .B2(n19686), .A(n19678), .ZN(n15518) );
  INV_X1 U18636 ( .A(n15543), .ZN(n15564) );
  AOI22_X1 U18637 ( .A1(n15565), .A2(n19644), .B1(n19659), .B2(n15564), .ZN(
        n15517) );
  INV_X1 U18638 ( .A(n15514), .ZN(n15515) );
  OAI221_X1 U18639 ( .B1(P1_REIP_REG_12__SCAN_IN), .B2(P1_REIP_REG_11__SCAN_IN), .C1(P1_REIP_REG_12__SCAN_IN), .C2(n15525), .A(n15515), .ZN(n15516) );
  NAND4_X1 U18640 ( .A1(n15519), .A2(n15518), .A3(n15517), .A4(n15516), .ZN(
        P1_U2828) );
  INV_X1 U18641 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15541) );
  INV_X1 U18642 ( .A(n15520), .ZN(n15521) );
  AOI21_X1 U18643 ( .B1(n15523), .B2(n15522), .A(n15521), .ZN(n15620) );
  INV_X1 U18644 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n15524) );
  AOI22_X1 U18645 ( .A1(n19686), .A2(n15620), .B1(n15525), .B2(n15524), .ZN(
        n15526) );
  OAI21_X1 U18646 ( .B1(n15541), .B2(n19662), .A(n15526), .ZN(n15527) );
  AOI211_X1 U18647 ( .C1(n19675), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n19678), .B(n15527), .ZN(n15532) );
  XNOR2_X1 U18648 ( .A(n15529), .B(n15528), .ZN(n15576) );
  AOI22_X1 U18649 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n15530), .B1(n19659), 
        .B2(n15576), .ZN(n15531) );
  OAI211_X1 U18650 ( .C1(n15579), .C2(n19690), .A(n15532), .B(n15531), .ZN(
        P1_U2829) );
  AOI22_X1 U18651 ( .A1(n15534), .A2(n19706), .B1(n19705), .B2(n15533), .ZN(
        n15535) );
  OAI21_X1 U18652 ( .B1(n19710), .B2(n15536), .A(n15535), .ZN(P1_U2851) );
  AOI22_X1 U18653 ( .A1(n15560), .A2(n19706), .B1(n19705), .B2(n15537), .ZN(
        n15538) );
  OAI21_X1 U18654 ( .B1(n19710), .B2(n15539), .A(n15538), .ZN(P1_U2857) );
  AOI22_X1 U18655 ( .A1(n15576), .A2(n19706), .B1(n19705), .B2(n15620), .ZN(
        n15540) );
  OAI21_X1 U18656 ( .B1(n19710), .B2(n15541), .A(n15540), .ZN(P1_U2861) );
  AOI22_X1 U18657 ( .A1(P1_EAX_REG_12__SCAN_IN), .A2(n15545), .B1(n15544), 
        .B2(n19758), .ZN(n15542) );
  OAI21_X1 U18658 ( .B1(n19714), .B2(n15543), .A(n15542), .ZN(P1_U2892) );
  INV_X1 U18659 ( .A(n15576), .ZN(n15547) );
  AOI22_X1 U18660 ( .A1(P1_EAX_REG_11__SCAN_IN), .A2(n15545), .B1(n15544), 
        .B2(n19756), .ZN(n15546) );
  OAI21_X1 U18661 ( .B1(n19714), .B2(n15547), .A(n15546), .ZN(P1_U2893) );
  AOI22_X1 U18662 ( .A1(n19782), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n19781), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15551) );
  AOI22_X1 U18663 ( .A1(n15549), .A2(n19788), .B1(n19787), .B2(n15548), .ZN(
        n15550) );
  OAI211_X1 U18664 ( .C1(n19793), .C2(n15552), .A(n15551), .B(n15550), .ZN(
        P1_U2980) );
  AOI22_X1 U18665 ( .A1(n19782), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n19781), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n15557) );
  INV_X1 U18666 ( .A(n15553), .ZN(n15555) );
  AOI22_X1 U18667 ( .A1(n15555), .A2(n19787), .B1(n15566), .B2(n15554), .ZN(
        n15556) );
  OAI211_X1 U18668 ( .C1(n15558), .C2(n19608), .A(n15557), .B(n15556), .ZN(
        P1_U2982) );
  AOI22_X1 U18669 ( .A1(n19782), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n19781), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n15562) );
  AOI22_X1 U18670 ( .A1(n15560), .A2(n19787), .B1(n15559), .B2(n15566), .ZN(
        n15561) );
  OAI211_X1 U18671 ( .C1(n15563), .C2(n19608), .A(n15562), .B(n15561), .ZN(
        P1_U2984) );
  AOI22_X1 U18672 ( .A1(n19782), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n19781), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15568) );
  AOI22_X1 U18673 ( .A1(n15566), .A2(n15565), .B1(n19787), .B2(n15564), .ZN(
        n15567) );
  OAI211_X1 U18674 ( .C1(n15569), .C2(n19608), .A(n15568), .B(n15567), .ZN(
        P1_U2987) );
  AOI22_X1 U18675 ( .A1(n19782), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n19781), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15578) );
  NOR2_X1 U18676 ( .A1(n15570), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15574) );
  NOR2_X1 U18677 ( .A1(n15571), .A2(n15629), .ZN(n15573) );
  MUX2_X1 U18678 ( .A(n15574), .B(n15573), .S(n15572), .Z(n15575) );
  XOR2_X1 U18679 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n15575), .Z(
        n15622) );
  AOI22_X1 U18680 ( .A1(n19788), .A2(n15622), .B1(n19787), .B2(n15576), .ZN(
        n15577) );
  OAI211_X1 U18681 ( .C1(n19793), .C2(n15579), .A(n15578), .B(n15577), .ZN(
        P1_U2988) );
  AOI22_X1 U18682 ( .A1(n19782), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n19781), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15585) );
  NAND2_X1 U18683 ( .A1(n15581), .A2(n15580), .ZN(n15582) );
  XNOR2_X1 U18684 ( .A(n15583), .B(n15582), .ZN(n15662) );
  AOI22_X1 U18685 ( .A1(n15662), .A2(n19788), .B1(n19787), .B2(n19638), .ZN(
        n15584) );
  OAI211_X1 U18686 ( .C1(n19793), .C2(n19642), .A(n15585), .B(n15584), .ZN(
        P1_U2992) );
  AOI22_X1 U18687 ( .A1(n19782), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n19781), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n15590) );
  XNOR2_X1 U18688 ( .A(n15586), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15587) );
  XNOR2_X1 U18689 ( .A(n15588), .B(n15587), .ZN(n15671) );
  AOI22_X1 U18690 ( .A1(n15671), .A2(n19788), .B1(n19787), .B2(n19707), .ZN(
        n15589) );
  OAI211_X1 U18691 ( .C1(n19793), .C2(n19656), .A(n15590), .B(n15589), .ZN(
        P1_U2993) );
  AOI22_X1 U18692 ( .A1(n19782), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n19781), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n15597) );
  OAI21_X1 U18693 ( .B1(n15593), .B2(n15592), .A(n15591), .ZN(n15594) );
  INV_X1 U18694 ( .A(n15594), .ZN(n15676) );
  INV_X1 U18695 ( .A(n15595), .ZN(n19670) );
  AOI22_X1 U18696 ( .A1(n15676), .A2(n19788), .B1(n19787), .B2(n19670), .ZN(
        n15596) );
  OAI211_X1 U18697 ( .C1(n19793), .C2(n19673), .A(n15597), .B(n15596), .ZN(
        P1_U2994) );
  NOR2_X1 U18698 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15598), .ZN(
        n15604) );
  NOR2_X1 U18699 ( .A1(n19798), .A2(n14178), .ZN(n15602) );
  OAI22_X1 U18700 ( .A1(n15600), .A2(n19820), .B1(n15599), .B2(n19823), .ZN(
        n15601) );
  AOI211_X1 U18701 ( .C1(n15604), .C2(n15603), .A(n15602), .B(n15601), .ZN(
        n15605) );
  OAI21_X1 U18702 ( .B1(n15607), .B2(n15606), .A(n15605), .ZN(P1_U3013) );
  NOR2_X1 U18703 ( .A1(n15609), .A2(n15608), .ZN(n15613) );
  NOR2_X1 U18704 ( .A1(n19798), .A2(n15610), .ZN(n15611) );
  AOI221_X1 U18705 ( .B1(n15613), .B2(n15618), .C1(n15612), .C2(n15618), .A(
        n15611), .ZN(n15617) );
  AOI22_X1 U18706 ( .A1(n15615), .A2(n19810), .B1(n19807), .B2(n15614), .ZN(
        n15616) );
  OAI211_X1 U18707 ( .C1(n15619), .C2(n15618), .A(n15617), .B(n15616), .ZN(
        P1_U3018) );
  AOI22_X1 U18708 ( .A1(n19807), .A2(n15620), .B1(n19781), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n15628) );
  AOI22_X1 U18709 ( .A1(n15622), .A2(n19810), .B1(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n15621), .ZN(n15627) );
  NAND3_X1 U18710 ( .A1(n15625), .A2(n15624), .A3(n15623), .ZN(n15626) );
  NAND3_X1 U18711 ( .A1(n15628), .A2(n15627), .A3(n15626), .ZN(P1_U3020) );
  INV_X1 U18712 ( .A(n15674), .ZN(n15654) );
  NAND2_X1 U18713 ( .A1(n15636), .A2(n15654), .ZN(n15647) );
  AOI22_X1 U18714 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n11134), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15629), .ZN(n15640) );
  AOI21_X1 U18715 ( .B1(n19807), .B2(n15631), .A(n15630), .ZN(n15639) );
  INV_X1 U18716 ( .A(n15632), .ZN(n15648) );
  AOI21_X1 U18717 ( .B1(n19818), .B2(n15633), .A(n15648), .ZN(n15635) );
  AOI21_X1 U18718 ( .B1(n15636), .B2(n15635), .A(n15634), .ZN(n15643) );
  AOI22_X1 U18719 ( .A1(n15637), .A2(n19810), .B1(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n15643), .ZN(n15638) );
  OAI211_X1 U18720 ( .C1(n15647), .C2(n15640), .A(n15639), .B(n15638), .ZN(
        P1_U3021) );
  INV_X1 U18721 ( .A(n15641), .ZN(n15642) );
  AOI21_X1 U18722 ( .B1(n19807), .B2(n19626), .A(n15642), .ZN(n15646) );
  AOI22_X1 U18723 ( .A1(n15644), .A2(n19810), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15643), .ZN(n15645) );
  OAI211_X1 U18724 ( .C1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n15647), .A(
        n15646), .B(n15645), .ZN(P1_U3022) );
  NOR2_X1 U18725 ( .A1(n19801), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15675) );
  INV_X1 U18726 ( .A(n15675), .ZN(n15650) );
  AOI221_X1 U18727 ( .B1(n15649), .B2(n19818), .C1(n19801), .C2(n19818), .A(
        n15648), .ZN(n15680) );
  OAI21_X1 U18728 ( .B1(n15651), .B2(n15650), .A(n15680), .ZN(n15670) );
  AOI21_X1 U18729 ( .B1(n12308), .B2(n15652), .A(n15670), .ZN(n15664) );
  INV_X1 U18730 ( .A(n15653), .ZN(n15659) );
  NAND2_X1 U18731 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15654), .ZN(
        n15666) );
  AOI221_X1 U18732 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n13212), .C2(n15665), .A(
        n15666), .ZN(n15658) );
  OAI22_X1 U18733 ( .A1(n19823), .A2(n15656), .B1(n15655), .B2(n19798), .ZN(
        n15657) );
  AOI211_X1 U18734 ( .C1(n15659), .C2(n19810), .A(n15658), .B(n15657), .ZN(
        n15660) );
  OAI21_X1 U18735 ( .B1(n15664), .B2(n13212), .A(n15660), .ZN(P1_U3023) );
  INV_X1 U18736 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n19650) );
  OAI22_X1 U18737 ( .A1(n19823), .A2(n19639), .B1(n19650), .B2(n19798), .ZN(
        n15661) );
  AOI21_X1 U18738 ( .B1(n15662), .B2(n19810), .A(n15661), .ZN(n15663) );
  OAI221_X1 U18739 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n15666), .C1(
        n15665), .C2(n15664), .A(n15663), .ZN(P1_U3024) );
  INV_X1 U18740 ( .A(n15667), .ZN(n15668) );
  XNOR2_X1 U18741 ( .A(n15669), .B(n15668), .ZN(n19704) );
  AOI22_X1 U18742 ( .A1(n19807), .A2(n19704), .B1(n19781), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n15673) );
  AOI22_X1 U18743 ( .A1(n15671), .A2(n19810), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15670), .ZN(n15672) );
  OAI211_X1 U18744 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n15674), .A(
        n15673), .B(n15672), .ZN(P1_U3025) );
  AOI22_X1 U18745 ( .A1(n19807), .A2(n19663), .B1(n19781), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n15678) );
  AOI22_X1 U18746 ( .A1(n15676), .A2(n19810), .B1(n19809), .B2(n15675), .ZN(
        n15677) );
  OAI211_X1 U18747 ( .C1(n15680), .C2(n15679), .A(n15678), .B(n15677), .ZN(
        P1_U3026) );
  NOR3_X1 U18748 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20446), .A3(n20445), 
        .ZN(n15681) );
  AOI22_X1 U18749 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n20547), .B1(n15681), 
        .B2(n20546), .ZN(n20447) );
  AOI21_X1 U18750 ( .B1(n20447), .B2(n15683), .A(n15682), .ZN(n15686) );
  AOI21_X1 U18751 ( .B1(n20270), .B2(n20546), .A(n15684), .ZN(n15685) );
  AOI211_X1 U18752 ( .C1(n20445), .C2(n15687), .A(n15686), .B(n15685), .ZN(
        P1_U3162) );
  OAI21_X1 U18753 ( .B1(n15689), .B2(n20270), .A(n15688), .ZN(P1_U3466) );
  OAI22_X1 U18754 ( .A1(n15691), .A2(n15690), .B1(n14828), .B2(n18601), .ZN(
        n15695) );
  INV_X1 U18755 ( .A(n15692), .ZN(n15693) );
  OAI22_X1 U18756 ( .A1(n15693), .A2(n18616), .B1(n18540), .B2(n11965), .ZN(
        n15694) );
  AOI211_X1 U18757 ( .C1(n18647), .C2(n18650), .A(n15695), .B(n15694), .ZN(
        n15699) );
  NAND4_X1 U18758 ( .A1(n18623), .A2(n15704), .A3(n15697), .A4(n15696), .ZN(
        n15698) );
  OAI211_X1 U18759 ( .C1(n15700), .C2(n18643), .A(n15699), .B(n15698), .ZN(
        P2_U2824) );
  AOI22_X1 U18760 ( .A1(P2_REIP_REG_29__SCAN_IN), .A2(n9772), .B1(n15701), 
        .B2(n18637), .ZN(n15710) );
  AOI22_X1 U18761 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18639), .B1(
        P2_EBX_REG_29__SCAN_IN), .B2(n18614), .ZN(n15709) );
  AOI22_X1 U18762 ( .A1(n15703), .A2(n18625), .B1(n15702), .B2(n18647), .ZN(
        n15708) );
  AOI21_X1 U18763 ( .B1(n15705), .B2(n9721), .A(n15704), .ZN(n15706) );
  NAND2_X1 U18764 ( .A1(n18623), .A2(n15706), .ZN(n15707) );
  NAND4_X1 U18765 ( .A1(n15710), .A2(n15709), .A3(n15708), .A4(n15707), .ZN(
        P2_U2826) );
  AOI22_X1 U18766 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18639), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n9772), .ZN(n15711) );
  OAI21_X1 U18767 ( .B1(n15712), .B2(n18616), .A(n15711), .ZN(n15713) );
  AOI21_X1 U18768 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n18614), .A(n15713), .ZN(
        n15720) );
  AOI21_X1 U18769 ( .B1(n15716), .B2(n15715), .A(n15714), .ZN(n15717) );
  AOI22_X1 U18770 ( .A1(n15718), .A2(n18647), .B1(n18623), .B2(n15717), .ZN(
        n15719) );
  OAI211_X1 U18771 ( .C1(n15721), .C2(n18643), .A(n15720), .B(n15719), .ZN(
        P2_U2827) );
  INV_X1 U18772 ( .A(n15722), .ZN(n15724) );
  AOI22_X1 U18773 ( .A1(n15724), .A2(n18625), .B1(n15723), .B2(n18647), .ZN(
        n15733) );
  AOI211_X1 U18774 ( .C1(n15727), .C2(n15726), .A(n15725), .B(n19437), .ZN(
        n15731) );
  AOI22_X1 U18775 ( .A1(P2_EBX_REG_27__SCAN_IN), .A2(n18614), .B1(
        P2_REIP_REG_27__SCAN_IN), .B2(n9772), .ZN(n15728) );
  OAI21_X1 U18776 ( .B1(n15729), .B2(n18616), .A(n15728), .ZN(n15730) );
  AOI211_X1 U18777 ( .C1(n18639), .C2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15731), .B(n15730), .ZN(n15732) );
  NAND2_X1 U18778 ( .A1(n15733), .A2(n15732), .ZN(P2_U2828) );
  AOI211_X1 U18779 ( .C1(n15736), .C2(n15735), .A(n15734), .B(n19437), .ZN(
        n15742) );
  AOI22_X1 U18780 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n18639), .B1(
        n15737), .B2(n18637), .ZN(n15739) );
  AOI22_X1 U18781 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n18614), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n9772), .ZN(n15738) );
  OAI211_X1 U18782 ( .C1(n15740), .C2(n18643), .A(n15739), .B(n15738), .ZN(
        n15741) );
  AOI211_X1 U18783 ( .C1(n18647), .C2(n15743), .A(n15742), .B(n15741), .ZN(
        n15744) );
  INV_X1 U18784 ( .A(n15744), .ZN(P2_U2829) );
  AOI22_X1 U18785 ( .A1(n15745), .A2(n18637), .B1(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n18639), .ZN(n15754) );
  AOI22_X1 U18786 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(n18614), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n9772), .ZN(n15753) );
  AOI22_X1 U18787 ( .A1(n15747), .A2(n18625), .B1(n15746), .B2(n18647), .ZN(
        n15752) );
  AOI21_X1 U18788 ( .B1(n15749), .B2(n10128), .A(n15748), .ZN(n15750) );
  NAND2_X1 U18789 ( .A1(n18623), .A2(n15750), .ZN(n15751) );
  NAND4_X1 U18790 ( .A1(n15754), .A2(n15753), .A3(n15752), .A4(n15751), .ZN(
        P2_U2830) );
  AOI22_X1 U18791 ( .A1(n15755), .A2(n18637), .B1(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n18639), .ZN(n15765) );
  AOI22_X1 U18792 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(n18614), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n9772), .ZN(n15764) );
  INV_X1 U18793 ( .A(n15756), .ZN(n15779) );
  AOI22_X1 U18794 ( .A1(n15757), .A2(n18625), .B1(n15779), .B2(n18647), .ZN(
        n15763) );
  AOI21_X1 U18795 ( .B1(n15760), .B2(n15759), .A(n15758), .ZN(n15761) );
  NAND2_X1 U18796 ( .A1(n18623), .A2(n15761), .ZN(n15762) );
  NAND4_X1 U18797 ( .A1(n15765), .A2(n15764), .A3(n15763), .A4(n15762), .ZN(
        P2_U2831) );
  AOI211_X1 U18798 ( .C1(n15768), .C2(n15767), .A(n15766), .B(n19437), .ZN(
        n15772) );
  AOI22_X1 U18799 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n18639), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n9772), .ZN(n15769) );
  OAI21_X1 U18800 ( .B1(n15770), .B2(n18616), .A(n15769), .ZN(n15771) );
  AOI211_X1 U18801 ( .C1(P2_EBX_REG_23__SCAN_IN), .C2(n18614), .A(n15772), .B(
        n15771), .ZN(n15777) );
  INV_X1 U18802 ( .A(n15773), .ZN(n15774) );
  AOI22_X1 U18803 ( .A1(n15775), .A2(n18625), .B1(n15774), .B2(n18647), .ZN(
        n15776) );
  NAND2_X1 U18804 ( .A1(n15777), .A2(n15776), .ZN(P2_U2832) );
  AOI22_X1 U18805 ( .A1(n15778), .A2(n18663), .B1(P2_EAX_REG_24__SCAN_IN), 
        .B2(n18691), .ZN(n15783) );
  AOI22_X1 U18806 ( .A1(n18651), .A2(BUF2_REG_24__SCAN_IN), .B1(n18652), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n15782) );
  AOI22_X1 U18807 ( .A1(n15780), .A2(n18694), .B1(n18692), .B2(n15779), .ZN(
        n15781) );
  NAND3_X1 U18808 ( .A1(n15783), .A2(n15782), .A3(n15781), .ZN(P2_U2895) );
  AOI22_X1 U18809 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n18850), .B1(n18829), 
        .B2(n15784), .ZN(n15789) );
  AOI222_X1 U18810 ( .A1(n15787), .A2(n18808), .B1(n18830), .B2(n15786), .C1(
        n18821), .C2(n15785), .ZN(n15788) );
  OAI211_X1 U18811 ( .C1(n15852), .C2(n10113), .A(n15789), .B(n15788), .ZN(
        P2_U2992) );
  AOI22_X1 U18812 ( .A1(n18820), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n18850), .ZN(n15798) );
  INV_X1 U18813 ( .A(n15790), .ZN(n15792) );
  AOI21_X1 U18814 ( .B1(n15792), .B2(n15861), .A(n15791), .ZN(n15860) );
  NAND2_X1 U18815 ( .A1(n15794), .A2(n15793), .ZN(n15795) );
  XNOR2_X1 U18816 ( .A(n15796), .B(n15795), .ZN(n15859) );
  AOI222_X1 U18817 ( .A1(n15860), .A2(n18821), .B1(n18808), .B2(n15859), .C1(
        n18830), .C2(n15858), .ZN(n15797) );
  OAI211_X1 U18818 ( .C1(n18816), .C2(n18511), .A(n15798), .B(n15797), .ZN(
        P2_U3000) );
  AOI22_X1 U18819 ( .A1(n18820), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n18850), .ZN(n15808) );
  OR2_X1 U18820 ( .A1(n15799), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15801) );
  NAND2_X1 U18821 ( .A1(n15801), .A2(n15800), .ZN(n15879) );
  INV_X1 U18822 ( .A(n15879), .ZN(n15806) );
  OR2_X1 U18823 ( .A1(n9737), .A2(n15802), .ZN(n15803) );
  XNOR2_X1 U18824 ( .A(n15804), .B(n15803), .ZN(n15876) );
  AOI222_X1 U18825 ( .A1(n15806), .A2(n18821), .B1(n18808), .B2(n15876), .C1(
        n18830), .C2(n15805), .ZN(n15807) );
  OAI211_X1 U18826 ( .C1(n18816), .C2(n18535), .A(n15808), .B(n15807), .ZN(
        P2_U3002) );
  AOI22_X1 U18827 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n18850), .B1(n18829), 
        .B2(n18548), .ZN(n15813) );
  OAI22_X1 U18828 ( .A1(n15810), .A2(n15838), .B1(n15809), .B2(n18833), .ZN(
        n15811) );
  AOI21_X1 U18829 ( .B1(n18830), .B2(n18545), .A(n15811), .ZN(n15812) );
  OAI211_X1 U18830 ( .C1(n15852), .C2(n18541), .A(n15813), .B(n15812), .ZN(
        P2_U3003) );
  AOI22_X1 U18831 ( .A1(n18820), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n18850), .ZN(n15818) );
  INV_X1 U18832 ( .A(n15814), .ZN(n15816) );
  AOI222_X1 U18833 ( .A1(n15816), .A2(n18808), .B1(n18830), .B2(n18562), .C1(
        n18821), .C2(n15815), .ZN(n15817) );
  OAI211_X1 U18834 ( .C1(n18816), .C2(n18559), .A(n15818), .B(n15817), .ZN(
        P2_U3004) );
  AOI22_X1 U18835 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n18850), .B1(n18829), 
        .B2(n18571), .ZN(n15823) );
  OAI22_X1 U18836 ( .A1(n15820), .A2(n15838), .B1(n18833), .B2(n15819), .ZN(
        n15821) );
  AOI21_X1 U18837 ( .B1(n18830), .B2(n18573), .A(n15821), .ZN(n15822) );
  OAI211_X1 U18838 ( .C1(n15852), .C2(n15824), .A(n15823), .B(n15822), .ZN(
        P2_U3005) );
  AOI22_X1 U18839 ( .A1(n18820), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n18850), .ZN(n15836) );
  AOI21_X1 U18840 ( .B1(n15827), .B2(n15826), .A(n15825), .ZN(n15832) );
  INV_X1 U18841 ( .A(n15828), .ZN(n15830) );
  NOR2_X1 U18842 ( .A1(n15830), .A2(n15829), .ZN(n15831) );
  XNOR2_X1 U18843 ( .A(n15832), .B(n15831), .ZN(n15891) );
  XOR2_X1 U18844 ( .A(n15834), .B(n15833), .Z(n15889) );
  AOI222_X1 U18845 ( .A1(n15891), .A2(n18808), .B1(n18830), .B2(n15890), .C1(
        n15889), .C2(n18821), .ZN(n15835) );
  OAI211_X1 U18846 ( .C1(n18816), .C2(n18582), .A(n15836), .B(n15835), .ZN(
        P2_U3006) );
  AOI22_X1 U18847 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n18850), .B1(n18829), 
        .B2(n18621), .ZN(n15842) );
  OAI22_X1 U18848 ( .A1(n15839), .A2(n15838), .B1(n15837), .B2(n18833), .ZN(
        n15840) );
  AOI21_X1 U18849 ( .B1(n18830), .B2(n18624), .A(n15840), .ZN(n15841) );
  OAI211_X1 U18850 ( .C1(n15852), .C2(n15843), .A(n15842), .B(n15841), .ZN(
        P2_U3009) );
  AOI22_X1 U18851 ( .A1(P2_REIP_REG_3__SCAN_IN), .A2(n18850), .B1(n18829), 
        .B2(n15844), .ZN(n15851) );
  XNOR2_X1 U18852 ( .A(n15845), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n15846) );
  XNOR2_X1 U18853 ( .A(n15847), .B(n15846), .ZN(n15900) );
  AOI222_X1 U18854 ( .A1(n18808), .A2(n15900), .B1(n9724), .B2(n18821), .C1(
        n15895), .C2(n18830), .ZN(n15850) );
  OAI211_X1 U18855 ( .C1(n15853), .C2(n15852), .A(n15851), .B(n15850), .ZN(
        P2_U3011) );
  AOI21_X1 U18856 ( .B1(n15856), .B2(n15855), .A(n15854), .ZN(n18655) );
  AOI22_X1 U18857 ( .A1(n15857), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n18875), .B2(n18655), .ZN(n15867) );
  AOI222_X1 U18858 ( .A1(n15860), .A2(n18849), .B1(n18846), .B2(n15859), .C1(
        n18868), .C2(n15858), .ZN(n15866) );
  NAND2_X1 U18859 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n18850), .ZN(n15865) );
  NAND3_X1 U18860 ( .A1(n15863), .A2(n15862), .A3(n15861), .ZN(n15864) );
  NAND4_X1 U18861 ( .A1(n15867), .A2(n15866), .A3(n15865), .A4(n15864), .ZN(
        P2_U3032) );
  AOI21_X1 U18862 ( .B1(n15870), .B2(n15869), .A(n15868), .ZN(n18659) );
  NAND2_X1 U18863 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n18850), .ZN(n15871) );
  OAI221_X1 U18864 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n15873), 
        .C1(n13774), .C2(n15872), .A(n15871), .ZN(n15874) );
  AOI21_X1 U18865 ( .B1(n18875), .B2(n18659), .A(n15874), .ZN(n15878) );
  NOR2_X1 U18866 ( .A1(n18839), .A2(n18538), .ZN(n15875) );
  AOI21_X1 U18867 ( .B1(n15876), .B2(n18846), .A(n15875), .ZN(n15877) );
  OAI211_X1 U18868 ( .C1(n18861), .C2(n15879), .A(n15878), .B(n15877), .ZN(
        P2_U3034) );
  INV_X1 U18869 ( .A(n15880), .ZN(n15882) );
  AOI211_X1 U18870 ( .C1(n13752), .C2(n15883), .A(n15882), .B(n15881), .ZN(
        n15888) );
  AOI21_X1 U18871 ( .B1(n15886), .B2(n15885), .A(n15884), .ZN(n18585) );
  INV_X1 U18872 ( .A(n18585), .ZN(n18665) );
  OAI22_X1 U18873 ( .A1(n15898), .A2(n18665), .B1(n12016), .B2(n18496), .ZN(
        n15887) );
  NOR2_X1 U18874 ( .A1(n15888), .A2(n15887), .ZN(n15893) );
  AOI222_X1 U18875 ( .A1(n15891), .A2(n18846), .B1(n18868), .B2(n15890), .C1(
        n15889), .C2(n18849), .ZN(n15892) );
  OAI211_X1 U18876 ( .C1(n15894), .C2(n13752), .A(n15893), .B(n15892), .ZN(
        P2_U3038) );
  NAND2_X1 U18877 ( .A1(n9724), .A2(n18849), .ZN(n15897) );
  AOI22_X1 U18878 ( .A1(n18868), .A2(n15895), .B1(P2_REIP_REG_3__SCAN_IN), 
        .B2(n13482), .ZN(n15896) );
  OAI211_X1 U18879 ( .C1(n19534), .C2(n15898), .A(n15897), .B(n15896), .ZN(
        n15899) );
  AOI21_X1 U18880 ( .B1(n18846), .B2(n15900), .A(n15899), .ZN(n15901) );
  OAI221_X1 U18881 ( .B1(n18841), .B2(n15903), .C1(n18841), .C2(n15902), .A(
        n15901), .ZN(P2_U3043) );
  INV_X1 U18882 ( .A(n15910), .ZN(n19434) );
  NOR2_X1 U18883 ( .A1(n19434), .A2(n19593), .ZN(n19436) );
  OAI21_X1 U18884 ( .B1(n15905), .B2(n19525), .A(n15904), .ZN(n15913) );
  INV_X1 U18885 ( .A(n15906), .ZN(n15908) );
  AOI211_X1 U18886 ( .C1(n19574), .C2(n15908), .A(n19435), .B(n15907), .ZN(
        n15912) );
  AOI22_X1 U18887 ( .A1(n15910), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n18699), 
        .B2(n15909), .ZN(n15911) );
  OAI211_X1 U18888 ( .C1(n19436), .C2(n15913), .A(n15912), .B(n15911), .ZN(
        P2_U3176) );
  INV_X1 U18889 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18349) );
  NAND3_X1 U18890 ( .A1(n18349), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15925) );
  INV_X1 U18891 ( .A(n15925), .ZN(n15961) );
  AOI21_X1 U18892 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15914), .A(
        n18349), .ZN(n15915) );
  AOI21_X1 U18893 ( .B1(n15974), .B2(n15961), .A(n15915), .ZN(n15963) );
  INV_X1 U18894 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16133) );
  NAND2_X1 U18895 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17314) );
  INV_X1 U18896 ( .A(n17314), .ZN(n17297) );
  NAND3_X1 U18897 ( .A1(n17297), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17226) );
  NOR2_X2 U18898 ( .A1(n16128), .A2(n15918), .ZN(n17186) );
  NAND3_X1 U18899 ( .A1(n10281), .A2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17153) );
  INV_X1 U18900 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17085) );
  INV_X1 U18901 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17098) );
  NOR2_X1 U18902 ( .A1(n17098), .A2(n17086), .ZN(n17083) );
  INV_X1 U18903 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16167) );
  NAND2_X1 U18904 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n15944), .ZN(
        n15920) );
  INV_X1 U18905 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18325) );
  NOR2_X1 U18906 ( .A1(n18325), .A2(n9746), .ZN(n15957) );
  NAND3_X1 U18907 ( .A1(n9766), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15949) );
  NOR2_X1 U18908 ( .A1(n16167), .A2(n15949), .ZN(n15921) );
  NAND2_X1 U18909 ( .A1(n18394), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18255) );
  OAI21_X2 U18910 ( .B1(n17402), .B2(n17070), .A(n18090), .ZN(n17261) );
  NAND2_X1 U18911 ( .A1(n15921), .A2(n17261), .ZN(n15935) );
  XNOR2_X1 U18912 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15922) );
  NOR2_X1 U18913 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17070), .ZN(
        n15946) );
  INV_X1 U18914 ( .A(n15945), .ZN(n16115) );
  OR2_X1 U18915 ( .A1(n18090), .A2(n15921), .ZN(n15950) );
  OAI211_X1 U18916 ( .C1(n16115), .C2(n18255), .A(n17408), .B(n15950), .ZN(
        n15955) );
  NOR2_X1 U18917 ( .A1(n15946), .A2(n15955), .ZN(n15934) );
  OAI22_X1 U18918 ( .A1(n15935), .A2(n15922), .B1(n15934), .B2(n16133), .ZN(
        n15923) );
  AOI211_X1 U18919 ( .C1(n17258), .C2(n10073), .A(n15957), .B(n15923), .ZN(
        n15930) );
  OAI21_X1 U18920 ( .B1(n15938), .B2(n15931), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15924) );
  OAI21_X1 U18921 ( .B1(n15925), .B2(n15976), .A(n15924), .ZN(n15959) );
  AOI22_X1 U18922 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17235), .B1(
        n17318), .B2(n18349), .ZN(n15928) );
  NOR2_X1 U18923 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18349), .ZN(
        n15958) );
  OAI211_X1 U18924 ( .C1(n15963), .C2(n17412), .A(n15930), .B(n15929), .ZN(
        P3_U2799) );
  INV_X1 U18925 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16156) );
  XNOR2_X1 U18926 ( .A(n16156), .B(n15944), .ZN(n16152) );
  NAND2_X1 U18927 ( .A1(n17309), .A2(n15931), .ZN(n15956) );
  NAND2_X1 U18928 ( .A1(n17401), .A2(n15932), .ZN(n15952) );
  AOI21_X1 U18929 ( .B1(n15956), .B2(n15952), .A(n15938), .ZN(n15937) );
  NAND2_X1 U18930 ( .A1(n17715), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n15933) );
  OAI221_X1 U18931 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n15935), .C1(
        n16156), .C2(n15934), .A(n15933), .ZN(n15936) );
  AOI211_X1 U18932 ( .C1(n17258), .C2(n16152), .A(n15937), .B(n15936), .ZN(
        n15942) );
  AOI22_X1 U18933 ( .A1(n17232), .A2(n17401), .B1(n17309), .B2(n17574), .ZN(
        n17303) );
  NOR2_X1 U18934 ( .A1(n17507), .A2(n17303), .ZN(n17195) );
  NAND2_X1 U18935 ( .A1(n15971), .A2(n17195), .ZN(n17108) );
  INV_X1 U18936 ( .A(n17108), .ZN(n17119) );
  NAND4_X1 U18937 ( .A1(n15940), .A2(n15939), .A3(n17119), .A4(n15938), .ZN(
        n15941) );
  OAI211_X1 U18938 ( .C1(n15943), .C2(n17322), .A(n15942), .B(n15941), .ZN(
        P3_U2800) );
  AOI21_X1 U18939 ( .B1(n16167), .B2(n15945), .A(n15944), .ZN(n16161) );
  OAI21_X1 U18940 ( .B1(n15946), .B2(n17258), .A(n16161), .ZN(n15947) );
  OAI211_X1 U18941 ( .C1(n15950), .C2(n15949), .A(n15948), .B(n15947), .ZN(
        n15954) );
  NOR2_X1 U18942 ( .A1(n15974), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15953) );
  AOI21_X1 U18943 ( .B1(n15958), .B2(n17631), .A(n15957), .ZN(n15967) );
  AOI22_X1 U18944 ( .A1(n15961), .A2(n15960), .B1(n17472), .B2(n15959), .ZN(
        n15962) );
  OAI22_X1 U18945 ( .A1(n15963), .A2(n17703), .B1(n15962), .B2(n17680), .ZN(
        n15964) );
  OAI211_X1 U18946 ( .C1(n18349), .C2(n15968), .A(n15967), .B(n15966), .ZN(
        P3_U2831) );
  AOI21_X1 U18947 ( .B1(n17318), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15969), .ZN(n17055) );
  NAND2_X1 U18948 ( .A1(n17061), .A2(n17613), .ZN(n15988) );
  AOI22_X1 U18949 ( .A1(n18217), .A2(n17232), .B1(n17574), .B2(n17472), .ZN(
        n17588) );
  OAI21_X1 U18950 ( .B1(n17588), .B2(n17507), .A(n15970), .ZN(n17466) );
  NAND2_X1 U18951 ( .A1(n15971), .A2(n17466), .ZN(n17458) );
  NOR2_X1 U18952 ( .A1(n17680), .A2(n17458), .ZN(n17444) );
  NOR2_X1 U18953 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n15972), .ZN(
        n17052) );
  OAI211_X1 U18954 ( .C1(n15974), .C2(n17468), .A(n15973), .B(n17705), .ZN(
        n15975) );
  AOI21_X1 U18955 ( .B1(n17472), .B2(n15976), .A(n15975), .ZN(n15982) );
  OAI21_X1 U18956 ( .B1(n17060), .B2(n17235), .A(n15977), .ZN(n17054) );
  NAND2_X1 U18957 ( .A1(n17055), .A2(n17054), .ZN(n17053) );
  NAND2_X1 U18958 ( .A1(n15985), .A2(n17060), .ZN(n15978) );
  NAND4_X1 U18959 ( .A1(n15980), .A2(n17053), .A3(n15979), .A4(n15978), .ZN(
        n15981) );
  AOI211_X1 U18960 ( .C1(n15982), .C2(n15981), .A(n17710), .B(n15984), .ZN(
        n15983) );
  INV_X1 U18961 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18322) );
  NOR2_X1 U18962 ( .A1(n9746), .A2(n18322), .ZN(n17051) );
  AOI211_X1 U18963 ( .C1(n17444), .C2(n17052), .A(n15983), .B(n17051), .ZN(
        n15987) );
  NAND4_X1 U18964 ( .A1(n15985), .A2(n17060), .A3(n17613), .A4(n15984), .ZN(
        n15986) );
  OAI211_X1 U18965 ( .C1(n17055), .C2(n15988), .A(n15987), .B(n15986), .ZN(
        P3_U2834) );
  NOR3_X1 U18966 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n15990) );
  NOR4_X1 U18967 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n15989) );
  NAND4_X1 U18968 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n15990), .A3(n15989), .A4(
        U215), .ZN(U213) );
  INV_X1 U18969 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n16081) );
  INV_X2 U18970 ( .A(U214), .ZN(n16045) );
  INV_X1 U18971 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16082) );
  OAI222_X1 U18972 ( .A1(U212), .A2(n16081), .B1(n16047), .B2(n15992), .C1(
        U214), .C2(n16082), .ZN(U216) );
  INV_X1 U18973 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n15994) );
  AOI22_X1 U18974 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16045), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16032), .ZN(n15993) );
  OAI21_X1 U18975 ( .B1(n15994), .B2(n16047), .A(n15993), .ZN(U217) );
  INV_X1 U18976 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20672) );
  AOI22_X1 U18977 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16045), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16032), .ZN(n15995) );
  OAI21_X1 U18978 ( .B1(n20672), .B2(n16047), .A(n15995), .ZN(U218) );
  INV_X1 U18979 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n15997) );
  AOI22_X1 U18980 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16045), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16032), .ZN(n15996) );
  OAI21_X1 U18981 ( .B1(n15997), .B2(n16047), .A(n15996), .ZN(U219) );
  AOI22_X1 U18982 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16045), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16032), .ZN(n15998) );
  OAI21_X1 U18983 ( .B1(n15999), .B2(n16047), .A(n15998), .ZN(U220) );
  INV_X1 U18984 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16001) );
  AOI22_X1 U18985 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16045), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16032), .ZN(n16000) );
  OAI21_X1 U18986 ( .B1(n16001), .B2(n16047), .A(n16000), .ZN(U221) );
  INV_X1 U18987 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16003) );
  AOI22_X1 U18988 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16045), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16032), .ZN(n16002) );
  OAI21_X1 U18989 ( .B1(n16003), .B2(n16047), .A(n16002), .ZN(U222) );
  AOI22_X1 U18990 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16045), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16032), .ZN(n16004) );
  OAI21_X1 U18991 ( .B1(n14042), .B2(n16047), .A(n16004), .ZN(U223) );
  INV_X1 U18992 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16006) );
  AOI22_X1 U18993 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16045), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16032), .ZN(n16005) );
  OAI21_X1 U18994 ( .B1(n16006), .B2(n16047), .A(n16005), .ZN(U224) );
  INV_X1 U18995 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n18918) );
  AOI22_X1 U18996 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16045), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16032), .ZN(n16007) );
  OAI21_X1 U18997 ( .B1(n18918), .B2(n16047), .A(n16007), .ZN(U225) );
  AOI22_X1 U18998 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16045), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16032), .ZN(n16008) );
  OAI21_X1 U18999 ( .B1(n16009), .B2(n16047), .A(n16008), .ZN(U226) );
  INV_X1 U19000 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16011) );
  AOI22_X1 U19001 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16045), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16032), .ZN(n16010) );
  OAI21_X1 U19002 ( .B1(n16011), .B2(n16047), .A(n16010), .ZN(U227) );
  AOI22_X1 U19003 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16045), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16032), .ZN(n16012) );
  OAI21_X1 U19004 ( .B1(n16013), .B2(n16047), .A(n16012), .ZN(U228) );
  AOI22_X1 U19005 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16045), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16032), .ZN(n16014) );
  OAI21_X1 U19006 ( .B1(n18899), .B2(n16047), .A(n16014), .ZN(U229) );
  INV_X1 U19007 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n18894) );
  AOI22_X1 U19008 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16045), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16032), .ZN(n16015) );
  OAI21_X1 U19009 ( .B1(n18894), .B2(n16047), .A(n16015), .ZN(U230) );
  INV_X1 U19010 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16017) );
  AOI22_X1 U19011 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16045), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16032), .ZN(n16016) );
  OAI21_X1 U19012 ( .B1(n16017), .B2(n16047), .A(n16016), .ZN(U231) );
  AOI22_X1 U19013 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16045), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16032), .ZN(n16018) );
  OAI21_X1 U19014 ( .B1(n12643), .B2(n16047), .A(n16018), .ZN(U232) );
  AOI22_X1 U19015 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16045), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16032), .ZN(n16019) );
  OAI21_X1 U19016 ( .B1(n12402), .B2(n16047), .A(n16019), .ZN(U233) );
  INV_X1 U19017 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16021) );
  AOI22_X1 U19018 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16045), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16032), .ZN(n16020) );
  OAI21_X1 U19019 ( .B1(n16021), .B2(n16047), .A(n16020), .ZN(U234) );
  AOI22_X1 U19020 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16045), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16032), .ZN(n16022) );
  OAI21_X1 U19021 ( .B1(n16023), .B2(n16047), .A(n16022), .ZN(U235) );
  INV_X1 U19022 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n16025) );
  AOI22_X1 U19023 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16045), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16032), .ZN(n16024) );
  OAI21_X1 U19024 ( .B1(n16025), .B2(n16047), .A(n16024), .ZN(U236) );
  INV_X1 U19025 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16027) );
  AOI22_X1 U19026 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16045), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16032), .ZN(n16026) );
  OAI21_X1 U19027 ( .B1(n16027), .B2(n16047), .A(n16026), .ZN(U237) );
  INV_X1 U19028 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16029) );
  AOI22_X1 U19029 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16045), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16032), .ZN(n16028) );
  OAI21_X1 U19030 ( .B1(n16029), .B2(n16047), .A(n16028), .ZN(U238) );
  AOI22_X1 U19031 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16045), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16032), .ZN(n16030) );
  OAI21_X1 U19032 ( .B1(n20584), .B2(n16047), .A(n16030), .ZN(U239) );
  INV_X1 U19033 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n20640) );
  AOI22_X1 U19034 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16045), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16032), .ZN(n16031) );
  OAI21_X1 U19035 ( .B1(n20640), .B2(n16047), .A(n16031), .ZN(U240) );
  INV_X1 U19036 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16034) );
  AOI22_X1 U19037 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16045), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16032), .ZN(n16033) );
  OAI21_X1 U19038 ( .B1(n16034), .B2(n16047), .A(n16033), .ZN(U241) );
  AOI22_X1 U19039 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16045), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16032), .ZN(n16035) );
  OAI21_X1 U19040 ( .B1(n16036), .B2(n16047), .A(n16035), .ZN(U242) );
  INV_X1 U19041 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16038) );
  AOI22_X1 U19042 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16045), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16032), .ZN(n16037) );
  OAI21_X1 U19043 ( .B1(n16038), .B2(n16047), .A(n16037), .ZN(U243) );
  INV_X1 U19044 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16040) );
  AOI22_X1 U19045 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16045), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16032), .ZN(n16039) );
  OAI21_X1 U19046 ( .B1(n16040), .B2(n16047), .A(n16039), .ZN(U244) );
  INV_X1 U19047 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16042) );
  AOI22_X1 U19048 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16045), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16032), .ZN(n16041) );
  OAI21_X1 U19049 ( .B1(n16042), .B2(n16047), .A(n16041), .ZN(U245) );
  INV_X1 U19050 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16044) );
  AOI22_X1 U19051 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16045), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16032), .ZN(n16043) );
  OAI21_X1 U19052 ( .B1(n16044), .B2(n16047), .A(n16043), .ZN(U246) );
  INV_X1 U19053 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16048) );
  AOI22_X1 U19054 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16045), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16032), .ZN(n16046) );
  OAI21_X1 U19055 ( .B1(n16048), .B2(n16047), .A(n16046), .ZN(U247) );
  OAI22_X1 U19056 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16079), .ZN(n16049) );
  INV_X1 U19057 ( .A(n16049), .ZN(U251) );
  OAI22_X1 U19058 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16079), .ZN(n16050) );
  INV_X1 U19059 ( .A(n16050), .ZN(U252) );
  OAI22_X1 U19060 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16079), .ZN(n16051) );
  INV_X1 U19061 ( .A(n16051), .ZN(U253) );
  OAI22_X1 U19062 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16079), .ZN(n16052) );
  INV_X1 U19063 ( .A(n16052), .ZN(U254) );
  OAI22_X1 U19064 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16079), .ZN(n16053) );
  INV_X1 U19065 ( .A(n16053), .ZN(U255) );
  OAI22_X1 U19066 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16079), .ZN(n16054) );
  INV_X1 U19067 ( .A(n16054), .ZN(U256) );
  OAI22_X1 U19068 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16079), .ZN(n16055) );
  INV_X1 U19069 ( .A(n16055), .ZN(U257) );
  INV_X1 U19070 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n20574) );
  INV_X1 U19071 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n17776) );
  AOI22_X1 U19072 ( .A1(n16079), .A2(n20574), .B1(n17776), .B2(U215), .ZN(U258) );
  OAI22_X1 U19073 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16079), .ZN(n16056) );
  INV_X1 U19074 ( .A(n16056), .ZN(U259) );
  OAI22_X1 U19075 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n16079), .ZN(n16057) );
  INV_X1 U19076 ( .A(n16057), .ZN(U260) );
  OAI22_X1 U19077 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16072), .ZN(n16058) );
  INV_X1 U19078 ( .A(n16058), .ZN(U261) );
  OAI22_X1 U19079 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16072), .ZN(n16059) );
  INV_X1 U19080 ( .A(n16059), .ZN(U262) );
  OAI22_X1 U19081 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16079), .ZN(n16060) );
  INV_X1 U19082 ( .A(n16060), .ZN(U263) );
  OAI22_X1 U19083 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16072), .ZN(n16061) );
  INV_X1 U19084 ( .A(n16061), .ZN(U264) );
  OAI22_X1 U19085 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16079), .ZN(n16062) );
  INV_X1 U19086 ( .A(n16062), .ZN(U265) );
  OAI22_X1 U19087 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16079), .ZN(n16063) );
  INV_X1 U19088 ( .A(n16063), .ZN(U266) );
  OAI22_X1 U19089 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16072), .ZN(n16064) );
  INV_X1 U19090 ( .A(n16064), .ZN(U267) );
  INV_X1 U19091 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n20655) );
  INV_X1 U19092 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n18893) );
  AOI22_X1 U19093 ( .A1(n16079), .A2(n20655), .B1(n18893), .B2(U215), .ZN(U268) );
  OAI22_X1 U19094 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16072), .ZN(n16065) );
  INV_X1 U19095 ( .A(n16065), .ZN(U269) );
  OAI22_X1 U19096 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16072), .ZN(n16066) );
  INV_X1 U19097 ( .A(n16066), .ZN(U270) );
  OAI22_X1 U19098 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16072), .ZN(n16067) );
  INV_X1 U19099 ( .A(n16067), .ZN(U271) );
  OAI22_X1 U19100 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16072), .ZN(n16068) );
  INV_X1 U19101 ( .A(n16068), .ZN(U272) );
  OAI22_X1 U19102 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16079), .ZN(n16069) );
  INV_X1 U19103 ( .A(n16069), .ZN(U273) );
  OAI22_X1 U19104 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16072), .ZN(n16070) );
  INV_X1 U19105 ( .A(n16070), .ZN(U274) );
  OAI22_X1 U19106 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16079), .ZN(n16071) );
  INV_X1 U19107 ( .A(n16071), .ZN(U275) );
  OAI22_X1 U19108 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16072), .ZN(n16073) );
  INV_X1 U19109 ( .A(n16073), .ZN(U276) );
  OAI22_X1 U19110 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16079), .ZN(n16074) );
  INV_X1 U19111 ( .A(n16074), .ZN(U277) );
  OAI22_X1 U19112 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16079), .ZN(n16075) );
  INV_X1 U19113 ( .A(n16075), .ZN(U278) );
  OAI22_X1 U19114 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16079), .ZN(n16076) );
  INV_X1 U19115 ( .A(n16076), .ZN(U279) );
  OAI22_X1 U19116 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16079), .ZN(n16077) );
  INV_X1 U19117 ( .A(n16077), .ZN(U280) );
  OAI22_X1 U19118 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16079), .ZN(n16078) );
  INV_X1 U19119 ( .A(n16078), .ZN(U281) );
  INV_X1 U19120 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n17780) );
  AOI22_X1 U19121 ( .A1(n16079), .A2(n16081), .B1(n17780), .B2(U215), .ZN(U282) );
  INV_X1 U19122 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16080) );
  AOI222_X1 U19123 ( .A1(n16082), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16081), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n16080), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16083) );
  INV_X2 U19124 ( .A(n16085), .ZN(n16084) );
  INV_X1 U19125 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18289) );
  INV_X1 U19126 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19474) );
  AOI22_X1 U19127 ( .A1(n16084), .A2(n18289), .B1(n19474), .B2(n16085), .ZN(
        U347) );
  INV_X1 U19128 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18287) );
  INV_X1 U19129 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19473) );
  AOI22_X1 U19130 ( .A1(n16084), .A2(n18287), .B1(n19473), .B2(n16085), .ZN(
        U348) );
  INV_X1 U19131 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18284) );
  INV_X1 U19132 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19472) );
  AOI22_X1 U19133 ( .A1(n16084), .A2(n18284), .B1(n19472), .B2(n16085), .ZN(
        U349) );
  INV_X1 U19134 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18283) );
  INV_X1 U19135 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19471) );
  AOI22_X1 U19136 ( .A1(n16084), .A2(n18283), .B1(n19471), .B2(n16085), .ZN(
        U350) );
  INV_X1 U19137 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18281) );
  INV_X1 U19138 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19469) );
  AOI22_X1 U19139 ( .A1(n16084), .A2(n18281), .B1(n19469), .B2(n16085), .ZN(
        U351) );
  INV_X1 U19140 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18279) );
  INV_X1 U19141 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19467) );
  AOI22_X1 U19142 ( .A1(n16084), .A2(n18279), .B1(n19467), .B2(n16085), .ZN(
        U352) );
  INV_X1 U19143 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18277) );
  INV_X1 U19144 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20626) );
  AOI22_X1 U19145 ( .A1(n16084), .A2(n18277), .B1(n20626), .B2(n16085), .ZN(
        U353) );
  INV_X1 U19146 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18275) );
  AOI22_X1 U19147 ( .A1(n16084), .A2(n18275), .B1(n19465), .B2(n16085), .ZN(
        U354) );
  INV_X1 U19148 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18326) );
  INV_X1 U19149 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19510) );
  AOI22_X1 U19150 ( .A1(n16084), .A2(n18326), .B1(n19510), .B2(n16085), .ZN(
        U355) );
  INV_X1 U19151 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18324) );
  INV_X1 U19152 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19507) );
  AOI22_X1 U19153 ( .A1(n16084), .A2(n18324), .B1(n19507), .B2(n16085), .ZN(
        U356) );
  INV_X1 U19154 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18321) );
  INV_X1 U19155 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19505) );
  AOI22_X1 U19156 ( .A1(n16084), .A2(n18321), .B1(n19505), .B2(n16085), .ZN(
        U357) );
  INV_X1 U19157 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18320) );
  INV_X1 U19158 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19502) );
  AOI22_X1 U19159 ( .A1(n16084), .A2(n18320), .B1(n19502), .B2(n16085), .ZN(
        U358) );
  INV_X1 U19160 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18317) );
  INV_X1 U19161 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19501) );
  AOI22_X1 U19162 ( .A1(n16084), .A2(n18317), .B1(n19501), .B2(n16085), .ZN(
        U359) );
  INV_X1 U19163 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18315) );
  INV_X1 U19164 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19499) );
  AOI22_X1 U19165 ( .A1(n16084), .A2(n18315), .B1(n19499), .B2(n16085), .ZN(
        U360) );
  INV_X1 U19166 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18312) );
  INV_X1 U19167 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19497) );
  AOI22_X1 U19168 ( .A1(n16084), .A2(n18312), .B1(n19497), .B2(n16085), .ZN(
        U361) );
  INV_X1 U19169 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18310) );
  INV_X1 U19170 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19495) );
  AOI22_X1 U19171 ( .A1(n16084), .A2(n18310), .B1(n19495), .B2(n16085), .ZN(
        U362) );
  INV_X1 U19172 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18309) );
  INV_X1 U19173 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19493) );
  AOI22_X1 U19174 ( .A1(n16084), .A2(n18309), .B1(n19493), .B2(n16085), .ZN(
        U363) );
  INV_X1 U19175 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18307) );
  INV_X1 U19176 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19491) );
  AOI22_X1 U19177 ( .A1(n16084), .A2(n18307), .B1(n19491), .B2(n16085), .ZN(
        U364) );
  INV_X1 U19178 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18273) );
  INV_X1 U19179 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19464) );
  AOI22_X1 U19180 ( .A1(n16084), .A2(n18273), .B1(n19464), .B2(n16085), .ZN(
        U365) );
  INV_X1 U19181 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18304) );
  INV_X1 U19182 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19489) );
  AOI22_X1 U19183 ( .A1(n16084), .A2(n18304), .B1(n19489), .B2(n16085), .ZN(
        U366) );
  INV_X1 U19184 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18303) );
  INV_X1 U19185 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19488) );
  AOI22_X1 U19186 ( .A1(n16084), .A2(n18303), .B1(n19488), .B2(n16085), .ZN(
        U367) );
  INV_X1 U19187 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18301) );
  INV_X1 U19188 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19486) );
  AOI22_X1 U19189 ( .A1(n16084), .A2(n18301), .B1(n19486), .B2(n16085), .ZN(
        U368) );
  INV_X1 U19190 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n20624) );
  INV_X1 U19191 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19484) );
  AOI22_X1 U19192 ( .A1(n16084), .A2(n20624), .B1(n19484), .B2(n16085), .ZN(
        U369) );
  INV_X1 U19193 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18298) );
  INV_X1 U19194 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19482) );
  AOI22_X1 U19195 ( .A1(n16084), .A2(n18298), .B1(n19482), .B2(n16085), .ZN(
        U370) );
  INV_X1 U19196 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18296) );
  INV_X1 U19197 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19481) );
  AOI22_X1 U19198 ( .A1(n16084), .A2(n18296), .B1(n19481), .B2(n16085), .ZN(
        U371) );
  INV_X1 U19199 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18294) );
  INV_X1 U19200 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19479) );
  AOI22_X1 U19201 ( .A1(n16084), .A2(n18294), .B1(n19479), .B2(n16085), .ZN(
        U372) );
  INV_X1 U19202 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n20707) );
  INV_X1 U19203 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19478) );
  AOI22_X1 U19204 ( .A1(n16084), .A2(n20707), .B1(n19478), .B2(n16085), .ZN(
        U373) );
  INV_X1 U19205 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18293) );
  INV_X1 U19206 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19476) );
  AOI22_X1 U19207 ( .A1(n16084), .A2(n18293), .B1(n19476), .B2(n16085), .ZN(
        U374) );
  INV_X1 U19208 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18291) );
  INV_X1 U19209 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19475) );
  AOI22_X1 U19210 ( .A1(n16084), .A2(n18291), .B1(n19475), .B2(n16085), .ZN(
        U375) );
  INV_X1 U19211 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18271) );
  INV_X1 U19212 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19461) );
  AOI22_X1 U19213 ( .A1(n16084), .A2(n18271), .B1(n19461), .B2(n16085), .ZN(
        U376) );
  INV_X1 U19214 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18270) );
  NAND2_X1 U19215 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18270), .ZN(n16086) );
  INV_X1 U19216 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n20611) );
  NAND2_X1 U19217 ( .A1(n20637), .A2(n20611), .ZN(n18257) );
  OAI21_X1 U19218 ( .B1(n16086), .B2(n20611), .A(n18257), .ZN(n18336) );
  AOI21_X1 U19219 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n18336), .ZN(n16087) );
  INV_X1 U19220 ( .A(n16087), .ZN(P3_U2633) );
  INV_X1 U19221 ( .A(P3_CODEFETCH_REG_SCAN_IN), .ZN(n16090) );
  NAND2_X1 U19222 ( .A1(n18222), .A2(n18235), .ZN(n16975) );
  NOR2_X1 U19223 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18394), .ZN(n18248) );
  NAND2_X1 U19224 ( .A1(n16088), .A2(n18248), .ZN(n16089) );
  OAI221_X1 U19225 ( .B1(n16090), .B2(n16974), .C1(n16090), .C2(n16094), .A(
        n16089), .ZN(P3_U2634) );
  NOR2_X1 U19226 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n16092) );
  AOI22_X1 U19227 ( .A1(P3_D_C_N_REG_SCAN_IN), .A2(n18401), .B1(n16092), .B2(
        n20637), .ZN(n16091) );
  OAI21_X1 U19228 ( .B1(P3_CODEFETCH_REG_SCAN_IN), .B2(n18401), .A(n16091), 
        .ZN(P3_U2635) );
  OAI21_X1 U19229 ( .B1(n16092), .B2(BS16), .A(n18336), .ZN(n18334) );
  OAI21_X1 U19230 ( .B1(n18336), .B2(n16113), .A(n18334), .ZN(P3_U2636) );
  AND3_X1 U19231 ( .A1(n16094), .A2(n18222), .A3(n16093), .ZN(n18225) );
  NOR2_X1 U19232 ( .A1(n18225), .A2(n18243), .ZN(n18382) );
  OAI21_X1 U19233 ( .B1(n18382), .B2(n17725), .A(n16095), .ZN(P3_U2637) );
  NOR4_X1 U19234 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16099) );
  NOR4_X1 U19235 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n16098) );
  NOR4_X1 U19236 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16097) );
  NOR4_X1 U19237 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16096) );
  NAND4_X1 U19238 ( .A1(n16099), .A2(n16098), .A3(n16097), .A4(n16096), .ZN(
        n16105) );
  NOR4_X1 U19239 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n16103) );
  AOI211_X1 U19240 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_19__SCAN_IN), .B(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n16102) );
  NOR4_X1 U19241 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n16101) );
  NOR4_X1 U19242 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n16100) );
  NAND4_X1 U19243 ( .A1(n16103), .A2(n16102), .A3(n16101), .A4(n16100), .ZN(
        n16104) );
  NOR2_X1 U19244 ( .A1(n16105), .A2(n16104), .ZN(n18375) );
  INV_X1 U19245 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16107) );
  NOR3_X1 U19246 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16108) );
  OAI21_X1 U19247 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16108), .A(n18375), .ZN(
        n16106) );
  OAI21_X1 U19248 ( .B1(n18375), .B2(n16107), .A(n16106), .ZN(P3_U2638) );
  INV_X1 U19249 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18371) );
  INV_X1 U19250 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18335) );
  AOI21_X1 U19251 ( .B1(n18371), .B2(n18335), .A(n16108), .ZN(n16110) );
  INV_X1 U19252 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16109) );
  INV_X1 U19253 ( .A(n18375), .ZN(n18378) );
  AOI22_X1 U19254 ( .A1(n18375), .A2(n16110), .B1(n16109), .B2(n18378), .ZN(
        P3_U2639) );
  NAND2_X1 U19255 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .ZN(n16141) );
  INV_X1 U19256 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18311) );
  INV_X1 U19257 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18305) );
  NAND3_X1 U19258 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .ZN(n16138) );
  INV_X1 U19259 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n20705) );
  INV_X1 U19260 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n20706) );
  NAND3_X1 U19261 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(P3_REIP_REG_10__SCAN_IN), 
        .A3(P3_REIP_REG_9__SCAN_IN), .ZN(n16137) );
  OAI211_X1 U19262 ( .C1(n18391), .C2(n18390), .A(n18385), .B(n16113), .ZN(
        n18237) );
  NOR2_X4 U19263 ( .A1(n18237), .A2(n16112), .ZN(n16470) );
  INV_X1 U19264 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18285) );
  INV_X1 U19265 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18280) );
  INV_X1 U19266 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18276) );
  NAND3_X1 U19267 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16429) );
  NOR2_X1 U19268 ( .A1(n18276), .A2(n16429), .ZN(n16416) );
  NAND2_X1 U19269 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16416), .ZN(n16414) );
  NOR2_X1 U19270 ( .A1(n18280), .A2(n16414), .ZN(n16388) );
  NAND2_X1 U19271 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n16388), .ZN(n16376) );
  NOR2_X1 U19272 ( .A1(n18285), .A2(n16376), .ZN(n16136) );
  NAND2_X1 U19273 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16335), .ZN(n16327) );
  NAND3_X1 U19274 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .A3(n16269), .ZN(n16254) );
  NAND3_X1 U19275 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .A3(n16241), .ZN(n16223) );
  NAND2_X1 U19276 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16140), .ZN(n16200) );
  NAND4_X1 U19277 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16185), .ZN(n16146) );
  NAND2_X1 U19278 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n18325), .ZN(n16145) );
  NAND2_X1 U19279 ( .A1(n16113), .A2(n18385), .ZN(n16114) );
  NOR2_X1 U19280 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n16464) );
  NAND2_X1 U19281 ( .A1(n16464), .A2(n16767), .ZN(n16453) );
  NOR2_X1 U19282 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n16453), .ZN(n16440) );
  NAND2_X1 U19283 ( .A1(n16440), .A2(n16759), .ZN(n16430) );
  NAND2_X1 U19284 ( .A1(n16411), .A2(n16756), .ZN(n16407) );
  INV_X1 U19285 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n16383) );
  NAND2_X1 U19286 ( .A1(n16387), .A2(n16383), .ZN(n16382) );
  NAND2_X1 U19287 ( .A1(n16367), .A2(n16701), .ZN(n16360) );
  NAND2_X1 U19288 ( .A1(n16345), .A2(n16337), .ZN(n16336) );
  NAND2_X1 U19289 ( .A1(n16320), .A2(n16308), .ZN(n16306) );
  NAND2_X1 U19290 ( .A1(n16297), .A2(n16647), .ZN(n16286) );
  NAND2_X1 U19291 ( .A1(n16274), .A2(n16604), .ZN(n16270) );
  INV_X1 U19292 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n16565) );
  NAND2_X1 U19293 ( .A1(n16257), .A2(n16565), .ZN(n16248) );
  INV_X1 U19294 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n16231) );
  NAND2_X1 U19295 ( .A1(n16236), .A2(n16231), .ZN(n16230) );
  INV_X1 U19296 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n20591) );
  NAND2_X1 U19297 ( .A1(n16217), .A2(n20591), .ZN(n16210) );
  INV_X1 U19298 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n16189) );
  NAND2_X1 U19299 ( .A1(n16198), .A2(n16189), .ZN(n16188) );
  NOR2_X1 U19300 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n16188), .ZN(n16180) );
  NAND2_X1 U19301 ( .A1(n16180), .A2(n16172), .ZN(n16171) );
  NOR2_X1 U19302 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16171), .ZN(n16147) );
  AND2_X1 U19303 ( .A1(n16466), .A2(n16147), .ZN(n16148) );
  INV_X1 U19304 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16492) );
  INV_X1 U19305 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16174) );
  NAND2_X1 U19306 ( .A1(n16117), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16116) );
  AOI21_X1 U19307 ( .B1(n16174), .B2(n16116), .A(n16115), .ZN(n17047) );
  OAI21_X1 U19308 ( .B1(n16117), .B2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16116), .ZN(n17069) );
  INV_X1 U19309 ( .A(n17069), .ZN(n16183) );
  INV_X1 U19310 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17140) );
  INV_X1 U19311 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17138) );
  NAND2_X1 U19312 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17124), .ZN(
        n16125) );
  NAND2_X1 U19313 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17084), .ZN(
        n16121) );
  INV_X1 U19314 ( .A(n16121), .ZN(n16120) );
  NAND2_X1 U19315 ( .A1(n17083), .A2(n16120), .ZN(n17046) );
  AOI21_X1 U19316 ( .B1(n10109), .B2(n17046), .A(n16117), .ZN(n17075) );
  NAND2_X1 U19317 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16120), .ZN(
        n16119) );
  INV_X1 U19318 ( .A(n17046), .ZN(n16118) );
  AOI21_X1 U19319 ( .B1(n17086), .B2(n16119), .A(n16118), .ZN(n17089) );
  AOI22_X1 U19320 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16120), .B1(
        n16121), .B2(n17098), .ZN(n17101) );
  OAI21_X1 U19321 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17084), .A(
        n16121), .ZN(n16122) );
  INV_X1 U19322 ( .A(n16122), .ZN(n17112) );
  INV_X1 U19323 ( .A(n16125), .ZN(n16124) );
  NAND2_X1 U19324 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16124), .ZN(
        n16123) );
  AOI21_X1 U19325 ( .B1(n17138), .B2(n16123), .A(n17084), .ZN(n17126) );
  AOI22_X1 U19326 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16124), .B1(
        n16125), .B2(n17140), .ZN(n17143) );
  INV_X1 U19327 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n20690) );
  INV_X1 U19328 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17166) );
  NAND3_X1 U19329 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17186), .A3(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17165) );
  NOR3_X1 U19330 ( .A1(n20690), .A2(n17166), .A3(n17165), .ZN(n17121) );
  OAI21_X1 U19331 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17121), .A(
        n16125), .ZN(n17155) );
  INV_X1 U19332 ( .A(n17155), .ZN(n16247) );
  INV_X1 U19333 ( .A(n17165), .ZN(n16127) );
  NAND2_X1 U19334 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16127), .ZN(
        n16126) );
  AOI21_X1 U19335 ( .B1(n17166), .B2(n16126), .A(n17121), .ZN(n17170) );
  XOR2_X1 U19336 ( .A(n20690), .B(n17165), .Z(n17178) );
  NAND2_X1 U19337 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17186), .ZN(
        n16129) );
  AOI21_X1 U19338 ( .B1(n17187), .B2(n16129), .A(n16127), .ZN(n17191) );
  INV_X1 U19339 ( .A(n16128), .ZN(n17202) );
  NAND2_X1 U19340 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17202), .ZN(
        n17203) );
  NOR2_X1 U19341 ( .A1(n17214), .A2(n17203), .ZN(n16294) );
  OAI21_X1 U19342 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16294), .A(
        n16129), .ZN(n16130) );
  INV_X1 U19343 ( .A(n16130), .ZN(n17205) );
  INV_X1 U19344 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16478) );
  NOR2_X1 U19345 ( .A1(n16276), .A2(n9609), .ZN(n16267) );
  NOR2_X1 U19346 ( .A1(n16245), .A2(n10079), .ZN(n16239) );
  NOR2_X1 U19347 ( .A1(n17143), .A2(n16239), .ZN(n16238) );
  NOR2_X1 U19348 ( .A1(n16216), .A2(n10079), .ZN(n16209) );
  NOR2_X1 U19349 ( .A1(n16208), .A2(n9609), .ZN(n16202) );
  NOR2_X1 U19350 ( .A1(n17089), .A2(n16202), .ZN(n16201) );
  NOR2_X1 U19351 ( .A1(n16182), .A2(n10079), .ZN(n16170) );
  NOR2_X1 U19352 ( .A1(n16169), .A2(n9609), .ZN(n16160) );
  NAND2_X1 U19353 ( .A1(n10073), .A2(n9771), .ZN(n16468) );
  NOR3_X1 U19354 ( .A1(n16152), .A2(n16151), .A3(n16468), .ZN(n16135) );
  NAND2_X1 U19355 ( .A1(n18403), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18246) );
  INV_X1 U19356 ( .A(n18246), .ZN(n18087) );
  NAND2_X1 U19357 ( .A1(n18087), .A2(n18248), .ZN(n18241) );
  NAND4_X1 U19358 ( .A1(n9746), .A2(n18384), .A3(n18251), .A4(n18241), .ZN(
        n16477) );
  INV_X1 U19359 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n16132) );
  OAI211_X1 U19360 ( .C1(n16132), .C2(n17741), .A(n18237), .B(n16131), .ZN(
        n16482) );
  OAI22_X1 U19361 ( .A1(n16133), .A2(n16467), .B1(n16132), .B2(n16482), .ZN(
        n16134) );
  AOI211_X1 U19362 ( .C1(n16148), .C2(n16492), .A(n16135), .B(n16134), .ZN(
        n16144) );
  NOR2_X1 U19363 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16146), .ZN(n16153) );
  INV_X1 U19364 ( .A(n16470), .ZN(n16450) );
  NAND2_X1 U19365 ( .A1(n16477), .A2(n16450), .ZN(n16485) );
  INV_X1 U19366 ( .A(n16485), .ZN(n16329) );
  INV_X1 U19367 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18323) );
  INV_X1 U19368 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18319) );
  NOR3_X1 U19369 ( .A1(n18322), .A2(n18323), .A3(n18319), .ZN(n16142) );
  NAND2_X1 U19370 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n16262) );
  NOR2_X1 U19371 ( .A1(n18305), .A2(n16262), .ZN(n16224) );
  NAND4_X1 U19372 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n16224), .A3(
        P3_REIP_REG_22__SCAN_IN), .A4(P3_REIP_REG_21__SCAN_IN), .ZN(n16139) );
  NAND2_X1 U19373 ( .A1(n16136), .A2(n16477), .ZN(n16358) );
  NOR2_X1 U19374 ( .A1(n16358), .A2(n16137), .ZN(n16328) );
  NAND2_X1 U19375 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16328), .ZN(n16316) );
  NOR2_X1 U19376 ( .A1(n20705), .A2(n16316), .ZN(n16311) );
  NAND2_X1 U19377 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16311), .ZN(n16283) );
  NOR2_X1 U19378 ( .A1(n16283), .A2(n16138), .ZN(n16225) );
  NOR2_X1 U19379 ( .A1(n16329), .A2(n16225), .ZN(n16280) );
  AOI21_X1 U19380 ( .B1(n16485), .B2(n16139), .A(n16280), .ZN(n16222) );
  INV_X1 U19381 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18313) );
  NAND2_X1 U19382 ( .A1(n16140), .A2(n18313), .ZN(n16214) );
  NAND2_X1 U19383 ( .A1(n16222), .A2(n16214), .ZN(n16204) );
  AOI21_X1 U19384 ( .B1(n16470), .B2(n16141), .A(n16204), .ZN(n16168) );
  OAI21_X1 U19385 ( .B1(n16329), .B2(n16142), .A(n16168), .ZN(n16163) );
  OAI21_X1 U19386 ( .B1(n16153), .B2(n16163), .A(P3_REIP_REG_31__SCAN_IN), 
        .ZN(n16143) );
  OAI211_X1 U19387 ( .C1(n16146), .C2(n16145), .A(n16144), .B(n16143), .ZN(
        P3_U2640) );
  NOR2_X1 U19388 ( .A1(n16147), .A2(n16481), .ZN(n16158) );
  INV_X1 U19389 ( .A(n16158), .ZN(n16150) );
  NOR2_X1 U19390 ( .A1(n16469), .A2(n16148), .ZN(n16149) );
  MUX2_X1 U19391 ( .A(n16150), .B(n16149), .S(P3_EBX_REG_30__SCAN_IN), .Z(
        n16155) );
  OAI211_X1 U19392 ( .C1(n16156), .C2(n16467), .A(n16155), .B(n16154), .ZN(
        P3_U2641) );
  NAND2_X1 U19393 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16171), .ZN(n16157) );
  AOI22_X1 U19394 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16469), .B1(n16158), 
        .B2(n16157), .ZN(n16166) );
  NAND2_X1 U19395 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16185), .ZN(n16179) );
  NOR2_X1 U19396 ( .A1(n18322), .A2(n16179), .ZN(n16164) );
  AOI211_X1 U19397 ( .C1(n16161), .C2(n16160), .A(n16159), .B(n18251), .ZN(
        n16162) );
  AOI221_X1 U19398 ( .B1(n16164), .B2(n18323), .C1(n16163), .C2(
        P3_REIP_REG_29__SCAN_IN), .A(n16162), .ZN(n16165) );
  OAI211_X1 U19399 ( .C1(n16167), .C2(n16467), .A(n16166), .B(n16165), .ZN(
        P3_U2642) );
  INV_X1 U19400 ( .A(n16168), .ZN(n16193) );
  AOI21_X1 U19401 ( .B1(n16185), .B2(n18319), .A(n16193), .ZN(n16178) );
  AOI211_X1 U19402 ( .C1(n17047), .C2(n16170), .A(n16169), .B(n18251), .ZN(
        n16176) );
  OAI21_X1 U19403 ( .B1(n16180), .B2(n16172), .A(n16171), .ZN(n16173) );
  OAI22_X1 U19404 ( .A1(n16174), .A2(n16467), .B1(n16481), .B2(n16173), .ZN(
        n16175) );
  AOI211_X1 U19405 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16469), .A(n16176), .B(
        n16175), .ZN(n16177) );
  OAI221_X1 U19406 ( .B1(P3_REIP_REG_28__SCAN_IN), .B2(n16179), .C1(n18322), 
        .C2(n16178), .A(n16177), .ZN(P3_U2643) );
  INV_X1 U19407 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n20580) );
  AOI211_X1 U19408 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n16188), .A(n16180), .B(
        n16481), .ZN(n16181) );
  AOI21_X1 U19409 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n16469), .A(n16181), .ZN(
        n16187) );
  AOI211_X1 U19410 ( .C1(n16183), .C2(n10094), .A(n16182), .B(n18251), .ZN(
        n16184) );
  AOI221_X1 U19411 ( .B1(n16185), .B2(n18319), .C1(n16193), .C2(
        P3_REIP_REG_27__SCAN_IN), .A(n16184), .ZN(n16186) );
  OAI211_X1 U19412 ( .C1(n20580), .C2(n16467), .A(n16187), .B(n16186), .ZN(
        P3_U2644) );
  OAI21_X1 U19413 ( .B1(n16198), .B2(n16189), .A(n16188), .ZN(n16197) );
  AOI22_X1 U19414 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n16443), .B1(
        n16469), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n16196) );
  INV_X1 U19415 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18314) );
  NOR2_X1 U19416 ( .A1(n18314), .A2(n16200), .ZN(n16194) );
  INV_X1 U19417 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18316) );
  AOI211_X1 U19418 ( .C1(n17075), .C2(n16191), .A(n16190), .B(n18251), .ZN(
        n16192) );
  AOI221_X1 U19419 ( .B1(n16194), .B2(n18316), .C1(n16193), .C2(
        P3_REIP_REG_26__SCAN_IN), .A(n16192), .ZN(n16195) );
  OAI211_X1 U19420 ( .C1(n16481), .C2(n16197), .A(n16196), .B(n16195), .ZN(
        P3_U2645) );
  AOI211_X1 U19421 ( .C1(P3_EBX_REG_25__SCAN_IN), .C2(n16210), .A(n16198), .B(
        n16481), .ZN(n16199) );
  AOI21_X1 U19422 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n16469), .A(n16199), .ZN(
        n16207) );
  INV_X1 U19423 ( .A(n16200), .ZN(n16205) );
  AOI211_X1 U19424 ( .C1(n17089), .C2(n16202), .A(n16201), .B(n18251), .ZN(
        n16203) );
  AOI221_X1 U19425 ( .B1(n16205), .B2(n18314), .C1(n16204), .C2(
        P3_REIP_REG_25__SCAN_IN), .A(n16203), .ZN(n16206) );
  OAI211_X1 U19426 ( .C1(n17086), .C2(n16467), .A(n16207), .B(n16206), .ZN(
        P3_U2646) );
  AOI211_X1 U19427 ( .C1(n17101), .C2(n16209), .A(n16208), .B(n18251), .ZN(
        n16213) );
  OAI21_X1 U19428 ( .B1(n16217), .B2(n20591), .A(n16210), .ZN(n16211) );
  OAI22_X1 U19429 ( .A1(n16482), .A2(n20591), .B1(n16481), .B2(n16211), .ZN(
        n16212) );
  AOI211_X1 U19430 ( .C1(n16443), .C2(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16213), .B(n16212), .ZN(n16215) );
  OAI211_X1 U19431 ( .C1(n16222), .C2(n18313), .A(n16215), .B(n16214), .ZN(
        P3_U2647) );
  AOI211_X1 U19432 ( .C1(n17112), .C2(n9742), .A(n16216), .B(n18251), .ZN(
        n16220) );
  AOI211_X1 U19433 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n16230), .A(n16217), .B(
        n16481), .ZN(n16219) );
  INV_X1 U19434 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16532) );
  OAI22_X1 U19435 ( .A1(n17085), .A2(n16467), .B1(n16482), .B2(n16532), .ZN(
        n16218) );
  NOR3_X1 U19436 ( .A1(n16220), .A2(n16219), .A3(n16218), .ZN(n16221) );
  OAI221_X1 U19437 ( .B1(P3_REIP_REG_23__SCAN_IN), .B2(n16223), .C1(n18311), 
        .C2(n16222), .A(n16221), .ZN(P3_U2648) );
  AOI22_X1 U19438 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n16443), .B1(
        n16469), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n16235) );
  AOI21_X1 U19439 ( .B1(n16225), .B2(n16224), .A(n16329), .ZN(n16244) );
  AOI211_X1 U19440 ( .C1(n17126), .C2(n16227), .A(n16226), .B(n18251), .ZN(
        n16228) );
  AOI21_X1 U19441 ( .B1(n16244), .B2(P3_REIP_REG_22__SCAN_IN), .A(n16228), 
        .ZN(n16234) );
  NAND2_X1 U19442 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .ZN(n16229) );
  OAI211_X1 U19443 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(P3_REIP_REG_21__SCAN_IN), .A(n16241), .B(n16229), .ZN(n16233) );
  OAI211_X1 U19444 ( .C1(n16236), .C2(n16231), .A(n16466), .B(n16230), .ZN(
        n16232) );
  NAND4_X1 U19445 ( .A1(n16235), .A2(n16234), .A3(n16233), .A4(n16232), .ZN(
        P3_U2649) );
  AOI211_X1 U19446 ( .C1(P3_EBX_REG_21__SCAN_IN), .C2(n16248), .A(n16236), .B(
        n16481), .ZN(n16237) );
  AOI21_X1 U19447 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n16469), .A(n16237), .ZN(
        n16243) );
  INV_X1 U19448 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18306) );
  AOI211_X1 U19449 ( .C1(n17143), .C2(n16239), .A(n16238), .B(n18251), .ZN(
        n16240) );
  AOI221_X1 U19450 ( .B1(n16244), .B2(P3_REIP_REG_21__SCAN_IN), .C1(n16241), 
        .C2(n18306), .A(n16240), .ZN(n16242) );
  OAI211_X1 U19451 ( .C1(n17140), .C2(n16467), .A(n16243), .B(n16242), .ZN(
        P3_U2650) );
  INV_X1 U19452 ( .A(n16244), .ZN(n16253) );
  AOI211_X1 U19453 ( .C1(n16247), .C2(n16246), .A(n16245), .B(n18251), .ZN(
        n16251) );
  OAI211_X1 U19454 ( .C1(n16257), .C2(n16565), .A(n16466), .B(n16248), .ZN(
        n16249) );
  OAI21_X1 U19455 ( .B1(n16565), .B2(n16482), .A(n16249), .ZN(n16250) );
  AOI211_X1 U19456 ( .C1(n16443), .C2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16251), .B(n16250), .ZN(n16252) );
  OAI221_X1 U19457 ( .B1(P3_REIP_REG_20__SCAN_IN), .B2(n16254), .C1(n18305), 
        .C2(n16253), .A(n16252), .ZN(P3_U2651) );
  INV_X1 U19458 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18302) );
  INV_X1 U19459 ( .A(n16280), .ZN(n16265) );
  AOI211_X1 U19460 ( .C1(n17170), .C2(n16256), .A(n16255), .B(n18251), .ZN(
        n16261) );
  AOI211_X1 U19461 ( .C1(P3_EBX_REG_19__SCAN_IN), .C2(n16270), .A(n16257), .B(
        n16481), .ZN(n16260) );
  AOI22_X1 U19462 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n16443), .B1(
        n16469), .B2(P3_EBX_REG_19__SCAN_IN), .ZN(n16258) );
  INV_X1 U19463 ( .A(n16258), .ZN(n16259) );
  NOR4_X1 U19464 ( .A1(n17710), .A2(n16261), .A3(n16260), .A4(n16259), .ZN(
        n16264) );
  OAI211_X1 U19465 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(P3_REIP_REG_18__SCAN_IN), .A(n16269), .B(n16262), .ZN(n16263) );
  OAI211_X1 U19466 ( .C1(n18302), .C2(n16265), .A(n16264), .B(n16263), .ZN(
        P3_U2652) );
  AOI22_X1 U19467 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16443), .B1(
        n16469), .B2(P3_EBX_REG_18__SCAN_IN), .ZN(n16273) );
  INV_X1 U19468 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18300) );
  AOI211_X1 U19469 ( .C1(n17178), .C2(n16267), .A(n16266), .B(n18251), .ZN(
        n16268) );
  AOI221_X1 U19470 ( .B1(n16280), .B2(P3_REIP_REG_18__SCAN_IN), .C1(n16269), 
        .C2(n18300), .A(n16268), .ZN(n16272) );
  OAI211_X1 U19471 ( .C1(n16274), .C2(n16604), .A(n16466), .B(n16270), .ZN(
        n16271) );
  NAND4_X1 U19472 ( .A1(n16273), .A2(n16272), .A3(n9746), .A4(n16271), .ZN(
        P3_U2653) );
  AOI211_X1 U19473 ( .C1(P3_EBX_REG_17__SCAN_IN), .C2(n16286), .A(n16274), .B(
        n16481), .ZN(n16275) );
  AOI211_X1 U19474 ( .C1(n16469), .C2(P3_EBX_REG_17__SCAN_IN), .A(n17710), .B(
        n16275), .ZN(n16282) );
  NAND2_X1 U19475 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16290) );
  NOR3_X1 U19476 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n16290), .A3(n16303), 
        .ZN(n16279) );
  AOI211_X1 U19477 ( .C1(n17191), .C2(n16277), .A(n16276), .B(n18251), .ZN(
        n16278) );
  AOI211_X1 U19478 ( .C1(n16280), .C2(P3_REIP_REG_17__SCAN_IN), .A(n16279), 
        .B(n16278), .ZN(n16281) );
  OAI211_X1 U19479 ( .C1(n17187), .C2(n16467), .A(n16282), .B(n16281), .ZN(
        P3_U2654) );
  NAND2_X1 U19480 ( .A1(n16485), .A2(n16283), .ZN(n16309) );
  INV_X1 U19481 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18297) );
  AOI211_X1 U19482 ( .C1(n17205), .C2(n16285), .A(n16284), .B(n18251), .ZN(
        n16289) );
  OAI211_X1 U19483 ( .C1(n16297), .C2(n16647), .A(n16466), .B(n16286), .ZN(
        n16287) );
  OAI211_X1 U19484 ( .C1(n16482), .C2(n16647), .A(n9746), .B(n16287), .ZN(
        n16288) );
  AOI211_X1 U19485 ( .C1(n16443), .C2(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n16289), .B(n16288), .ZN(n16293) );
  OAI211_X1 U19486 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(P3_REIP_REG_15__SCAN_IN), .A(n16291), .B(n16290), .ZN(n16292) );
  OAI211_X1 U19487 ( .C1(n16309), .C2(n18297), .A(n16293), .B(n16292), .ZN(
        P3_U2655) );
  INV_X1 U19488 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18295) );
  AOI21_X1 U19489 ( .B1(n17214), .B2(n17203), .A(n16294), .ZN(n17217) );
  NOR2_X1 U19490 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17402), .ZN(
        n16460) );
  AOI21_X1 U19491 ( .B1(n17202), .B2(n16460), .A(n9609), .ZN(n16296) );
  OAI21_X1 U19492 ( .B1(n17217), .B2(n16296), .A(n9771), .ZN(n16295) );
  AOI21_X1 U19493 ( .B1(n17217), .B2(n16296), .A(n16295), .ZN(n16301) );
  AOI211_X1 U19494 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n16306), .A(n16297), .B(
        n16481), .ZN(n16300) );
  AOI22_X1 U19495 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n16443), .B1(
        n16469), .B2(P3_EBX_REG_15__SCAN_IN), .ZN(n16298) );
  INV_X1 U19496 ( .A(n16298), .ZN(n16299) );
  NOR4_X1 U19497 ( .A1(n17710), .A2(n16301), .A3(n16300), .A4(n16299), .ZN(
        n16302) );
  OAI221_X1 U19498 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n16303), .C1(n18295), 
        .C2(n16309), .A(n16302), .ZN(P3_U2656) );
  AOI21_X1 U19499 ( .B1(n17260), .B2(n16460), .A(n9609), .ZN(n16333) );
  AOI21_X1 U19500 ( .B1(n10073), .B2(n17228), .A(n16333), .ZN(n16305) );
  INV_X1 U19501 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17227) );
  NAND2_X1 U19502 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16343), .ZN(
        n16357) );
  INV_X1 U19503 ( .A(n16357), .ZN(n16342) );
  NAND2_X1 U19504 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n16342), .ZN(
        n16341) );
  INV_X1 U19505 ( .A(n16341), .ZN(n17246) );
  NAND2_X1 U19506 ( .A1(n17250), .A2(n17246), .ZN(n16317) );
  INV_X1 U19507 ( .A(n17203), .ZN(n16304) );
  AOI21_X1 U19508 ( .B1(n17227), .B2(n16317), .A(n16304), .ZN(n17229) );
  XOR2_X1 U19509 ( .A(n16305), .B(n17229), .Z(n16315) );
  OAI211_X1 U19510 ( .C1(n16320), .C2(n16308), .A(n16466), .B(n16306), .ZN(
        n16307) );
  OAI211_X1 U19511 ( .C1(n16482), .C2(n16308), .A(n9746), .B(n16307), .ZN(
        n16313) );
  OAI22_X1 U19512 ( .A1(n16311), .A2(n16310), .B1(n20705), .B2(n16309), .ZN(
        n16312) );
  AOI211_X1 U19513 ( .C1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .C2(n16443), .A(
        n16313), .B(n16312), .ZN(n16314) );
  OAI21_X1 U19514 ( .B1(n16315), .B2(n18251), .A(n16314), .ZN(P3_U2657) );
  NAND2_X1 U19515 ( .A1(n16485), .A2(n16316), .ZN(n16326) );
  INV_X1 U19516 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17267) );
  AOI21_X1 U19517 ( .B1(n10073), .B2(n17267), .A(n16333), .ZN(n16319) );
  NOR2_X1 U19518 ( .A1(n17267), .A2(n16341), .ZN(n16330) );
  OAI21_X1 U19519 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16330), .A(
        n16317), .ZN(n17248) );
  OAI21_X1 U19520 ( .B1(n16319), .B2(n17248), .A(n9771), .ZN(n16318) );
  AOI21_X1 U19521 ( .B1(n16319), .B2(n17248), .A(n16318), .ZN(n16324) );
  AOI211_X1 U19522 ( .C1(P3_EBX_REG_13__SCAN_IN), .C2(n16336), .A(n16320), .B(
        n16481), .ZN(n16323) );
  AOI22_X1 U19523 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n16443), .B1(
        n16469), .B2(P3_EBX_REG_13__SCAN_IN), .ZN(n16321) );
  INV_X1 U19524 ( .A(n16321), .ZN(n16322) );
  NOR4_X1 U19525 ( .A1(n17710), .A2(n16324), .A3(n16323), .A4(n16322), .ZN(
        n16325) );
  OAI221_X1 U19526 ( .B1(P3_REIP_REG_13__SCAN_IN), .B2(n16327), .C1(n20706), 
        .C2(n16326), .A(n16325), .ZN(P3_U2658) );
  AOI22_X1 U19527 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16443), .B1(
        n16469), .B2(P3_EBX_REG_12__SCAN_IN), .ZN(n16340) );
  NOR2_X1 U19528 ( .A1(n16329), .A2(n16328), .ZN(n16346) );
  INV_X1 U19529 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18292) );
  AOI21_X1 U19530 ( .B1(n17267), .B2(n16341), .A(n16330), .ZN(n17257) );
  INV_X1 U19531 ( .A(n17257), .ZN(n16332) );
  INV_X1 U19532 ( .A(n16333), .ZN(n16331) );
  AOI221_X1 U19533 ( .B1(n17257), .B2(n16333), .C1(n16332), .C2(n16331), .A(
        n18251), .ZN(n16334) );
  AOI221_X1 U19534 ( .B1(n16346), .B2(P3_REIP_REG_12__SCAN_IN), .C1(n16335), 
        .C2(n18292), .A(n16334), .ZN(n16339) );
  OAI211_X1 U19535 ( .C1(n16345), .C2(n16337), .A(n16466), .B(n16336), .ZN(
        n16338) );
  NAND4_X1 U19536 ( .A1(n16340), .A2(n16339), .A3(n9746), .A4(n16338), .ZN(
        P3_U2659) );
  OAI21_X1 U19537 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16342), .A(
        n16341), .ZN(n17277) );
  AOI21_X1 U19538 ( .B1(n16343), .B2(n16460), .A(n9609), .ZN(n16344) );
  XOR2_X1 U19539 ( .A(n17277), .B(n16344), .Z(n16352) );
  AOI211_X1 U19540 ( .C1(P3_EBX_REG_11__SCAN_IN), .C2(n16360), .A(n16345), .B(
        n16481), .ZN(n16350) );
  INV_X1 U19541 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18288) );
  INV_X1 U19542 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18286) );
  NOR2_X1 U19543 ( .A1(n18288), .A2(n18286), .ZN(n16354) );
  INV_X1 U19544 ( .A(n16353), .ZN(n16366) );
  OAI221_X1 U19545 ( .B1(P3_REIP_REG_11__SCAN_IN), .B2(n16354), .C1(
        P3_REIP_REG_11__SCAN_IN), .C2(n16366), .A(n16346), .ZN(n16347) );
  OAI211_X1 U19546 ( .C1(n16482), .C2(n16348), .A(n9746), .B(n16347), .ZN(
        n16349) );
  AOI211_X1 U19547 ( .C1(n16443), .C2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n16350), .B(n16349), .ZN(n16351) );
  OAI21_X1 U19548 ( .B1(n18251), .B2(n16352), .A(n16351), .ZN(P3_U2660) );
  AOI211_X1 U19549 ( .C1(n18288), .C2(n18286), .A(n16354), .B(n16353), .ZN(
        n16355) );
  AOI211_X1 U19550 ( .C1(n16469), .C2(P3_EBX_REG_10__SCAN_IN), .A(n17715), .B(
        n16355), .ZN(n16364) );
  INV_X1 U19551 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17287) );
  INV_X1 U19552 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17331) );
  NOR3_X1 U19553 ( .A1(n17402), .A2(n17313), .A3(n17331), .ZN(n16393) );
  NAND2_X1 U19554 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16393), .ZN(
        n16375) );
  NOR2_X1 U19555 ( .A1(n17287), .A2(n16375), .ZN(n16365) );
  AOI21_X1 U19556 ( .B1(n16365), .B2(n16478), .A(n9609), .ZN(n16356) );
  INV_X1 U19557 ( .A(n16356), .ZN(n16368) );
  OAI21_X1 U19558 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16365), .A(
        n16357), .ZN(n17288) );
  XOR2_X1 U19559 ( .A(n16368), .B(n17288), .Z(n16359) );
  AND2_X1 U19560 ( .A1(n16485), .A2(n16358), .ZN(n16381) );
  AOI22_X1 U19561 ( .A1(n9771), .A2(n16359), .B1(P3_REIP_REG_10__SCAN_IN), 
        .B2(n16381), .ZN(n16363) );
  OAI211_X1 U19562 ( .C1(n16367), .C2(n16701), .A(n16466), .B(n16360), .ZN(
        n16362) );
  NAND2_X1 U19563 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n16443), .ZN(
        n16361) );
  NAND4_X1 U19564 ( .A1(n16364), .A2(n16363), .A3(n16362), .A4(n16361), .ZN(
        P3_U2661) );
  AOI22_X1 U19565 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16443), .B1(
        n16469), .B2(P3_EBX_REG_9__SCAN_IN), .ZN(n16374) );
  NAND2_X1 U19566 ( .A1(n9609), .A2(n9771), .ZN(n16463) );
  INV_X1 U19567 ( .A(n16463), .ZN(n16396) );
  AOI21_X1 U19568 ( .B1(n17287), .B2(n16375), .A(n16365), .ZN(n17306) );
  AOI22_X1 U19569 ( .A1(n16396), .A2(n17306), .B1(n16366), .B2(n18286), .ZN(
        n16373) );
  AOI211_X1 U19570 ( .C1(P3_EBX_REG_9__SCAN_IN), .C2(n16382), .A(n16367), .B(
        n16481), .ZN(n16371) );
  INV_X1 U19571 ( .A(n17313), .ZN(n17312) );
  NAND3_X1 U19572 ( .A1(n17312), .A2(n17297), .A3(n16460), .ZN(n16369) );
  AOI211_X1 U19573 ( .C1(n17306), .C2(n16369), .A(n18251), .B(n16368), .ZN(
        n16370) );
  AOI211_X1 U19574 ( .C1(n16381), .C2(P3_REIP_REG_9__SCAN_IN), .A(n16371), .B(
        n16370), .ZN(n16372) );
  NAND4_X1 U19575 ( .A1(n16374), .A2(n16373), .A3(n16372), .A4(n9746), .ZN(
        P3_U2662) );
  INV_X1 U19576 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16386) );
  AOI21_X1 U19577 ( .B1(n16393), .B2(n16478), .A(n9609), .ZN(n16397) );
  OAI21_X1 U19578 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16393), .A(
        n16375), .ZN(n17317) );
  XOR2_X1 U19579 ( .A(n16397), .B(n17317), .Z(n16379) );
  NOR2_X1 U19580 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16376), .ZN(n16377) );
  AOI22_X1 U19581 ( .A1(n16470), .A2(n16377), .B1(n16469), .B2(
        P3_EBX_REG_8__SCAN_IN), .ZN(n16378) );
  OAI211_X1 U19582 ( .C1(n18251), .C2(n16379), .A(n16378), .B(n9746), .ZN(
        n16380) );
  AOI21_X1 U19583 ( .B1(P3_REIP_REG_8__SCAN_IN), .B2(n16381), .A(n16380), .ZN(
        n16385) );
  OAI211_X1 U19584 ( .C1(n16387), .C2(n16383), .A(n16466), .B(n16382), .ZN(
        n16384) );
  OAI211_X1 U19585 ( .C1(n16467), .C2(n16386), .A(n16385), .B(n16384), .ZN(
        P3_U2663) );
  AOI211_X1 U19586 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n16407), .A(n16387), .B(
        n16481), .ZN(n16392) );
  NAND2_X1 U19587 ( .A1(n16470), .A2(n16388), .ZN(n16390) );
  INV_X1 U19588 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18282) );
  AOI221_X1 U19589 ( .B1(n18280), .B2(n16470), .C1(n16414), .C2(n16470), .A(
        n16479), .ZN(n16389) );
  OAI221_X1 U19590 ( .B1(P3_REIP_REG_7__SCAN_IN), .B2(n16390), .C1(n18282), 
        .C2(n16389), .A(n9746), .ZN(n16391) );
  AOI211_X1 U19591 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n16469), .A(n16392), .B(
        n16391), .ZN(n16399) );
  NOR2_X1 U19592 ( .A1(n17402), .A2(n17313), .ZN(n16400) );
  INV_X1 U19593 ( .A(n16400), .ZN(n16394) );
  AOI21_X1 U19594 ( .B1(n17331), .B2(n16394), .A(n16393), .ZN(n17336) );
  NAND2_X1 U19595 ( .A1(n17312), .A2(n16460), .ZN(n16401) );
  AOI21_X1 U19596 ( .B1(n17336), .B2(n16401), .A(n18251), .ZN(n16395) );
  OAI22_X1 U19597 ( .A1(n17336), .A2(n16397), .B1(n16396), .B2(n16395), .ZN(
        n16398) );
  OAI211_X1 U19598 ( .C1(n16467), .C2(n17331), .A(n16399), .B(n16398), .ZN(
        P3_U2664) );
  INV_X1 U19599 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n16410) );
  NOR3_X1 U19600 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n16450), .A3(n16414), .ZN(
        n16406) );
  AOI21_X1 U19601 ( .B1(n16470), .B2(n16414), .A(n16479), .ZN(n16422) );
  NAND2_X1 U19602 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17354), .ZN(
        n16412) );
  AOI21_X1 U19603 ( .B1(n16410), .B2(n16412), .A(n16400), .ZN(n17347) );
  AOI221_X1 U19604 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n10073), .C1(
        n16412), .C2(n10073), .A(n18251), .ZN(n16403) );
  NOR2_X1 U19605 ( .A1(n17347), .A2(n16468), .ZN(n16402) );
  AOI22_X1 U19606 ( .A1(n17347), .A2(n16403), .B1(n16402), .B2(n16401), .ZN(
        n16404) );
  OAI211_X1 U19607 ( .C1(n16422), .C2(n18280), .A(n16404), .B(n9746), .ZN(
        n16405) );
  AOI211_X1 U19608 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16469), .A(n16406), .B(
        n16405), .ZN(n16409) );
  OAI211_X1 U19609 ( .C1(n16411), .C2(n16756), .A(n16466), .B(n16407), .ZN(
        n16408) );
  OAI211_X1 U19610 ( .C1(n16467), .C2(n16410), .A(n16409), .B(n16408), .ZN(
        P3_U2665) );
  INV_X1 U19611 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18278) );
  AOI211_X1 U19612 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n16430), .A(n16411), .B(
        n16481), .ZN(n16420) );
  NOR2_X1 U19613 ( .A1(n17402), .A2(n17352), .ZN(n16413) );
  OAI21_X1 U19614 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n16413), .A(
        n16412), .ZN(n17359) );
  AOI21_X1 U19615 ( .B1(n10090), .B2(n16460), .A(n9609), .ZN(n16425) );
  XOR2_X1 U19616 ( .A(n17359), .B(n16425), .Z(n16418) );
  AND2_X1 U19617 ( .A1(n16414), .A2(n16470), .ZN(n16415) );
  AOI22_X1 U19618 ( .A1(n16416), .A2(n16415), .B1(n16469), .B2(
        P3_EBX_REG_5__SCAN_IN), .ZN(n16417) );
  OAI211_X1 U19619 ( .C1(n18251), .C2(n16418), .A(n16417), .B(n9746), .ZN(
        n16419) );
  AOI211_X1 U19620 ( .C1(n16443), .C2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n16420), .B(n16419), .ZN(n16421) );
  OAI21_X1 U19621 ( .B1(n16422), .B2(n18278), .A(n16421), .ZN(P3_U2666) );
  NAND2_X1 U19622 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16424) );
  NOR2_X1 U19623 ( .A1(n17402), .A2(n16424), .ZN(n16436) );
  OAI22_X1 U19624 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n16436), .B1(
        n17402), .B2(n17352), .ZN(n17371) );
  OAI22_X1 U19625 ( .A1(n16482), .A2(n16759), .B1(n17371), .B2(n16463), .ZN(
        n16423) );
  INV_X1 U19626 ( .A(n16423), .ZN(n16434) );
  NOR2_X1 U19627 ( .A1(n17736), .A2(n18384), .ZN(n18408) );
  INV_X1 U19628 ( .A(n18408), .ZN(n16487) );
  OAI221_X1 U19629 ( .B1(n16487), .B2(n9683), .C1(n16487), .C2(n18228), .A(
        n9746), .ZN(n16428) );
  AOI21_X1 U19630 ( .B1(n16470), .B2(n16429), .A(n16479), .ZN(n16447) );
  NOR2_X1 U19631 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n16424), .ZN(
        n17366) );
  AOI22_X1 U19632 ( .A1(n16460), .A2(n17366), .B1(n16425), .B2(n17371), .ZN(
        n16426) );
  OAI22_X1 U19633 ( .A1(n16447), .A2(n18276), .B1(n16426), .B2(n18251), .ZN(
        n16427) );
  AOI211_X1 U19634 ( .C1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .C2(n16443), .A(
        n16428), .B(n16427), .ZN(n16433) );
  OR3_X1 U19635 ( .A1(n16450), .A2(n16429), .A3(P3_REIP_REG_4__SCAN_IN), .ZN(
        n16432) );
  OAI211_X1 U19636 ( .C1(n16440), .C2(n16759), .A(n16466), .B(n16430), .ZN(
        n16431) );
  NAND4_X1 U19637 ( .A1(n16434), .A2(n16433), .A3(n16432), .A4(n16431), .ZN(
        P3_U2667) );
  INV_X1 U19638 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18272) );
  NOR2_X1 U19639 ( .A1(n18371), .A2(n18272), .ZN(n16451) );
  AOI21_X1 U19640 ( .B1(n16470), .B2(n16451), .A(P3_REIP_REG_3__SCAN_IN), .ZN(
        n16446) );
  NOR2_X1 U19641 ( .A1(n18355), .A2(n18362), .ZN(n18201) );
  NAND2_X1 U19642 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18201), .ZN(
        n18204) );
  INV_X1 U19643 ( .A(n18204), .ZN(n16452) );
  OAI21_X1 U19644 ( .B1(n16452), .B2(n18345), .A(n16435), .ZN(n18340) );
  AOI22_X1 U19645 ( .A1(n16469), .A2(P3_EBX_REG_3__SCAN_IN), .B1(n18408), .B2(
        n18340), .ZN(n16445) );
  INV_X1 U19646 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17395) );
  NOR2_X1 U19647 ( .A1(n17402), .A2(n17395), .ZN(n16448) );
  INV_X1 U19648 ( .A(n16436), .ZN(n16437) );
  OAI21_X1 U19649 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n16448), .A(
        n16437), .ZN(n17381) );
  AOI21_X1 U19650 ( .B1(n16478), .B2(n16448), .A(n9609), .ZN(n16458) );
  INV_X1 U19651 ( .A(n16458), .ZN(n16439) );
  OAI21_X1 U19652 ( .B1(n17381), .B2(n16439), .A(n9771), .ZN(n16438) );
  AOI21_X1 U19653 ( .B1(n17381), .B2(n16439), .A(n16438), .ZN(n16442) );
  AOI211_X1 U19654 ( .C1(P3_EBX_REG_3__SCAN_IN), .C2(n16453), .A(n16440), .B(
        n16481), .ZN(n16441) );
  AOI211_X1 U19655 ( .C1(n16443), .C2(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n16442), .B(n16441), .ZN(n16444) );
  OAI211_X1 U19656 ( .C1(n16447), .C2(n16446), .A(n16445), .B(n16444), .ZN(
        P3_U2668) );
  AOI21_X1 U19657 ( .B1(n17402), .B2(n17395), .A(n16448), .ZN(n16449) );
  INV_X1 U19658 ( .A(n16449), .ZN(n17392) );
  AOI211_X1 U19659 ( .C1(n18371), .C2(n18272), .A(n16451), .B(n16450), .ZN(
        n16457) );
  AOI21_X1 U19660 ( .B1(n18355), .B2(n18205), .A(n16452), .ZN(n18351) );
  AOI22_X1 U19661 ( .A1(n16479), .A2(P3_REIP_REG_2__SCAN_IN), .B1(n18351), 
        .B2(n18408), .ZN(n16455) );
  OAI211_X1 U19662 ( .C1(n16464), .C2(n16767), .A(n16466), .B(n16453), .ZN(
        n16454) );
  OAI211_X1 U19663 ( .C1(n16467), .C2(n17395), .A(n16455), .B(n16454), .ZN(
        n16456) );
  AOI211_X1 U19664 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16469), .A(n16457), .B(
        n16456), .ZN(n16462) );
  OAI211_X1 U19665 ( .C1(n16460), .C2(n17392), .A(n9771), .B(n16458), .ZN(
        n16461) );
  OAI211_X1 U19666 ( .C1(n16463), .C2(n17392), .A(n16462), .B(n16461), .ZN(
        P3_U2669) );
  AOI21_X1 U19667 ( .B1(P3_EBX_REG_1__SCAN_IN), .B2(P3_EBX_REG_0__SCAN_IN), 
        .A(n16464), .ZN(n16771) );
  AND2_X1 U19668 ( .A1(n16465), .A2(n18205), .ZN(n18359) );
  AOI22_X1 U19669 ( .A1(n16466), .A2(n16771), .B1(n18359), .B2(n18408), .ZN(
        n16476) );
  OAI21_X1 U19670 ( .B1(n16478), .B2(n16468), .A(n16467), .ZN(n16474) );
  AOI21_X1 U19671 ( .B1(n10073), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n18251), .ZN(n16473) );
  AOI22_X1 U19672 ( .A1(n18371), .A2(n16470), .B1(n16469), .B2(
        P3_EBX_REG_1__SCAN_IN), .ZN(n16471) );
  INV_X1 U19673 ( .A(n16471), .ZN(n16472) );
  AOI221_X1 U19674 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16474), .C1(
        n17402), .C2(n16473), .A(n16472), .ZN(n16475) );
  OAI211_X1 U19675 ( .C1(n16477), .C2(n18371), .A(n16476), .B(n16475), .ZN(
        P3_U2670) );
  NOR3_X1 U19676 ( .A1(n18404), .A2(n16479), .A3(n16478), .ZN(n16484) );
  AOI21_X1 U19677 ( .B1(n16482), .B2(n16481), .A(n16480), .ZN(n16483) );
  AOI211_X1 U19678 ( .C1(P3_REIP_REG_0__SCAN_IN), .C2(n16485), .A(n16484), .B(
        n16483), .ZN(n16486) );
  OAI21_X1 U19679 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n16487), .A(
        n16486), .ZN(P3_U2671) );
  NOR4_X1 U19680 ( .A1(n16565), .A2(n16602), .A3(n16523), .A4(n16522), .ZN(
        n16488) );
  NAND4_X1 U19681 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(P3_EBX_REG_21__SCAN_IN), .A4(n16488), .ZN(n16491) );
  NOR2_X1 U19682 ( .A1(n16492), .A2(n16491), .ZN(n16518) );
  NAND2_X1 U19683 ( .A1(n16774), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16490) );
  NAND2_X1 U19684 ( .A1(n16518), .A2(n17778), .ZN(n16489) );
  OAI22_X1 U19685 ( .A1(n16518), .A2(n16490), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n16489), .ZN(P3_U2672) );
  NAND2_X1 U19686 ( .A1(n16492), .A2(n16491), .ZN(n16493) );
  NAND2_X1 U19687 ( .A1(n16493), .A2(n16774), .ZN(n16517) );
  AOI22_X1 U19688 ( .A1(n9630), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n16634), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16497) );
  AOI22_X1 U19689 ( .A1(n9616), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16496) );
  AOI22_X1 U19690 ( .A1(n9622), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9640), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16495) );
  AOI22_X1 U19691 ( .A1(n16740), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9611), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16494) );
  NAND4_X1 U19692 ( .A1(n16497), .A2(n16496), .A3(n16495), .A4(n16494), .ZN(
        n16503) );
  AOI22_X1 U19693 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n16508), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16501) );
  AOI22_X1 U19694 ( .A1(n16739), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n15269), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16500) );
  AOI22_X1 U19695 ( .A1(n9629), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n16721), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16499) );
  AOI22_X1 U19696 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n16741), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16498) );
  NAND4_X1 U19697 ( .A1(n16501), .A2(n16500), .A3(n16499), .A4(n16498), .ZN(
        n16502) );
  NOR2_X1 U19698 ( .A1(n16503), .A2(n16502), .ZN(n16516) );
  AOI22_X1 U19699 ( .A1(n9616), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16721), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16507) );
  AOI22_X1 U19700 ( .A1(n16741), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16506) );
  AOI22_X1 U19701 ( .A1(n9613), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n16716), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16505) );
  AOI22_X1 U19702 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9642), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16504) );
  NAND4_X1 U19703 ( .A1(n16507), .A2(n16506), .A3(n16505), .A4(n16504), .ZN(
        n16514) );
  AOI22_X1 U19704 ( .A1(n16740), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9629), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16512) );
  AOI22_X1 U19705 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n16508), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16511) );
  AOI22_X1 U19706 ( .A1(n16739), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n15241), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16510) );
  AOI22_X1 U19707 ( .A1(n9630), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n16610), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16509) );
  NAND4_X1 U19708 ( .A1(n16512), .A2(n16511), .A3(n16510), .A4(n16509), .ZN(
        n16513) );
  NOR2_X1 U19709 ( .A1(n16514), .A2(n16513), .ZN(n16520) );
  NOR3_X1 U19710 ( .A1(n16520), .A2(n16528), .A3(n16519), .ZN(n16515) );
  XOR2_X1 U19711 ( .A(n16516), .B(n16515), .Z(n16785) );
  OAI22_X1 U19712 ( .A1(n16518), .A2(n16517), .B1(n16785), .B2(n16774), .ZN(
        P3_U2673) );
  INV_X1 U19713 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16526) );
  NOR2_X1 U19714 ( .A1(n16528), .A2(n16519), .ZN(n16521) );
  XNOR2_X1 U19715 ( .A(n16521), .B(n16520), .ZN(n16789) );
  NOR4_X1 U19716 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16546), .A3(n16523), .A4(
        n16522), .ZN(n16524) );
  AOI21_X1 U19717 ( .B1(n16765), .B2(n16789), .A(n16524), .ZN(n16525) );
  OAI21_X1 U19718 ( .B1(n16527), .B2(n16526), .A(n16525), .ZN(P3_U2674) );
  OAI21_X1 U19719 ( .B1(n16533), .B2(n16529), .A(n16528), .ZN(n16802) );
  INV_X1 U19720 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16530) );
  AOI22_X1 U19721 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n16535), .B1(n16537), 
        .B2(n16530), .ZN(n16531) );
  OAI21_X1 U19722 ( .B1(n16774), .B2(n16802), .A(n16531), .ZN(P3_U2676) );
  NOR2_X2 U19723 ( .A1(n16532), .A2(n16546), .ZN(n16551) );
  NAND2_X1 U19724 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n16545), .ZN(n16541) );
  AOI21_X1 U19725 ( .B1(n16534), .B2(n16538), .A(n16533), .ZN(n16803) );
  AOI22_X1 U19726 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16535), .B1(n16765), 
        .B2(n16803), .ZN(n16536) );
  OAI21_X1 U19727 ( .B1(n16537), .B2(n16541), .A(n16536), .ZN(P3_U2677) );
  OAI21_X1 U19728 ( .B1(n16540), .B2(n16539), .A(n16538), .ZN(n16811) );
  OAI211_X1 U19729 ( .C1(n16545), .C2(P3_EBX_REG_25__SCAN_IN), .A(n16774), .B(
        n16541), .ZN(n16542) );
  OAI21_X1 U19730 ( .B1(n16811), .B2(n16774), .A(n16542), .ZN(P3_U2678) );
  AOI21_X1 U19731 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n16774), .A(n16551), .ZN(
        n16544) );
  XNOR2_X1 U19732 ( .A(n16543), .B(n16547), .ZN(n16817) );
  OAI22_X1 U19733 ( .A1(n16545), .A2(n16544), .B1(n16774), .B2(n16817), .ZN(
        P3_U2679) );
  INV_X1 U19734 ( .A(n16546), .ZN(n16564) );
  AOI21_X1 U19735 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n16774), .A(n16564), .ZN(
        n16550) );
  OAI21_X1 U19736 ( .B1(n16549), .B2(n16548), .A(n16547), .ZN(n16823) );
  OAI22_X1 U19737 ( .A1(n16551), .A2(n16550), .B1(n16774), .B2(n16823), .ZN(
        P3_U2680) );
  AOI21_X1 U19738 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n16774), .A(n16552), .ZN(
        n16563) );
  AOI22_X1 U19739 ( .A1(n16740), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n16723), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16556) );
  AOI22_X1 U19740 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n16668), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16555) );
  AOI22_X1 U19741 ( .A1(n9629), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(n9642), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16554) );
  AOI22_X1 U19742 ( .A1(n16738), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16553) );
  NAND4_X1 U19743 ( .A1(n16556), .A2(n16555), .A3(n16554), .A4(n16553), .ZN(
        n16562) );
  AOI22_X1 U19744 ( .A1(n16623), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9613), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16560) );
  AOI22_X1 U19745 ( .A1(n16733), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9622), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16559) );
  AOI22_X1 U19746 ( .A1(n9616), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(n9620), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16558) );
  AOI22_X1 U19747 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n16610), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16557) );
  NAND4_X1 U19748 ( .A1(n16560), .A2(n16559), .A3(n16558), .A4(n16557), .ZN(
        n16561) );
  NOR2_X1 U19749 ( .A1(n16562), .A2(n16561), .ZN(n16824) );
  OAI22_X1 U19750 ( .A1(n16564), .A2(n16563), .B1(n16824), .B2(n16774), .ZN(
        P3_U2681) );
  OAI21_X1 U19751 ( .B1(n16565), .B2(n16602), .A(n16774), .ZN(n16590) );
  AOI22_X1 U19752 ( .A1(n16739), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9629), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16575) );
  AOI22_X1 U19753 ( .A1(n16740), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n16634), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n16574) );
  INV_X1 U19754 ( .A(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n20578) );
  AOI22_X1 U19755 ( .A1(n16716), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16566) );
  OAI21_X1 U19756 ( .B1(n9679), .B2(n20578), .A(n16566), .ZN(n16572) );
  AOI22_X1 U19757 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(n9630), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16570) );
  AOI22_X1 U19758 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n16721), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16569) );
  AOI22_X1 U19759 ( .A1(n16733), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n16723), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16568) );
  AOI22_X1 U19760 ( .A1(n9622), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9642), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16567) );
  NAND4_X1 U19761 ( .A1(n16570), .A2(n16569), .A3(n16568), .A4(n16567), .ZN(
        n16571) );
  AOI211_X1 U19762 ( .C1(n9613), .C2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A(
        n16572), .B(n16571), .ZN(n16573) );
  NAND3_X1 U19763 ( .A1(n16575), .A2(n16574), .A3(n16573), .ZN(n16831) );
  NAND2_X1 U19764 ( .A1(n16765), .A2(n16831), .ZN(n16576) );
  OAI221_X1 U19765 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n16578), .C1(n16577), 
        .C2(n16590), .A(n16576), .ZN(P3_U2682) );
  AOI22_X1 U19766 ( .A1(n16739), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n16721), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16582) );
  AOI22_X1 U19767 ( .A1(n16682), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9622), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16581) );
  AOI22_X1 U19768 ( .A1(n15219), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9620), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16580) );
  AOI22_X1 U19769 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9640), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16579) );
  NAND4_X1 U19770 ( .A1(n16582), .A2(n16581), .A3(n16580), .A4(n16579), .ZN(
        n16588) );
  AOI22_X1 U19771 ( .A1(n9611), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n16723), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16586) );
  AOI22_X1 U19772 ( .A1(n16733), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16585) );
  AOI22_X1 U19773 ( .A1(n9616), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(n9629), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n16584) );
  AOI22_X1 U19774 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n16634), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16583) );
  NAND4_X1 U19775 ( .A1(n16586), .A2(n16585), .A3(n16584), .A4(n16583), .ZN(
        n16587) );
  NOR2_X1 U19776 ( .A1(n16588), .A2(n16587), .ZN(n16839) );
  NOR2_X1 U19777 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16589), .ZN(n16591) );
  OAI22_X1 U19778 ( .A1(n16839), .A2(n16774), .B1(n16591), .B2(n16590), .ZN(
        P3_U2683) );
  AOI22_X1 U19779 ( .A1(n16733), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n15241), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n16595) );
  AOI22_X1 U19780 ( .A1(n9616), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15097), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n16594) );
  AOI22_X1 U19781 ( .A1(n9629), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(n9620), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n16593) );
  AOI22_X1 U19782 ( .A1(n16741), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9640), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16592) );
  NAND4_X1 U19783 ( .A1(n16595), .A2(n16594), .A3(n16593), .A4(n16592), .ZN(
        n16601) );
  AOI22_X1 U19784 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9621), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16599) );
  AOI22_X1 U19785 ( .A1(n16739), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9612), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16598) );
  AOI22_X1 U19786 ( .A1(n9630), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n16597) );
  AOI22_X1 U19787 ( .A1(n15219), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n16610), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n16596) );
  NAND4_X1 U19788 ( .A1(n16599), .A2(n16598), .A3(n16597), .A4(n16596), .ZN(
        n16600) );
  NOR2_X1 U19789 ( .A1(n16601), .A2(n16600), .ZN(n16844) );
  OAI21_X1 U19790 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n16618), .A(n16602), .ZN(
        n16603) );
  AOI22_X1 U19791 ( .A1(n16765), .A2(n16844), .B1(n16603), .B2(n16774), .ZN(
        P3_U2684) );
  AOI21_X1 U19792 ( .B1(n16604), .B2(n16631), .A(n16765), .ZN(n16605) );
  INV_X1 U19793 ( .A(n16605), .ZN(n16617) );
  AOI22_X1 U19794 ( .A1(n9611), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n16721), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n16609) );
  AOI22_X1 U19795 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(n9622), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n16608) );
  AOI22_X1 U19796 ( .A1(n16623), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n16607) );
  AOI22_X1 U19797 ( .A1(n16733), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9641), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n16606) );
  NAND4_X1 U19798 ( .A1(n16609), .A2(n16608), .A3(n16607), .A4(n16606), .ZN(
        n16616) );
  AOI22_X1 U19799 ( .A1(n15219), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9629), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n16614) );
  AOI22_X1 U19800 ( .A1(n9616), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n16610), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n16613) );
  AOI22_X1 U19801 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n16668), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n16612) );
  AOI22_X1 U19802 ( .A1(n16723), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n15269), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n16611) );
  NAND4_X1 U19803 ( .A1(n16614), .A2(n16613), .A3(n16612), .A4(n16611), .ZN(
        n16615) );
  NOR2_X1 U19804 ( .A1(n16616), .A2(n16615), .ZN(n16848) );
  OAI22_X1 U19805 ( .A1(n16618), .A2(n16617), .B1(n16848), .B2(n16774), .ZN(
        P3_U2685) );
  AOI22_X1 U19806 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n9612), .B1(
        n16668), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n16622) );
  AOI22_X1 U19807 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9616), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n16621) );
  AOI22_X1 U19808 ( .A1(n9629), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n15241), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n16620) );
  AOI22_X1 U19809 ( .A1(n15219), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9642), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n16619) );
  NAND4_X1 U19810 ( .A1(n16622), .A2(n16621), .A3(n16620), .A4(n16619), .ZN(
        n16630) );
  AOI22_X1 U19811 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n9630), .ZN(n16628) );
  AOI22_X1 U19812 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n15217), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n16634), .ZN(n16627) );
  AOI22_X1 U19813 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n16721), .B1(
        n16733), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n16626) );
  AOI22_X1 U19814 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n16723), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n16716), .ZN(n16625) );
  NAND4_X1 U19815 ( .A1(n16628), .A2(n16627), .A3(n16626), .A4(n16625), .ZN(
        n16629) );
  NOR2_X1 U19816 ( .A1(n16630), .A2(n16629), .ZN(n16855) );
  OAI21_X1 U19817 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n16632), .A(n16631), .ZN(
        n16633) );
  AOI22_X1 U19818 ( .A1(n16765), .A2(n16855), .B1(n16633), .B2(n16774), .ZN(
        P3_U2686) );
  AOI22_X1 U19819 ( .A1(n9622), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9620), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n16638) );
  AOI22_X1 U19820 ( .A1(n16623), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n16741), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n16637) );
  AOI22_X1 U19821 ( .A1(n9629), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(n9641), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n16636) );
  AOI22_X1 U19822 ( .A1(n16739), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n16634), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n16635) );
  NAND4_X1 U19823 ( .A1(n16638), .A2(n16637), .A3(n16636), .A4(n16635), .ZN(
        n16644) );
  AOI22_X1 U19824 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n16642) );
  AOI22_X1 U19825 ( .A1(n15219), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9612), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n16641) );
  AOI22_X1 U19826 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n16733), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n16640) );
  AOI22_X1 U19827 ( .A1(n9616), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n16721), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n16639) );
  NAND4_X1 U19828 ( .A1(n16642), .A2(n16641), .A3(n16640), .A4(n16639), .ZN(
        n16643) );
  NOR2_X1 U19829 ( .A1(n16644), .A2(n16643), .ZN(n16862) );
  AND3_X1 U19830 ( .A1(n17778), .A2(n16646), .A3(n16645), .ZN(n16662) );
  NAND4_X1 U19831 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .A3(n16662), .A4(n16647), .ZN(n16649) );
  NAND3_X1 U19832 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16774), .A3(n16660), 
        .ZN(n16648) );
  OAI211_X1 U19833 ( .C1(n16862), .C2(n16774), .A(n16649), .B(n16648), .ZN(
        P3_U2687) );
  AOI22_X1 U19834 ( .A1(n9616), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(n9620), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16653) );
  AOI22_X1 U19835 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n16668), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16652) );
  AOI22_X1 U19836 ( .A1(n9630), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n16634), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16651) );
  AOI22_X1 U19837 ( .A1(n16741), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9642), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16650) );
  NAND4_X1 U19838 ( .A1(n16653), .A2(n16652), .A3(n16651), .A4(n16650), .ZN(
        n16659) );
  AOI22_X1 U19839 ( .A1(n16738), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16657) );
  AOI22_X1 U19840 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9629), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16656) );
  AOI22_X1 U19841 ( .A1(n15219), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9611), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16655) );
  AOI22_X1 U19842 ( .A1(n16733), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n15241), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16654) );
  NAND4_X1 U19843 ( .A1(n16657), .A2(n16656), .A3(n16655), .A4(n16654), .ZN(
        n16658) );
  NOR2_X1 U19844 ( .A1(n16659), .A2(n16658), .ZN(n16866) );
  OAI211_X1 U19845 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n16676), .A(n16660), .B(
        n16774), .ZN(n16661) );
  OAI21_X1 U19846 ( .B1(n16866), .B2(n16774), .A(n16661), .ZN(P3_U2688) );
  OAI21_X1 U19847 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n16662), .A(n16774), .ZN(
        n16675) );
  AOI22_X1 U19848 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9616), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16667) );
  AOI22_X1 U19849 ( .A1(n9630), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n16721), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16666) );
  AOI22_X1 U19850 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n16723), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16665) );
  AOI22_X1 U19851 ( .A1(n9629), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(n9642), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16664) );
  NAND4_X1 U19852 ( .A1(n16667), .A2(n16666), .A3(n16665), .A4(n16664), .ZN(
        n16674) );
  AOI22_X1 U19853 ( .A1(n16733), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n16716), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16672) );
  AOI22_X1 U19854 ( .A1(n15219), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16668), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16671) );
  AOI22_X1 U19855 ( .A1(n15241), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16670) );
  AOI22_X1 U19856 ( .A1(n9613), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n16634), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16669) );
  NAND4_X1 U19857 ( .A1(n16672), .A2(n16671), .A3(n16670), .A4(n16669), .ZN(
        n16673) );
  NOR2_X1 U19858 ( .A1(n16674), .A2(n16673), .ZN(n16871) );
  OAI22_X1 U19859 ( .A1(n16676), .A2(n16675), .B1(n16871), .B2(n16774), .ZN(
        P3_U2689) );
  AOI21_X1 U19860 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n16774), .A(n16677), .ZN(
        n16689) );
  AOI22_X1 U19861 ( .A1(n9616), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(n9629), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n16681) );
  AOI22_X1 U19862 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n16733), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16680) );
  AOI22_X1 U19863 ( .A1(n16634), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n16679) );
  AOI22_X1 U19864 ( .A1(n15219), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9642), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16678) );
  NAND4_X1 U19865 ( .A1(n16681), .A2(n16680), .A3(n16679), .A4(n16678), .ZN(
        n16688) );
  AOI22_X1 U19866 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n16716), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16686) );
  AOI22_X1 U19867 ( .A1(n16682), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9612), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16685) );
  AOI22_X1 U19868 ( .A1(n16738), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n16723), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16684) );
  AOI22_X1 U19869 ( .A1(n16739), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9622), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16683) );
  NAND4_X1 U19870 ( .A1(n16686), .A2(n16685), .A3(n16684), .A4(n16683), .ZN(
        n16687) );
  NOR2_X1 U19871 ( .A1(n16688), .A2(n16687), .ZN(n16878) );
  OAI22_X1 U19872 ( .A1(n16690), .A2(n16689), .B1(n16878), .B2(n16774), .ZN(
        P3_U2691) );
  AOI22_X1 U19873 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n15241), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n16694) );
  AOI22_X1 U19874 ( .A1(n16739), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9612), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n16693) );
  AOI22_X1 U19875 ( .A1(n15219), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n16721), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n16692) );
  AOI22_X1 U19876 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9641), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16691) );
  NAND4_X1 U19877 ( .A1(n16694), .A2(n16693), .A3(n16692), .A4(n16691), .ZN(
        n16700) );
  AOI22_X1 U19878 ( .A1(n16733), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9616), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n16698) );
  AOI22_X1 U19879 ( .A1(n16741), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n16634), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16697) );
  AOI22_X1 U19880 ( .A1(n16682), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9629), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n16696) );
  AOI22_X1 U19881 ( .A1(n16716), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n16695) );
  NAND4_X1 U19882 ( .A1(n16698), .A2(n16697), .A3(n16696), .A4(n16695), .ZN(
        n16699) );
  NOR2_X1 U19883 ( .A1(n16700), .A2(n16699), .ZN(n16882) );
  NOR2_X1 U19884 ( .A1(n16701), .A2(n16730), .ZN(n16715) );
  OAI21_X1 U19885 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n16715), .A(n16702), .ZN(
        n16703) );
  AOI22_X1 U19886 ( .A1(n16765), .A2(n16882), .B1(n16703), .B2(n16774), .ZN(
        P3_U2692) );
  OAI21_X1 U19887 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n16646), .A(n16774), .ZN(
        n16714) );
  AOI22_X1 U19888 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(n9629), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n16707) );
  AOI22_X1 U19889 ( .A1(n16733), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n16739), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n16706) );
  AOI22_X1 U19890 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n16723), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n16705) );
  AOI22_X1 U19891 ( .A1(n15241), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9641), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n16704) );
  NAND4_X1 U19892 ( .A1(n16707), .A2(n16706), .A3(n16705), .A4(n16704), .ZN(
        n16713) );
  AOI22_X1 U19893 ( .A1(n15219), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n16716), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n16711) );
  AOI22_X1 U19894 ( .A1(n9616), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n16634), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n16710) );
  AOI22_X1 U19895 ( .A1(n16623), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n16709) );
  AOI22_X1 U19896 ( .A1(n9611), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n16721), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n16708) );
  NAND4_X1 U19897 ( .A1(n16711), .A2(n16710), .A3(n16709), .A4(n16708), .ZN(
        n16712) );
  NOR2_X1 U19898 ( .A1(n16713), .A2(n16712), .ZN(n16886) );
  OAI22_X1 U19899 ( .A1(n16715), .A2(n16714), .B1(n16886), .B2(n16774), .ZN(
        P3_U2693) );
  AOI22_X1 U19900 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n16716), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n15217), .ZN(n16720) );
  AOI22_X1 U19901 ( .A1(n15219), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n9616), .ZN(n16719) );
  AOI22_X1 U19902 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n9613), .B1(
        n16739), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n16718) );
  AOI22_X1 U19903 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n9642), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n15241), .ZN(n16717) );
  NAND4_X1 U19904 ( .A1(n16720), .A2(n16719), .A3(n16718), .A4(n16717), .ZN(
        n16729) );
  AOI22_X1 U19905 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n16721), .ZN(n16727) );
  AOI22_X1 U19906 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n16634), .B1(
        n16723), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n16726) );
  AOI22_X1 U19907 ( .A1(n9630), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9629), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n16725) );
  AOI22_X1 U19908 ( .A1(n9621), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n16733), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n16724) );
  NAND4_X1 U19909 ( .A1(n16727), .A2(n16726), .A3(n16725), .A4(n16724), .ZN(
        n16728) );
  NOR2_X1 U19910 ( .A1(n16729), .A2(n16728), .ZN(n16892) );
  OAI21_X1 U19911 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n16731), .A(n16730), .ZN(
        n16732) );
  AOI22_X1 U19912 ( .A1(n16765), .A2(n16892), .B1(n16732), .B2(n16774), .ZN(
        P3_U2694) );
  AOI22_X1 U19913 ( .A1(n16733), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n15269), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n16737) );
  AOI22_X1 U19914 ( .A1(n16722), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9621), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n16736) );
  AOI22_X1 U19915 ( .A1(n9613), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9642), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n16735) );
  AOI22_X1 U19916 ( .A1(n9622), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n15217), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n16734) );
  NAND4_X1 U19917 ( .A1(n16737), .A2(n16736), .A3(n16735), .A4(n16734), .ZN(
        n16747) );
  AOI22_X1 U19918 ( .A1(n16738), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n16634), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n16745) );
  AOI22_X1 U19919 ( .A1(n16739), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9629), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n16744) );
  AOI22_X1 U19920 ( .A1(n16740), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9616), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n16743) );
  AOI22_X1 U19921 ( .A1(n9630), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n16741), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n16742) );
  NAND4_X1 U19922 ( .A1(n16745), .A2(n16744), .A3(n16743), .A4(n16742), .ZN(
        n16746) );
  NOR2_X1 U19923 ( .A1(n16747), .A2(n16746), .ZN(n16900) );
  NOR3_X1 U19924 ( .A1(n16890), .A2(n16756), .A3(n16753), .ZN(n16750) );
  OAI221_X1 U19925 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(P3_EBX_REG_7__SCAN_IN), 
        .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16750), .A(n16748), .ZN(n16749) );
  AOI22_X1 U19926 ( .A1(n16765), .A2(n16900), .B1(n16749), .B2(n16774), .ZN(
        P3_U2695) );
  AOI21_X1 U19927 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n16774), .A(n16750), .ZN(
        n16751) );
  INV_X1 U19928 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17784) );
  OAI22_X1 U19929 ( .A1(n16752), .A2(n16751), .B1(n17784), .B2(n16774), .ZN(
        P3_U2696) );
  NAND2_X1 U19930 ( .A1(n16774), .A2(n16753), .ZN(n16757) );
  NOR2_X1 U19931 ( .A1(n16890), .A2(n16753), .ZN(n16754) );
  AOI22_X1 U19932 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n16765), .B1(
        n16754), .B2(n16756), .ZN(n16755) );
  OAI21_X1 U19933 ( .B1(n16756), .B2(n16757), .A(n16755), .ZN(P3_U2697) );
  NOR2_X1 U19934 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n16762), .ZN(n16758) );
  INV_X1 U19935 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17769) );
  OAI22_X1 U19936 ( .A1(n16758), .A2(n16757), .B1(n17769), .B2(n16774), .ZN(
        P3_U2698) );
  AOI21_X1 U19937 ( .B1(n16759), .B2(n16763), .A(n16765), .ZN(n16760) );
  INV_X1 U19938 ( .A(n16760), .ZN(n16761) );
  INV_X1 U19939 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17763) );
  OAI22_X1 U19940 ( .A1(n16762), .A2(n16761), .B1(n17763), .B2(n16774), .ZN(
        P3_U2699) );
  INV_X1 U19941 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17757) );
  OAI21_X1 U19942 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n16770), .A(n16763), .ZN(
        n16764) );
  AOI22_X1 U19943 ( .A1(n16765), .A2(n17757), .B1(n16764), .B2(n16774), .ZN(
        P3_U2700) );
  AOI21_X1 U19944 ( .B1(n16767), .B2(n16766), .A(n16765), .ZN(n16768) );
  INV_X1 U19945 ( .A(n16768), .ZN(n16769) );
  INV_X1 U19946 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17751) );
  OAI22_X1 U19947 ( .A1(n16770), .A2(n16769), .B1(n17751), .B2(n16774), .ZN(
        P3_U2701) );
  INV_X1 U19948 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17745) );
  AOI22_X1 U19949 ( .A1(P3_EBX_REG_1__SCAN_IN), .A2(n16772), .B1(n16775), .B2(
        n16771), .ZN(n16773) );
  OAI21_X1 U19950 ( .B1(n17745), .B2(n16774), .A(n16773), .ZN(P3_U2702) );
  NOR2_X1 U19951 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n16775), .ZN(n16776) );
  INV_X1 U19952 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17739) );
  OAI22_X1 U19953 ( .A1(n16777), .A2(n16776), .B1(n17739), .B2(n16774), .ZN(
        P3_U2703) );
  INV_X1 U19954 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17001) );
  INV_X1 U19955 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n16997) );
  INV_X1 U19956 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n16995) );
  INV_X1 U19957 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n16993) );
  INV_X1 U19958 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n16979) );
  INV_X1 U19959 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17011) );
  NAND4_X1 U19960 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n16778) );
  NOR3_X1 U19961 ( .A1(n17011), .A2(n17009), .A3(n16778), .ZN(n16779) );
  NAND3_X1 U19962 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(P3_EAX_REG_7__SCAN_IN), 
        .A3(n16779), .ZN(n16901) );
  NOR2_X1 U19963 ( .A1(n16929), .A2(n16901), .ZN(n16897) );
  NAND2_X1 U19964 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n16897), .ZN(n16896) );
  INV_X1 U19965 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17032) );
  INV_X1 U19966 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17029) );
  NAND4_X1 U19967 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(P3_EAX_REG_13__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(P3_EAX_REG_9__SCAN_IN), .ZN(n16780)
         );
  NAND2_X1 U19968 ( .A1(P3_EAX_REG_15__SCAN_IN), .A2(n16867), .ZN(n16863) );
  INV_X1 U19969 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n16991) );
  INV_X1 U19970 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n16985) );
  INV_X1 U19971 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n16983) );
  INV_X1 U19972 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n16981) );
  NOR4_X1 U19973 ( .A1(n16991), .A2(n16985), .A3(n16983), .A4(n16981), .ZN(
        n16781) );
  NOR2_X1 U19974 ( .A1(P3_EAX_REG_31__SCAN_IN), .A2(n16790), .ZN(n16782) );
  OAI21_X1 U19975 ( .B1(n17780), .B2(n16825), .A(n16783), .ZN(P3_U2704) );
  INV_X1 U19976 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17007) );
  NOR2_X2 U19977 ( .A1(n16784), .A2(n16922), .ZN(n16857) );
  INV_X1 U19978 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n17770) );
  OAI22_X1 U19979 ( .A1(n16785), .A2(n16924), .B1(n17770), .B2(n16825), .ZN(
        n16786) );
  AOI21_X1 U19980 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n16857), .A(n16786), .ZN(
        n16787) );
  OAI221_X1 U19981 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n16790), .C1(n17007), 
        .C2(n16788), .A(n16787), .ZN(P3_U2705) );
  INV_X1 U19982 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n17765) );
  AOI22_X1 U19983 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n16857), .B1(n16789), .B2(
        n16931), .ZN(n16793) );
  OAI211_X1 U19984 ( .C1(n16791), .C2(P3_EAX_REG_29__SCAN_IN), .A(n16922), .B(
        n16790), .ZN(n16792) );
  OAI211_X1 U19985 ( .C1(n16825), .C2(n17765), .A(n16793), .B(n16792), .ZN(
        P3_U2706) );
  INV_X1 U19986 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n17759) );
  AOI22_X1 U19987 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n16857), .B1(n16794), .B2(
        n16931), .ZN(n16797) );
  OAI211_X1 U19988 ( .C1(n16798), .C2(P3_EAX_REG_28__SCAN_IN), .A(n16922), .B(
        n16795), .ZN(n16796) );
  OAI211_X1 U19989 ( .C1(n16825), .C2(n17759), .A(n16797), .B(n16796), .ZN(
        P3_U2707) );
  AOI22_X1 U19990 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n16857), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16856), .ZN(n16801) );
  AOI211_X1 U19991 ( .C1(n17001), .C2(n16804), .A(n16798), .B(n16868), .ZN(
        n16799) );
  INV_X1 U19992 ( .A(n16799), .ZN(n16800) );
  OAI211_X1 U19993 ( .C1(n16924), .C2(n16802), .A(n16801), .B(n16800), .ZN(
        P3_U2708) );
  INV_X1 U19994 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n17747) );
  AOI22_X1 U19995 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n16857), .B1(n16803), .B2(
        n16931), .ZN(n16806) );
  OAI211_X1 U19996 ( .C1(n16807), .C2(P3_EAX_REG_26__SCAN_IN), .A(n16922), .B(
        n16804), .ZN(n16805) );
  OAI211_X1 U19997 ( .C1(n16825), .C2(n17747), .A(n16806), .B(n16805), .ZN(
        P3_U2709) );
  AOI22_X1 U19998 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n16857), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16856), .ZN(n16810) );
  AOI211_X1 U19999 ( .C1(n16997), .C2(n16813), .A(n16807), .B(n16868), .ZN(
        n16808) );
  INV_X1 U20000 ( .A(n16808), .ZN(n16809) );
  OAI211_X1 U20001 ( .C1(n16924), .C2(n16811), .A(n16810), .B(n16809), .ZN(
        P3_U2710) );
  AOI22_X1 U20002 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n16857), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16856), .ZN(n16816) );
  OAI21_X1 U20003 ( .B1(n16995), .B2(n16868), .A(n16812), .ZN(n16814) );
  NAND2_X1 U20004 ( .A1(n16814), .A2(n16813), .ZN(n16815) );
  OAI211_X1 U20005 ( .C1(n16924), .C2(n16817), .A(n16816), .B(n16815), .ZN(
        P3_U2711) );
  AOI211_X1 U20006 ( .C1(n16993), .C2(n16819), .A(n16868), .B(n16818), .ZN(
        n16820) );
  AOI21_X1 U20007 ( .B1(n16856), .B2(BUF2_REG_23__SCAN_IN), .A(n16820), .ZN(
        n16822) );
  NAND2_X1 U20008 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n16857), .ZN(n16821) );
  OAI211_X1 U20009 ( .C1(n16924), .C2(n16823), .A(n16822), .B(n16821), .ZN(
        P3_U2712) );
  NAND2_X1 U20010 ( .A1(n17778), .A2(n16858), .ZN(n16849) );
  NAND2_X1 U20011 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n16850), .ZN(n16845) );
  NAND3_X1 U20012 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .A3(n16840), .ZN(n16830) );
  INV_X1 U20013 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n18916) );
  OAI22_X1 U20014 ( .A1(n18916), .A2(n16825), .B1(n16924), .B2(n16824), .ZN(
        n16826) );
  INV_X1 U20015 ( .A(n16826), .ZN(n16829) );
  NAND2_X1 U20016 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n16840), .ZN(n16836) );
  NAND2_X1 U20017 ( .A1(n16922), .A2(n16836), .ZN(n16832) );
  OAI21_X1 U20018 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n16928), .A(n16832), .ZN(
        n16827) );
  AOI22_X1 U20019 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n16857), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n16827), .ZN(n16828) );
  OAI211_X1 U20020 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n16830), .A(n16829), .B(
        n16828), .ZN(P3_U2713) );
  AOI22_X1 U20021 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n16856), .B1(n16931), .B2(
        n16831), .ZN(n16835) );
  INV_X1 U20022 ( .A(n16832), .ZN(n16833) );
  AOI22_X1 U20023 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n16857), .B1(
        P3_EAX_REG_21__SCAN_IN), .B2(n16833), .ZN(n16834) );
  OAI211_X1 U20024 ( .C1(P3_EAX_REG_21__SCAN_IN), .C2(n16836), .A(n16835), .B(
        n16834), .ZN(P3_U2714) );
  AOI22_X1 U20025 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n16857), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16856), .ZN(n16838) );
  OAI211_X1 U20026 ( .C1(n16840), .C2(P3_EAX_REG_20__SCAN_IN), .A(n16922), .B(
        n16836), .ZN(n16837) );
  OAI211_X1 U20027 ( .C1(n16839), .C2(n16924), .A(n16838), .B(n16837), .ZN(
        P3_U2715) );
  AOI22_X1 U20028 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n16857), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16856), .ZN(n16843) );
  AOI211_X1 U20029 ( .C1(n16985), .C2(n16845), .A(n16840), .B(n16868), .ZN(
        n16841) );
  INV_X1 U20030 ( .A(n16841), .ZN(n16842) );
  OAI211_X1 U20031 ( .C1(n16844), .C2(n16924), .A(n16843), .B(n16842), .ZN(
        P3_U2716) );
  AOI22_X1 U20032 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n16857), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16856), .ZN(n16847) );
  OAI211_X1 U20033 ( .C1(n16850), .C2(P3_EAX_REG_18__SCAN_IN), .A(n16922), .B(
        n16845), .ZN(n16846) );
  OAI211_X1 U20034 ( .C1(n16848), .C2(n16924), .A(n16847), .B(n16846), .ZN(
        P3_U2717) );
  AOI22_X1 U20035 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n16857), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16856), .ZN(n16854) );
  OAI21_X1 U20036 ( .B1(n16981), .B2(n16868), .A(n16849), .ZN(n16852) );
  INV_X1 U20037 ( .A(n16850), .ZN(n16851) );
  NAND2_X1 U20038 ( .A1(n16852), .A2(n16851), .ZN(n16853) );
  OAI211_X1 U20039 ( .C1(n16855), .C2(n16924), .A(n16854), .B(n16853), .ZN(
        P3_U2718) );
  AOI22_X1 U20040 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n16857), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16856), .ZN(n16861) );
  AOI211_X1 U20041 ( .C1(n16979), .C2(n16863), .A(n16868), .B(n16858), .ZN(
        n16859) );
  INV_X1 U20042 ( .A(n16859), .ZN(n16860) );
  OAI211_X1 U20043 ( .C1(n16862), .C2(n16924), .A(n16861), .B(n16860), .ZN(
        P3_U2719) );
  OAI211_X1 U20044 ( .C1(P3_EAX_REG_15__SCAN_IN), .C2(n16867), .A(n16922), .B(
        n16863), .ZN(n16865) );
  NAND2_X1 U20045 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n16932), .ZN(n16864) );
  OAI211_X1 U20046 ( .C1(n16866), .C2(n16924), .A(n16865), .B(n16864), .ZN(
        P3_U2720) );
  INV_X1 U20047 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17034) );
  INV_X1 U20048 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17025) );
  NOR3_X1 U20049 ( .A1(n16890), .A2(n16896), .A3(n17025), .ZN(n16894) );
  NAND2_X1 U20050 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n16894), .ZN(n16885) );
  NOR2_X1 U20051 ( .A1(n17029), .A2(n16885), .ZN(n16877) );
  NAND2_X1 U20052 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n16877), .ZN(n16872) );
  NOR2_X1 U20053 ( .A1(n17034), .A2(n16872), .ZN(n16875) );
  INV_X1 U20054 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17036) );
  AOI22_X1 U20055 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n16932), .B1(n16875), .B2(
        n17036), .ZN(n16870) );
  OR3_X1 U20056 ( .A1(n17036), .A2(n16868), .A3(n16867), .ZN(n16869) );
  OAI211_X1 U20057 ( .C1(n16871), .C2(n16924), .A(n16870), .B(n16869), .ZN(
        P3_U2721) );
  INV_X1 U20058 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n16876) );
  INV_X1 U20059 ( .A(n16872), .ZN(n16880) );
  AOI21_X1 U20060 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n16922), .A(n16880), .ZN(
        n16874) );
  OAI222_X1 U20061 ( .A1(n16927), .A2(n16876), .B1(n16875), .B2(n16874), .C1(
        n16924), .C2(n16873), .ZN(P3_U2722) );
  INV_X1 U20062 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n16881) );
  AOI21_X1 U20063 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n16922), .A(n16877), .ZN(
        n16879) );
  OAI222_X1 U20064 ( .A1(n16927), .A2(n16881), .B1(n16880), .B2(n16879), .C1(
        n16924), .C2(n16878), .ZN(P3_U2723) );
  NAND2_X1 U20065 ( .A1(n16922), .A2(n16885), .ZN(n16888) );
  INV_X1 U20066 ( .A(n16882), .ZN(n16883) );
  AOI22_X1 U20067 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n16932), .B1(n16931), .B2(
        n16883), .ZN(n16884) );
  OAI221_X1 U20068 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n16885), .C1(n17029), 
        .C2(n16888), .A(n16884), .ZN(P3_U2724) );
  INV_X1 U20069 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n16889) );
  NOR2_X1 U20070 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n16894), .ZN(n16887) );
  OAI222_X1 U20071 ( .A1(n16927), .A2(n16889), .B1(n16888), .B2(n16887), .C1(
        n16924), .C2(n16886), .ZN(P3_U2725) );
  INV_X1 U20072 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n16895) );
  NOR2_X1 U20073 ( .A1(n16890), .A2(n16896), .ZN(n16891) );
  AOI21_X1 U20074 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n16922), .A(n16891), .ZN(
        n16893) );
  OAI222_X1 U20075 ( .A1(n16927), .A2(n16895), .B1(n16894), .B2(n16893), .C1(
        n16924), .C2(n16892), .ZN(P3_U2726) );
  NAND2_X1 U20076 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n16932), .ZN(n16899) );
  OAI211_X1 U20077 ( .C1(P3_EAX_REG_8__SCAN_IN), .C2(n16897), .A(n16922), .B(
        n16896), .ZN(n16898) );
  OAI211_X1 U20078 ( .C1(n16900), .C2(n16924), .A(n16899), .B(n16898), .ZN(
        P3_U2727) );
  INV_X1 U20079 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n20610) );
  INV_X1 U20080 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17017) );
  INV_X1 U20081 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17013) );
  NOR4_X1 U20082 ( .A1(n17013), .A2(n17011), .A3(n17009), .A4(n16928), .ZN(
        n16926) );
  NAND2_X1 U20083 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n16926), .ZN(n16913) );
  NOR2_X1 U20084 ( .A1(n17017), .A2(n16913), .ZN(n16917) );
  NAND2_X1 U20085 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n16917), .ZN(n16905) );
  NOR2_X1 U20086 ( .A1(n20610), .A2(n16905), .ZN(n16909) );
  AOI21_X1 U20087 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n16922), .A(n16909), .ZN(
        n16904) );
  NOR2_X1 U20088 ( .A1(n16901), .A2(n16928), .ZN(n16903) );
  OAI222_X1 U20089 ( .A1(n17776), .A2(n16927), .B1(n16904), .B2(n16903), .C1(
        n16924), .C2(n16902), .ZN(P3_U2728) );
  INV_X1 U20090 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n17771) );
  INV_X1 U20091 ( .A(n16905), .ZN(n16912) );
  AOI21_X1 U20092 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n16922), .A(n16912), .ZN(
        n16908) );
  INV_X1 U20093 ( .A(n16906), .ZN(n16907) );
  OAI222_X1 U20094 ( .A1(n17771), .A2(n16927), .B1(n16909), .B2(n16908), .C1(
        n16924), .C2(n16907), .ZN(P3_U2729) );
  AOI21_X1 U20095 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n16922), .A(n16917), .ZN(
        n16911) );
  OAI222_X1 U20096 ( .A1(n17764), .A2(n16927), .B1(n16912), .B2(n16911), .C1(
        n16924), .C2(n16910), .ZN(P3_U2730) );
  INV_X1 U20097 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n17758) );
  INV_X1 U20098 ( .A(n16913), .ZN(n16920) );
  AOI21_X1 U20099 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n16922), .A(n16920), .ZN(
        n16916) );
  INV_X1 U20100 ( .A(n16914), .ZN(n16915) );
  OAI222_X1 U20101 ( .A1(n17758), .A2(n16927), .B1(n16917), .B2(n16916), .C1(
        n16924), .C2(n16915), .ZN(P3_U2731) );
  INV_X1 U20102 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n17752) );
  AOI21_X1 U20103 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n16922), .A(n16926), .ZN(
        n16919) );
  OAI222_X1 U20104 ( .A1(n17752), .A2(n16927), .B1(n16920), .B2(n16919), .C1(
        n16924), .C2(n16918), .ZN(P3_U2732) );
  INV_X1 U20105 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n17746) );
  NOR3_X1 U20106 ( .A1(n17011), .A2(n17009), .A3(n16928), .ZN(n16921) );
  AOI21_X1 U20107 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n16922), .A(n16921), .ZN(
        n16925) );
  OAI222_X1 U20108 ( .A1(n17746), .A2(n16927), .B1(n16926), .B2(n16925), .C1(
        n16924), .C2(n16923), .ZN(P3_U2733) );
  OR2_X1 U20109 ( .A1(n17009), .A2(n16928), .ZN(n16935) );
  AOI21_X1 U20110 ( .B1(n17778), .B2(n17009), .A(n16929), .ZN(n16934) );
  AOI22_X1 U20111 ( .A1(n16932), .A2(BUF2_REG_1__SCAN_IN), .B1(n16931), .B2(
        n16930), .ZN(n16933) );
  OAI221_X1 U20112 ( .B1(P3_EAX_REG_1__SCAN_IN), .B2(n16935), .C1(n17011), 
        .C2(n16934), .A(n16933), .ZN(P3_U2734) );
  AND2_X1 U20113 ( .A1(n16963), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NAND2_X1 U20114 ( .A1(n16953), .A2(n17736), .ZN(n16952) );
  AOI22_X1 U20115 ( .A1(n18386), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n16970), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n16937) );
  OAI21_X1 U20116 ( .B1(n17007), .B2(n16952), .A(n16937), .ZN(P3_U2737) );
  INV_X1 U20117 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17005) );
  AOI22_X1 U20118 ( .A1(n18386), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n16970), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n16938) );
  OAI21_X1 U20119 ( .B1(n17005), .B2(n16952), .A(n16938), .ZN(P3_U2738) );
  INV_X1 U20120 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17003) );
  AOI22_X1 U20121 ( .A1(n18386), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n16970), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n16939) );
  OAI21_X1 U20122 ( .B1(n17003), .B2(n16952), .A(n16939), .ZN(P3_U2739) );
  AOI22_X1 U20123 ( .A1(n18386), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n16963), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n16940) );
  OAI21_X1 U20124 ( .B1(n17001), .B2(n16952), .A(n16940), .ZN(P3_U2740) );
  INV_X1 U20125 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n16999) );
  AOI22_X1 U20126 ( .A1(n18386), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n16963), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n16941) );
  OAI21_X1 U20127 ( .B1(n16999), .B2(n16952), .A(n16941), .ZN(P3_U2741) );
  AOI22_X1 U20128 ( .A1(n18386), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n16963), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n16942) );
  OAI21_X1 U20129 ( .B1(n16997), .B2(n16952), .A(n16942), .ZN(P3_U2742) );
  AOI22_X1 U20130 ( .A1(n18386), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n16963), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n16943) );
  OAI21_X1 U20131 ( .B1(n16995), .B2(n16952), .A(n16943), .ZN(P3_U2743) );
  CLKBUF_X1 U20132 ( .A(n18386), .Z(n16971) );
  AOI22_X1 U20133 ( .A1(n16971), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n16970), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n16944) );
  OAI21_X1 U20134 ( .B1(n16993), .B2(n16952), .A(n16944), .ZN(P3_U2744) );
  AOI22_X1 U20135 ( .A1(n16971), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n16970), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n16945) );
  OAI21_X1 U20136 ( .B1(n16991), .B2(n16952), .A(n16945), .ZN(P3_U2745) );
  INV_X1 U20137 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n16989) );
  AOI22_X1 U20138 ( .A1(n16971), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n16970), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n16946) );
  OAI21_X1 U20139 ( .B1(n16989), .B2(n16952), .A(n16946), .ZN(P3_U2746) );
  INV_X1 U20140 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n16987) );
  AOI22_X1 U20141 ( .A1(n16971), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n16970), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n16947) );
  OAI21_X1 U20142 ( .B1(n16987), .B2(n16952), .A(n16947), .ZN(P3_U2747) );
  AOI22_X1 U20143 ( .A1(n16971), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n16970), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n16948) );
  OAI21_X1 U20144 ( .B1(n16985), .B2(n16952), .A(n16948), .ZN(P3_U2748) );
  AOI22_X1 U20145 ( .A1(n16971), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n16970), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n16949) );
  OAI21_X1 U20146 ( .B1(n16983), .B2(n16952), .A(n16949), .ZN(P3_U2749) );
  AOI22_X1 U20147 ( .A1(n16971), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n16970), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n16950) );
  OAI21_X1 U20148 ( .B1(n16981), .B2(n16952), .A(n16950), .ZN(P3_U2750) );
  AOI22_X1 U20149 ( .A1(n16971), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n16970), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n16951) );
  OAI21_X1 U20150 ( .B1(n16979), .B2(n16952), .A(n16951), .ZN(P3_U2751) );
  INV_X1 U20151 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17041) );
  AOI22_X1 U20152 ( .A1(n16971), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n16970), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n16954) );
  OAI21_X1 U20153 ( .B1(n17041), .B2(n16973), .A(n16954), .ZN(P3_U2752) );
  AOI22_X1 U20154 ( .A1(n16971), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n16970), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n16955) );
  OAI21_X1 U20155 ( .B1(n17036), .B2(n16973), .A(n16955), .ZN(P3_U2753) );
  AOI22_X1 U20156 ( .A1(n16971), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n16970), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n16956) );
  OAI21_X1 U20157 ( .B1(n17034), .B2(n16973), .A(n16956), .ZN(P3_U2754) );
  AOI22_X1 U20158 ( .A1(n16971), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n16970), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n16957) );
  OAI21_X1 U20159 ( .B1(n17032), .B2(n16973), .A(n16957), .ZN(P3_U2755) );
  AOI22_X1 U20160 ( .A1(n16971), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n16963), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n16958) );
  OAI21_X1 U20161 ( .B1(n17029), .B2(n16973), .A(n16958), .ZN(P3_U2756) );
  INV_X1 U20162 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17027) );
  AOI22_X1 U20163 ( .A1(n16971), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n16963), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n16959) );
  OAI21_X1 U20164 ( .B1(n17027), .B2(n16973), .A(n16959), .ZN(P3_U2757) );
  AOI22_X1 U20165 ( .A1(n16971), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n16963), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n16960) );
  OAI21_X1 U20166 ( .B1(n17025), .B2(n16973), .A(n16960), .ZN(P3_U2758) );
  INV_X1 U20167 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n20659) );
  AOI22_X1 U20168 ( .A1(n16971), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n16963), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n16961) );
  OAI21_X1 U20169 ( .B1(n20659), .B2(n16973), .A(n16961), .ZN(P3_U2759) );
  INV_X1 U20170 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17022) );
  AOI22_X1 U20171 ( .A1(n16971), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n16963), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n16962) );
  OAI21_X1 U20172 ( .B1(n17022), .B2(n16973), .A(n16962), .ZN(P3_U2760) );
  AOI22_X1 U20173 ( .A1(n16971), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n16963), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n16964) );
  OAI21_X1 U20174 ( .B1(n20610), .B2(n16973), .A(n16964), .ZN(P3_U2761) );
  INV_X1 U20175 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17019) );
  AOI22_X1 U20176 ( .A1(n16971), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n16970), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n16965) );
  OAI21_X1 U20177 ( .B1(n17019), .B2(n16973), .A(n16965), .ZN(P3_U2762) );
  AOI22_X1 U20178 ( .A1(n16971), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n16970), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n16966) );
  OAI21_X1 U20179 ( .B1(n17017), .B2(n16973), .A(n16966), .ZN(P3_U2763) );
  INV_X1 U20180 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17015) );
  AOI22_X1 U20181 ( .A1(n16971), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n16970), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n16967) );
  OAI21_X1 U20182 ( .B1(n17015), .B2(n16973), .A(n16967), .ZN(P3_U2764) );
  AOI22_X1 U20183 ( .A1(n16971), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n16970), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n16968) );
  OAI21_X1 U20184 ( .B1(n17013), .B2(n16973), .A(n16968), .ZN(P3_U2765) );
  AOI22_X1 U20185 ( .A1(n16971), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n16970), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n16969) );
  OAI21_X1 U20186 ( .B1(n17011), .B2(n16973), .A(n16969), .ZN(P3_U2766) );
  AOI22_X1 U20187 ( .A1(n16971), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n16970), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n16972) );
  OAI21_X1 U20188 ( .B1(n17009), .B2(n16973), .A(n16972), .ZN(P3_U2767) );
  NOR2_X1 U20189 ( .A1(n18391), .A2(n16976), .ZN(n18234) );
  INV_X1 U20190 ( .A(n18385), .ZN(n18392) );
  AOI211_X1 U20191 ( .C1(n18391), .C2(n18392), .A(n16976), .B(n16975), .ZN(
        n16977) );
  AOI22_X1 U20192 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17038), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17037), .ZN(n16978) );
  OAI21_X1 U20193 ( .B1(n16979), .B2(n17040), .A(n16978), .ZN(P3_U2768) );
  AOI22_X1 U20194 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17038), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17037), .ZN(n16980) );
  OAI21_X1 U20195 ( .B1(n16981), .B2(n17040), .A(n16980), .ZN(P3_U2769) );
  AOI22_X1 U20196 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17038), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17037), .ZN(n16982) );
  OAI21_X1 U20197 ( .B1(n16983), .B2(n17040), .A(n16982), .ZN(P3_U2770) );
  AOI22_X1 U20198 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17030), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17037), .ZN(n16984) );
  OAI21_X1 U20199 ( .B1(n16985), .B2(n17040), .A(n16984), .ZN(P3_U2771) );
  AOI22_X1 U20200 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17030), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17037), .ZN(n16986) );
  OAI21_X1 U20201 ( .B1(n16987), .B2(n17040), .A(n16986), .ZN(P3_U2772) );
  AOI22_X1 U20202 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17030), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17037), .ZN(n16988) );
  OAI21_X1 U20203 ( .B1(n16989), .B2(n17040), .A(n16988), .ZN(P3_U2773) );
  AOI22_X1 U20204 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17030), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17037), .ZN(n16990) );
  OAI21_X1 U20205 ( .B1(n16991), .B2(n17040), .A(n16990), .ZN(P3_U2774) );
  AOI22_X1 U20206 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17030), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17037), .ZN(n16992) );
  OAI21_X1 U20207 ( .B1(n16993), .B2(n17040), .A(n16992), .ZN(P3_U2775) );
  AOI22_X1 U20208 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17030), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17037), .ZN(n16994) );
  OAI21_X1 U20209 ( .B1(n16995), .B2(n17040), .A(n16994), .ZN(P3_U2776) );
  AOI22_X1 U20210 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17030), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17037), .ZN(n16996) );
  OAI21_X1 U20211 ( .B1(n16997), .B2(n17040), .A(n16996), .ZN(P3_U2777) );
  AOI22_X1 U20212 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17030), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17037), .ZN(n16998) );
  OAI21_X1 U20213 ( .B1(n16999), .B2(n17040), .A(n16998), .ZN(P3_U2778) );
  AOI22_X1 U20214 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17030), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17037), .ZN(n17000) );
  OAI21_X1 U20215 ( .B1(n17001), .B2(n17040), .A(n17000), .ZN(P3_U2779) );
  AOI22_X1 U20216 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17038), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17037), .ZN(n17002) );
  OAI21_X1 U20217 ( .B1(n17003), .B2(n17040), .A(n17002), .ZN(P3_U2780) );
  AOI22_X1 U20218 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17038), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17037), .ZN(n17004) );
  OAI21_X1 U20219 ( .B1(n17005), .B2(n17040), .A(n17004), .ZN(P3_U2781) );
  AOI22_X1 U20220 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17038), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17037), .ZN(n17006) );
  OAI21_X1 U20221 ( .B1(n17007), .B2(n17040), .A(n17006), .ZN(P3_U2782) );
  AOI22_X1 U20222 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17038), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17037), .ZN(n17008) );
  OAI21_X1 U20223 ( .B1(n17009), .B2(n17040), .A(n17008), .ZN(P3_U2783) );
  AOI22_X1 U20224 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17038), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17037), .ZN(n17010) );
  OAI21_X1 U20225 ( .B1(n17011), .B2(n17040), .A(n17010), .ZN(P3_U2784) );
  AOI22_X1 U20226 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17038), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17037), .ZN(n17012) );
  OAI21_X1 U20227 ( .B1(n17013), .B2(n17040), .A(n17012), .ZN(P3_U2785) );
  AOI22_X1 U20228 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17038), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17037), .ZN(n17014) );
  OAI21_X1 U20229 ( .B1(n17015), .B2(n17040), .A(n17014), .ZN(P3_U2786) );
  AOI22_X1 U20230 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17038), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17037), .ZN(n17016) );
  OAI21_X1 U20231 ( .B1(n17017), .B2(n17040), .A(n17016), .ZN(P3_U2787) );
  AOI22_X1 U20232 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17038), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17037), .ZN(n17018) );
  OAI21_X1 U20233 ( .B1(n17019), .B2(n17040), .A(n17018), .ZN(P3_U2788) );
  AOI22_X1 U20234 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17038), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17037), .ZN(n17020) );
  OAI21_X1 U20235 ( .B1(n20610), .B2(n17040), .A(n17020), .ZN(P3_U2789) );
  AOI22_X1 U20236 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17038), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17037), .ZN(n17021) );
  OAI21_X1 U20237 ( .B1(n17022), .B2(n17040), .A(n17021), .ZN(P3_U2790) );
  AOI22_X1 U20238 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17038), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17037), .ZN(n17023) );
  OAI21_X1 U20239 ( .B1(n20659), .B2(n17040), .A(n17023), .ZN(P3_U2791) );
  AOI22_X1 U20240 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17038), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17037), .ZN(n17024) );
  OAI21_X1 U20241 ( .B1(n17025), .B2(n17040), .A(n17024), .ZN(P3_U2792) );
  AOI22_X1 U20242 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17030), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17037), .ZN(n17026) );
  OAI21_X1 U20243 ( .B1(n17027), .B2(n17040), .A(n17026), .ZN(P3_U2793) );
  AOI22_X1 U20244 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17038), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17037), .ZN(n17028) );
  OAI21_X1 U20245 ( .B1(n17029), .B2(n17040), .A(n17028), .ZN(P3_U2794) );
  AOI22_X1 U20246 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17030), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17037), .ZN(n17031) );
  OAI21_X1 U20247 ( .B1(n17032), .B2(n17040), .A(n17031), .ZN(P3_U2795) );
  AOI22_X1 U20248 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17038), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17037), .ZN(n17033) );
  OAI21_X1 U20249 ( .B1(n17034), .B2(n17040), .A(n17033), .ZN(P3_U2796) );
  AOI22_X1 U20250 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17038), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17037), .ZN(n17035) );
  OAI21_X1 U20251 ( .B1(n17036), .B2(n17040), .A(n17035), .ZN(P3_U2797) );
  AOI22_X1 U20252 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17038), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17037), .ZN(n17039) );
  OAI21_X1 U20253 ( .B1(n17041), .B2(n17040), .A(n17039), .ZN(P3_U2798) );
  INV_X1 U20254 ( .A(n17309), .ZN(n17240) );
  NAND2_X1 U20255 ( .A1(n17412), .A2(n17240), .ZN(n17132) );
  INV_X1 U20256 ( .A(n17132), .ZN(n17160) );
  INV_X1 U20257 ( .A(n17042), .ZN(n17414) );
  AOI22_X1 U20258 ( .A1(n17401), .A2(n17415), .B1(n17309), .B2(n17414), .ZN(
        n17080) );
  NAND2_X1 U20259 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17080), .ZN(
        n17066) );
  NAND2_X1 U20260 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17066), .ZN(
        n17058) );
  NAND4_X1 U20261 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n9765), .A3(
        n17083), .A4(n17261), .ZN(n17063) );
  OAI21_X1 U20262 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17043), .ZN(n17049) );
  INV_X1 U20263 ( .A(n18255), .ZN(n17204) );
  INV_X1 U20264 ( .A(n17044), .ZN(n17311) );
  OAI21_X1 U20265 ( .B1(n9766), .B2(n17311), .A(n17408), .ZN(n17045) );
  AOI21_X1 U20266 ( .B1(n17204), .B2(n17046), .A(n17045), .ZN(n17071) );
  OAI21_X1 U20267 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17070), .A(
        n17071), .ZN(n17059) );
  AOI22_X1 U20268 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17059), .B1(
        n17258), .B2(n17047), .ZN(n17048) );
  OAI21_X1 U20269 ( .B1(n17063), .B2(n17049), .A(n17048), .ZN(n17050) );
  AOI211_X1 U20270 ( .C1(n17052), .C2(n17119), .A(n17051), .B(n17050), .ZN(
        n17057) );
  OAI211_X1 U20271 ( .C1(n17055), .C2(n17054), .A(n17293), .B(n17053), .ZN(
        n17056) );
  OAI211_X1 U20272 ( .C1(n17160), .C2(n17058), .A(n17057), .B(n17056), .ZN(
        P3_U2802) );
  AOI22_X1 U20273 ( .A1(n17715), .A2(P3_REIP_REG_27__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n17059), .ZN(n17068) );
  NOR2_X1 U20274 ( .A1(n17413), .A2(n17108), .ZN(n17065) );
  NOR2_X1 U20275 ( .A1(n17061), .A2(n17060), .ZN(n17062) );
  XOR2_X1 U20276 ( .A(n17062), .B(n17318), .Z(n17421) );
  OAI22_X1 U20277 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17063), .B1(
        n17421), .B2(n17322), .ZN(n17064) );
  AOI221_X1 U20278 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17066), 
        .C1(n17065), .C2(n17066), .A(n17064), .ZN(n17067) );
  OAI211_X1 U20279 ( .C1(n17247), .C2(n17069), .A(n17068), .B(n17067), .ZN(
        P3_U2803) );
  NAND2_X1 U20280 ( .A1(n17247), .A2(n17070), .ZN(n17185) );
  NAND3_X1 U20281 ( .A1(n9765), .A2(n17083), .A3(n18121), .ZN(n17072) );
  AOI21_X1 U20282 ( .B1(n10109), .B2(n17072), .A(n17071), .ZN(n17074) );
  NAND2_X1 U20283 ( .A1(n17715), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17426) );
  INV_X1 U20284 ( .A(n17426), .ZN(n17073) );
  AOI211_X1 U20285 ( .C1(n17075), .C2(n17185), .A(n17074), .B(n17073), .ZN(
        n17079) );
  OAI21_X1 U20286 ( .B1(n17077), .B2(n17418), .A(n17076), .ZN(n17423) );
  NOR3_X1 U20287 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17435), .A3(
        n17431), .ZN(n17422) );
  AOI22_X1 U20288 ( .A1(n17293), .A2(n17423), .B1(n17119), .B2(n17422), .ZN(
        n17078) );
  OAI211_X1 U20289 ( .C1(n17080), .C2(n17418), .A(n17079), .B(n17078), .ZN(
        P3_U2804) );
  OAI21_X1 U20290 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17082), .A(
        n17081), .ZN(n17442) );
  NAND2_X1 U20291 ( .A1(n9765), .A2(n17261), .ZN(n17099) );
  AOI211_X1 U20292 ( .C1(n17098), .C2(n17086), .A(n17083), .B(n17099), .ZN(
        n17088) );
  OR2_X1 U20293 ( .A1(n18090), .A2(n9765), .ZN(n17116) );
  OAI211_X1 U20294 ( .C1(n17084), .C2(n18255), .A(n17408), .B(n17116), .ZN(
        n17113) );
  AOI21_X1 U20295 ( .B1(n17154), .B2(n17085), .A(n17113), .ZN(n17097) );
  OAI22_X1 U20296 ( .A1(n17097), .A2(n17086), .B1(n9746), .B2(n18314), .ZN(
        n17087) );
  AOI211_X1 U20297 ( .C1(n17089), .C2(n17258), .A(n17088), .B(n17087), .ZN(
        n17096) );
  AOI21_X1 U20298 ( .B1(n17435), .B2(n17091), .A(n17090), .ZN(n17439) );
  AOI21_X1 U20299 ( .B1(n17318), .B2(n17093), .A(n17092), .ZN(n17094) );
  XOR2_X1 U20300 ( .A(n17094), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17438) );
  AOI22_X1 U20301 ( .A1(n17401), .A2(n17439), .B1(n17293), .B2(n17438), .ZN(
        n17095) );
  OAI211_X1 U20302 ( .C1(n17240), .C2(n17442), .A(n17096), .B(n17095), .ZN(
        P3_U2805) );
  NOR2_X1 U20303 ( .A1(n17451), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17443) );
  INV_X1 U20304 ( .A(n17443), .ZN(n17107) );
  NAND2_X1 U20305 ( .A1(n17715), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n17456) );
  OAI221_X1 U20306 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n17099), .C1(
        n17098), .C2(n17097), .A(n17456), .ZN(n17100) );
  AOI21_X1 U20307 ( .B1(n17258), .B2(n17101), .A(n17100), .ZN(n17106) );
  OAI22_X1 U20308 ( .A1(n17450), .A2(n17412), .B1(n15358), .B2(n17240), .ZN(
        n17118) );
  OAI21_X1 U20309 ( .B1(n17104), .B2(n17103), .A(n17102), .ZN(n17445) );
  AOI22_X1 U20310 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17118), .B1(
        n17293), .B2(n17445), .ZN(n17105) );
  OAI211_X1 U20311 ( .C1(n17108), .C2(n17107), .A(n17106), .B(n17105), .ZN(
        P3_U2806) );
  OAI22_X1 U20312 ( .A1(n17318), .A2(n17480), .B1(n17127), .B2(n17109), .ZN(
        n17110) );
  NOR2_X1 U20313 ( .A1(n17110), .A2(n17150), .ZN(n17111) );
  XOR2_X1 U20314 ( .A(n17111), .B(n17451), .Z(n17463) );
  AOI22_X1 U20315 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17113), .B1(
        n17112), .B2(n17185), .ZN(n17114) );
  NAND2_X1 U20316 ( .A1(n17715), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17462) );
  OAI211_X1 U20317 ( .C1(n17116), .C2(n17115), .A(n17114), .B(n17462), .ZN(
        n17117) );
  AOI221_X1 U20318 ( .B1(n17119), .B2(n17451), .C1(n17118), .C2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n17117), .ZN(n17120) );
  OAI21_X1 U20319 ( .B1(n17322), .B2(n17463), .A(n17120), .ZN(P3_U2807) );
  INV_X1 U20320 ( .A(n17121), .ZN(n17122) );
  NAND2_X1 U20321 ( .A1(n17204), .A2(n17122), .ZN(n17123) );
  OAI211_X1 U20322 ( .C1(n17124), .C2(n17311), .A(n17408), .B(n17123), .ZN(
        n17158) );
  AOI21_X1 U20323 ( .B1(n17154), .B2(n17152), .A(n17158), .ZN(n17139) );
  INV_X1 U20324 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18308) );
  NOR2_X1 U20325 ( .A1(n9746), .A2(n18308), .ZN(n17464) );
  NAND2_X1 U20326 ( .A1(n17124), .A2(n17261), .ZN(n17141) );
  AOI221_X1 U20327 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C1(n17140), .C2(n17138), .A(
        n17141), .ZN(n17125) );
  AOI211_X1 U20328 ( .C1(n17126), .C2(n17258), .A(n17464), .B(n17125), .ZN(
        n17137) );
  INV_X1 U20329 ( .A(n17127), .ZN(n17128) );
  AOI21_X1 U20330 ( .B1(n17129), .B2(n17128), .A(n17150), .ZN(n17130) );
  XOR2_X1 U20331 ( .A(n17130), .B(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(
        n17465) );
  INV_X1 U20332 ( .A(n17195), .ZN(n17212) );
  NOR2_X1 U20333 ( .A1(n17473), .A2(n17212), .ZN(n17134) );
  NAND2_X1 U20334 ( .A1(n17401), .A2(n17131), .ZN(n17225) );
  OAI21_X1 U20335 ( .B1(n17541), .B2(n17240), .A(n17225), .ZN(n17159) );
  AOI21_X1 U20336 ( .B1(n17473), .B2(n17132), .A(n17159), .ZN(n17149) );
  INV_X1 U20337 ( .A(n17149), .ZN(n17133) );
  MUX2_X1 U20338 ( .A(n17134), .B(n17133), .S(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(n17135) );
  AOI21_X1 U20339 ( .B1(n17293), .B2(n17465), .A(n17135), .ZN(n17136) );
  OAI211_X1 U20340 ( .C1(n17139), .C2(n17138), .A(n17137), .B(n17136), .ZN(
        P3_U2808) );
  NAND2_X1 U20341 ( .A1(n17715), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n17488) );
  OAI221_X1 U20342 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n17141), .C1(
        n17140), .C2(n17139), .A(n17488), .ZN(n17142) );
  AOI21_X1 U20343 ( .B1(n17258), .B2(n17143), .A(n17142), .ZN(n17148) );
  OAI22_X1 U20344 ( .A1(n17482), .A2(n17163), .B1(n17145), .B2(n17182), .ZN(
        n17146) );
  XOR2_X1 U20345 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17146), .Z(
        n17487) );
  NOR2_X1 U20346 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17482), .ZN(
        n17486) );
  NOR2_X1 U20347 ( .A1(n17484), .A2(n17212), .ZN(n17171) );
  AOI22_X1 U20348 ( .A1(n17293), .A2(n17487), .B1(n17486), .B2(n17171), .ZN(
        n17147) );
  OAI211_X1 U20349 ( .C1(n17149), .C2(n17491), .A(n17148), .B(n17147), .ZN(
        P3_U2809) );
  INV_X1 U20350 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17502) );
  AOI221_X1 U20351 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17163), 
        .C1(n17502), .C2(n17179), .A(n17150), .ZN(n17151) );
  XOR2_X1 U20352 ( .A(n17474), .B(n17151), .Z(n17500) );
  OAI21_X1 U20353 ( .B1(n17153), .B2(n18090), .A(n17152), .ZN(n17157) );
  AOI21_X1 U20354 ( .B1(n17247), .B2(n17070), .A(n17155), .ZN(n17156) );
  NOR2_X1 U20355 ( .A1(n9746), .A2(n18305), .ZN(n17492) );
  AOI211_X1 U20356 ( .C1(n17158), .C2(n17157), .A(n17156), .B(n17492), .ZN(
        n17162) );
  NOR2_X1 U20357 ( .A1(n17484), .A2(n17502), .ZN(n17496) );
  INV_X1 U20358 ( .A(n17159), .ZN(n17211) );
  OAI21_X1 U20359 ( .B1(n17160), .B2(n17496), .A(n17211), .ZN(n17172) );
  NOR2_X1 U20360 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17502), .ZN(
        n17493) );
  AOI22_X1 U20361 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17172), .B1(
        n17171), .B2(n17493), .ZN(n17161) );
  OAI211_X1 U20362 ( .C1(n17322), .C2(n17500), .A(n17162), .B(n17161), .ZN(
        P3_U2810) );
  OAI21_X1 U20363 ( .B1(n17182), .B2(n17179), .A(n17163), .ZN(n17164) );
  XOR2_X1 U20364 ( .A(n17164), .B(n17502), .Z(n17506) );
  NOR2_X1 U20365 ( .A1(n9746), .A2(n18302), .ZN(n17501) );
  NOR2_X1 U20366 ( .A1(n20690), .A2(n17166), .ZN(n17168) );
  OAI211_X1 U20367 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n10281), .B(n17261), .ZN(n17167) );
  OAI21_X1 U20368 ( .B1(n10281), .B2(n17311), .A(n17408), .ZN(n17190) );
  AOI21_X1 U20369 ( .B1(n17204), .B2(n17165), .A(n17190), .ZN(n17175) );
  OAI22_X1 U20370 ( .A1(n17168), .A2(n17167), .B1(n17175), .B2(n17166), .ZN(
        n17169) );
  AOI211_X1 U20371 ( .C1(n17170), .C2(n17258), .A(n17501), .B(n17169), .ZN(
        n17174) );
  AOI22_X1 U20372 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17172), .B1(
        n17171), .B2(n17502), .ZN(n17173) );
  OAI211_X1 U20373 ( .C1(n17506), .C2(n17322), .A(n17174), .B(n17173), .ZN(
        P3_U2811) );
  NAND2_X1 U20374 ( .A1(n17513), .A2(n17180), .ZN(n17521) );
  NAND2_X1 U20375 ( .A1(n10281), .A2(n17261), .ZN(n17176) );
  NAND2_X1 U20376 ( .A1(n17715), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n17519) );
  OAI221_X1 U20377 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17176), .C1(
        n20690), .C2(n17175), .A(n17519), .ZN(n17177) );
  AOI21_X1 U20378 ( .B1(n17258), .B2(n17178), .A(n17177), .ZN(n17184) );
  OAI21_X1 U20379 ( .B1(n17513), .B2(n17212), .A(n17211), .ZN(n17194) );
  OAI21_X1 U20380 ( .B1(n17180), .B2(n17235), .A(n17179), .ZN(n17181) );
  XOR2_X1 U20381 ( .A(n17182), .B(n17181), .Z(n17517) );
  AOI22_X1 U20382 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17194), .B1(
        n17293), .B2(n17517), .ZN(n17183) );
  OAI211_X1 U20383 ( .C1(n17212), .C2(n17521), .A(n17184), .B(n17183), .ZN(
        P3_U2812) );
  INV_X1 U20384 ( .A(n17185), .ZN(n17393) );
  OAI21_X1 U20385 ( .B1(n17188), .B2(n18090), .A(n17187), .ZN(n17189) );
  AOI22_X1 U20386 ( .A1(n17191), .A2(n17185), .B1(n17190), .B2(n17189), .ZN(
        n17198) );
  OAI21_X1 U20387 ( .B1(n17193), .B2(n17522), .A(n17192), .ZN(n17525) );
  AOI22_X1 U20388 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17194), .B1(
        n17293), .B2(n17525), .ZN(n17197) );
  NAND3_X1 U20389 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17195), .A3(
        n17522), .ZN(n17196) );
  NAND2_X1 U20390 ( .A1(n17710), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n17526) );
  NAND4_X1 U20391 ( .A1(n17198), .A2(n17197), .A3(n17196), .A4(n17526), .ZN(
        P3_U2813) );
  AOI21_X1 U20392 ( .B1(n17318), .B2(n17200), .A(n17199), .ZN(n17201) );
  XOR2_X1 U20393 ( .A(n17201), .B(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .Z(
        n17536) );
  NAND2_X1 U20394 ( .A1(n17202), .A2(n17261), .ZN(n17215) );
  AOI221_X1 U20395 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C1(n17214), .C2(n17207), .A(
        n17215), .ZN(n17209) );
  OAI21_X1 U20396 ( .B1(n17202), .B2(n17311), .A(n17408), .ZN(n17231) );
  AOI21_X1 U20397 ( .B1(n17204), .B2(n17203), .A(n17231), .ZN(n17213) );
  AOI22_X1 U20398 ( .A1(n17715), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n17258), 
        .B2(n17205), .ZN(n17206) );
  OAI21_X1 U20399 ( .B1(n17213), .B2(n17207), .A(n17206), .ZN(n17208) );
  AOI211_X1 U20400 ( .C1(n17536), .C2(n17293), .A(n17209), .B(n17208), .ZN(
        n17210) );
  OAI221_X1 U20401 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17212), 
        .C1(n17539), .C2(n17211), .A(n17210), .ZN(P3_U2814) );
  NOR3_X1 U20402 ( .A1(n17576), .A2(n17556), .A3(n17562), .ZN(n17233) );
  NOR2_X1 U20403 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17233), .ZN(
        n17547) );
  NAND2_X1 U20404 ( .A1(n17715), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n17549) );
  OAI221_X1 U20405 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17215), .C1(
        n17214), .C2(n17213), .A(n17549), .ZN(n17216) );
  AOI21_X1 U20406 ( .B1(n17258), .B2(n17217), .A(n17216), .ZN(n17224) );
  INV_X1 U20407 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17550) );
  NAND3_X1 U20408 ( .A1(n17597), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n17574), .ZN(n17219) );
  INV_X1 U20409 ( .A(n17262), .ZN(n17218) );
  AOI22_X1 U20410 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17219), .B1(
        n17218), .B2(n17559), .ZN(n17220) );
  OAI221_X1 U20411 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n17562), 
        .C1(n17591), .C2(n17318), .A(n17220), .ZN(n17221) );
  XOR2_X1 U20412 ( .A(n17550), .B(n17221), .Z(n17553) );
  NOR2_X1 U20413 ( .A1(n17541), .A2(n17240), .ZN(n17222) );
  INV_X1 U20414 ( .A(n17533), .ZN(n17542) );
  OAI21_X1 U20415 ( .B1(n17542), .B2(n17310), .A(n17550), .ZN(n17545) );
  AOI22_X1 U20416 ( .A1(n17293), .A2(n17553), .B1(n17222), .B2(n17545), .ZN(
        n17223) );
  OAI211_X1 U20417 ( .C1(n17547), .C2(n17225), .A(n17224), .B(n17223), .ZN(
        P3_U2815) );
  NOR2_X1 U20418 ( .A1(n17313), .A2(n18090), .ZN(n17345) );
  INV_X1 U20419 ( .A(n17345), .ZN(n17286) );
  NOR2_X1 U20420 ( .A1(n17226), .A2(n17286), .ZN(n17290) );
  NAND2_X1 U20421 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n17290), .ZN(
        n17274) );
  OAI21_X1 U20422 ( .B1(n17228), .B2(n17274), .A(n17227), .ZN(n17230) );
  AOI22_X1 U20423 ( .A1(n17231), .A2(n17230), .B1(n17229), .B2(n17185), .ZN(
        n17243) );
  NAND2_X1 U20424 ( .A1(n17239), .A2(n17232), .ZN(n17234) );
  AOI21_X1 U20425 ( .B1(n17562), .B2(n17234), .A(n17233), .ZN(n17569) );
  NOR2_X1 U20426 ( .A1(n17235), .A2(n17310), .ZN(n17284) );
  AOI21_X1 U20427 ( .B1(n17284), .B2(n17239), .A(n17236), .ZN(n17237) );
  XOR2_X1 U20428 ( .A(n17237), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(
        n17567) );
  NAND2_X1 U20429 ( .A1(n17533), .A2(n17574), .ZN(n17238) );
  OAI221_X1 U20430 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17239), 
        .C1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n17574), .A(n17238), .ZN(
        n17565) );
  OAI22_X1 U20431 ( .A1(n17567), .A2(n17322), .B1(n17240), .B2(n17565), .ZN(
        n17241) );
  AOI21_X1 U20432 ( .B1(n17401), .B2(n17569), .A(n17241), .ZN(n17242) );
  OAI211_X1 U20433 ( .C1(n9746), .C2(n20705), .A(n17243), .B(n17242), .ZN(
        P3_U2816) );
  INV_X1 U20434 ( .A(n17303), .ZN(n17279) );
  AOI22_X1 U20435 ( .A1(n17310), .A2(n17309), .B1(n17401), .B2(n17576), .ZN(
        n17308) );
  INV_X1 U20436 ( .A(n17308), .ZN(n17280) );
  AOI21_X1 U20437 ( .B1(n17580), .B2(n17279), .A(n17280), .ZN(n17265) );
  INV_X1 U20438 ( .A(n17367), .ZN(n17403) );
  OAI21_X1 U20439 ( .B1(n17396), .B2(n17244), .A(n17403), .ZN(n17245) );
  OAI21_X1 U20440 ( .B1(n17246), .B2(n18255), .A(n17245), .ZN(n17259) );
  NOR2_X1 U20441 ( .A1(n9746), .A2(n20706), .ZN(n17252) );
  OAI211_X1 U20442 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17260), .B(n17261), .ZN(n17249) );
  OAI22_X1 U20443 ( .A1(n17250), .A2(n17249), .B1(n17248), .B2(n17247), .ZN(
        n17251) );
  AOI211_X1 U20444 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17259), .A(
        n17252), .B(n17251), .ZN(n17256) );
  INV_X1 U20445 ( .A(n17284), .ZN(n17301) );
  OAI21_X1 U20446 ( .B1(n17580), .B2(n17301), .A(n17253), .ZN(n17254) );
  XOR2_X1 U20447 ( .A(n17254), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .Z(
        n17583) );
  NOR2_X1 U20448 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17580), .ZN(
        n17582) );
  AOI22_X1 U20449 ( .A1(n17293), .A2(n17583), .B1(n17582), .B2(n17279), .ZN(
        n17255) );
  OAI211_X1 U20450 ( .C1(n17265), .C2(n17559), .A(n17256), .B(n17255), .ZN(
        P3_U2817) );
  AOI22_X1 U20451 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17259), .B1(
        n17258), .B2(n17257), .ZN(n17270) );
  AND2_X1 U20452 ( .A1(n17261), .A2(n17260), .ZN(n17268) );
  AOI21_X1 U20453 ( .B1(n17284), .B2(n17597), .A(n17262), .ZN(n17263) );
  XOR2_X1 U20454 ( .A(n17263), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n17595) );
  AOI21_X1 U20455 ( .B1(n17597), .B2(n17279), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17264) );
  OAI22_X1 U20456 ( .A1(n17595), .A2(n17322), .B1(n17265), .B2(n17264), .ZN(
        n17266) );
  AOI21_X1 U20457 ( .B1(n17268), .B2(n17267), .A(n17266), .ZN(n17269) );
  OAI211_X1 U20458 ( .C1(n9746), .C2(n18292), .A(n17270), .B(n17269), .ZN(
        P3_U2818) );
  INV_X1 U20459 ( .A(n17604), .ZN(n17273) );
  OAI21_X1 U20460 ( .B1(n17273), .B2(n17301), .A(n17271), .ZN(n17272) );
  XNOR2_X1 U20461 ( .A(n17272), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17608) );
  NOR2_X1 U20462 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17273), .ZN(
        n17596) );
  OAI211_X1 U20463 ( .C1(n17290), .C2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n17403), .B(n17274), .ZN(n17276) );
  NAND2_X1 U20464 ( .A1(n17710), .A2(P3_REIP_REG_11__SCAN_IN), .ZN(n17275) );
  OAI211_X1 U20465 ( .C1(n17393), .C2(n17277), .A(n17276), .B(n17275), .ZN(
        n17278) );
  AOI21_X1 U20466 ( .B1(n17596), .B2(n17279), .A(n17278), .ZN(n17282) );
  NOR2_X1 U20467 ( .A1(n17604), .A2(n17303), .ZN(n17294) );
  OAI21_X1 U20468 ( .B1(n17294), .B2(n17280), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17281) );
  OAI211_X1 U20469 ( .C1(n17608), .C2(n17322), .A(n17282), .B(n17281), .ZN(
        P3_U2819) );
  AOI21_X1 U20470 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17284), .A(
        n17283), .ZN(n17285) );
  XOR2_X1 U20471 ( .A(n17616), .B(n17285), .Z(n17612) );
  NOR2_X1 U20472 ( .A1(n9746), .A2(n18288), .ZN(n17292) );
  NOR3_X1 U20473 ( .A1(n17314), .A2(n17287), .A3(n17286), .ZN(n17299) );
  AOI21_X1 U20474 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17403), .A(
        n17299), .ZN(n17289) );
  OAI22_X1 U20475 ( .A1(n17290), .A2(n17289), .B1(n17393), .B2(n17288), .ZN(
        n17291) );
  AOI211_X1 U20476 ( .C1(n17293), .C2(n17612), .A(n17292), .B(n17291), .ZN(
        n17296) );
  OAI21_X1 U20477 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n17294), .ZN(n17295) );
  OAI211_X1 U20478 ( .C1(n17308), .C2(n17616), .A(n17296), .B(n17295), .ZN(
        P3_U2820) );
  AOI22_X1 U20479 ( .A1(n17297), .A2(n17345), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17403), .ZN(n17298) );
  NAND2_X1 U20480 ( .A1(n17715), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n17621) );
  OAI21_X1 U20481 ( .B1(n17299), .B2(n17298), .A(n17621), .ZN(n17305) );
  NAND2_X1 U20482 ( .A1(n17301), .A2(n17300), .ZN(n17302) );
  XOR2_X1 U20483 ( .A(n17302), .B(n17609), .Z(n17623) );
  OAI22_X1 U20484 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17303), .B1(
        n17623), .B2(n17322), .ZN(n17304) );
  AOI211_X1 U20485 ( .C1(n17306), .C2(n17185), .A(n17305), .B(n17304), .ZN(
        n17307) );
  OAI21_X1 U20486 ( .B1(n17308), .B2(n17609), .A(n17307), .ZN(P3_U2821) );
  NAND2_X1 U20487 ( .A1(n17310), .A2(n17309), .ZN(n17326) );
  OAI21_X1 U20488 ( .B1(n17312), .B2(n17311), .A(n17408), .ZN(n17330) );
  NOR2_X1 U20489 ( .A1(n17313), .A2(n17331), .ZN(n17315) );
  OAI211_X1 U20490 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17315), .A(
        n18121), .B(n17314), .ZN(n17316) );
  NAND2_X1 U20491 ( .A1(n17710), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n17632) );
  OAI211_X1 U20492 ( .C1(n17393), .C2(n17317), .A(n17316), .B(n17632), .ZN(
        n17324) );
  NOR2_X1 U20493 ( .A1(n17327), .A2(n17574), .ZN(n17319) );
  XOR2_X1 U20494 ( .A(n17319), .B(n17318), .Z(n17640) );
  OAI21_X1 U20495 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17321), .A(
        n17320), .ZN(n17642) );
  OAI22_X1 U20496 ( .A1(n17640), .A2(n17322), .B1(n17412), .B2(n17642), .ZN(
        n17323) );
  AOI211_X1 U20497 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17330), .A(
        n17324), .B(n17323), .ZN(n17325) );
  OAI21_X1 U20498 ( .B1(n17327), .B2(n17326), .A(n17325), .ZN(P3_U2822) );
  OAI21_X1 U20499 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17329), .A(
        n17328), .ZN(n17651) );
  NOR2_X1 U20500 ( .A1(n9746), .A2(n18282), .ZN(n17643) );
  AOI221_X1 U20501 ( .B1(n17345), .B2(n17331), .C1(n17330), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n17643), .ZN(n17338) );
  AOI21_X1 U20502 ( .B1(n17334), .B2(n17333), .A(n17332), .ZN(n17335) );
  XOR2_X1 U20503 ( .A(n17335), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n17648) );
  AOI22_X1 U20504 ( .A1(n17401), .A2(n17648), .B1(n17336), .B2(n17185), .ZN(
        n17337) );
  OAI211_X1 U20505 ( .C1(n17411), .C2(n17651), .A(n17338), .B(n17337), .ZN(
        P3_U2823) );
  OAI21_X1 U20506 ( .B1(n17341), .B2(n17340), .A(n17339), .ZN(n17654) );
  AOI22_X1 U20507 ( .A1(n17354), .A2(n18121), .B1(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17403), .ZN(n17344) );
  OAI21_X1 U20508 ( .B1(n17343), .B2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n17342), .ZN(n17655) );
  OAI22_X1 U20509 ( .A1(n17345), .A2(n17344), .B1(n17412), .B2(n17655), .ZN(
        n17346) );
  AOI21_X1 U20510 ( .B1(n17347), .B2(n17185), .A(n17346), .ZN(n17348) );
  NAND2_X1 U20511 ( .A1(n17710), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n17658) );
  OAI211_X1 U20512 ( .C1(n17411), .C2(n17654), .A(n17348), .B(n17658), .ZN(
        P3_U2824) );
  OAI21_X1 U20513 ( .B1(n17351), .B2(n17350), .A(n17349), .ZN(n17662) );
  AOI221_X1 U20514 ( .B1(n17396), .B2(n17353), .C1(n17352), .C2(n17353), .A(
        n17367), .ZN(n17362) );
  NAND2_X1 U20515 ( .A1(n17354), .A2(n18121), .ZN(n17361) );
  OAI21_X1 U20516 ( .B1(n17357), .B2(n17356), .A(n17355), .ZN(n17358) );
  XOR2_X1 U20517 ( .A(n17358), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(
        n17661) );
  OAI22_X1 U20518 ( .A1(n17393), .A2(n17359), .B1(n17411), .B2(n17661), .ZN(
        n17360) );
  AOI21_X1 U20519 ( .B1(n17362), .B2(n17361), .A(n17360), .ZN(n17363) );
  NAND2_X1 U20520 ( .A1(n17710), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n17665) );
  OAI211_X1 U20521 ( .C1(n17412), .C2(n17662), .A(n17363), .B(n17665), .ZN(
        P3_U2825) );
  OAI21_X1 U20522 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n17365), .A(
        n17364), .ZN(n17673) );
  AOI22_X1 U20523 ( .A1(n17715), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18121), 
        .B2(n17366), .ZN(n17374) );
  NOR2_X1 U20524 ( .A1(n17396), .A2(n17395), .ZN(n17383) );
  AOI21_X1 U20525 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17383), .A(
        n17367), .ZN(n17384) );
  OAI21_X1 U20526 ( .B1(n17370), .B2(n17369), .A(n17368), .ZN(n17679) );
  OAI22_X1 U20527 ( .A1(n17393), .A2(n17371), .B1(n17411), .B2(n17679), .ZN(
        n17372) );
  AOI21_X1 U20528 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17384), .A(
        n17372), .ZN(n17373) );
  OAI211_X1 U20529 ( .C1(n17412), .C2(n17673), .A(n17374), .B(n17373), .ZN(
        P3_U2826) );
  OAI21_X1 U20530 ( .B1(n17377), .B2(n17376), .A(n17375), .ZN(n17689) );
  OAI21_X1 U20531 ( .B1(n17380), .B2(n17379), .A(n17378), .ZN(n17685) );
  OAI22_X1 U20532 ( .A1(n17393), .A2(n17381), .B1(n17411), .B2(n17685), .ZN(
        n17382) );
  AOI221_X1 U20533 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17384), .C1(
        n17383), .C2(n17384), .A(n17382), .ZN(n17385) );
  NAND2_X1 U20534 ( .A1(n17715), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n17684) );
  OAI211_X1 U20535 ( .C1(n17412), .C2(n17689), .A(n17385), .B(n17684), .ZN(
        P3_U2827) );
  OAI21_X1 U20536 ( .B1(n17388), .B2(n17387), .A(n17386), .ZN(n17702) );
  OAI21_X1 U20537 ( .B1(n17391), .B2(n17390), .A(n17389), .ZN(n17697) );
  OAI22_X1 U20538 ( .A1(n17393), .A2(n17392), .B1(n17411), .B2(n17697), .ZN(
        n17394) );
  AOI221_X1 U20539 ( .B1(n17396), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C1(
        n18121), .C2(n17395), .A(n17394), .ZN(n17397) );
  NAND2_X1 U20540 ( .A1(n17715), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n17700) );
  OAI211_X1 U20541 ( .C1(n17412), .C2(n17702), .A(n17397), .B(n17700), .ZN(
        P3_U2828) );
  OAI21_X1 U20542 ( .B1(n17399), .B2(n17406), .A(n17398), .ZN(n17714) );
  NAND2_X1 U20543 ( .A1(n18366), .A2(n17407), .ZN(n17400) );
  XNOR2_X1 U20544 ( .A(n17400), .B(n17399), .ZN(n17709) );
  AOI22_X1 U20545 ( .A1(n17401), .A2(n17709), .B1(n17710), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17405) );
  AOI22_X1 U20546 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17403), .B1(
        n17185), .B2(n17402), .ZN(n17404) );
  OAI211_X1 U20547 ( .C1(n17411), .C2(n17714), .A(n17405), .B(n17404), .ZN(
        P3_U2829) );
  AOI21_X1 U20548 ( .B1(n17407), .B2(n18366), .A(n17406), .ZN(n17720) );
  INV_X1 U20549 ( .A(n17720), .ZN(n17718) );
  NAND3_X1 U20550 ( .A1(n18348), .A2(n18255), .A3(n17408), .ZN(n17409) );
  AOI22_X1 U20551 ( .A1(n17715), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17409), .ZN(n17410) );
  OAI221_X1 U20552 ( .B1(n17720), .B2(n17412), .C1(n17718), .C2(n17411), .A(
        n17410), .ZN(P3_U2830) );
  NOR2_X1 U20553 ( .A1(n17413), .A2(n17458), .ZN(n17420) );
  NOR2_X1 U20554 ( .A1(n18190), .A2(n17602), .ZN(n17627) );
  NAND2_X1 U20555 ( .A1(n17602), .A2(n18366), .ZN(n17510) );
  INV_X1 U20556 ( .A(n17510), .ZN(n17669) );
  AOI221_X1 U20557 ( .B1(n17431), .B2(n17671), .C1(n17446), .C2(n17671), .A(
        n17669), .ZN(n17429) );
  AOI22_X1 U20558 ( .A1(n17602), .A2(n17418), .B1(n17435), .B2(n17671), .ZN(
        n17417) );
  AOI21_X1 U20559 ( .B1(n18190), .B2(n17418), .A(n17424), .ZN(n17419) );
  AOI22_X1 U20560 ( .A1(n17613), .A2(n17423), .B1(n17444), .B2(n17422), .ZN(
        n17427) );
  OAI211_X1 U20561 ( .C1(n17680), .C2(n17424), .A(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n9746), .ZN(n17425) );
  NAND3_X1 U20562 ( .A1(n17427), .A2(n17426), .A3(n17425), .ZN(P3_U2836) );
  NOR2_X1 U20563 ( .A1(n17428), .A2(n17431), .ZN(n17434) );
  INV_X1 U20564 ( .A(n17429), .ZN(n17430) );
  AOI221_X1 U20565 ( .B1(n17431), .B2(n18218), .C1(n17452), .C2(n18218), .A(
        n17430), .ZN(n17432) );
  INV_X1 U20566 ( .A(n17432), .ZN(n17433) );
  MUX2_X1 U20567 ( .A(n17434), .B(n17433), .S(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(n17437) );
  OAI22_X1 U20568 ( .A1(n17435), .A2(n17705), .B1(n9746), .B2(n18314), .ZN(
        n17436) );
  AOI21_X1 U20569 ( .B1(n17716), .B2(n17437), .A(n17436), .ZN(n17441) );
  AOI22_X1 U20570 ( .A1(n17719), .A2(n17439), .B1(n17613), .B2(n17438), .ZN(
        n17440) );
  OAI211_X1 U20571 ( .C1(n17566), .C2(n17442), .A(n17441), .B(n17440), .ZN(
        P3_U2837) );
  AOI22_X1 U20572 ( .A1(n17613), .A2(n17445), .B1(n17444), .B2(n17443), .ZN(
        n17457) );
  AOI21_X1 U20573 ( .B1(n17671), .B2(n17446), .A(n17669), .ZN(n17449) );
  AOI21_X1 U20574 ( .B1(n17472), .B2(n17447), .A(n17699), .ZN(n17448) );
  OAI211_X1 U20575 ( .C1(n17450), .C2(n17468), .A(n17449), .B(n17448), .ZN(
        n17454) );
  AOI211_X1 U20576 ( .C1(n18218), .C2(n17452), .A(n17451), .B(n17454), .ZN(
        n17453) );
  NOR2_X1 U20577 ( .A1(n17710), .A2(n17453), .ZN(n17459) );
  OAI211_X1 U20578 ( .C1(n17534), .C2(n17454), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n17459), .ZN(n17455) );
  NAND3_X1 U20579 ( .A1(n17457), .A2(n17456), .A3(n17455), .ZN(P3_U2838) );
  INV_X1 U20580 ( .A(n17458), .ZN(n17460) );
  OAI221_X1 U20581 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17460), 
        .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n17705), .A(n17459), .ZN(
        n17461) );
  OAI211_X1 U20582 ( .C1(n17463), .C2(n17636), .A(n17462), .B(n17461), .ZN(
        P3_U2839) );
  AOI21_X1 U20583 ( .B1(n17465), .B2(n17613), .A(n17464), .ZN(n17479) );
  INV_X1 U20584 ( .A(n17466), .ZN(n17485) );
  NOR2_X1 U20585 ( .A1(n17485), .A2(n17473), .ZN(n17477) );
  AOI21_X1 U20586 ( .B1(n17467), .B2(n17512), .A(n18185), .ZN(n17471) );
  NOR3_X1 U20587 ( .A1(n18366), .A2(n17507), .A3(n17557), .ZN(n17530) );
  AOI21_X1 U20588 ( .B1(n17467), .B2(n17530), .A(n18188), .ZN(n17470) );
  AOI21_X1 U20589 ( .B1(n17511), .B2(n17496), .A(n18202), .ZN(n17469) );
  OAI22_X1 U20590 ( .A1(n17548), .A2(n17468), .B1(n17541), .B2(n17573), .ZN(
        n17514) );
  NOR4_X1 U20591 ( .A1(n17471), .A2(n17470), .A3(n17469), .A4(n17514), .ZN(
        n17494) );
  NOR2_X1 U20592 ( .A1(n18217), .A2(n17472), .ZN(n17603) );
  INV_X1 U20593 ( .A(n17603), .ZN(n17579) );
  AOI22_X1 U20594 ( .A1(n18190), .A2(n17474), .B1(n17473), .B2(n17579), .ZN(
        n17481) );
  OAI211_X1 U20595 ( .C1(n17630), .C2(n17475), .A(n17494), .B(n17481), .ZN(
        n17476) );
  OAI221_X1 U20596 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n17477), 
        .C1(n17480), .C2(n17476), .A(n17716), .ZN(n17478) );
  OAI211_X1 U20597 ( .C1(n17705), .C2(n17480), .A(n17479), .B(n17478), .ZN(
        P3_U2840) );
  NAND3_X1 U20598 ( .A1(n17716), .A2(n17494), .A3(n17481), .ZN(n17483) );
  NAND2_X1 U20599 ( .A1(n18188), .A2(n18185), .ZN(n17704) );
  OAI221_X1 U20600 ( .B1(n17483), .B2(n17482), .C1(n17483), .C2(n17704), .A(
        n9746), .ZN(n17490) );
  NOR3_X1 U20601 ( .A1(n17485), .A2(n17680), .A3(n17484), .ZN(n17503) );
  AOI22_X1 U20602 ( .A1(n17613), .A2(n17487), .B1(n17486), .B2(n17503), .ZN(
        n17489) );
  OAI211_X1 U20603 ( .C1(n17491), .C2(n17490), .A(n17489), .B(n17488), .ZN(
        P3_U2841) );
  AOI21_X1 U20604 ( .B1(n17493), .B2(n17503), .A(n17492), .ZN(n17499) );
  AND2_X1 U20605 ( .A1(n17716), .A2(n17494), .ZN(n17495) );
  AOI221_X1 U20606 ( .B1(n17496), .B2(n17495), .C1(n17603), .C2(n17495), .A(
        n17715), .ZN(n17504) );
  AND3_X1 U20607 ( .A1(n17502), .A2(n17704), .A3(P3_STATE2_REG_2__SCAN_IN), 
        .ZN(n17497) );
  OAI21_X1 U20608 ( .B1(n17504), .B2(n17497), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17498) );
  OAI211_X1 U20609 ( .C1(n17500), .C2(n17636), .A(n17499), .B(n17498), .ZN(
        P3_U2842) );
  AOI221_X1 U20610 ( .B1(n17504), .B2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), 
        .C1(n17503), .C2(n17502), .A(n17501), .ZN(n17505) );
  OAI21_X1 U20611 ( .B1(n17506), .B2(n17636), .A(n17505), .ZN(P3_U2843) );
  OAI22_X1 U20612 ( .A1(n17692), .A2(n18185), .B1(n17690), .B2(n17670), .ZN(
        n17624) );
  INV_X1 U20613 ( .A(n17624), .ZN(n17683) );
  NOR2_X1 U20614 ( .A1(n17683), .A2(n17508), .ZN(n17644) );
  NAND2_X1 U20615 ( .A1(n17509), .A2(n17644), .ZN(n17587) );
  AOI21_X1 U20616 ( .B1(n17588), .B2(n17587), .A(n17680), .ZN(n17620) );
  NAND2_X1 U20617 ( .A1(n9802), .A2(n17620), .ZN(n17540) );
  NAND3_X1 U20618 ( .A1(n17511), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n17510), .ZN(n17516) );
  AOI222_X1 U20619 ( .A1(n17513), .A2(n18185), .B1(n17513), .B2(n17512), .C1(
        n18185), .C2(n17603), .ZN(n17515) );
  OR2_X1 U20620 ( .A1(n17680), .A2(n17514), .ZN(n17535) );
  AOI211_X1 U20621 ( .C1(n17671), .C2(n17516), .A(n17515), .B(n17535), .ZN(
        n17523) );
  AOI221_X1 U20622 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17523), 
        .C1(n17627), .C2(n17523), .A(n17715), .ZN(n17518) );
  AOI22_X1 U20623 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17518), .B1(
        n17613), .B2(n17517), .ZN(n17520) );
  OAI211_X1 U20624 ( .C1(n17521), .C2(n17540), .A(n17520), .B(n17519), .ZN(
        P3_U2844) );
  NAND2_X1 U20625 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17522), .ZN(
        n17528) );
  NOR3_X1 U20626 ( .A1(n17715), .A2(n17523), .A3(n17522), .ZN(n17524) );
  AOI21_X1 U20627 ( .B1(n17613), .B2(n17525), .A(n17524), .ZN(n17527) );
  OAI211_X1 U20628 ( .C1(n17528), .C2(n17540), .A(n17527), .B(n17526), .ZN(
        P3_U2845) );
  INV_X1 U20629 ( .A(n17610), .ZN(n17598) );
  AOI22_X1 U20630 ( .A1(n18218), .A2(n17529), .B1(n18190), .B2(n17557), .ZN(
        n17572) );
  AOI21_X1 U20631 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18188), .A(
        n17530), .ZN(n17531) );
  INV_X1 U20632 ( .A(n17531), .ZN(n17532) );
  OAI211_X1 U20633 ( .C1(n17598), .C2(n17533), .A(n17572), .B(n17532), .ZN(
        n17544) );
  OAI221_X1 U20634 ( .B1(n17535), .B2(n17534), .C1(n17535), .C2(n17544), .A(
        n9746), .ZN(n17538) );
  AOI22_X1 U20635 ( .A1(n17715), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n17613), 
        .B2(n17536), .ZN(n17537) );
  OAI221_X1 U20636 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17540), 
        .C1(n17539), .C2(n17538), .A(n17537), .ZN(P3_U2846) );
  NOR2_X1 U20637 ( .A1(n17541), .A2(n17573), .ZN(n17546) );
  OAI21_X1 U20638 ( .B1(n17542), .B2(n17587), .A(n17550), .ZN(n17543) );
  AOI22_X1 U20639 ( .A1(n17546), .A2(n17545), .B1(n17544), .B2(n17543), .ZN(
        n17555) );
  NOR3_X1 U20640 ( .A1(n17548), .A2(n17547), .A3(n17703), .ZN(n17552) );
  OAI21_X1 U20641 ( .B1(n17705), .B2(n17550), .A(n17549), .ZN(n17551) );
  AOI211_X1 U20642 ( .C1(n17553), .C2(n17613), .A(n17552), .B(n17551), .ZN(
        n17554) );
  OAI21_X1 U20643 ( .B1(n17555), .B2(n17680), .A(n17554), .ZN(P3_U2847) );
  NOR2_X1 U20644 ( .A1(n17556), .A2(n17587), .ZN(n17564) );
  AOI22_X1 U20645 ( .A1(n18218), .A2(n17580), .B1(n18190), .B2(n17556), .ZN(
        n17558) );
  OR2_X1 U20646 ( .A1(n18366), .A2(n17557), .ZN(n17601) );
  OAI21_X1 U20647 ( .B1(n17580), .B2(n17601), .A(n17602), .ZN(n17577) );
  NAND4_X1 U20648 ( .A1(n17572), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n17558), .A4(n17577), .ZN(n17560) );
  OAI221_X1 U20649 ( .B1(n17560), .B2(n17559), .C1(n17560), .C2(n17704), .A(
        n17716), .ZN(n17561) );
  OAI21_X1 U20650 ( .B1(n17705), .B2(n17562), .A(n17561), .ZN(n17563) );
  OAI21_X1 U20651 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17564), .A(
        n17563), .ZN(n17571) );
  OAI22_X1 U20652 ( .A1(n17567), .A2(n17636), .B1(n17566), .B2(n17565), .ZN(
        n17568) );
  AOI21_X1 U20653 ( .B1(n17719), .B2(n17569), .A(n17568), .ZN(n17570) );
  OAI211_X1 U20654 ( .C1(n9746), .C2(n20705), .A(n17571), .B(n17570), .ZN(
        P3_U2848) );
  OAI21_X1 U20655 ( .B1(n17574), .B2(n17573), .A(n17572), .ZN(n17575) );
  AOI21_X1 U20656 ( .B1(n18217), .B2(n17576), .A(n17575), .ZN(n17599) );
  OAI211_X1 U20657 ( .C1(n17598), .C2(n17597), .A(n17599), .B(n17577), .ZN(
        n17578) );
  AOI21_X1 U20658 ( .B1(n17580), .B2(n17579), .A(n17578), .ZN(n17589) );
  OAI211_X1 U20659 ( .C1(n17598), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n17716), .B(n17589), .ZN(n17581) );
  NAND2_X1 U20660 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17581), .ZN(
        n17585) );
  AOI22_X1 U20661 ( .A1(n17613), .A2(n17583), .B1(n17620), .B2(n17582), .ZN(
        n17584) );
  OAI221_X1 U20662 ( .B1(n17710), .B2(n17585), .C1(n9746), .C2(n20706), .A(
        n17584), .ZN(P3_U2849) );
  AOI22_X1 U20663 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17699), .B1(
        n17710), .B2(P3_REIP_REG_12__SCAN_IN), .ZN(n17594) );
  AOI21_X1 U20664 ( .B1(n17588), .B2(n17587), .A(n17586), .ZN(n17592) );
  INV_X1 U20665 ( .A(n17589), .ZN(n17590) );
  OAI221_X1 U20666 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n17592), 
        .C1(n17591), .C2(n17590), .A(n17716), .ZN(n17593) );
  OAI211_X1 U20667 ( .C1(n17595), .C2(n17636), .A(n17594), .B(n17593), .ZN(
        P3_U2850) );
  AOI22_X1 U20668 ( .A1(n17715), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n17620), 
        .B2(n17596), .ZN(n17607) );
  NOR2_X1 U20669 ( .A1(n17598), .A2(n17597), .ZN(n17605) );
  INV_X1 U20670 ( .A(n17599), .ZN(n17600) );
  AOI211_X1 U20671 ( .C1(n17602), .C2(n17601), .A(n17680), .B(n17600), .ZN(
        n17618) );
  OAI221_X1 U20672 ( .B1(n17604), .B2(n18188), .C1(n17604), .C2(n17603), .A(
        n17618), .ZN(n17611) );
  OAI211_X1 U20673 ( .C1(n17605), .C2(n17611), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n9746), .ZN(n17606) );
  OAI211_X1 U20674 ( .C1(n17608), .C2(n17636), .A(n17607), .B(n17606), .ZN(
        P3_U2851) );
  NAND2_X1 U20675 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17620), .ZN(
        n17617) );
  OAI221_X1 U20676 ( .B1(n17611), .B2(n17610), .C1(n17611), .C2(n17609), .A(
        n9746), .ZN(n17615) );
  AOI22_X1 U20677 ( .A1(n17715), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n17613), 
        .B2(n17612), .ZN(n17614) );
  OAI221_X1 U20678 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n17617), 
        .C1(n17616), .C2(n17615), .A(n17614), .ZN(P3_U2852) );
  OAI21_X1 U20679 ( .B1(n17710), .B2(n17618), .A(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17619) );
  OAI21_X1 U20680 ( .B1(n17620), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17619), .ZN(n17622) );
  OAI211_X1 U20681 ( .C1(n17623), .C2(n17636), .A(n17622), .B(n17621), .ZN(
        P3_U2853) );
  INV_X1 U20682 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n17625) );
  NAND3_X1 U20683 ( .A1(n17716), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n17624), .ZN(n17674) );
  NOR3_X1 U20684 ( .A1(n17667), .A2(n17625), .A3(n17674), .ZN(n17657) );
  NAND3_X1 U20685 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n17657), .ZN(n17635) );
  OAI22_X1 U20686 ( .A1(n17628), .A2(n18185), .B1(n17627), .B2(n17626), .ZN(
        n17629) );
  NOR2_X1 U20687 ( .A1(n17669), .A2(n17629), .ZN(n17652) );
  OAI211_X1 U20688 ( .C1(n17630), .C2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B(n17652), .ZN(n17646) );
  AOI21_X1 U20689 ( .B1(n17631), .B2(n17646), .A(n17699), .ZN(n17633) );
  OAI221_X1 U20690 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17635), .C1(
        n17634), .C2(n17633), .A(n17632), .ZN(n17638) );
  NOR2_X1 U20691 ( .A1(n17636), .A2(n17640), .ZN(n17637) );
  AOI211_X1 U20692 ( .C1(n17640), .C2(n17639), .A(n17638), .B(n17637), .ZN(
        n17641) );
  OAI21_X1 U20693 ( .B1(n17703), .B2(n17642), .A(n17641), .ZN(P3_U2854) );
  INV_X1 U20694 ( .A(n17721), .ZN(n17713) );
  AOI21_X1 U20695 ( .B1(n17699), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n17643), .ZN(n17650) );
  AOI21_X1 U20696 ( .B1(n17644), .B2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17645) );
  NOR2_X1 U20697 ( .A1(n17645), .A2(n17680), .ZN(n17647) );
  AOI22_X1 U20698 ( .A1(n17719), .A2(n17648), .B1(n17647), .B2(n17646), .ZN(
        n17649) );
  OAI211_X1 U20699 ( .C1(n17713), .C2(n17651), .A(n17650), .B(n17649), .ZN(
        P3_U2855) );
  OAI21_X1 U20700 ( .B1(n17680), .B2(n17652), .A(n17705), .ZN(n17653) );
  INV_X1 U20701 ( .A(n17653), .ZN(n17668) );
  OAI22_X1 U20702 ( .A1(n17703), .A2(n17655), .B1(n17713), .B2(n17654), .ZN(
        n17656) );
  AOI21_X1 U20703 ( .B1(n17657), .B2(n17660), .A(n17656), .ZN(n17659) );
  OAI211_X1 U20704 ( .C1(n17668), .C2(n17660), .A(n17659), .B(n17658), .ZN(
        P3_U2856) );
  NOR2_X1 U20705 ( .A1(n17674), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17664) );
  OAI22_X1 U20706 ( .A1(n17703), .A2(n17662), .B1(n17713), .B2(n17661), .ZN(
        n17663) );
  AOI21_X1 U20707 ( .B1(n17664), .B2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n17663), .ZN(n17666) );
  OAI211_X1 U20708 ( .C1(n17668), .C2(n17667), .A(n17666), .B(n17665), .ZN(
        P3_U2857) );
  AOI21_X1 U20709 ( .B1(n17671), .B2(n17670), .A(n17669), .ZN(n17672) );
  INV_X1 U20710 ( .A(n17672), .ZN(n17694) );
  AOI211_X1 U20711 ( .C1(n18218), .C2(n17692), .A(n17682), .B(n17694), .ZN(
        n17681) );
  OAI21_X1 U20712 ( .B1(n17681), .B2(n17706), .A(n17705), .ZN(n17676) );
  OAI22_X1 U20713 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n17674), .B1(
        n17673), .B2(n17703), .ZN(n17675) );
  AOI21_X1 U20714 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n17676), .A(
        n17675), .ZN(n17678) );
  NAND2_X1 U20715 ( .A1(n17710), .A2(P3_REIP_REG_4__SCAN_IN), .ZN(n17677) );
  OAI211_X1 U20716 ( .C1(n17679), .C2(n17713), .A(n17678), .B(n17677), .ZN(
        P3_U2858) );
  AOI211_X1 U20717 ( .C1(n17683), .C2(n17682), .A(n17681), .B(n17680), .ZN(
        n17687) );
  OAI21_X1 U20718 ( .B1(n17685), .B2(n17713), .A(n17684), .ZN(n17686) );
  AOI211_X1 U20719 ( .C1(n17699), .C2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n17687), .B(n17686), .ZN(n17688) );
  OAI21_X1 U20720 ( .B1(n17703), .B2(n17689), .A(n17688), .ZN(P3_U2859) );
  NOR2_X1 U20721 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n17690), .ZN(
        n17691) );
  AOI22_X1 U20722 ( .A1(n18218), .A2(n17692), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n17691), .ZN(n17696) );
  INV_X1 U20723 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18350) );
  NOR2_X1 U20724 ( .A1(n18366), .A2(n18350), .ZN(n17693) );
  OAI221_X1 U20725 ( .B1(n17694), .B2(n18218), .C1(n17694), .C2(n17693), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n17695) );
  OAI211_X1 U20726 ( .C1(n17697), .C2(n18224), .A(n17696), .B(n17695), .ZN(
        n17698) );
  AOI22_X1 U20727 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n17699), .B1(
        n17716), .B2(n17698), .ZN(n17701) );
  OAI211_X1 U20728 ( .C1(n17703), .C2(n17702), .A(n17701), .B(n17700), .ZN(
        P3_U2860) );
  NAND3_X1 U20729 ( .A1(n17716), .A2(n18366), .A3(n17704), .ZN(n17722) );
  AOI21_X1 U20730 ( .B1(n17705), .B2(n17722), .A(n18350), .ZN(n17708) );
  AOI211_X1 U20731 ( .C1(n18202), .C2(n18366), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n17706), .ZN(n17707) );
  AOI211_X1 U20732 ( .C1(n17719), .C2(n17709), .A(n17708), .B(n17707), .ZN(
        n17712) );
  NAND2_X1 U20733 ( .A1(n17710), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n17711) );
  OAI211_X1 U20734 ( .C1(n17714), .C2(n17713), .A(n17712), .B(n17711), .ZN(
        P3_U2861) );
  INV_X1 U20735 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n18377) );
  AOI211_X1 U20736 ( .C1(n18202), .C2(n17716), .A(n17715), .B(n18366), .ZN(
        n17717) );
  AOI221_X1 U20737 ( .B1(n17721), .B2(n17720), .C1(n17719), .C2(n17718), .A(
        n17717), .ZN(n17723) );
  OAI211_X1 U20738 ( .C1(n18377), .C2(n9746), .A(n17723), .B(n17722), .ZN(
        P3_U2862) );
  AOI211_X1 U20739 ( .C1(n17725), .C2(n17724), .A(n18403), .B(n18348), .ZN(
        n18238) );
  OAI21_X1 U20740 ( .B1(n18238), .B2(n17785), .A(n17730), .ZN(n17726) );
  OAI221_X1 U20741 ( .B1(n17988), .B2(n18388), .C1(n17988), .C2(n17730), .A(
        n17726), .ZN(P3_U2863) );
  NAND2_X1 U20742 ( .A1(n18209), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n17986) );
  INV_X1 U20743 ( .A(n17986), .ZN(n18013) );
  NAND2_X1 U20744 ( .A1(n18196), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n17872) );
  INV_X1 U20745 ( .A(n17872), .ZN(n17920) );
  NOR2_X1 U20746 ( .A1(n18013), .A2(n17920), .ZN(n17728) );
  OAI22_X1 U20747 ( .A1(n17729), .A2(n18196), .B1(n17728), .B2(n17727), .ZN(
        P3_U2866) );
  INV_X1 U20748 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18195) );
  NOR2_X1 U20749 ( .A1(n18195), .A2(n17730), .ZN(P3_U2867) );
  NOR2_X1 U20750 ( .A1(n18196), .A2(n17895), .ZN(n18119) );
  NAND2_X1 U20751 ( .A1(n17988), .A2(n18119), .ZN(n18115) );
  NAND3_X1 U20752 ( .A1(n17987), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18059) );
  INV_X1 U20753 ( .A(n18059), .ZN(n18120) );
  NAND2_X1 U20754 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18120), .ZN(
        n18149) );
  INV_X1 U20755 ( .A(n18149), .ZN(n18167) );
  OAI21_X1 U20756 ( .B1(n18106), .B2(n18167), .A(n18037), .ZN(n18089) );
  NOR2_X1 U20757 ( .A1(n17987), .A2(n17988), .ZN(n18191) );
  NAND3_X1 U20758 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n18191), .ZN(n18174) );
  INV_X1 U20759 ( .A(n18174), .ZN(n18159) );
  NOR2_X1 U20760 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18192) );
  NAND2_X1 U20761 ( .A1(n18209), .A2(n18196), .ZN(n17807) );
  INV_X1 U20762 ( .A(n17807), .ZN(n17829) );
  NAND2_X1 U20763 ( .A1(n18192), .A2(n17829), .ZN(n17836) );
  NOR2_X1 U20764 ( .A1(n18159), .A2(n17846), .ZN(n17808) );
  AOI211_X1 U20765 ( .C1(P3_STATE2_REG_3__SCAN_IN), .C2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n17896), .B(n17808), .ZN(
        n17731) );
  INV_X1 U20766 ( .A(n17731), .ZN(n17732) );
  OAI21_X1 U20767 ( .B1(n18035), .B2(n18089), .A(n17732), .ZN(n17783) );
  INV_X1 U20768 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n17733) );
  NOR2_X2 U20769 ( .A1(n17733), .A2(n18090), .ZN(n18088) );
  AND2_X1 U20770 ( .A1(n18037), .A2(BUF2_REG_0__SCAN_IN), .ZN(n18116) );
  NOR2_X1 U20771 ( .A1(n18087), .A2(n17808), .ZN(n17777) );
  AOI22_X1 U20772 ( .A1(n18088), .A2(n18167), .B1(n18116), .B2(n17777), .ZN(
        n17738) );
  NOR2_X1 U20773 ( .A1(n17735), .A2(n17734), .ZN(n17740) );
  NAND2_X1 U20774 ( .A1(n17736), .A2(n17740), .ZN(n18095) );
  INV_X1 U20775 ( .A(n18095), .ZN(n18122) );
  AND2_X1 U20776 ( .A1(n18121), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18117) );
  AOI22_X1 U20777 ( .A1(n18122), .A2(n17846), .B1(n18117), .B2(n18106), .ZN(
        n17737) );
  OAI211_X1 U20778 ( .C1(n17739), .C2(n17783), .A(n17738), .B(n17737), .ZN(
        P3_U2868) );
  NOR2_X2 U20779 ( .A1(n18090), .A2(n18893), .ZN(n18128) );
  AND2_X1 U20780 ( .A1(n18037), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18126) );
  AOI22_X1 U20781 ( .A1(n18128), .A2(n18106), .B1(n18126), .B2(n17777), .ZN(
        n17744) );
  INV_X1 U20782 ( .A(n17740), .ZN(n17779) );
  NOR2_X1 U20783 ( .A1(n17779), .A2(n17741), .ZN(n17788) );
  INV_X1 U20784 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n17742) );
  NOR2_X2 U20785 ( .A1(n17742), .A2(n18090), .ZN(n18127) );
  AOI22_X1 U20786 ( .A1(n17788), .A2(n17846), .B1(n18127), .B2(n18167), .ZN(
        n17743) );
  OAI211_X1 U20787 ( .C1(n17745), .C2(n17783), .A(n17744), .B(n17743), .ZN(
        P3_U2869) );
  NAND2_X1 U20788 ( .A1(n18121), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18137) );
  INV_X1 U20789 ( .A(n18137), .ZN(n18065) );
  NOR2_X2 U20790 ( .A1(n17896), .A2(n17746), .ZN(n18132) );
  AOI22_X1 U20791 ( .A1(n18065), .A2(n18106), .B1(n18132), .B2(n17777), .ZN(
        n17750) );
  NOR2_X1 U20792 ( .A1(n17747), .A2(n18090), .ZN(n18133) );
  NOR2_X2 U20793 ( .A1(n17748), .A2(n17779), .ZN(n18134) );
  AOI22_X1 U20794 ( .A1(n18133), .A2(n18167), .B1(n18134), .B2(n17846), .ZN(
        n17749) );
  OAI211_X1 U20795 ( .C1(n17751), .C2(n17783), .A(n17750), .B(n17749), .ZN(
        P3_U2870) );
  NOR2_X2 U20796 ( .A1(n17896), .A2(n17752), .ZN(n18138) );
  NAND2_X1 U20797 ( .A1(n18121), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18143) );
  INV_X1 U20798 ( .A(n18143), .ZN(n18069) );
  AOI22_X1 U20799 ( .A1(n18138), .A2(n17777), .B1(n18069), .B2(n18106), .ZN(
        n17756) );
  INV_X1 U20800 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n17753) );
  NOR2_X1 U20801 ( .A1(n17753), .A2(n18090), .ZN(n18139) );
  NOR2_X2 U20802 ( .A1(n17754), .A2(n17779), .ZN(n18140) );
  AOI22_X1 U20803 ( .A1(n18139), .A2(n18167), .B1(n18140), .B2(n17846), .ZN(
        n17755) );
  OAI211_X1 U20804 ( .C1(n17757), .C2(n17783), .A(n17756), .B(n17755), .ZN(
        P3_U2871) );
  NAND2_X1 U20805 ( .A1(n18121), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18150) );
  INV_X1 U20806 ( .A(n18150), .ZN(n18073) );
  NOR2_X2 U20807 ( .A1(n17896), .A2(n17758), .ZN(n18144) );
  AOI22_X1 U20808 ( .A1(n18073), .A2(n18106), .B1(n18144), .B2(n17777), .ZN(
        n17762) );
  NOR2_X1 U20809 ( .A1(n17759), .A2(n18090), .ZN(n18145) );
  NOR2_X2 U20810 ( .A1(n17760), .A2(n17779), .ZN(n18146) );
  AOI22_X1 U20811 ( .A1(n18145), .A2(n18167), .B1(n18146), .B2(n17846), .ZN(
        n17761) );
  OAI211_X1 U20812 ( .C1(n17763), .C2(n17783), .A(n17762), .B(n17761), .ZN(
        P3_U2872) );
  NOR2_X2 U20813 ( .A1(n17896), .A2(n17764), .ZN(n18151) );
  NOR2_X2 U20814 ( .A1(n17765), .A2(n18090), .ZN(n18152) );
  AOI22_X1 U20815 ( .A1(n18151), .A2(n17777), .B1(n18152), .B2(n18167), .ZN(
        n17768) );
  AND2_X1 U20816 ( .A1(n18121), .A2(BUF2_REG_21__SCAN_IN), .ZN(n18153) );
  NOR2_X1 U20817 ( .A1(n17779), .A2(n17766), .ZN(n17797) );
  AOI22_X1 U20818 ( .A1(n18153), .A2(n18106), .B1(n17797), .B2(n17846), .ZN(
        n17767) );
  OAI211_X1 U20819 ( .C1(n17769), .C2(n17783), .A(n17768), .B(n17767), .ZN(
        P3_U2873) );
  INV_X1 U20820 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17775) );
  NOR2_X1 U20821 ( .A1(n17770), .A2(n18090), .ZN(n18004) );
  NOR2_X2 U20822 ( .A1(n17896), .A2(n17771), .ZN(n18158) );
  AOI22_X1 U20823 ( .A1(n18004), .A2(n18167), .B1(n18158), .B2(n17777), .ZN(
        n17774) );
  NOR2_X2 U20824 ( .A1(n17772), .A2(n17779), .ZN(n18160) );
  NAND2_X1 U20825 ( .A1(n18121), .A2(BUF2_REG_22__SCAN_IN), .ZN(n18007) );
  INV_X1 U20826 ( .A(n18007), .ZN(n18157) );
  AOI22_X1 U20827 ( .A1(n18160), .A2(n17846), .B1(n18157), .B2(n18106), .ZN(
        n17773) );
  OAI211_X1 U20828 ( .C1(n17775), .C2(n17783), .A(n17774), .B(n17773), .ZN(
        P3_U2874) );
  AND2_X1 U20829 ( .A1(n18121), .A2(BUF2_REG_23__SCAN_IN), .ZN(n18168) );
  NOR2_X2 U20830 ( .A1(n17896), .A2(n17776), .ZN(n18166) );
  AOI22_X1 U20831 ( .A1(n18168), .A2(n18106), .B1(n18166), .B2(n17777), .ZN(
        n17782) );
  NOR2_X1 U20832 ( .A1(n17779), .A2(n17778), .ZN(n17802) );
  NOR2_X2 U20833 ( .A1(n18090), .A2(n17780), .ZN(n18169) );
  AOI22_X1 U20834 ( .A1(n17802), .A2(n17846), .B1(n18169), .B2(n18167), .ZN(
        n17781) );
  OAI211_X1 U20835 ( .C1(n17784), .C2(n17783), .A(n17782), .B(n17781), .ZN(
        P3_U2875) );
  INV_X1 U20836 ( .A(n18088), .ZN(n18125) );
  NAND2_X1 U20837 ( .A1(n17987), .A2(n18246), .ZN(n17964) );
  NOR2_X1 U20838 ( .A1(n17807), .A2(n17964), .ZN(n17803) );
  AOI22_X1 U20839 ( .A1(n18117), .A2(n18159), .B1(n18116), .B2(n17803), .ZN(
        n17787) );
  NOR2_X1 U20840 ( .A1(n17896), .A2(n17785), .ZN(n18118) );
  INV_X1 U20841 ( .A(n18118), .ZN(n17828) );
  NOR2_X1 U20842 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n17828), .ZN(
        n17873) );
  AOI22_X1 U20843 ( .A1(n18121), .A2(n18119), .B1(n17829), .B2(n17873), .ZN(
        n17804) );
  NAND2_X1 U20844 ( .A1(n17987), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n17963) );
  NOR2_X2 U20845 ( .A1(n17963), .A2(n17807), .ZN(n17868) );
  AOI22_X1 U20846 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n17804), .B1(
        n18122), .B2(n17868), .ZN(n17786) );
  OAI211_X1 U20847 ( .C1(n18125), .C2(n18115), .A(n17787), .B(n17786), .ZN(
        P3_U2876) );
  INV_X1 U20848 ( .A(n17868), .ZN(n17862) );
  AOI22_X1 U20849 ( .A1(n18127), .A2(n18106), .B1(n18126), .B2(n17803), .ZN(
        n17790) );
  AOI22_X1 U20850 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n17804), .B1(
        n18128), .B2(n18159), .ZN(n17789) );
  OAI211_X1 U20851 ( .C1(n18131), .C2(n17862), .A(n17790), .B(n17789), .ZN(
        P3_U2877) );
  AOI22_X1 U20852 ( .A1(n18133), .A2(n18106), .B1(n18132), .B2(n17803), .ZN(
        n17792) );
  AOI22_X1 U20853 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n17804), .B1(
        n18134), .B2(n17868), .ZN(n17791) );
  OAI211_X1 U20854 ( .C1(n18137), .C2(n18174), .A(n17792), .B(n17791), .ZN(
        P3_U2878) );
  AOI22_X1 U20855 ( .A1(n18139), .A2(n18106), .B1(n18138), .B2(n17803), .ZN(
        n17794) );
  AOI22_X1 U20856 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n17804), .B1(
        n18140), .B2(n17868), .ZN(n17793) );
  OAI211_X1 U20857 ( .C1(n18143), .C2(n18174), .A(n17794), .B(n17793), .ZN(
        P3_U2879) );
  AOI22_X1 U20858 ( .A1(n18145), .A2(n18106), .B1(n18144), .B2(n17803), .ZN(
        n17796) );
  AOI22_X1 U20859 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n17804), .B1(
        n18146), .B2(n17868), .ZN(n17795) );
  OAI211_X1 U20860 ( .C1(n18150), .C2(n18174), .A(n17796), .B(n17795), .ZN(
        P3_U2880) );
  AOI22_X1 U20861 ( .A1(n18153), .A2(n18159), .B1(n18151), .B2(n17803), .ZN(
        n17799) );
  AOI22_X1 U20862 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n17804), .B1(
        n18152), .B2(n18106), .ZN(n17798) );
  OAI211_X1 U20863 ( .C1(n18156), .C2(n17862), .A(n17799), .B(n17798), .ZN(
        P3_U2881) );
  AOI22_X1 U20864 ( .A1(n18004), .A2(n18106), .B1(n18158), .B2(n17803), .ZN(
        n17801) );
  AOI22_X1 U20865 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n17804), .B1(
        n18160), .B2(n17868), .ZN(n17800) );
  OAI211_X1 U20866 ( .C1(n18007), .C2(n18174), .A(n17801), .B(n17800), .ZN(
        P3_U2882) );
  INV_X1 U20867 ( .A(n17802), .ZN(n18175) );
  AOI22_X1 U20868 ( .A1(n18169), .A2(n18106), .B1(n18166), .B2(n17803), .ZN(
        n17806) );
  AOI22_X1 U20869 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n17804), .B1(
        n18168), .B2(n18159), .ZN(n17805) );
  OAI211_X1 U20870 ( .C1(n18175), .C2(n17862), .A(n17806), .B(n17805), .ZN(
        P3_U2883) );
  NOR2_X1 U20871 ( .A1(n17987), .A2(n17807), .ZN(n17874) );
  NAND2_X1 U20872 ( .A1(n17988), .A2(n17874), .ZN(n17881) );
  NOR2_X1 U20873 ( .A1(n17868), .A2(n17891), .ZN(n17850) );
  NOR2_X1 U20874 ( .A1(n18087), .A2(n17850), .ZN(n17824) );
  AOI22_X1 U20875 ( .A1(n18117), .A2(n17846), .B1(n18116), .B2(n17824), .ZN(
        n17811) );
  OAI21_X1 U20876 ( .B1(n17808), .B2(n18035), .A(n17850), .ZN(n17809) );
  OAI211_X1 U20877 ( .C1(n17891), .C2(n18339), .A(n18037), .B(n17809), .ZN(
        n17825) );
  AOI22_X1 U20878 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n17825), .B1(
        n18122), .B2(n17891), .ZN(n17810) );
  OAI211_X1 U20879 ( .C1(n18125), .C2(n18174), .A(n17811), .B(n17810), .ZN(
        P3_U2884) );
  AOI22_X1 U20880 ( .A1(n18128), .A2(n17846), .B1(n18126), .B2(n17824), .ZN(
        n17813) );
  AOI22_X1 U20881 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17825), .B1(
        n18127), .B2(n18159), .ZN(n17812) );
  OAI211_X1 U20882 ( .C1(n18131), .C2(n17881), .A(n17813), .B(n17812), .ZN(
        P3_U2885) );
  INV_X1 U20883 ( .A(n18133), .ZN(n18068) );
  AOI22_X1 U20884 ( .A1(n18065), .A2(n17846), .B1(n18132), .B2(n17824), .ZN(
        n17815) );
  AOI22_X1 U20885 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n17825), .B1(
        n18134), .B2(n17891), .ZN(n17814) );
  OAI211_X1 U20886 ( .C1(n18068), .C2(n18174), .A(n17815), .B(n17814), .ZN(
        P3_U2886) );
  INV_X1 U20887 ( .A(n18139), .ZN(n18072) );
  AOI22_X1 U20888 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n17825), .B1(
        n18138), .B2(n17824), .ZN(n17817) );
  AOI22_X1 U20889 ( .A1(n18140), .A2(n17891), .B1(n18069), .B2(n17846), .ZN(
        n17816) );
  OAI211_X1 U20890 ( .C1(n18072), .C2(n18174), .A(n17817), .B(n17816), .ZN(
        P3_U2887) );
  INV_X1 U20891 ( .A(n18145), .ZN(n18076) );
  AOI22_X1 U20892 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n17825), .B1(
        n18144), .B2(n17824), .ZN(n17819) );
  AOI22_X1 U20893 ( .A1(n18146), .A2(n17891), .B1(n18073), .B2(n17846), .ZN(
        n17818) );
  OAI211_X1 U20894 ( .C1(n18076), .C2(n18174), .A(n17819), .B(n17818), .ZN(
        P3_U2888) );
  AOI22_X1 U20895 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n17825), .B1(
        n18151), .B2(n17824), .ZN(n17821) );
  AOI22_X1 U20896 ( .A1(n18153), .A2(n17846), .B1(n18152), .B2(n18159), .ZN(
        n17820) );
  OAI211_X1 U20897 ( .C1(n18156), .C2(n17881), .A(n17821), .B(n17820), .ZN(
        P3_U2889) );
  AOI22_X1 U20898 ( .A1(n18004), .A2(n18159), .B1(n18158), .B2(n17824), .ZN(
        n17823) );
  AOI22_X1 U20899 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n17825), .B1(
        n18160), .B2(n17891), .ZN(n17822) );
  OAI211_X1 U20900 ( .C1(n18007), .C2(n17836), .A(n17823), .B(n17822), .ZN(
        P3_U2890) );
  AOI22_X1 U20901 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n17825), .B1(
        n18166), .B2(n17824), .ZN(n17827) );
  AOI22_X1 U20902 ( .A1(n18168), .A2(n17846), .B1(n18169), .B2(n18159), .ZN(
        n17826) );
  OAI211_X1 U20903 ( .C1(n18175), .C2(n17881), .A(n17827), .B(n17826), .ZN(
        P3_U2891) );
  NAND2_X1 U20904 ( .A1(n18191), .A2(n17829), .ZN(n17914) );
  AND2_X1 U20905 ( .A1(n18246), .A2(n17874), .ZN(n17845) );
  AOI22_X1 U20906 ( .A1(n18088), .A2(n17846), .B1(n18116), .B2(n17845), .ZN(
        n17831) );
  AOI21_X1 U20907 ( .B1(n17987), .B2(n18035), .A(n17828), .ZN(n17921) );
  NAND2_X1 U20908 ( .A1(n17829), .A2(n17921), .ZN(n17847) );
  AOI22_X1 U20909 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n17847), .B1(
        n18117), .B2(n17868), .ZN(n17830) );
  OAI211_X1 U20910 ( .C1(n18095), .C2(n17914), .A(n17831), .B(n17830), .ZN(
        P3_U2892) );
  AOI22_X1 U20911 ( .A1(n18128), .A2(n17868), .B1(n18126), .B2(n17845), .ZN(
        n17833) );
  AOI22_X1 U20912 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n17847), .B1(
        n18127), .B2(n17846), .ZN(n17832) );
  OAI211_X1 U20913 ( .C1(n18131), .C2(n17914), .A(n17833), .B(n17832), .ZN(
        P3_U2893) );
  AOI22_X1 U20914 ( .A1(n18065), .A2(n17868), .B1(n18132), .B2(n17845), .ZN(
        n17835) );
  INV_X1 U20915 ( .A(n17914), .ZN(n17916) );
  AOI22_X1 U20916 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n17847), .B1(
        n18134), .B2(n17916), .ZN(n17834) );
  OAI211_X1 U20917 ( .C1(n18068), .C2(n17836), .A(n17835), .B(n17834), .ZN(
        P3_U2894) );
  AOI22_X1 U20918 ( .A1(n18139), .A2(n17846), .B1(n18138), .B2(n17845), .ZN(
        n17838) );
  AOI22_X1 U20919 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n17847), .B1(
        n18140), .B2(n17916), .ZN(n17837) );
  OAI211_X1 U20920 ( .C1(n18143), .C2(n17862), .A(n17838), .B(n17837), .ZN(
        P3_U2895) );
  AOI22_X1 U20921 ( .A1(n18145), .A2(n17846), .B1(n18144), .B2(n17845), .ZN(
        n17840) );
  AOI22_X1 U20922 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n17847), .B1(
        n18146), .B2(n17916), .ZN(n17839) );
  OAI211_X1 U20923 ( .C1(n18150), .C2(n17862), .A(n17840), .B(n17839), .ZN(
        P3_U2896) );
  AOI22_X1 U20924 ( .A1(n18153), .A2(n17868), .B1(n18151), .B2(n17845), .ZN(
        n17842) );
  AOI22_X1 U20925 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n17847), .B1(
        n18152), .B2(n17846), .ZN(n17841) );
  OAI211_X1 U20926 ( .C1(n18156), .C2(n17914), .A(n17842), .B(n17841), .ZN(
        P3_U2897) );
  AOI22_X1 U20927 ( .A1(n18004), .A2(n17846), .B1(n18158), .B2(n17845), .ZN(
        n17844) );
  AOI22_X1 U20928 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n17847), .B1(
        n18160), .B2(n17916), .ZN(n17843) );
  OAI211_X1 U20929 ( .C1(n18007), .C2(n17862), .A(n17844), .B(n17843), .ZN(
        P3_U2898) );
  AOI22_X1 U20930 ( .A1(n18169), .A2(n17846), .B1(n18166), .B2(n17845), .ZN(
        n17849) );
  AOI22_X1 U20931 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n17847), .B1(
        n18168), .B2(n17868), .ZN(n17848) );
  OAI211_X1 U20932 ( .C1(n18175), .C2(n17914), .A(n17849), .B(n17848), .ZN(
        P3_U2899) );
  NAND2_X1 U20933 ( .A1(n18192), .A2(n17920), .ZN(n17905) );
  NOR2_X1 U20934 ( .A1(n17916), .A2(n17937), .ZN(n17897) );
  NOR2_X1 U20935 ( .A1(n18087), .A2(n17897), .ZN(n17867) );
  AOI22_X1 U20936 ( .A1(n18088), .A2(n17868), .B1(n18116), .B2(n17867), .ZN(
        n17853) );
  OAI22_X1 U20937 ( .A1(n17850), .A2(n18090), .B1(n17897), .B2(n17896), .ZN(
        n17851) );
  OAI21_X1 U20938 ( .B1(n17937), .B2(n18339), .A(n17851), .ZN(n17869) );
  AOI22_X1 U20939 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n17869), .B1(
        n18117), .B2(n17891), .ZN(n17852) );
  OAI211_X1 U20940 ( .C1(n18095), .C2(n17905), .A(n17853), .B(n17852), .ZN(
        P3_U2900) );
  AOI22_X1 U20941 ( .A1(n18128), .A2(n17891), .B1(n18126), .B2(n17867), .ZN(
        n17855) );
  AOI22_X1 U20942 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n17869), .B1(
        n18127), .B2(n17868), .ZN(n17854) );
  OAI211_X1 U20943 ( .C1(n18131), .C2(n17905), .A(n17855), .B(n17854), .ZN(
        P3_U2901) );
  AOI22_X1 U20944 ( .A1(n18133), .A2(n17868), .B1(n18132), .B2(n17867), .ZN(
        n17857) );
  AOI22_X1 U20945 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n17869), .B1(
        n18134), .B2(n17937), .ZN(n17856) );
  OAI211_X1 U20946 ( .C1(n18137), .C2(n17881), .A(n17857), .B(n17856), .ZN(
        P3_U2902) );
  AOI22_X1 U20947 ( .A1(n18138), .A2(n17867), .B1(n18069), .B2(n17891), .ZN(
        n17859) );
  AOI22_X1 U20948 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n17869), .B1(
        n18140), .B2(n17937), .ZN(n17858) );
  OAI211_X1 U20949 ( .C1(n18072), .C2(n17862), .A(n17859), .B(n17858), .ZN(
        P3_U2903) );
  AOI22_X1 U20950 ( .A1(n18073), .A2(n17891), .B1(n18144), .B2(n17867), .ZN(
        n17861) );
  AOI22_X1 U20951 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n17869), .B1(
        n18146), .B2(n17937), .ZN(n17860) );
  OAI211_X1 U20952 ( .C1(n18076), .C2(n17862), .A(n17861), .B(n17860), .ZN(
        P3_U2904) );
  AOI22_X1 U20953 ( .A1(n18153), .A2(n17891), .B1(n18151), .B2(n17867), .ZN(
        n17864) );
  AOI22_X1 U20954 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n17869), .B1(
        n18152), .B2(n17868), .ZN(n17863) );
  OAI211_X1 U20955 ( .C1(n18156), .C2(n17905), .A(n17864), .B(n17863), .ZN(
        P3_U2905) );
  AOI22_X1 U20956 ( .A1(n18004), .A2(n17868), .B1(n18158), .B2(n17867), .ZN(
        n17866) );
  AOI22_X1 U20957 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n17869), .B1(
        n18160), .B2(n17937), .ZN(n17865) );
  OAI211_X1 U20958 ( .C1(n18007), .C2(n17881), .A(n17866), .B(n17865), .ZN(
        P3_U2906) );
  AOI22_X1 U20959 ( .A1(n18168), .A2(n17891), .B1(n18166), .B2(n17867), .ZN(
        n17871) );
  AOI22_X1 U20960 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n17869), .B1(
        n18169), .B2(n17868), .ZN(n17870) );
  OAI211_X1 U20961 ( .C1(n18175), .C2(n17905), .A(n17871), .B(n17870), .ZN(
        P3_U2907) );
  NOR2_X2 U20962 ( .A1(n17963), .A2(n17872), .ZN(n17959) );
  INV_X1 U20963 ( .A(n17959), .ZN(n17957) );
  NOR2_X1 U20964 ( .A1(n17964), .A2(n17872), .ZN(n17890) );
  AOI22_X1 U20965 ( .A1(n18117), .A2(n17916), .B1(n18116), .B2(n17890), .ZN(
        n17876) );
  AOI22_X1 U20966 ( .A1(n18121), .A2(n17874), .B1(n17873), .B2(n17920), .ZN(
        n17892) );
  AOI22_X1 U20967 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n17892), .B1(
        n18088), .B2(n17891), .ZN(n17875) );
  OAI211_X1 U20968 ( .C1(n18095), .C2(n17957), .A(n17876), .B(n17875), .ZN(
        P3_U2908) );
  AOI22_X1 U20969 ( .A1(n18127), .A2(n17891), .B1(n18126), .B2(n17890), .ZN(
        n17878) );
  AOI22_X1 U20970 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n17892), .B1(
        n18128), .B2(n17916), .ZN(n17877) );
  OAI211_X1 U20971 ( .C1(n18131), .C2(n17957), .A(n17878), .B(n17877), .ZN(
        P3_U2909) );
  AOI22_X1 U20972 ( .A1(n18065), .A2(n17916), .B1(n18132), .B2(n17890), .ZN(
        n17880) );
  AOI22_X1 U20973 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n17892), .B1(
        n18134), .B2(n17959), .ZN(n17879) );
  OAI211_X1 U20974 ( .C1(n18068), .C2(n17881), .A(n17880), .B(n17879), .ZN(
        P3_U2910) );
  AOI22_X1 U20975 ( .A1(n18139), .A2(n17891), .B1(n18138), .B2(n17890), .ZN(
        n17883) );
  AOI22_X1 U20976 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n17892), .B1(
        n18140), .B2(n17959), .ZN(n17882) );
  OAI211_X1 U20977 ( .C1(n18143), .C2(n17914), .A(n17883), .B(n17882), .ZN(
        P3_U2911) );
  AOI22_X1 U20978 ( .A1(n18145), .A2(n17891), .B1(n18144), .B2(n17890), .ZN(
        n17885) );
  AOI22_X1 U20979 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n17892), .B1(
        n18146), .B2(n17959), .ZN(n17884) );
  OAI211_X1 U20980 ( .C1(n18150), .C2(n17914), .A(n17885), .B(n17884), .ZN(
        P3_U2912) );
  AOI22_X1 U20981 ( .A1(n18153), .A2(n17916), .B1(n18151), .B2(n17890), .ZN(
        n17887) );
  AOI22_X1 U20982 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n17892), .B1(
        n18152), .B2(n17891), .ZN(n17886) );
  OAI211_X1 U20983 ( .C1(n18156), .C2(n17957), .A(n17887), .B(n17886), .ZN(
        P3_U2913) );
  AOI22_X1 U20984 ( .A1(n18004), .A2(n17891), .B1(n18158), .B2(n17890), .ZN(
        n17889) );
  AOI22_X1 U20985 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n17892), .B1(
        n18160), .B2(n17959), .ZN(n17888) );
  OAI211_X1 U20986 ( .C1(n18007), .C2(n17914), .A(n17889), .B(n17888), .ZN(
        P3_U2914) );
  AOI22_X1 U20987 ( .A1(n18169), .A2(n17891), .B1(n18166), .B2(n17890), .ZN(
        n17894) );
  AOI22_X1 U20988 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n17892), .B1(
        n18168), .B2(n17916), .ZN(n17893) );
  OAI211_X1 U20989 ( .C1(n18175), .C2(n17957), .A(n17894), .B(n17893), .ZN(
        P3_U2915) );
  NOR2_X1 U20990 ( .A1(n17895), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n17965) );
  NAND2_X1 U20991 ( .A1(n17988), .A2(n17965), .ZN(n17980) );
  NOR2_X1 U20992 ( .A1(n17959), .A2(n17982), .ZN(n17941) );
  NOR2_X1 U20993 ( .A1(n18087), .A2(n17941), .ZN(n17915) );
  AOI22_X1 U20994 ( .A1(n18117), .A2(n17937), .B1(n18116), .B2(n17915), .ZN(
        n17900) );
  OAI22_X1 U20995 ( .A1(n17897), .A2(n18090), .B1(n17941), .B2(n17896), .ZN(
        n17898) );
  OAI21_X1 U20996 ( .B1(n17982), .B2(n18339), .A(n17898), .ZN(n17917) );
  AOI22_X1 U20997 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n17917), .B1(
        n18122), .B2(n17982), .ZN(n17899) );
  OAI211_X1 U20998 ( .C1(n18125), .C2(n17914), .A(n17900), .B(n17899), .ZN(
        P3_U2916) );
  AOI22_X1 U20999 ( .A1(n18127), .A2(n17916), .B1(n18126), .B2(n17915), .ZN(
        n17902) );
  AOI22_X1 U21000 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17917), .B1(
        n18128), .B2(n17937), .ZN(n17901) );
  OAI211_X1 U21001 ( .C1(n18131), .C2(n17980), .A(n17902), .B(n17901), .ZN(
        P3_U2917) );
  AOI22_X1 U21002 ( .A1(n18133), .A2(n17916), .B1(n18132), .B2(n17915), .ZN(
        n17904) );
  AOI22_X1 U21003 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n17917), .B1(
        n18134), .B2(n17982), .ZN(n17903) );
  OAI211_X1 U21004 ( .C1(n18137), .C2(n17905), .A(n17904), .B(n17903), .ZN(
        P3_U2918) );
  AOI22_X1 U21005 ( .A1(n18138), .A2(n17915), .B1(n18069), .B2(n17937), .ZN(
        n17907) );
  AOI22_X1 U21006 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n17917), .B1(
        n18140), .B2(n17982), .ZN(n17906) );
  OAI211_X1 U21007 ( .C1(n18072), .C2(n17914), .A(n17907), .B(n17906), .ZN(
        P3_U2919) );
  AOI22_X1 U21008 ( .A1(n18073), .A2(n17937), .B1(n18144), .B2(n17915), .ZN(
        n17909) );
  AOI22_X1 U21009 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n17917), .B1(
        n18146), .B2(n17982), .ZN(n17908) );
  OAI211_X1 U21010 ( .C1(n18076), .C2(n17914), .A(n17909), .B(n17908), .ZN(
        P3_U2920) );
  AOI22_X1 U21011 ( .A1(n18151), .A2(n17915), .B1(n18152), .B2(n17916), .ZN(
        n17911) );
  AOI22_X1 U21012 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n17917), .B1(
        n18153), .B2(n17937), .ZN(n17910) );
  OAI211_X1 U21013 ( .C1(n18156), .C2(n17980), .A(n17911), .B(n17910), .ZN(
        P3_U2921) );
  INV_X1 U21014 ( .A(n18004), .ZN(n18163) );
  AOI22_X1 U21015 ( .A1(n18158), .A2(n17915), .B1(n18157), .B2(n17937), .ZN(
        n17913) );
  AOI22_X1 U21016 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n17917), .B1(
        n18160), .B2(n17982), .ZN(n17912) );
  OAI211_X1 U21017 ( .C1(n18163), .C2(n17914), .A(n17913), .B(n17912), .ZN(
        P3_U2922) );
  AOI22_X1 U21018 ( .A1(n18168), .A2(n17937), .B1(n18166), .B2(n17915), .ZN(
        n17919) );
  AOI22_X1 U21019 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n17917), .B1(
        n18169), .B2(n17916), .ZN(n17918) );
  OAI211_X1 U21020 ( .C1(n18175), .C2(n17980), .A(n17919), .B(n17918), .ZN(
        P3_U2923) );
  NAND2_X1 U21021 ( .A1(n18191), .A2(n17920), .ZN(n18001) );
  AND2_X1 U21022 ( .A1(n18246), .A2(n17965), .ZN(n17936) );
  AOI22_X1 U21023 ( .A1(n18088), .A2(n17937), .B1(n18116), .B2(n17936), .ZN(
        n17923) );
  NAND2_X1 U21024 ( .A1(n17921), .A2(n17920), .ZN(n17938) );
  AOI22_X1 U21025 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n17938), .B1(
        n18117), .B2(n17959), .ZN(n17922) );
  OAI211_X1 U21026 ( .C1(n18095), .C2(n18001), .A(n17923), .B(n17922), .ZN(
        P3_U2924) );
  AOI22_X1 U21027 ( .A1(n18128), .A2(n17959), .B1(n18126), .B2(n17936), .ZN(
        n17925) );
  AOI22_X1 U21028 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n17938), .B1(
        n18127), .B2(n17937), .ZN(n17924) );
  OAI211_X1 U21029 ( .C1(n18131), .C2(n18001), .A(n17925), .B(n17924), .ZN(
        P3_U2925) );
  AOI22_X1 U21030 ( .A1(n18133), .A2(n17937), .B1(n18132), .B2(n17936), .ZN(
        n17927) );
  INV_X1 U21031 ( .A(n18001), .ZN(n18009) );
  AOI22_X1 U21032 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n17938), .B1(
        n18134), .B2(n18009), .ZN(n17926) );
  OAI211_X1 U21033 ( .C1(n18137), .C2(n17957), .A(n17927), .B(n17926), .ZN(
        P3_U2926) );
  AOI22_X1 U21034 ( .A1(n18139), .A2(n17937), .B1(n18138), .B2(n17936), .ZN(
        n17929) );
  AOI22_X1 U21035 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n17938), .B1(
        n18140), .B2(n18009), .ZN(n17928) );
  OAI211_X1 U21036 ( .C1(n18143), .C2(n17957), .A(n17929), .B(n17928), .ZN(
        P3_U2927) );
  AOI22_X1 U21037 ( .A1(n18145), .A2(n17937), .B1(n18144), .B2(n17936), .ZN(
        n17931) );
  AOI22_X1 U21038 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n17938), .B1(
        n18146), .B2(n18009), .ZN(n17930) );
  OAI211_X1 U21039 ( .C1(n18150), .C2(n17957), .A(n17931), .B(n17930), .ZN(
        P3_U2928) );
  AOI22_X1 U21040 ( .A1(n18151), .A2(n17936), .B1(n18152), .B2(n17937), .ZN(
        n17933) );
  AOI22_X1 U21041 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n17938), .B1(
        n18153), .B2(n17959), .ZN(n17932) );
  OAI211_X1 U21042 ( .C1(n18156), .C2(n18001), .A(n17933), .B(n17932), .ZN(
        P3_U2929) );
  AOI22_X1 U21043 ( .A1(n18004), .A2(n17937), .B1(n18158), .B2(n17936), .ZN(
        n17935) );
  AOI22_X1 U21044 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n17938), .B1(
        n18160), .B2(n18009), .ZN(n17934) );
  OAI211_X1 U21045 ( .C1(n18007), .C2(n17957), .A(n17935), .B(n17934), .ZN(
        P3_U2930) );
  AOI22_X1 U21046 ( .A1(n18169), .A2(n17937), .B1(n18166), .B2(n17936), .ZN(
        n17940) );
  AOI22_X1 U21047 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n17938), .B1(
        n18168), .B2(n17959), .ZN(n17939) );
  OAI211_X1 U21048 ( .C1(n18175), .C2(n18001), .A(n17940), .B(n17939), .ZN(
        P3_U2931) );
  NAND2_X1 U21049 ( .A1(n18192), .A2(n18013), .ZN(n18029) );
  NOR2_X1 U21050 ( .A1(n18009), .A2(n18031), .ZN(n17989) );
  NOR2_X1 U21051 ( .A1(n18087), .A2(n17989), .ZN(n17958) );
  AOI22_X1 U21052 ( .A1(n18088), .A2(n17959), .B1(n18116), .B2(n17958), .ZN(
        n17944) );
  OAI21_X1 U21053 ( .B1(n17941), .B2(n18035), .A(n17989), .ZN(n17942) );
  OAI211_X1 U21054 ( .C1(n18031), .C2(n18339), .A(n18037), .B(n17942), .ZN(
        n17960) );
  AOI22_X1 U21055 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n17960), .B1(
        n18117), .B2(n17982), .ZN(n17943) );
  OAI211_X1 U21056 ( .C1(n18095), .C2(n18029), .A(n17944), .B(n17943), .ZN(
        P3_U2932) );
  AOI22_X1 U21057 ( .A1(n18128), .A2(n17982), .B1(n18126), .B2(n17958), .ZN(
        n17946) );
  AOI22_X1 U21058 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n17960), .B1(
        n18127), .B2(n17959), .ZN(n17945) );
  OAI211_X1 U21059 ( .C1(n18131), .C2(n18029), .A(n17946), .B(n17945), .ZN(
        P3_U2933) );
  AOI22_X1 U21060 ( .A1(n18065), .A2(n17982), .B1(n18132), .B2(n17958), .ZN(
        n17948) );
  AOI22_X1 U21061 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n17960), .B1(
        n18134), .B2(n18031), .ZN(n17947) );
  OAI211_X1 U21062 ( .C1(n18068), .C2(n17957), .A(n17948), .B(n17947), .ZN(
        P3_U2934) );
  AOI22_X1 U21063 ( .A1(n18138), .A2(n17958), .B1(n18069), .B2(n17982), .ZN(
        n17950) );
  AOI22_X1 U21064 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n17960), .B1(
        n18140), .B2(n18031), .ZN(n17949) );
  OAI211_X1 U21065 ( .C1(n18072), .C2(n17957), .A(n17950), .B(n17949), .ZN(
        P3_U2935) );
  AOI22_X1 U21066 ( .A1(n18073), .A2(n17982), .B1(n18144), .B2(n17958), .ZN(
        n17952) );
  AOI22_X1 U21067 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n17960), .B1(
        n18146), .B2(n18031), .ZN(n17951) );
  OAI211_X1 U21068 ( .C1(n18076), .C2(n17957), .A(n17952), .B(n17951), .ZN(
        P3_U2936) );
  AOI22_X1 U21069 ( .A1(n18151), .A2(n17958), .B1(n18152), .B2(n17959), .ZN(
        n17954) );
  AOI22_X1 U21070 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n17960), .B1(
        n18153), .B2(n17982), .ZN(n17953) );
  OAI211_X1 U21071 ( .C1(n18156), .C2(n18029), .A(n17954), .B(n17953), .ZN(
        P3_U2937) );
  AOI22_X1 U21072 ( .A1(n18158), .A2(n17958), .B1(n18157), .B2(n17982), .ZN(
        n17956) );
  AOI22_X1 U21073 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n17960), .B1(
        n18160), .B2(n18031), .ZN(n17955) );
  OAI211_X1 U21074 ( .C1(n18163), .C2(n17957), .A(n17956), .B(n17955), .ZN(
        P3_U2938) );
  AOI22_X1 U21075 ( .A1(n18169), .A2(n17959), .B1(n18166), .B2(n17958), .ZN(
        n17962) );
  AOI22_X1 U21076 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n17960), .B1(
        n18168), .B2(n17982), .ZN(n17961) );
  OAI211_X1 U21077 ( .C1(n18175), .C2(n18029), .A(n17962), .B(n17961), .ZN(
        P3_U2939) );
  NOR2_X2 U21078 ( .A1(n17986), .A2(n17963), .ZN(n18055) );
  INV_X1 U21079 ( .A(n18055), .ZN(n18053) );
  NOR2_X1 U21080 ( .A1(n17986), .A2(n17964), .ZN(n17981) );
  AOI22_X1 U21081 ( .A1(n18088), .A2(n17982), .B1(n18116), .B2(n17981), .ZN(
        n17967) );
  NOR2_X1 U21082 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n17986), .ZN(
        n18014) );
  AOI22_X1 U21083 ( .A1(n18121), .A2(n17965), .B1(n18118), .B2(n18014), .ZN(
        n17983) );
  AOI22_X1 U21084 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n17983), .B1(
        n18117), .B2(n18009), .ZN(n17966) );
  OAI211_X1 U21085 ( .C1(n18053), .C2(n18095), .A(n17967), .B(n17966), .ZN(
        P3_U2940) );
  AOI22_X1 U21086 ( .A1(n18127), .A2(n17982), .B1(n18126), .B2(n17981), .ZN(
        n17969) );
  AOI22_X1 U21087 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n17983), .B1(
        n18128), .B2(n18009), .ZN(n17968) );
  OAI211_X1 U21088 ( .C1(n18053), .C2(n18131), .A(n17969), .B(n17968), .ZN(
        P3_U2941) );
  AOI22_X1 U21089 ( .A1(n18065), .A2(n18009), .B1(n18132), .B2(n17981), .ZN(
        n17971) );
  AOI22_X1 U21090 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n17983), .B1(
        n18055), .B2(n18134), .ZN(n17970) );
  OAI211_X1 U21091 ( .C1(n18068), .C2(n17980), .A(n17971), .B(n17970), .ZN(
        P3_U2942) );
  AOI22_X1 U21092 ( .A1(n18138), .A2(n17981), .B1(n18069), .B2(n18009), .ZN(
        n17973) );
  AOI22_X1 U21093 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n17983), .B1(
        n18055), .B2(n18140), .ZN(n17972) );
  OAI211_X1 U21094 ( .C1(n18072), .C2(n17980), .A(n17973), .B(n17972), .ZN(
        P3_U2943) );
  AOI22_X1 U21095 ( .A1(n18145), .A2(n17982), .B1(n18144), .B2(n17981), .ZN(
        n17975) );
  AOI22_X1 U21096 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n17983), .B1(
        n18055), .B2(n18146), .ZN(n17974) );
  OAI211_X1 U21097 ( .C1(n18150), .C2(n18001), .A(n17975), .B(n17974), .ZN(
        P3_U2944) );
  AOI22_X1 U21098 ( .A1(n18151), .A2(n17981), .B1(n18152), .B2(n17982), .ZN(
        n17977) );
  AOI22_X1 U21099 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n17983), .B1(
        n18153), .B2(n18009), .ZN(n17976) );
  OAI211_X1 U21100 ( .C1(n18053), .C2(n18156), .A(n17977), .B(n17976), .ZN(
        P3_U2945) );
  AOI22_X1 U21101 ( .A1(n18158), .A2(n17981), .B1(n18157), .B2(n18009), .ZN(
        n17979) );
  AOI22_X1 U21102 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n17983), .B1(
        n18055), .B2(n18160), .ZN(n17978) );
  OAI211_X1 U21103 ( .C1(n18163), .C2(n17980), .A(n17979), .B(n17978), .ZN(
        P3_U2946) );
  AOI22_X1 U21104 ( .A1(n18169), .A2(n17982), .B1(n18166), .B2(n17981), .ZN(
        n17985) );
  AOI22_X1 U21105 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n17983), .B1(
        n18168), .B2(n18009), .ZN(n17984) );
  OAI211_X1 U21106 ( .C1(n18053), .C2(n18175), .A(n17985), .B(n17984), .ZN(
        P3_U2947) );
  NOR2_X1 U21107 ( .A1(n17987), .A2(n17986), .ZN(n18060) );
  NAND2_X1 U21108 ( .A1(n17988), .A2(n18060), .ZN(n18081) );
  NOR2_X1 U21109 ( .A1(n18055), .A2(n18083), .ZN(n18036) );
  NOR2_X1 U21110 ( .A1(n18087), .A2(n18036), .ZN(n18008) );
  AOI22_X1 U21111 ( .A1(n18088), .A2(n18009), .B1(n18116), .B2(n18008), .ZN(
        n17992) );
  OAI21_X1 U21112 ( .B1(n17989), .B2(n18035), .A(n18036), .ZN(n17990) );
  OAI211_X1 U21113 ( .C1(n18083), .C2(n18339), .A(n18037), .B(n17990), .ZN(
        n18010) );
  AOI22_X1 U21114 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18010), .B1(
        n18117), .B2(n18031), .ZN(n17991) );
  OAI211_X1 U21115 ( .C1(n18081), .C2(n18095), .A(n17992), .B(n17991), .ZN(
        P3_U2948) );
  AOI22_X1 U21116 ( .A1(n18127), .A2(n18009), .B1(n18126), .B2(n18008), .ZN(
        n17994) );
  AOI22_X1 U21117 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18010), .B1(
        n18128), .B2(n18031), .ZN(n17993) );
  OAI211_X1 U21118 ( .C1(n18081), .C2(n18131), .A(n17994), .B(n17993), .ZN(
        P3_U2949) );
  AOI22_X1 U21119 ( .A1(n18065), .A2(n18031), .B1(n18132), .B2(n18008), .ZN(
        n17996) );
  AOI22_X1 U21120 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18010), .B1(
        n18083), .B2(n18134), .ZN(n17995) );
  OAI211_X1 U21121 ( .C1(n18068), .C2(n18001), .A(n17996), .B(n17995), .ZN(
        P3_U2950) );
  AOI22_X1 U21122 ( .A1(n18139), .A2(n18009), .B1(n18138), .B2(n18008), .ZN(
        n17998) );
  AOI22_X1 U21123 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18010), .B1(
        n18083), .B2(n18140), .ZN(n17997) );
  OAI211_X1 U21124 ( .C1(n18143), .C2(n18029), .A(n17998), .B(n17997), .ZN(
        P3_U2951) );
  AOI22_X1 U21125 ( .A1(n18073), .A2(n18031), .B1(n18144), .B2(n18008), .ZN(
        n18000) );
  AOI22_X1 U21126 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18010), .B1(
        n18083), .B2(n18146), .ZN(n17999) );
  OAI211_X1 U21127 ( .C1(n18076), .C2(n18001), .A(n18000), .B(n17999), .ZN(
        P3_U2952) );
  AOI22_X1 U21128 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18010), .B1(
        n18151), .B2(n18008), .ZN(n18003) );
  AOI22_X1 U21129 ( .A1(n18153), .A2(n18031), .B1(n18152), .B2(n18009), .ZN(
        n18002) );
  OAI211_X1 U21130 ( .C1(n18081), .C2(n18156), .A(n18003), .B(n18002), .ZN(
        P3_U2953) );
  AOI22_X1 U21131 ( .A1(n18004), .A2(n18009), .B1(n18158), .B2(n18008), .ZN(
        n18006) );
  AOI22_X1 U21132 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18010), .B1(
        n18083), .B2(n18160), .ZN(n18005) );
  OAI211_X1 U21133 ( .C1(n18007), .C2(n18029), .A(n18006), .B(n18005), .ZN(
        P3_U2954) );
  AOI22_X1 U21134 ( .A1(n18168), .A2(n18031), .B1(n18166), .B2(n18008), .ZN(
        n18012) );
  AOI22_X1 U21135 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18010), .B1(
        n18169), .B2(n18009), .ZN(n18011) );
  OAI211_X1 U21136 ( .C1(n18081), .C2(n18175), .A(n18012), .B(n18011), .ZN(
        P3_U2955) );
  NAND2_X1 U21137 ( .A1(n18191), .A2(n18013), .ZN(n18109) );
  AND2_X1 U21138 ( .A1(n18246), .A2(n18060), .ZN(n18030) );
  AOI22_X1 U21139 ( .A1(n18088), .A2(n18031), .B1(n18116), .B2(n18030), .ZN(
        n18016) );
  AOI22_X1 U21140 ( .A1(n18121), .A2(n18014), .B1(n18060), .B2(n18118), .ZN(
        n18032) );
  AOI22_X1 U21141 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18032), .B1(
        n18055), .B2(n18117), .ZN(n18015) );
  OAI211_X1 U21142 ( .C1(n18109), .C2(n18095), .A(n18016), .B(n18015), .ZN(
        P3_U2956) );
  AOI22_X1 U21143 ( .A1(n18127), .A2(n18031), .B1(n18126), .B2(n18030), .ZN(
        n18018) );
  AOI22_X1 U21144 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18032), .B1(
        n18055), .B2(n18128), .ZN(n18017) );
  OAI211_X1 U21145 ( .C1(n18109), .C2(n18131), .A(n18018), .B(n18017), .ZN(
        P3_U2957) );
  AOI22_X1 U21146 ( .A1(n18133), .A2(n18031), .B1(n18132), .B2(n18030), .ZN(
        n18020) );
  INV_X1 U21147 ( .A(n18109), .ZN(n18111) );
  AOI22_X1 U21148 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18032), .B1(
        n18111), .B2(n18134), .ZN(n18019) );
  OAI211_X1 U21149 ( .C1(n18053), .C2(n18137), .A(n18020), .B(n18019), .ZN(
        P3_U2958) );
  AOI22_X1 U21150 ( .A1(n18055), .A2(n18069), .B1(n18138), .B2(n18030), .ZN(
        n18022) );
  AOI22_X1 U21151 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18032), .B1(
        n18111), .B2(n18140), .ZN(n18021) );
  OAI211_X1 U21152 ( .C1(n18072), .C2(n18029), .A(n18022), .B(n18021), .ZN(
        P3_U2959) );
  AOI22_X1 U21153 ( .A1(n18055), .A2(n18073), .B1(n18144), .B2(n18030), .ZN(
        n18024) );
  AOI22_X1 U21154 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18032), .B1(
        n18111), .B2(n18146), .ZN(n18023) );
  OAI211_X1 U21155 ( .C1(n18076), .C2(n18029), .A(n18024), .B(n18023), .ZN(
        P3_U2960) );
  AOI22_X1 U21156 ( .A1(n18055), .A2(n18153), .B1(n18151), .B2(n18030), .ZN(
        n18026) );
  AOI22_X1 U21157 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18032), .B1(
        n18152), .B2(n18031), .ZN(n18025) );
  OAI211_X1 U21158 ( .C1(n18109), .C2(n18156), .A(n18026), .B(n18025), .ZN(
        P3_U2961) );
  AOI22_X1 U21159 ( .A1(n18055), .A2(n18157), .B1(n18158), .B2(n18030), .ZN(
        n18028) );
  AOI22_X1 U21160 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18032), .B1(
        n18111), .B2(n18160), .ZN(n18027) );
  OAI211_X1 U21161 ( .C1(n18163), .C2(n18029), .A(n18028), .B(n18027), .ZN(
        P3_U2962) );
  AOI22_X1 U21162 ( .A1(n18169), .A2(n18031), .B1(n18166), .B2(n18030), .ZN(
        n18034) );
  AOI22_X1 U21163 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18032), .B1(
        n18055), .B2(n18168), .ZN(n18033) );
  OAI211_X1 U21164 ( .C1(n18109), .C2(n18175), .A(n18034), .B(n18033), .ZN(
        P3_U2963) );
  NOR2_X2 U21165 ( .A1(n18059), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18170) );
  INV_X1 U21166 ( .A(n18170), .ZN(n18164) );
  AOI21_X1 U21167 ( .B1(n18164), .B2(n18109), .A(n18087), .ZN(n18054) );
  AOI22_X1 U21168 ( .A1(n18083), .A2(n18117), .B1(n18116), .B2(n18054), .ZN(
        n18040) );
  AOI221_X1 U21169 ( .B1(n18036), .B2(n18109), .C1(n18035), .C2(n18109), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18038) );
  OAI21_X1 U21170 ( .B1(n18170), .B2(n18038), .A(n18037), .ZN(n18056) );
  AOI22_X1 U21171 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18056), .B1(
        n18170), .B2(n18122), .ZN(n18039) );
  OAI211_X1 U21172 ( .C1(n18125), .C2(n18053), .A(n18040), .B(n18039), .ZN(
        P3_U2964) );
  AOI22_X1 U21173 ( .A1(n18055), .A2(n18127), .B1(n18054), .B2(n18126), .ZN(
        n18042) );
  AOI22_X1 U21174 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18056), .B1(
        n18083), .B2(n18128), .ZN(n18041) );
  OAI211_X1 U21175 ( .C1(n18164), .C2(n18131), .A(n18042), .B(n18041), .ZN(
        P3_U2965) );
  AOI22_X1 U21176 ( .A1(n18083), .A2(n18065), .B1(n18054), .B2(n18132), .ZN(
        n18044) );
  AOI22_X1 U21177 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18056), .B1(
        n18170), .B2(n18134), .ZN(n18043) );
  OAI211_X1 U21178 ( .C1(n18053), .C2(n18068), .A(n18044), .B(n18043), .ZN(
        P3_U2966) );
  AOI22_X1 U21179 ( .A1(n18083), .A2(n18069), .B1(n18054), .B2(n18138), .ZN(
        n18046) );
  AOI22_X1 U21180 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18056), .B1(
        n18170), .B2(n18140), .ZN(n18045) );
  OAI211_X1 U21181 ( .C1(n18053), .C2(n18072), .A(n18046), .B(n18045), .ZN(
        P3_U2967) );
  AOI22_X1 U21182 ( .A1(n18083), .A2(n18073), .B1(n18054), .B2(n18144), .ZN(
        n18048) );
  AOI22_X1 U21183 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18056), .B1(
        n18170), .B2(n18146), .ZN(n18047) );
  OAI211_X1 U21184 ( .C1(n18053), .C2(n18076), .A(n18048), .B(n18047), .ZN(
        P3_U2968) );
  AOI22_X1 U21185 ( .A1(n18055), .A2(n18152), .B1(n18054), .B2(n18151), .ZN(
        n18050) );
  AOI22_X1 U21186 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18056), .B1(
        n18083), .B2(n18153), .ZN(n18049) );
  OAI211_X1 U21187 ( .C1(n18164), .C2(n18156), .A(n18050), .B(n18049), .ZN(
        P3_U2969) );
  AOI22_X1 U21188 ( .A1(n18083), .A2(n18157), .B1(n18054), .B2(n18158), .ZN(
        n18052) );
  AOI22_X1 U21189 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18056), .B1(
        n18170), .B2(n18160), .ZN(n18051) );
  OAI211_X1 U21190 ( .C1(n18053), .C2(n18163), .A(n18052), .B(n18051), .ZN(
        P3_U2970) );
  AOI22_X1 U21191 ( .A1(n18055), .A2(n18169), .B1(n18054), .B2(n18166), .ZN(
        n18058) );
  AOI22_X1 U21192 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18056), .B1(
        n18083), .B2(n18168), .ZN(n18057) );
  OAI211_X1 U21193 ( .C1(n18164), .C2(n18175), .A(n18058), .B(n18057), .ZN(
        P3_U2971) );
  NOR2_X1 U21194 ( .A1(n18087), .A2(n18059), .ZN(n18082) );
  AOI22_X1 U21195 ( .A1(n18088), .A2(n18083), .B1(n18116), .B2(n18082), .ZN(
        n18062) );
  AOI22_X1 U21196 ( .A1(n18121), .A2(n18060), .B1(n18120), .B2(n18118), .ZN(
        n18084) );
  AOI22_X1 U21197 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18084), .B1(
        n18111), .B2(n18117), .ZN(n18061) );
  OAI211_X1 U21198 ( .C1(n18095), .C2(n18149), .A(n18062), .B(n18061), .ZN(
        P3_U2972) );
  AOI22_X1 U21199 ( .A1(n18083), .A2(n18127), .B1(n18126), .B2(n18082), .ZN(
        n18064) );
  AOI22_X1 U21200 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18084), .B1(
        n18111), .B2(n18128), .ZN(n18063) );
  OAI211_X1 U21201 ( .C1(n18131), .C2(n18149), .A(n18064), .B(n18063), .ZN(
        P3_U2973) );
  AOI22_X1 U21202 ( .A1(n18111), .A2(n18065), .B1(n18132), .B2(n18082), .ZN(
        n18067) );
  AOI22_X1 U21203 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18084), .B1(
        n18134), .B2(n18167), .ZN(n18066) );
  OAI211_X1 U21204 ( .C1(n18081), .C2(n18068), .A(n18067), .B(n18066), .ZN(
        P3_U2974) );
  AOI22_X1 U21205 ( .A1(n18111), .A2(n18069), .B1(n18138), .B2(n18082), .ZN(
        n18071) );
  AOI22_X1 U21206 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18084), .B1(
        n18140), .B2(n18167), .ZN(n18070) );
  OAI211_X1 U21207 ( .C1(n18081), .C2(n18072), .A(n18071), .B(n18070), .ZN(
        P3_U2975) );
  AOI22_X1 U21208 ( .A1(n18111), .A2(n18073), .B1(n18144), .B2(n18082), .ZN(
        n18075) );
  AOI22_X1 U21209 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18084), .B1(
        n18146), .B2(n18167), .ZN(n18074) );
  OAI211_X1 U21210 ( .C1(n18081), .C2(n18076), .A(n18075), .B(n18074), .ZN(
        P3_U2976) );
  AOI22_X1 U21211 ( .A1(n18111), .A2(n18153), .B1(n18151), .B2(n18082), .ZN(
        n18078) );
  AOI22_X1 U21212 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18084), .B1(
        n18083), .B2(n18152), .ZN(n18077) );
  OAI211_X1 U21213 ( .C1(n18156), .C2(n18149), .A(n18078), .B(n18077), .ZN(
        P3_U2977) );
  AOI22_X1 U21214 ( .A1(n18111), .A2(n18157), .B1(n18158), .B2(n18082), .ZN(
        n18080) );
  AOI22_X1 U21215 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18084), .B1(
        n18160), .B2(n18167), .ZN(n18079) );
  OAI211_X1 U21216 ( .C1(n18081), .C2(n18163), .A(n18080), .B(n18079), .ZN(
        P3_U2978) );
  AOI22_X1 U21217 ( .A1(n18083), .A2(n18169), .B1(n18166), .B2(n18082), .ZN(
        n18086) );
  AOI22_X1 U21218 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18084), .B1(
        n18111), .B2(n18168), .ZN(n18085) );
  OAI211_X1 U21219 ( .C1(n18175), .C2(n18149), .A(n18086), .B(n18085), .ZN(
        P3_U2979) );
  AOI21_X1 U21220 ( .B1(n18115), .B2(n18149), .A(n18087), .ZN(n18110) );
  AOI22_X1 U21221 ( .A1(n18088), .A2(n18111), .B1(n18116), .B2(n18110), .ZN(
        n18094) );
  NOR2_X1 U21222 ( .A1(n18170), .A2(n18111), .ZN(n18091) );
  OAI21_X1 U21223 ( .B1(n18091), .B2(n18090), .A(n18089), .ZN(n18092) );
  OAI21_X1 U21224 ( .B1(n18106), .B2(n18339), .A(n18092), .ZN(n18112) );
  AOI22_X1 U21225 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18112), .B1(
        n18170), .B2(n18117), .ZN(n18093) );
  OAI211_X1 U21226 ( .C1(n18095), .C2(n18115), .A(n18094), .B(n18093), .ZN(
        P3_U2980) );
  AOI22_X1 U21227 ( .A1(n18111), .A2(n18127), .B1(n18126), .B2(n18110), .ZN(
        n18097) );
  AOI22_X1 U21228 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18112), .B1(
        n18170), .B2(n18128), .ZN(n18096) );
  OAI211_X1 U21229 ( .C1(n18131), .C2(n18115), .A(n18097), .B(n18096), .ZN(
        P3_U2981) );
  AOI22_X1 U21230 ( .A1(n18111), .A2(n18133), .B1(n18132), .B2(n18110), .ZN(
        n18099) );
  AOI22_X1 U21231 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18112), .B1(
        n18134), .B2(n18106), .ZN(n18098) );
  OAI211_X1 U21232 ( .C1(n18164), .C2(n18137), .A(n18099), .B(n18098), .ZN(
        P3_U2982) );
  AOI22_X1 U21233 ( .A1(n18111), .A2(n18139), .B1(n18138), .B2(n18110), .ZN(
        n18101) );
  AOI22_X1 U21234 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18112), .B1(
        n18140), .B2(n18106), .ZN(n18100) );
  OAI211_X1 U21235 ( .C1(n18164), .C2(n18143), .A(n18101), .B(n18100), .ZN(
        P3_U2983) );
  AOI22_X1 U21236 ( .A1(n18111), .A2(n18145), .B1(n18144), .B2(n18110), .ZN(
        n18103) );
  AOI22_X1 U21237 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18112), .B1(
        n18146), .B2(n18106), .ZN(n18102) );
  OAI211_X1 U21238 ( .C1(n18164), .C2(n18150), .A(n18103), .B(n18102), .ZN(
        P3_U2984) );
  AOI22_X1 U21239 ( .A1(n18170), .A2(n18153), .B1(n18151), .B2(n18110), .ZN(
        n18105) );
  AOI22_X1 U21240 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18112), .B1(
        n18111), .B2(n18152), .ZN(n18104) );
  OAI211_X1 U21241 ( .C1(n18156), .C2(n18115), .A(n18105), .B(n18104), .ZN(
        P3_U2985) );
  AOI22_X1 U21242 ( .A1(n18170), .A2(n18157), .B1(n18158), .B2(n18110), .ZN(
        n18108) );
  AOI22_X1 U21243 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18112), .B1(
        n18160), .B2(n18106), .ZN(n18107) );
  OAI211_X1 U21244 ( .C1(n18109), .C2(n18163), .A(n18108), .B(n18107), .ZN(
        P3_U2986) );
  AOI22_X1 U21245 ( .A1(n18170), .A2(n18168), .B1(n18166), .B2(n18110), .ZN(
        n18114) );
  AOI22_X1 U21246 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18112), .B1(
        n18111), .B2(n18169), .ZN(n18113) );
  OAI211_X1 U21247 ( .C1(n18175), .C2(n18115), .A(n18114), .B(n18113), .ZN(
        P3_U2987) );
  AND2_X1 U21248 ( .A1(n18246), .A2(n18119), .ZN(n18165) );
  AOI22_X1 U21249 ( .A1(n18117), .A2(n18167), .B1(n18116), .B2(n18165), .ZN(
        n18124) );
  AOI22_X1 U21250 ( .A1(n18121), .A2(n18120), .B1(n18119), .B2(n18118), .ZN(
        n18171) );
  AOI22_X1 U21251 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18171), .B1(
        n18122), .B2(n18159), .ZN(n18123) );
  OAI211_X1 U21252 ( .C1(n18125), .C2(n18164), .A(n18124), .B(n18123), .ZN(
        P3_U2988) );
  AOI22_X1 U21253 ( .A1(n18170), .A2(n18127), .B1(n18126), .B2(n18165), .ZN(
        n18130) );
  AOI22_X1 U21254 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18171), .B1(
        n18128), .B2(n18167), .ZN(n18129) );
  OAI211_X1 U21255 ( .C1(n18131), .C2(n18174), .A(n18130), .B(n18129), .ZN(
        P3_U2989) );
  AOI22_X1 U21256 ( .A1(n18170), .A2(n18133), .B1(n18132), .B2(n18165), .ZN(
        n18136) );
  AOI22_X1 U21257 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18171), .B1(
        n18134), .B2(n18159), .ZN(n18135) );
  OAI211_X1 U21258 ( .C1(n18137), .C2(n18149), .A(n18136), .B(n18135), .ZN(
        P3_U2990) );
  AOI22_X1 U21259 ( .A1(n18170), .A2(n18139), .B1(n18138), .B2(n18165), .ZN(
        n18142) );
  AOI22_X1 U21260 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18171), .B1(
        n18140), .B2(n18159), .ZN(n18141) );
  OAI211_X1 U21261 ( .C1(n18143), .C2(n18149), .A(n18142), .B(n18141), .ZN(
        P3_U2991) );
  AOI22_X1 U21262 ( .A1(n18170), .A2(n18145), .B1(n18144), .B2(n18165), .ZN(
        n18148) );
  AOI22_X1 U21263 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18171), .B1(
        n18146), .B2(n18159), .ZN(n18147) );
  OAI211_X1 U21264 ( .C1(n18150), .C2(n18149), .A(n18148), .B(n18147), .ZN(
        P3_U2992) );
  AOI22_X1 U21265 ( .A1(n18170), .A2(n18152), .B1(n18151), .B2(n18165), .ZN(
        n18155) );
  AOI22_X1 U21266 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18171), .B1(
        n18153), .B2(n18167), .ZN(n18154) );
  OAI211_X1 U21267 ( .C1(n18156), .C2(n18174), .A(n18155), .B(n18154), .ZN(
        P3_U2993) );
  AOI22_X1 U21268 ( .A1(n18158), .A2(n18165), .B1(n18157), .B2(n18167), .ZN(
        n18162) );
  AOI22_X1 U21269 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18171), .B1(
        n18160), .B2(n18159), .ZN(n18161) );
  OAI211_X1 U21270 ( .C1(n18164), .C2(n18163), .A(n18162), .B(n18161), .ZN(
        P3_U2994) );
  AOI22_X1 U21271 ( .A1(n18168), .A2(n18167), .B1(n18166), .B2(n18165), .ZN(
        n18173) );
  AOI22_X1 U21272 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18171), .B1(
        n18170), .B2(n18169), .ZN(n18172) );
  OAI211_X1 U21273 ( .C1(n18175), .C2(n18174), .A(n18173), .B(n18172), .ZN(
        P3_U2995) );
  OAI21_X1 U21274 ( .B1(n18188), .B2(n18369), .A(n18176), .ZN(n18178) );
  NAND2_X1 U21275 ( .A1(n18362), .A2(n18355), .ZN(n18177) );
  OAI221_X1 U21276 ( .B1(n18362), .B2(n18355), .C1(n18216), .C2(n18178), .A(
        n18177), .ZN(n18184) );
  AOI21_X1 U21277 ( .B1(n18181), .B2(n18180), .A(n18179), .ZN(n18200) );
  INV_X1 U21278 ( .A(n18200), .ZN(n18182) );
  NAND3_X1 U21279 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18205), .A3(
        n18182), .ZN(n18183) );
  OAI211_X1 U21280 ( .C1(n18351), .C2(n18185), .A(n18184), .B(n18183), .ZN(
        n18353) );
  INV_X1 U21281 ( .A(n18186), .ZN(n18229) );
  AOI22_X1 U21282 ( .A1(n18186), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n18353), .B2(n18229), .ZN(n18214) );
  NAND2_X1 U21283 ( .A1(n18188), .A2(n18187), .ZN(n18189) );
  NAND2_X1 U21284 ( .A1(n18202), .A2(n18369), .ZN(n18197) );
  AOI22_X1 U21285 ( .A1(n18359), .A2(n18189), .B1(n18362), .B2(n18197), .ZN(
        n18356) );
  AOI22_X1 U21286 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18190), .B1(
        n18189), .B2(n18369), .ZN(n18363) );
  AOI222_X1 U21287 ( .A1(n18356), .A2(n18363), .B1(n18356), .B2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C1(n18363), .C2(n18191), .ZN(
        n18193) );
  AOI21_X1 U21288 ( .B1(n18193), .B2(n18229), .A(n18192), .ZN(n18194) );
  AOI21_X1 U21289 ( .B1(n18214), .B2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n18194), .ZN(n18210) );
  OAI21_X1 U21290 ( .B1(n18210), .B2(n18196), .A(n18195), .ZN(n18213) );
  NAND2_X1 U21291 ( .A1(n18355), .A2(n18205), .ZN(n18198) );
  AOI22_X1 U21292 ( .A1(n18218), .A2(n18198), .B1(n18201), .B2(n18197), .ZN(
        n18199) );
  NOR2_X1 U21293 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18199), .ZN(
        n18341) );
  OAI21_X1 U21294 ( .B1(n18202), .B2(n18201), .A(n18200), .ZN(n18203) );
  AOI22_X1 U21295 ( .A1(n18355), .A2(n18205), .B1(n18204), .B2(n18203), .ZN(
        n18342) );
  AOI21_X1 U21296 ( .B1(n18342), .B2(n18229), .A(n18345), .ZN(n18206) );
  AOI21_X1 U21297 ( .B1(n18229), .B2(n18341), .A(n18206), .ZN(n18212) );
  INV_X1 U21298 ( .A(n18214), .ZN(n18208) );
  NOR2_X1 U21299 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18207) );
  OAI221_X1 U21300 ( .B1(n18210), .B2(n18209), .C1(n18210), .C2(n18208), .A(
        n18207), .ZN(n18211) );
  AOI22_X1 U21301 ( .A1(n18214), .A2(n18213), .B1(n18212), .B2(n18211), .ZN(
        n18232) );
  NOR2_X1 U21302 ( .A1(n18216), .A2(n18215), .ZN(n18221) );
  NOR2_X1 U21303 ( .A1(n18218), .A2(n18217), .ZN(n18220) );
  OAI222_X1 U21304 ( .A1(n18224), .A2(n18223), .B1(n18222), .B2(n18221), .C1(
        n18220), .C2(n18219), .ZN(n18383) );
  OAI21_X1 U21305 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18225), .ZN(n18226) );
  OAI211_X1 U21306 ( .C1(n18229), .C2(n18228), .A(n18227), .B(n18226), .ZN(
        n18230) );
  NOR4_X1 U21307 ( .A1(n18232), .A2(n18383), .A3(n18231), .A4(n18230), .ZN(
        n18244) );
  AOI22_X1 U21308 ( .A1(n18364), .A2(n18397), .B1(n18392), .B2(n18386), .ZN(
        n18233) );
  INV_X1 U21309 ( .A(n18233), .ZN(n18240) );
  INV_X1 U21310 ( .A(n18234), .ZN(n18236) );
  OAI211_X1 U21311 ( .C1(n18237), .C2(n18236), .A(n18235), .B(n18244), .ZN(
        n18338) );
  OAI21_X1 U21312 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18385), .A(n18338), 
        .ZN(n18245) );
  NOR2_X1 U21313 ( .A1(n18238), .A2(n18245), .ZN(n18239) );
  MUX2_X1 U21314 ( .A(n18240), .B(n18239), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18242) );
  OAI211_X1 U21315 ( .C1(n18244), .C2(n18243), .A(n18242), .B(n18241), .ZN(
        P3_U2996) );
  NAND2_X1 U21316 ( .A1(n18392), .A2(n18386), .ZN(n18250) );
  NAND4_X1 U21317 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(n18392), .A4(n18403), .ZN(n18252) );
  INV_X1 U21318 ( .A(n18245), .ZN(n18247) );
  NAND3_X1 U21319 ( .A1(n18248), .A2(n18247), .A3(n18246), .ZN(n18249) );
  NAND4_X1 U21320 ( .A1(n18251), .A2(n18250), .A3(n18252), .A4(n18249), .ZN(
        P3_U2997) );
  OAI211_X1 U21321 ( .C1(P3_STATE2_REG_0__SCAN_IN), .C2(
        P3_STATEBS16_REG_SCAN_IN), .A(n18253), .B(n18252), .ZN(n18254) );
  NAND2_X1 U21322 ( .A1(n18255), .A2(n18254), .ZN(P3_U2998) );
  AND2_X1 U21323 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18256), .ZN(
        P3_U2999) );
  AND2_X1 U21324 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18256), .ZN(
        P3_U3000) );
  AND2_X1 U21325 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18256), .ZN(
        P3_U3001) );
  AND2_X1 U21326 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18256), .ZN(
        P3_U3002) );
  AND2_X1 U21327 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18256), .ZN(
        P3_U3003) );
  AND2_X1 U21328 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18256), .ZN(
        P3_U3004) );
  AND2_X1 U21329 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18256), .ZN(
        P3_U3005) );
  AND2_X1 U21330 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18256), .ZN(
        P3_U3006) );
  AND2_X1 U21331 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18256), .ZN(
        P3_U3007) );
  AND2_X1 U21332 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18256), .ZN(
        P3_U3008) );
  AND2_X1 U21333 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18256), .ZN(
        P3_U3009) );
  AND2_X1 U21334 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18256), .ZN(
        P3_U3010) );
  INV_X1 U21335 ( .A(P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20636) );
  NOR2_X1 U21336 ( .A1(n20636), .A2(n18336), .ZN(P3_U3011) );
  AND2_X1 U21337 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18256), .ZN(
        P3_U3012) );
  AND2_X1 U21338 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18256), .ZN(
        P3_U3013) );
  AND2_X1 U21339 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18256), .ZN(
        P3_U3014) );
  AND2_X1 U21340 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18256), .ZN(
        P3_U3015) );
  AND2_X1 U21341 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18256), .ZN(
        P3_U3016) );
  AND2_X1 U21342 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18256), .ZN(
        P3_U3017) );
  AND2_X1 U21343 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18256), .ZN(
        P3_U3018) );
  AND2_X1 U21344 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18256), .ZN(
        P3_U3019) );
  AND2_X1 U21345 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18256), .ZN(
        P3_U3020) );
  AND2_X1 U21346 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18256), .ZN(P3_U3021) );
  AND2_X1 U21347 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18256), .ZN(P3_U3022) );
  AND2_X1 U21348 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18256), .ZN(P3_U3023) );
  AND2_X1 U21349 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18256), .ZN(P3_U3024) );
  AND2_X1 U21350 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18256), .ZN(P3_U3025) );
  AND2_X1 U21351 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18256), .ZN(P3_U3026) );
  AND2_X1 U21352 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18256), .ZN(P3_U3027) );
  AND2_X1 U21353 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18256), .ZN(P3_U3028) );
  NOR2_X1 U21354 ( .A1(n20611), .A2(n19451), .ZN(n18260) );
  NAND2_X1 U21355 ( .A1(HOLD), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18261) );
  INV_X1 U21356 ( .A(n18261), .ZN(n18266) );
  INV_X1 U21357 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18399) );
  NOR3_X1 U21358 ( .A1(n18260), .A2(n18266), .A3(n18399), .ZN(n18259) );
  NAND2_X1 U21359 ( .A1(n18392), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18264) );
  AND2_X1 U21360 ( .A1(n18264), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n18269) );
  INV_X1 U21361 ( .A(NA), .ZN(n20458) );
  OAI21_X1 U21362 ( .B1(n20458), .B2(n18257), .A(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18268) );
  INV_X1 U21363 ( .A(n18268), .ZN(n18258) );
  OAI22_X1 U21364 ( .A1(n18380), .A2(n18259), .B1(n18269), .B2(n18258), .ZN(
        P3_U3029) );
  AOI22_X1 U21365 ( .A1(P3_REQUESTPENDING_REG_SCAN_IN), .A2(n18261), .B1(
        n18260), .B2(n18270), .ZN(n18263) );
  OAI211_X1 U21366 ( .C1(n18263), .C2(n20637), .A(n18264), .B(n18262), .ZN(
        P3_U3030) );
  OAI22_X1 U21367 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18264), .ZN(n18265) );
  OAI22_X1 U21368 ( .A1(n18266), .A2(n18265), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18267) );
  OAI22_X1 U21369 ( .A1(n18269), .A2(n18268), .B1(n20637), .B2(n18267), .ZN(
        P3_U3031) );
  OAI222_X1 U21370 ( .A1(n18371), .A2(n18328), .B1(n18271), .B2(n18380), .C1(
        n18272), .C2(n18318), .ZN(P3_U3032) );
  INV_X1 U21371 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18274) );
  OAI222_X1 U21372 ( .A1(n18318), .A2(n18274), .B1(n18273), .B2(n18380), .C1(
        n18272), .C2(n18328), .ZN(P3_U3033) );
  OAI222_X1 U21373 ( .A1(n18318), .A2(n18276), .B1(n18275), .B2(n18380), .C1(
        n18274), .C2(n18328), .ZN(P3_U3034) );
  OAI222_X1 U21374 ( .A1(n18318), .A2(n18278), .B1(n18277), .B2(n18380), .C1(
        n18276), .C2(n18328), .ZN(P3_U3035) );
  OAI222_X1 U21375 ( .A1(n18318), .A2(n18280), .B1(n18279), .B2(n18380), .C1(
        n18278), .C2(n18328), .ZN(P3_U3036) );
  OAI222_X1 U21376 ( .A1(n18318), .A2(n18282), .B1(n18281), .B2(n18380), .C1(
        n18280), .C2(n18328), .ZN(P3_U3037) );
  OAI222_X1 U21377 ( .A1(n18318), .A2(n18285), .B1(n18283), .B2(n18380), .C1(
        n18282), .C2(n18328), .ZN(P3_U3038) );
  OAI222_X1 U21378 ( .A1(n18285), .A2(n18328), .B1(n18284), .B2(n18380), .C1(
        n18286), .C2(n18318), .ZN(P3_U3039) );
  OAI222_X1 U21379 ( .A1(n18318), .A2(n18288), .B1(n18287), .B2(n18380), .C1(
        n18286), .C2(n18328), .ZN(P3_U3040) );
  INV_X1 U21380 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18290) );
  OAI222_X1 U21381 ( .A1(n18318), .A2(n18290), .B1(n18289), .B2(n18380), .C1(
        n18288), .C2(n18328), .ZN(P3_U3041) );
  OAI222_X1 U21382 ( .A1(n18318), .A2(n18292), .B1(n18291), .B2(n18380), .C1(
        n18290), .C2(n18328), .ZN(P3_U3042) );
  OAI222_X1 U21383 ( .A1(n18318), .A2(n20706), .B1(n18293), .B2(n18380), .C1(
        n18292), .C2(n18328), .ZN(P3_U3043) );
  OAI222_X1 U21384 ( .A1(n20705), .A2(n18328), .B1(n18294), .B2(n18380), .C1(
        n18295), .C2(n18318), .ZN(P3_U3045) );
  OAI222_X1 U21385 ( .A1(n18318), .A2(n18297), .B1(n18296), .B2(n18380), .C1(
        n18295), .C2(n18328), .ZN(P3_U3046) );
  INV_X1 U21386 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18299) );
  OAI222_X1 U21387 ( .A1(n18318), .A2(n18299), .B1(n18298), .B2(n18380), .C1(
        n18297), .C2(n18328), .ZN(P3_U3047) );
  OAI222_X1 U21388 ( .A1(n18299), .A2(n18328), .B1(n20624), .B2(n18380), .C1(
        n18300), .C2(n18318), .ZN(P3_U3048) );
  OAI222_X1 U21389 ( .A1(n18318), .A2(n18302), .B1(n18301), .B2(n18380), .C1(
        n18300), .C2(n18328), .ZN(P3_U3049) );
  OAI222_X1 U21390 ( .A1(n18318), .A2(n18305), .B1(n18303), .B2(n18380), .C1(
        n18302), .C2(n18328), .ZN(P3_U3050) );
  OAI222_X1 U21391 ( .A1(n18305), .A2(n18328), .B1(n18304), .B2(n18380), .C1(
        n18306), .C2(n18318), .ZN(P3_U3051) );
  OAI222_X1 U21392 ( .A1(n18318), .A2(n18308), .B1(n18307), .B2(n18380), .C1(
        n18306), .C2(n18328), .ZN(P3_U3052) );
  OAI222_X1 U21393 ( .A1(n18318), .A2(n18311), .B1(n18309), .B2(n18380), .C1(
        n18308), .C2(n18328), .ZN(P3_U3053) );
  OAI222_X1 U21394 ( .A1(n18311), .A2(n18328), .B1(n18310), .B2(n18380), .C1(
        n18313), .C2(n18318), .ZN(P3_U3054) );
  OAI222_X1 U21395 ( .A1(n18313), .A2(n18328), .B1(n18312), .B2(n18380), .C1(
        n18314), .C2(n18318), .ZN(P3_U3055) );
  OAI222_X1 U21396 ( .A1(n18318), .A2(n18316), .B1(n18315), .B2(n18380), .C1(
        n18314), .C2(n18328), .ZN(P3_U3056) );
  OAI222_X1 U21397 ( .A1(n18318), .A2(n18319), .B1(n18317), .B2(n18380), .C1(
        n18316), .C2(n18328), .ZN(P3_U3057) );
  OAI222_X1 U21398 ( .A1(n18318), .A2(n18322), .B1(n18320), .B2(n18380), .C1(
        n18319), .C2(n18328), .ZN(P3_U3058) );
  OAI222_X1 U21399 ( .A1(n18322), .A2(n18328), .B1(n18321), .B2(n18380), .C1(
        n18323), .C2(n18318), .ZN(P3_U3059) );
  INV_X1 U21400 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18327) );
  OAI222_X1 U21401 ( .A1(n18318), .A2(n18327), .B1(n18324), .B2(n18380), .C1(
        n18323), .C2(n18328), .ZN(P3_U3060) );
  OAI222_X1 U21402 ( .A1(n18328), .A2(n18327), .B1(n18326), .B2(n18380), .C1(
        n18325), .C2(n18318), .ZN(P3_U3061) );
  OAI22_X1 U21403 ( .A1(n18401), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n18380), .ZN(n18329) );
  INV_X1 U21404 ( .A(n18329), .ZN(P3_U3274) );
  OAI22_X1 U21405 ( .A1(n18401), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n18380), .ZN(n18330) );
  INV_X1 U21406 ( .A(n18330), .ZN(P3_U3275) );
  OAI22_X1 U21407 ( .A1(n18401), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18380), .ZN(n18331) );
  INV_X1 U21408 ( .A(n18331), .ZN(P3_U3276) );
  OAI22_X1 U21409 ( .A1(n18401), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n18380), .ZN(n18332) );
  INV_X1 U21410 ( .A(n18332), .ZN(P3_U3277) );
  OAI21_X1 U21411 ( .B1(n18336), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n18334), 
        .ZN(n18333) );
  INV_X1 U21412 ( .A(n18333), .ZN(P3_U3280) );
  OAI21_X1 U21413 ( .B1(n18336), .B2(n18335), .A(n18334), .ZN(P3_U3281) );
  OAI221_X1 U21414 ( .B1(n18339), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18339), 
        .C2(n18338), .A(n18337), .ZN(P3_U3282) );
  AOI22_X1 U21415 ( .A1(n18404), .A2(n18341), .B1(n18364), .B2(n18340), .ZN(
        n18347) );
  OAI21_X1 U21416 ( .B1(n18343), .B2(n18342), .A(n18367), .ZN(n18344) );
  INV_X1 U21417 ( .A(n18344), .ZN(n18346) );
  OAI22_X1 U21418 ( .A1(n18370), .A2(n18347), .B1(n18346), .B2(n18345), .ZN(
        P3_U3285) );
  NOR2_X1 U21419 ( .A1(n18348), .A2(n18366), .ZN(n18357) );
  OAI22_X1 U21420 ( .A1(n18350), .A2(n18349), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18358) );
  INV_X1 U21421 ( .A(n18358), .ZN(n18352) );
  AOI222_X1 U21422 ( .A1(n18353), .A2(n18404), .B1(n18357), .B2(n18352), .C1(
        n18364), .C2(n18351), .ZN(n18354) );
  AOI22_X1 U21423 ( .A1(n18370), .A2(n18355), .B1(n18354), .B2(n18367), .ZN(
        P3_U3288) );
  INV_X1 U21424 ( .A(n18356), .ZN(n18360) );
  AOI222_X1 U21425 ( .A1(n18360), .A2(n18404), .B1(n18364), .B2(n18359), .C1(
        n18358), .C2(n18357), .ZN(n18361) );
  AOI22_X1 U21426 ( .A1(n18370), .A2(n18362), .B1(n18361), .B2(n18367), .ZN(
        P3_U3289) );
  INV_X1 U21427 ( .A(n18363), .ZN(n18365) );
  AOI222_X1 U21428 ( .A1(n18366), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18404), 
        .B2(n18365), .C1(n18369), .C2(n18364), .ZN(n18368) );
  AOI22_X1 U21429 ( .A1(n18370), .A2(n18369), .B1(n18368), .B2(n18367), .ZN(
        P3_U3290) );
  AOI21_X1 U21430 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18372) );
  AOI22_X1 U21431 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18372), .B2(n18371), .ZN(n18374) );
  INV_X1 U21432 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18373) );
  AOI22_X1 U21433 ( .A1(n18375), .A2(n18374), .B1(n18373), .B2(n18378), .ZN(
        P3_U3292) );
  INV_X1 U21434 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18379) );
  NOR2_X1 U21435 ( .A1(n18378), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18376) );
  AOI22_X1 U21436 ( .A1(n18379), .A2(n18378), .B1(n18377), .B2(n18376), .ZN(
        P3_U3293) );
  INV_X1 U21437 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18405) );
  OAI22_X1 U21438 ( .A1(n18401), .A2(n18405), .B1(P3_W_R_N_REG_SCAN_IN), .B2(
        n18380), .ZN(n18381) );
  INV_X1 U21439 ( .A(n18381), .ZN(P3_U3294) );
  MUX2_X1 U21440 ( .A(P3_MORE_REG_SCAN_IN), .B(n18383), .S(n18382), .Z(
        P3_U3295) );
  NOR2_X1 U21441 ( .A1(n18403), .A2(n18394), .ZN(n18389) );
  INV_X1 U21442 ( .A(n18384), .ZN(n18406) );
  AOI21_X1 U21443 ( .B1(n18386), .B2(n18385), .A(n18406), .ZN(n18387) );
  OAI21_X1 U21444 ( .B1(n18389), .B2(n18388), .A(n18387), .ZN(n18400) );
  OAI21_X1 U21445 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n18391), .A(n18390), 
        .ZN(n18393) );
  AOI211_X1 U21446 ( .C1(n18407), .C2(n18393), .A(n18392), .B(n18403), .ZN(
        n18395) );
  NOR2_X1 U21447 ( .A1(n18395), .A2(n18394), .ZN(n18396) );
  OAI21_X1 U21448 ( .B1(n18397), .B2(n18396), .A(n18400), .ZN(n18398) );
  OAI21_X1 U21449 ( .B1(n18400), .B2(n18399), .A(n18398), .ZN(P3_U3296) );
  OAI22_X1 U21450 ( .A1(n18401), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18380), .ZN(n18402) );
  INV_X1 U21451 ( .A(n18402), .ZN(P3_U3297) );
  AOI21_X1 U21452 ( .B1(n18404), .B2(n18403), .A(n18406), .ZN(n18410) );
  AOI22_X1 U21453 ( .A1(n18407), .A2(n18406), .B1(n18410), .B2(n18405), .ZN(
        P3_U3298) );
  INV_X1 U21454 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18409) );
  AOI21_X1 U21455 ( .B1(n18410), .B2(n18409), .A(n18408), .ZN(P3_U3299) );
  INV_X1 U21456 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19442) );
  NAND2_X1 U21457 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20627), .ZN(n19450) );
  NAND2_X1 U21458 ( .A1(n19442), .A2(n18411), .ZN(n19447) );
  OAI21_X1 U21459 ( .B1(n19442), .B2(n19450), .A(n19447), .ZN(n19518) );
  AOI21_X1 U21460 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n19518), .ZN(n18412) );
  INV_X1 U21461 ( .A(n18412), .ZN(P2_U2815) );
  INV_X1 U21462 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18413) );
  OAI22_X1 U21463 ( .A1(n18414), .A2(n18413), .B1(n19440), .B2(n19533), .ZN(
        P2_U2816) );
  NAND2_X1 U21464 ( .A1(n19442), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19597) );
  INV_X2 U21465 ( .A(n19597), .ZN(n19509) );
  AOI21_X1 U21466 ( .B1(n19442), .B2(n20627), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n18415) );
  AOI22_X1 U21467 ( .A1(n19509), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n18415), 
        .B2(n19597), .ZN(P2_U2817) );
  OAI21_X1 U21468 ( .B1(n19454), .B2(BS16), .A(n19518), .ZN(n19516) );
  OAI21_X1 U21469 ( .B1(n19518), .B2(n19263), .A(n19516), .ZN(P2_U2818) );
  NOR2_X1 U21470 ( .A1(n18417), .A2(n18416), .ZN(n19581) );
  OAI21_X1 U21471 ( .B1(n19581), .B2(n12450), .A(n18418), .ZN(P2_U2819) );
  NOR4_X1 U21472 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18422) );
  NOR4_X1 U21473 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18421) );
  NOR4_X1 U21474 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18420) );
  NOR4_X1 U21475 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n18419) );
  NAND4_X1 U21476 ( .A1(n18422), .A2(n18421), .A3(n18420), .A4(n18419), .ZN(
        n18428) );
  NOR4_X1 U21477 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18426) );
  AOI211_X1 U21478 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_30__SCAN_IN), .B(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18425) );
  NOR4_X1 U21479 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18424) );
  NOR4_X1 U21480 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18423) );
  NAND4_X1 U21481 ( .A1(n18426), .A2(n18425), .A3(n18424), .A4(n18423), .ZN(
        n18427) );
  NOR2_X1 U21482 ( .A1(n18428), .A2(n18427), .ZN(n18439) );
  INV_X1 U21483 ( .A(n18439), .ZN(n18437) );
  NOR2_X1 U21484 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18437), .ZN(n18431) );
  INV_X1 U21485 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18429) );
  AOI22_X1 U21486 ( .A1(n18431), .A2(n18432), .B1(n18437), .B2(n18429), .ZN(
        P2_U2820) );
  OR3_X1 U21487 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18436) );
  INV_X1 U21488 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18430) );
  AOI22_X1 U21489 ( .A1(n18431), .A2(n18436), .B1(n18437), .B2(n18430), .ZN(
        P2_U2821) );
  INV_X1 U21490 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19517) );
  NAND2_X1 U21491 ( .A1(n18431), .A2(n19517), .ZN(n18435) );
  OAI21_X1 U21492 ( .B1(n18432), .B2(n19462), .A(n18439), .ZN(n18433) );
  OAI21_X1 U21493 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18439), .A(n18433), 
        .ZN(n18434) );
  OAI221_X1 U21494 ( .B1(n18435), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18435), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18434), .ZN(P2_U2822) );
  INV_X1 U21495 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18438) );
  OAI221_X1 U21496 ( .B1(n18439), .B2(n18438), .C1(n18437), .C2(n18436), .A(
        n18435), .ZN(P2_U2823) );
  AOI22_X1 U21497 ( .A1(n18440), .A2(n18625), .B1(n9725), .B2(n18647), .ZN(
        n18449) );
  AOI211_X1 U21498 ( .C1(n18443), .C2(n18442), .A(n19437), .B(n18441), .ZN(
        n18447) );
  AOI22_X1 U21499 ( .A1(P2_EBX_REG_20__SCAN_IN), .A2(n18614), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n9772), .ZN(n18444) );
  OAI21_X1 U21500 ( .B1(n18445), .B2(n18616), .A(n18444), .ZN(n18446) );
  AOI211_X1 U21501 ( .C1(n18639), .C2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n18447), .B(n18446), .ZN(n18448) );
  NAND2_X1 U21502 ( .A1(n18449), .A2(n18448), .ZN(P2_U2835) );
  AOI211_X1 U21503 ( .C1(n18452), .C2(n18451), .A(n19437), .B(n18450), .ZN(
        n18458) );
  OAI22_X1 U21504 ( .A1(n18642), .A2(n11918), .B1(n18453), .B2(n18616), .ZN(
        n18454) );
  AOI211_X1 U21505 ( .C1(P2_REIP_REG_19__SCAN_IN), .C2(n9772), .A(n18850), .B(
        n18454), .ZN(n18455) );
  OAI21_X1 U21506 ( .B1(n18456), .B2(n18540), .A(n18455), .ZN(n18457) );
  AOI211_X1 U21507 ( .C1(n18625), .C2(n18459), .A(n18458), .B(n18457), .ZN(
        n18460) );
  OAI21_X1 U21508 ( .B1(n18461), .B2(n18628), .A(n18460), .ZN(P2_U2836) );
  AOI211_X1 U21509 ( .C1(n18464), .C2(n18463), .A(n19437), .B(n18462), .ZN(
        n18469) );
  AOI21_X1 U21510 ( .B1(P2_REIP_REG_18__SCAN_IN), .B2(n9772), .A(n18850), .ZN(
        n18466) );
  AOI22_X1 U21511 ( .A1(P2_EBX_REG_18__SCAN_IN), .A2(n18614), .B1(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18639), .ZN(n18465) );
  OAI211_X1 U21512 ( .C1(n18467), .C2(n18616), .A(n18466), .B(n18465), .ZN(
        n18468) );
  AOI211_X1 U21513 ( .C1(n18647), .C2(n18470), .A(n18469), .B(n18468), .ZN(
        n18471) );
  OAI21_X1 U21514 ( .B1(n18472), .B2(n18643), .A(n18471), .ZN(P2_U2837) );
  AOI211_X1 U21515 ( .C1(n18475), .C2(n18474), .A(n18473), .B(n19437), .ZN(
        n18481) );
  OAI22_X1 U21516 ( .A1(n18642), .A2(n11911), .B1(n18476), .B2(n18616), .ZN(
        n18477) );
  AOI211_X1 U21517 ( .C1(P2_REIP_REG_17__SCAN_IN), .C2(n9772), .A(n18850), .B(
        n18477), .ZN(n18478) );
  OAI21_X1 U21518 ( .B1(n18479), .B2(n18540), .A(n18478), .ZN(n18480) );
  AOI211_X1 U21519 ( .C1(n18625), .C2(n18482), .A(n18481), .B(n18480), .ZN(
        n18483) );
  OAI21_X1 U21520 ( .B1(n18484), .B2(n18628), .A(n18483), .ZN(P2_U2838) );
  XNOR2_X1 U21521 ( .A(n18486), .B(n18485), .ZN(n18494) );
  AOI22_X1 U21522 ( .A1(P2_EBX_REG_16__SCAN_IN), .A2(n18614), .B1(n18487), 
        .B2(n18637), .ZN(n18488) );
  OAI211_X1 U21523 ( .C1(n12178), .C2(n18601), .A(n18488), .B(n18496), .ZN(
        n18489) );
  AOI21_X1 U21524 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n18639), .A(
        n18489), .ZN(n18493) );
  AOI22_X1 U21525 ( .A1(n18491), .A2(n18647), .B1(n18490), .B2(n18625), .ZN(
        n18492) );
  OAI211_X1 U21526 ( .C1(n19437), .C2(n18494), .A(n18493), .B(n18492), .ZN(
        P2_U2839) );
  AOI22_X1 U21527 ( .A1(P2_EBX_REG_15__SCAN_IN), .A2(n18614), .B1(n18495), 
        .B2(n18637), .ZN(n18497) );
  OAI211_X1 U21528 ( .C1(n19480), .C2(n18601), .A(n18497), .B(n18496), .ZN(
        n18498) );
  AOI21_X1 U21529 ( .B1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18639), .A(
        n18498), .ZN(n18505) );
  NAND2_X1 U21530 ( .A1(n15696), .A2(n18499), .ZN(n18500) );
  XNOR2_X1 U21531 ( .A(n18501), .B(n18500), .ZN(n18502) );
  AOI22_X1 U21532 ( .A1(n18625), .A2(n18503), .B1(n18623), .B2(n18502), .ZN(
        n18504) );
  OAI211_X1 U21533 ( .C1(n18628), .C2(n18506), .A(n18505), .B(n18504), .ZN(
        P2_U2840) );
  AOI22_X1 U21534 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n18639), .B1(
        n18507), .B2(n18637), .ZN(n18508) );
  OAI21_X1 U21535 ( .B1(n18642), .B2(n11860), .A(n18508), .ZN(n18509) );
  AOI211_X1 U21536 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n9772), .A(n18850), .B(
        n18509), .ZN(n18515) );
  NOR2_X1 U21537 ( .A1(n18630), .A2(n18510), .ZN(n18512) );
  XNOR2_X1 U21538 ( .A(n18512), .B(n18511), .ZN(n18513) );
  AOI22_X1 U21539 ( .A1(n18647), .A2(n18655), .B1(n18623), .B2(n18513), .ZN(
        n18514) );
  OAI211_X1 U21540 ( .C1(n18643), .C2(n18516), .A(n18515), .B(n18514), .ZN(
        P2_U2841) );
  OAI21_X1 U21541 ( .B1(n19477), .B2(n18601), .A(n18600), .ZN(n18520) );
  OAI22_X1 U21542 ( .A1(n18518), .A2(n18540), .B1(n18517), .B2(n18616), .ZN(
        n18519) );
  AOI211_X1 U21543 ( .C1(P2_EBX_REG_13__SCAN_IN), .C2(n18614), .A(n18520), .B(
        n18519), .ZN(n18527) );
  NAND2_X1 U21544 ( .A1(n15696), .A2(n18521), .ZN(n18522) );
  XNOR2_X1 U21545 ( .A(n18523), .B(n18522), .ZN(n18524) );
  AOI22_X1 U21546 ( .A1(n18625), .A2(n18525), .B1(n18623), .B2(n18524), .ZN(
        n18526) );
  OAI211_X1 U21547 ( .C1(n18628), .C2(n18528), .A(n18527), .B(n18526), .ZN(
        P2_U2842) );
  NOR2_X1 U21548 ( .A1(n18630), .A2(n18534), .ZN(n18529) );
  NOR3_X1 U21549 ( .A1(n18529), .A2(n18535), .A3(n19437), .ZN(n18533) );
  AOI22_X1 U21550 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18639), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n9772), .ZN(n18530) );
  OAI211_X1 U21551 ( .C1(n18531), .C2(n18616), .A(n18530), .B(n18600), .ZN(
        n18532) );
  AOI211_X1 U21552 ( .C1(P2_EBX_REG_12__SCAN_IN), .C2(n18614), .A(n18533), .B(
        n18532), .ZN(n18537) );
  NOR3_X1 U21553 ( .A1(n18630), .A2(n18534), .A3(n19437), .ZN(n18546) );
  AOI22_X1 U21554 ( .A1(n18647), .A2(n18659), .B1(n18546), .B2(n18535), .ZN(
        n18536) );
  OAI211_X1 U21555 ( .C1(n18643), .C2(n18538), .A(n18537), .B(n18536), .ZN(
        P2_U2843) );
  INV_X1 U21556 ( .A(n18539), .ZN(n18543) );
  OAI22_X1 U21557 ( .A1(n18541), .A2(n18540), .B1(n12161), .B2(n18601), .ZN(
        n18542) );
  AOI211_X1 U21558 ( .C1(n18647), .C2(n18543), .A(n18850), .B(n18542), .ZN(
        n18554) );
  AOI22_X1 U21559 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n18614), .B1(n10282), 
        .B2(n18637), .ZN(n18553) );
  AOI22_X1 U21560 ( .A1(n18625), .A2(n18545), .B1(n18548), .B2(n18544), .ZN(
        n18552) );
  INV_X1 U21561 ( .A(n18546), .ZN(n18547) );
  AOI21_X1 U21562 ( .B1(n18549), .B2(n18548), .A(n18547), .ZN(n18550) );
  INV_X1 U21563 ( .A(n18550), .ZN(n18551) );
  NAND4_X1 U21564 ( .A1(n18554), .A2(n18553), .A3(n18552), .A4(n18551), .ZN(
        P2_U2844) );
  OAI21_X1 U21565 ( .B1(n12159), .B2(n18601), .A(n18600), .ZN(n18557) );
  OAI22_X1 U21566 ( .A1(n18642), .A2(n10071), .B1(n18555), .B2(n18616), .ZN(
        n18556) );
  AOI211_X1 U21567 ( .C1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n18639), .A(
        n18557), .B(n18556), .ZN(n18564) );
  NOR2_X1 U21568 ( .A1(n18630), .A2(n18558), .ZN(n18560) );
  XNOR2_X1 U21569 ( .A(n18560), .B(n18559), .ZN(n18561) );
  AOI22_X1 U21570 ( .A1(n18625), .A2(n18562), .B1(n18623), .B2(n18561), .ZN(
        n18563) );
  OAI211_X1 U21571 ( .C1(n18628), .C2(n18565), .A(n18564), .B(n18563), .ZN(
        P2_U2845) );
  AOI22_X1 U21572 ( .A1(P2_EBX_REG_9__SCAN_IN), .A2(n18614), .B1(n18637), .B2(
        n18566), .ZN(n18567) );
  OAI211_X1 U21573 ( .C1(n12156), .C2(n18601), .A(n18567), .B(n18600), .ZN(
        n18568) );
  AOI21_X1 U21574 ( .B1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18639), .A(
        n18568), .ZN(n18575) );
  NAND2_X1 U21575 ( .A1(n15696), .A2(n18569), .ZN(n18570) );
  XNOR2_X1 U21576 ( .A(n18571), .B(n18570), .ZN(n18572) );
  AOI22_X1 U21577 ( .A1(n18625), .A2(n18573), .B1(n18623), .B2(n18572), .ZN(
        n18574) );
  OAI211_X1 U21578 ( .C1(n18628), .C2(n18576), .A(n18575), .B(n18574), .ZN(
        P2_U2846) );
  OAI21_X1 U21579 ( .B1(n12016), .B2(n18601), .A(n18600), .ZN(n18580) );
  OAI22_X1 U21580 ( .A1(n18642), .A2(n18578), .B1(n18577), .B2(n18616), .ZN(
        n18579) );
  AOI211_X1 U21581 ( .C1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n18639), .A(
        n18580), .B(n18579), .ZN(n18587) );
  NOR2_X1 U21582 ( .A1(n18630), .A2(n18581), .ZN(n18583) );
  XNOR2_X1 U21583 ( .A(n18583), .B(n18582), .ZN(n18584) );
  AOI22_X1 U21584 ( .A1(n18647), .A2(n18585), .B1(n18623), .B2(n18584), .ZN(
        n18586) );
  OAI211_X1 U21585 ( .C1(n18643), .C2(n18588), .A(n18587), .B(n18586), .ZN(
        P2_U2847) );
  AOI22_X1 U21586 ( .A1(P2_EBX_REG_7__SCAN_IN), .A2(n18614), .B1(n18589), .B2(
        n18637), .ZN(n18590) );
  OAI211_X1 U21587 ( .C1(n19470), .C2(n18601), .A(n18590), .B(n18600), .ZN(
        n18591) );
  AOI21_X1 U21588 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18639), .A(
        n18591), .ZN(n18598) );
  NAND2_X1 U21589 ( .A1(n15696), .A2(n18592), .ZN(n18593) );
  XNOR2_X1 U21590 ( .A(n18594), .B(n18593), .ZN(n18595) );
  AOI22_X1 U21591 ( .A1(n18625), .A2(n18596), .B1(n18623), .B2(n18595), .ZN(
        n18597) );
  OAI211_X1 U21592 ( .C1(n18628), .C2(n18599), .A(n18598), .B(n18597), .ZN(
        P2_U2848) );
  OAI21_X1 U21593 ( .B1(n19468), .B2(n18601), .A(n18600), .ZN(n18605) );
  AOI22_X1 U21594 ( .A1(n18614), .A2(P2_EBX_REG_6__SCAN_IN), .B1(n18602), .B2(
        n18637), .ZN(n18603) );
  INV_X1 U21595 ( .A(n18603), .ZN(n18604) );
  AOI211_X1 U21596 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n18639), .A(
        n18605), .B(n18604), .ZN(n18612) );
  NOR2_X1 U21597 ( .A1(n18630), .A2(n18606), .ZN(n18608) );
  XNOR2_X1 U21598 ( .A(n18608), .B(n18607), .ZN(n18609) );
  AOI22_X1 U21599 ( .A1(n18625), .A2(n18610), .B1(n18623), .B2(n18609), .ZN(
        n18611) );
  OAI211_X1 U21600 ( .C1(n18628), .C2(n18613), .A(n18612), .B(n18611), .ZN(
        P2_U2849) );
  AOI22_X1 U21601 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n18639), .B1(
        P2_EBX_REG_5__SCAN_IN), .B2(n18614), .ZN(n18615) );
  OAI21_X1 U21602 ( .B1(n18617), .B2(n18616), .A(n18615), .ZN(n18618) );
  AOI211_X1 U21603 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n9772), .A(n18850), .B(
        n18618), .ZN(n18627) );
  NAND2_X1 U21604 ( .A1(n15696), .A2(n18619), .ZN(n18620) );
  XNOR2_X1 U21605 ( .A(n18621), .B(n18620), .ZN(n18622) );
  AOI22_X1 U21606 ( .A1(n18625), .A2(n18624), .B1(n18623), .B2(n18622), .ZN(
        n18626) );
  OAI211_X1 U21607 ( .C1(n18628), .C2(n18674), .A(n18627), .B(n18626), .ZN(
        P2_U2850) );
  NOR2_X1 U21608 ( .A1(n18630), .A2(n18629), .ZN(n18631) );
  XOR2_X1 U21609 ( .A(n18815), .B(n18631), .Z(n18649) );
  NAND2_X1 U21610 ( .A1(n18633), .A2(n18632), .ZN(n18635) );
  AND2_X1 U21611 ( .A1(n18635), .A2(n10179), .ZN(n18843) );
  AOI21_X1 U21612 ( .B1(P2_REIP_REG_4__SCAN_IN), .B2(n9772), .A(n18850), .ZN(
        n18641) );
  AOI22_X1 U21613 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18639), .B1(
        n18638), .B2(n18637), .ZN(n18640) );
  OAI211_X1 U21614 ( .C1(n18642), .C2(n12671), .A(n18641), .B(n18640), .ZN(
        n18646) );
  OAI22_X1 U21615 ( .A1(n18677), .A2(n18644), .B1(n18838), .B2(n18643), .ZN(
        n18645) );
  AOI211_X1 U21616 ( .C1(n18647), .C2(n18843), .A(n18646), .B(n18645), .ZN(
        n18648) );
  OAI21_X1 U21617 ( .B1(n19437), .B2(n18649), .A(n18648), .ZN(P2_U2851) );
  AOI22_X1 U21618 ( .A1(n18651), .A2(BUF2_REG_31__SCAN_IN), .B1(n18692), .B2(
        n18650), .ZN(n18654) );
  AOI22_X1 U21619 ( .A1(n18652), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n18691), .ZN(n18653) );
  NAND2_X1 U21620 ( .A1(n18654), .A2(n18653), .ZN(P2_U2888) );
  INV_X1 U21621 ( .A(n18655), .ZN(n18658) );
  AOI22_X1 U21622 ( .A1(n18667), .A2(n18656), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n18691), .ZN(n18657) );
  OAI21_X1 U21623 ( .B1(n18675), .B2(n18658), .A(n18657), .ZN(P2_U2905) );
  INV_X1 U21624 ( .A(n18659), .ZN(n18662) );
  AOI22_X1 U21625 ( .A1(n18667), .A2(n18660), .B1(P2_EAX_REG_12__SCAN_IN), 
        .B2(n18691), .ZN(n18661) );
  OAI21_X1 U21626 ( .B1(n18675), .B2(n18662), .A(n18661), .ZN(P2_U2907) );
  AOI22_X1 U21627 ( .A1(n18667), .A2(n18663), .B1(P2_EAX_REG_8__SCAN_IN), .B2(
        n18691), .ZN(n18664) );
  OAI21_X1 U21628 ( .B1(n18675), .B2(n18665), .A(n18664), .ZN(P2_U2911) );
  AOI22_X1 U21629 ( .A1(n18667), .A2(n18666), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n18691), .ZN(n18673) );
  NAND2_X1 U21630 ( .A1(n19534), .A2(n19540), .ZN(n18670) );
  XOR2_X1 U21631 ( .A(n19540), .B(n19534), .Z(n18683) );
  NAND2_X1 U21632 ( .A1(n19546), .A2(n18863), .ZN(n18669) );
  NAND2_X1 U21633 ( .A1(n18669), .A2(n18668), .ZN(n18682) );
  NAND2_X1 U21634 ( .A1(n18683), .A2(n18682), .ZN(n18681) );
  AOI21_X1 U21635 ( .B1(n18670), .B2(n18681), .A(n18843), .ZN(n18676) );
  OR3_X1 U21636 ( .A1(n18676), .A2(n18677), .A3(n18671), .ZN(n18672) );
  OAI211_X1 U21637 ( .C1(n18675), .C2(n18674), .A(n18673), .B(n18672), .ZN(
        P2_U2914) );
  AOI22_X1 U21638 ( .A1(n18692), .A2(n18843), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n18691), .ZN(n18680) );
  XOR2_X1 U21639 ( .A(n18677), .B(n18676), .Z(n18678) );
  NAND2_X1 U21640 ( .A1(n18678), .A2(n18694), .ZN(n18679) );
  OAI211_X1 U21641 ( .C1(n18908), .C2(n18698), .A(n18680), .B(n18679), .ZN(
        P2_U2915) );
  OAI21_X1 U21642 ( .B1(n18683), .B2(n18682), .A(n18681), .ZN(n18684) );
  NAND2_X1 U21643 ( .A1(n18684), .A2(n18694), .ZN(n18690) );
  INV_X1 U21644 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n18685) );
  OAI22_X1 U21645 ( .A1(n19534), .A2(n18687), .B1(n18686), .B2(n18685), .ZN(
        n18688) );
  INV_X1 U21646 ( .A(n18688), .ZN(n18689) );
  OAI211_X1 U21647 ( .C1(n18904), .C2(n18698), .A(n18690), .B(n18689), .ZN(
        P2_U2916) );
  AOI22_X1 U21648 ( .A1(n18692), .A2(n18695), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n18691), .ZN(n18697) );
  OAI211_X1 U21649 ( .C1(n19128), .C2(n18695), .A(n18694), .B(n18693), .ZN(
        n18696) );
  OAI211_X1 U21650 ( .C1(n18785), .C2(n18698), .A(n18697), .B(n18696), .ZN(
        P2_U2919) );
  NAND3_X1 U21651 ( .A1(n18701), .A2(n18700), .A3(n18699), .ZN(n18703) );
  NAND2_X1 U21652 ( .A1(n18703), .A2(n18702), .ZN(n18704) );
  NOR2_X1 U21653 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19563), .ZN(n18767) );
  CLKBUF_X2 U21654 ( .A(n18767), .Z(n19594) );
  NOR2_X4 U21655 ( .A1(n18737), .A2(n19594), .ZN(n18755) );
  AND2_X1 U21656 ( .A1(n18755), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  AOI22_X1 U21657 ( .A1(n19594), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n18755), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n18706) );
  OAI21_X1 U21658 ( .B1(n18707), .B2(n18735), .A(n18706), .ZN(P2_U2921) );
  AOI22_X1 U21659 ( .A1(n19594), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n18755), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n18708) );
  OAI21_X1 U21660 ( .B1(n18709), .B2(n18735), .A(n18708), .ZN(P2_U2922) );
  AOI22_X1 U21661 ( .A1(n19594), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n18755), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n18710) );
  OAI21_X1 U21662 ( .B1(n18711), .B2(n18735), .A(n18710), .ZN(P2_U2923) );
  AOI22_X1 U21663 ( .A1(n19594), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n18755), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n18712) );
  OAI21_X1 U21664 ( .B1(n18713), .B2(n18735), .A(n18712), .ZN(P2_U2924) );
  AOI22_X1 U21665 ( .A1(n19594), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n18755), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n18714) );
  OAI21_X1 U21666 ( .B1(n18715), .B2(n18735), .A(n18714), .ZN(P2_U2925) );
  INV_X1 U21667 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n18717) );
  AOI22_X1 U21668 ( .A1(n19594), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n18755), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n18716) );
  OAI21_X1 U21669 ( .B1(n18717), .B2(n18735), .A(n18716), .ZN(P2_U2926) );
  AOI22_X1 U21670 ( .A1(n19594), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n18755), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n18718) );
  OAI21_X1 U21671 ( .B1(n18719), .B2(n18735), .A(n18718), .ZN(P2_U2927) );
  INV_X1 U21672 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n18721) );
  AOI22_X1 U21673 ( .A1(n19594), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n18755), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n18720) );
  OAI21_X1 U21674 ( .B1(n18721), .B2(n18735), .A(n18720), .ZN(P2_U2928) );
  INV_X1 U21675 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n18723) );
  AOI22_X1 U21676 ( .A1(n19594), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n18755), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n18722) );
  OAI21_X1 U21677 ( .B1(n18723), .B2(n18735), .A(n18722), .ZN(P2_U2929) );
  AOI22_X1 U21678 ( .A1(n19594), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n18755), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n18724) );
  OAI21_X1 U21679 ( .B1(n18725), .B2(n18735), .A(n18724), .ZN(P2_U2930) );
  INV_X1 U21680 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n18727) );
  AOI22_X1 U21681 ( .A1(n19594), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n18755), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n18726) );
  OAI21_X1 U21682 ( .B1(n18727), .B2(n18735), .A(n18726), .ZN(P2_U2931) );
  INV_X1 U21683 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n18729) );
  AOI22_X1 U21684 ( .A1(n19594), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n18755), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n18728) );
  OAI21_X1 U21685 ( .B1(n18729), .B2(n18735), .A(n18728), .ZN(P2_U2932) );
  INV_X1 U21686 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n18731) );
  AOI22_X1 U21687 ( .A1(n19594), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n18755), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n18730) );
  OAI21_X1 U21688 ( .B1(n18731), .B2(n18735), .A(n18730), .ZN(P2_U2933) );
  INV_X1 U21689 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n18733) );
  AOI22_X1 U21690 ( .A1(n19594), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n18755), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n18732) );
  OAI21_X1 U21691 ( .B1(n18733), .B2(n18735), .A(n18732), .ZN(P2_U2934) );
  INV_X1 U21692 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n18736) );
  AOI22_X1 U21693 ( .A1(n19594), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n18755), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n18734) );
  OAI21_X1 U21694 ( .B1(n18736), .B2(n18735), .A(n18734), .ZN(P2_U2935) );
  AOI22_X1 U21695 ( .A1(n19594), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n18755), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n18738) );
  OAI21_X1 U21696 ( .B1(n18739), .B2(n18769), .A(n18738), .ZN(P2_U2936) );
  AOI22_X1 U21697 ( .A1(n19594), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n18755), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n18740) );
  OAI21_X1 U21698 ( .B1(n18741), .B2(n18769), .A(n18740), .ZN(P2_U2937) );
  AOI22_X1 U21699 ( .A1(n19594), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n18755), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n18742) );
  OAI21_X1 U21700 ( .B1(n18743), .B2(n18769), .A(n18742), .ZN(P2_U2938) );
  AOI22_X1 U21701 ( .A1(n19594), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n18755), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n18744) );
  OAI21_X1 U21702 ( .B1(n18745), .B2(n18769), .A(n18744), .ZN(P2_U2939) );
  AOI22_X1 U21703 ( .A1(n19594), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n18755), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n18746) );
  OAI21_X1 U21704 ( .B1(n18747), .B2(n18769), .A(n18746), .ZN(P2_U2940) );
  AOI22_X1 U21705 ( .A1(n19594), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n18755), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n18748) );
  OAI21_X1 U21706 ( .B1(n20620), .B2(n18769), .A(n18748), .ZN(P2_U2941) );
  AOI22_X1 U21707 ( .A1(n18767), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n18755), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n18749) );
  OAI21_X1 U21708 ( .B1(n18750), .B2(n18769), .A(n18749), .ZN(P2_U2942) );
  AOI22_X1 U21709 ( .A1(n18767), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n18755), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n18751) );
  OAI21_X1 U21710 ( .B1(n18752), .B2(n18769), .A(n18751), .ZN(P2_U2943) );
  AOI22_X1 U21711 ( .A1(n18767), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n18755), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n18753) );
  OAI21_X1 U21712 ( .B1(n18754), .B2(n18769), .A(n18753), .ZN(P2_U2944) );
  AOI22_X1 U21713 ( .A1(n18767), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n18755), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n18756) );
  OAI21_X1 U21714 ( .B1(n18757), .B2(n18769), .A(n18756), .ZN(P2_U2945) );
  INV_X1 U21715 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n18759) );
  AOI22_X1 U21716 ( .A1(n18767), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n18755), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n18758) );
  OAI21_X1 U21717 ( .B1(n18759), .B2(n18769), .A(n18758), .ZN(P2_U2946) );
  INV_X1 U21718 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n18761) );
  AOI22_X1 U21719 ( .A1(n18767), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n18755), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n18760) );
  OAI21_X1 U21720 ( .B1(n18761), .B2(n18769), .A(n18760), .ZN(P2_U2947) );
  AOI22_X1 U21721 ( .A1(n18767), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n18755), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n18762) );
  OAI21_X1 U21722 ( .B1(n18685), .B2(n18769), .A(n18762), .ZN(P2_U2948) );
  INV_X1 U21723 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n18764) );
  AOI22_X1 U21724 ( .A1(n18767), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n18755), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n18763) );
  OAI21_X1 U21725 ( .B1(n18764), .B2(n18769), .A(n18763), .ZN(P2_U2949) );
  INV_X1 U21726 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n18766) );
  AOI22_X1 U21727 ( .A1(n18767), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n18755), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n18765) );
  OAI21_X1 U21728 ( .B1(n18766), .B2(n18769), .A(n18765), .ZN(P2_U2950) );
  INV_X1 U21729 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n18770) );
  AOI22_X1 U21730 ( .A1(n18767), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n18755), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n18768) );
  OAI21_X1 U21731 ( .B1(n18770), .B2(n18769), .A(n18768), .ZN(P2_U2951) );
  AOI22_X1 U21732 ( .A1(n18773), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_16__SCAN_IN), .B2(n18801), .ZN(n18771) );
  OAI21_X1 U21733 ( .B1(n18785), .B2(n18804), .A(n18771), .ZN(P2_U2952) );
  AOI22_X1 U21734 ( .A1(n18773), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n18801), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n18772) );
  OAI21_X1 U21735 ( .B1(n18896), .B2(n18804), .A(n18772), .ZN(P2_U2953) );
  AOI22_X1 U21736 ( .A1(n18773), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n18801), .ZN(n18774) );
  OAI21_X1 U21737 ( .B1(n18901), .B2(n18804), .A(n18774), .ZN(P2_U2954) );
  AOI22_X1 U21738 ( .A1(n18802), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n18801), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n18775) );
  OAI21_X1 U21739 ( .B1(n18904), .B2(n18804), .A(n18775), .ZN(P2_U2955) );
  AOI22_X1 U21740 ( .A1(n18802), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n18801), .ZN(n18776) );
  OAI21_X1 U21741 ( .B1(n18908), .B2(n18804), .A(n18776), .ZN(P2_U2956) );
  AOI22_X1 U21742 ( .A1(n18802), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n18801), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n18777) );
  OAI21_X1 U21743 ( .B1(n18912), .B2(n18804), .A(n18777), .ZN(P2_U2957) );
  AOI22_X1 U21744 ( .A1(n18802), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n18801), .ZN(n18778) );
  OAI21_X1 U21745 ( .B1(n18920), .B2(n18804), .A(n18778), .ZN(P2_U2958) );
  AOI22_X1 U21746 ( .A1(n18802), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n18801), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n18779) );
  OAI21_X1 U21747 ( .B1(n18928), .B2(n18804), .A(n18779), .ZN(P2_U2959) );
  AOI22_X1 U21748 ( .A1(n18802), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n18801), 
        .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n18780) );
  OAI21_X1 U21749 ( .B1(n18794), .B2(n18804), .A(n18780), .ZN(P2_U2961) );
  AOI22_X1 U21750 ( .A1(n18802), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(
        P2_EAX_REG_26__SCAN_IN), .B2(n18801), .ZN(n18781) );
  OAI21_X1 U21751 ( .B1(n18796), .B2(n18804), .A(n18781), .ZN(P2_U2962) );
  AOI22_X1 U21752 ( .A1(n18802), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n18801), .ZN(n18782) );
  OAI21_X1 U21753 ( .B1(n18798), .B2(n18804), .A(n18782), .ZN(P2_U2963) );
  AOI22_X1 U21754 ( .A1(n18802), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n18801), .ZN(n18783) );
  OAI21_X1 U21755 ( .B1(n18800), .B2(n18804), .A(n18783), .ZN(P2_U2965) );
  AOI22_X1 U21756 ( .A1(n18802), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_0__SCAN_IN), .B2(n18801), .ZN(n18784) );
  OAI21_X1 U21757 ( .B1(n18785), .B2(n18804), .A(n18784), .ZN(P2_U2967) );
  AOI22_X1 U21758 ( .A1(n18802), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n18801), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n18786) );
  OAI21_X1 U21759 ( .B1(n18896), .B2(n18804), .A(n18786), .ZN(P2_U2968) );
  AOI22_X1 U21760 ( .A1(n18802), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n18801), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n18787) );
  OAI21_X1 U21761 ( .B1(n18901), .B2(n18804), .A(n18787), .ZN(P2_U2969) );
  AOI22_X1 U21762 ( .A1(n18802), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n18801), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n18788) );
  OAI21_X1 U21763 ( .B1(n18904), .B2(n18804), .A(n18788), .ZN(P2_U2970) );
  AOI22_X1 U21764 ( .A1(n18802), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n18801), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n18789) );
  OAI21_X1 U21765 ( .B1(n18908), .B2(n18804), .A(n18789), .ZN(P2_U2971) );
  AOI22_X1 U21766 ( .A1(n18802), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n18801), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n18790) );
  OAI21_X1 U21767 ( .B1(n18912), .B2(n18804), .A(n18790), .ZN(P2_U2972) );
  AOI22_X1 U21768 ( .A1(n18802), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n18801), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n18791) );
  OAI21_X1 U21769 ( .B1(n18920), .B2(n18804), .A(n18791), .ZN(P2_U2973) );
  AOI22_X1 U21770 ( .A1(n18802), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n18801), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n18792) );
  OAI21_X1 U21771 ( .B1(n18928), .B2(n18804), .A(n18792), .ZN(P2_U2974) );
  AOI22_X1 U21772 ( .A1(n18802), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_9__SCAN_IN), .B2(n18801), .ZN(n18793) );
  OAI21_X1 U21773 ( .B1(n18794), .B2(n18804), .A(n18793), .ZN(P2_U2976) );
  AOI22_X1 U21774 ( .A1(n18802), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(
        P2_EAX_REG_10__SCAN_IN), .B2(n18801), .ZN(n18795) );
  OAI21_X1 U21775 ( .B1(n18796), .B2(n18804), .A(n18795), .ZN(P2_U2977) );
  AOI22_X1 U21776 ( .A1(n18802), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n18801), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n18797) );
  OAI21_X1 U21777 ( .B1(n18798), .B2(n18804), .A(n18797), .ZN(P2_U2978) );
  AOI22_X1 U21778 ( .A1(n18802), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_13__SCAN_IN), .B2(n18801), .ZN(n18799) );
  OAI21_X1 U21779 ( .B1(n18800), .B2(n18804), .A(n18799), .ZN(P2_U2980) );
  AOI22_X1 U21780 ( .A1(n18802), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n18801), 
        .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n18803) );
  OAI21_X1 U21781 ( .B1(n18805), .B2(n18804), .A(n18803), .ZN(P2_U2982) );
  AOI22_X1 U21782 ( .A1(n18820), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n18850), .ZN(n18814) );
  XNOR2_X1 U21783 ( .A(n18806), .B(n18844), .ZN(n18848) );
  NAND2_X1 U21784 ( .A1(n18848), .A2(n18821), .ZN(n18810) );
  XNOR2_X1 U21785 ( .A(n18807), .B(n9749), .ZN(n18847) );
  NAND2_X1 U21786 ( .A1(n18847), .A2(n18808), .ZN(n18809) );
  OAI211_X1 U21787 ( .C1(n18811), .C2(n18838), .A(n18810), .B(n18809), .ZN(
        n18812) );
  INV_X1 U21788 ( .A(n18812), .ZN(n18813) );
  OAI211_X1 U21789 ( .C1(n18816), .C2(n18815), .A(n18814), .B(n18813), .ZN(
        P2_U3010) );
  AOI21_X1 U21790 ( .B1(n18819), .B2(n18818), .A(n18817), .ZN(n18857) );
  AOI22_X1 U21791 ( .A1(n18857), .A2(n18821), .B1(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18820), .ZN(n18836) );
  NAND2_X1 U21792 ( .A1(n18823), .A2(n18822), .ZN(n18824) );
  NAND2_X1 U21793 ( .A1(n18825), .A2(n18824), .ZN(n18858) );
  INV_X1 U21794 ( .A(n18826), .ZN(n18828) );
  NAND2_X1 U21795 ( .A1(n13482), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n18871) );
  INV_X1 U21796 ( .A(n18871), .ZN(n18827) );
  AOI21_X1 U21797 ( .B1(n18829), .B2(n18828), .A(n18827), .ZN(n18832) );
  NAND2_X1 U21798 ( .A1(n13260), .A2(n18830), .ZN(n18831) );
  OAI211_X1 U21799 ( .C1(n18858), .C2(n18833), .A(n18832), .B(n18831), .ZN(
        n18834) );
  INV_X1 U21800 ( .A(n18834), .ZN(n18835) );
  NAND2_X1 U21801 ( .A1(n18836), .A2(n18835), .ZN(P2_U3012) );
  NAND2_X1 U21802 ( .A1(n18837), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18840) );
  OAI22_X1 U21803 ( .A1(n18841), .A2(n18840), .B1(n18839), .B2(n18838), .ZN(
        n18842) );
  INV_X1 U21804 ( .A(n18842), .ZN(n18854) );
  AOI22_X1 U21805 ( .A1(n18845), .A2(n18844), .B1(n18843), .B2(n18875), .ZN(
        n18853) );
  AOI22_X1 U21806 ( .A1(n18849), .A2(n18848), .B1(n18847), .B2(n18846), .ZN(
        n18852) );
  NAND2_X1 U21807 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n18850), .ZN(n18851) );
  NAND4_X1 U21808 ( .A1(n18854), .A2(n18853), .A3(n18852), .A4(n18851), .ZN(
        P2_U3042) );
  AOI21_X1 U21809 ( .B1(n18856), .B2(n18869), .A(n18855), .ZN(n18879) );
  INV_X1 U21810 ( .A(n18857), .ZN(n18860) );
  OAI22_X1 U21811 ( .A1(n18861), .A2(n18860), .B1(n18859), .B2(n18858), .ZN(
        n18862) );
  INV_X1 U21812 ( .A(n18862), .ZN(n18877) );
  INV_X1 U21813 ( .A(n18863), .ZN(n19548) );
  AOI21_X1 U21814 ( .B1(n18866), .B2(n18865), .A(n18864), .ZN(n18867) );
  AOI21_X1 U21815 ( .B1(n18868), .B2(n13233), .A(n18867), .ZN(n18873) );
  OR3_X1 U21816 ( .A1(n18870), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A3(
        n18869), .ZN(n18872) );
  NAND3_X1 U21817 ( .A1(n18873), .A2(n18872), .A3(n18871), .ZN(n18874) );
  AOI21_X1 U21818 ( .B1(n18875), .B2(n19548), .A(n18874), .ZN(n18876) );
  OAI211_X1 U21819 ( .C1(n18879), .C2(n18878), .A(n18877), .B(n18876), .ZN(
        P2_U3044) );
  NAND2_X1 U21820 ( .A1(n12827), .A2(n19550), .ZN(n18987) );
  INV_X1 U21821 ( .A(n18987), .ZN(n18988) );
  NAND2_X1 U21822 ( .A1(n18988), .A2(n19560), .ZN(n18936) );
  NOR2_X1 U21823 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18936), .ZN(
        n18927) );
  AOI22_X1 U21824 ( .A1(n19303), .A2(n19427), .B1(n19370), .B2(n18927), .ZN(
        n18892) );
  INV_X1 U21825 ( .A(n18958), .ZN(n18880) );
  OAI21_X1 U21826 ( .B1(n19427), .B2(n18880), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n18881) );
  NAND2_X1 U21827 ( .A1(n18881), .A2(n19333), .ZN(n18890) );
  NOR2_X1 U21828 ( .A1(n18882), .A2(n12827), .ZN(n19422) );
  NOR2_X1 U21829 ( .A1(n19422), .A2(n18927), .ZN(n18889) );
  INV_X1 U21830 ( .A(n18889), .ZN(n18886) );
  INV_X1 U21831 ( .A(n18927), .ZN(n18883) );
  OAI211_X1 U21832 ( .C1(n18884), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n18883), 
        .B(n19533), .ZN(n18885) );
  OAI211_X1 U21833 ( .C1(n18890), .C2(n18886), .A(n19377), .B(n18885), .ZN(
        n18930) );
  OAI21_X1 U21834 ( .B1(n18887), .B2(n18927), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n18888) );
  AOI22_X1 U21835 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18930), .B1(
        n19371), .B2(n18929), .ZN(n18891) );
  OAI211_X1 U21836 ( .C1(n19306), .C2(n18958), .A(n18892), .B(n18891), .ZN(
        P2_U3048) );
  AOI22_X1 U21837 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n18924), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n18923), .ZN(n19389) );
  INV_X1 U21838 ( .A(n19389), .ZN(n19236) );
  NOR2_X2 U21839 ( .A1(n18895), .A2(n18925), .ZN(n19384) );
  AOI22_X1 U21840 ( .A1(n19236), .A2(n19427), .B1(n19384), .B2(n18927), .ZN(
        n18898) );
  NOR2_X2 U21841 ( .A1(n18896), .A2(n19104), .ZN(n19385) );
  AOI22_X1 U21842 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18930), .B1(
        n19385), .B2(n18929), .ZN(n18897) );
  OAI211_X1 U21843 ( .C1(n19239), .C2(n18958), .A(n18898), .B(n18897), .ZN(
        P2_U3049) );
  INV_X1 U21844 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n20604) );
  INV_X1 U21845 ( .A(n19392), .ZN(n19243) );
  AOI22_X1 U21846 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n18924), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n18923), .ZN(n19395) );
  INV_X1 U21847 ( .A(n19395), .ZN(n19240) );
  NOR2_X2 U21848 ( .A1(n18900), .A2(n18925), .ZN(n19390) );
  AOI22_X1 U21849 ( .A1(n19240), .A2(n19427), .B1(n19390), .B2(n18927), .ZN(
        n18903) );
  NOR2_X2 U21850 ( .A1(n18901), .A2(n19104), .ZN(n19391) );
  AOI22_X1 U21851 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18930), .B1(
        n19391), .B2(n18929), .ZN(n18902) );
  OAI211_X1 U21852 ( .C1(n19243), .C2(n18958), .A(n18903), .B(n18902), .ZN(
        P2_U3050) );
  AOI22_X1 U21853 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n18924), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n18923), .ZN(n19315) );
  NOR2_X2 U21854 ( .A1(n9808), .A2(n18925), .ZN(n19396) );
  AOI22_X1 U21855 ( .A1(n19398), .A2(n19427), .B1(n19396), .B2(n18927), .ZN(
        n18906) );
  NOR2_X2 U21856 ( .A1(n18904), .A2(n19104), .ZN(n19397) );
  AOI22_X1 U21857 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18930), .B1(
        n19397), .B2(n18929), .ZN(n18905) );
  OAI211_X1 U21858 ( .C1(n19401), .C2(n18958), .A(n18906), .B(n18905), .ZN(
        P2_U3051) );
  AOI22_X1 U21859 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n18924), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n18923), .ZN(n19319) );
  AOI22_X1 U21860 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n18924), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n18923), .ZN(n19407) );
  INV_X1 U21861 ( .A(n19407), .ZN(n19316) );
  NOR2_X2 U21862 ( .A1(n18907), .A2(n18925), .ZN(n19402) );
  AOI22_X1 U21863 ( .A1(n19316), .A2(n19427), .B1(n19402), .B2(n18927), .ZN(
        n18910) );
  NOR2_X2 U21864 ( .A1(n18908), .A2(n19104), .ZN(n19403) );
  AOI22_X1 U21865 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18930), .B1(
        n19403), .B2(n18929), .ZN(n18909) );
  OAI211_X1 U21866 ( .C1(n19319), .C2(n18958), .A(n18910), .B(n18909), .ZN(
        P2_U3052) );
  AOI22_X2 U21867 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n18924), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n18923), .ZN(n19415) );
  AOI22_X1 U21868 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18923), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n18924), .ZN(n19283) );
  NOR2_X2 U21869 ( .A1(n18911), .A2(n18925), .ZN(n19408) );
  AOI22_X1 U21870 ( .A1(n19410), .A2(n19427), .B1(n19408), .B2(n18927), .ZN(
        n18914) );
  NOR2_X2 U21871 ( .A1(n18912), .A2(n19104), .ZN(n19409) );
  AOI22_X1 U21872 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18930), .B1(
        n19409), .B2(n18929), .ZN(n18913) );
  OAI211_X1 U21873 ( .C1(n19415), .C2(n18958), .A(n18914), .B(n18913), .ZN(
        P2_U3053) );
  AOI22_X1 U21874 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18923), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n18924), .ZN(n19421) );
  INV_X1 U21875 ( .A(n19421), .ZN(n19357) );
  AOI22_X1 U21876 ( .A1(n19357), .A2(n19427), .B1(n9773), .B2(n18927), .ZN(
        n18922) );
  NOR2_X2 U21877 ( .A1(n18920), .A2(n19104), .ZN(n19417) );
  AOI22_X1 U21878 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18930), .B1(
        n19417), .B2(n18929), .ZN(n18921) );
  OAI211_X1 U21879 ( .C1(n19360), .C2(n18958), .A(n18922), .B(n18921), .ZN(
        P2_U3054) );
  AOI22_X1 U21880 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n18924), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n18923), .ZN(n19330) );
  AOI22_X1 U21881 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n18924), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n18923), .ZN(n19432) );
  AOI22_X1 U21882 ( .A1(n19325), .A2(n19427), .B1(n19423), .B2(n18927), .ZN(
        n18932) );
  NOR2_X2 U21883 ( .A1(n18928), .A2(n19104), .ZN(n19424) );
  AOI22_X1 U21884 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18930), .B1(
        n19424), .B2(n18929), .ZN(n18931) );
  OAI211_X1 U21885 ( .C1(n19330), .C2(n18958), .A(n18932), .B(n18931), .ZN(
        P2_U3055) );
  INV_X1 U21886 ( .A(n18933), .ZN(n18934) );
  NAND2_X1 U21887 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19560), .ZN(
        n19160) );
  NOR2_X1 U21888 ( .A1(n19160), .A2(n18987), .ZN(n18953) );
  NOR3_X1 U21889 ( .A1(n18934), .A2(n18953), .A3(n19586), .ZN(n18935) );
  AOI211_X2 U21890 ( .C1(n18936), .C2(n19586), .A(n19101), .B(n18935), .ZN(
        n18954) );
  AOI22_X1 U21891 ( .A1(n18954), .A2(n19371), .B1(n19370), .B2(n18953), .ZN(
        n18940) );
  NAND2_X1 U21892 ( .A1(n19540), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19049) );
  INV_X1 U21893 ( .A(n19049), .ZN(n19103) );
  NAND2_X1 U21894 ( .A1(n19103), .A2(n19161), .ZN(n18937) );
  AOI21_X1 U21895 ( .B1(n18937), .B2(n18936), .A(n18935), .ZN(n18938) );
  OAI211_X1 U21896 ( .C1(n18953), .C2(n19535), .A(n18938), .B(n19377), .ZN(
        n18955) );
  NOR2_X2 U21897 ( .A1(n19159), .A2(n19108), .ZN(n18983) );
  AOI22_X1 U21898 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18955), .B1(
        n18983), .B2(n19380), .ZN(n18939) );
  OAI211_X1 U21899 ( .C1(n19383), .C2(n18958), .A(n18940), .B(n18939), .ZN(
        P2_U3056) );
  AOI22_X1 U21900 ( .A1(n18954), .A2(n19385), .B1(n19384), .B2(n18953), .ZN(
        n18942) );
  AOI22_X1 U21901 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18955), .B1(
        n18983), .B2(n19386), .ZN(n18941) );
  OAI211_X1 U21902 ( .C1(n19389), .C2(n18958), .A(n18942), .B(n18941), .ZN(
        P2_U3057) );
  AOI22_X1 U21903 ( .A1(n18954), .A2(n19391), .B1(n19390), .B2(n18953), .ZN(
        n18944) );
  AOI22_X1 U21904 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18955), .B1(
        n18983), .B2(n19392), .ZN(n18943) );
  OAI211_X1 U21905 ( .C1(n19395), .C2(n18958), .A(n18944), .B(n18943), .ZN(
        P2_U3058) );
  AOI22_X1 U21906 ( .A1(n18954), .A2(n19397), .B1(n19396), .B2(n18953), .ZN(
        n18946) );
  INV_X1 U21907 ( .A(n19401), .ZN(n19311) );
  AOI22_X1 U21908 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18955), .B1(
        n18983), .B2(n19311), .ZN(n18945) );
  OAI211_X1 U21909 ( .C1(n19315), .C2(n18958), .A(n18946), .B(n18945), .ZN(
        P2_U3059) );
  AOI22_X1 U21910 ( .A1(n18954), .A2(n19403), .B1(n19402), .B2(n18953), .ZN(
        n18948) );
  INV_X1 U21911 ( .A(n19319), .ZN(n19404) );
  AOI22_X1 U21912 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18955), .B1(
        n18983), .B2(n19404), .ZN(n18947) );
  OAI211_X1 U21913 ( .C1(n19407), .C2(n18958), .A(n18948), .B(n18947), .ZN(
        P2_U3060) );
  AOI22_X1 U21914 ( .A1(n18954), .A2(n19409), .B1(n19408), .B2(n18953), .ZN(
        n18950) );
  INV_X1 U21915 ( .A(n19415), .ZN(n19280) );
  AOI22_X1 U21916 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18955), .B1(
        n18983), .B2(n19280), .ZN(n18949) );
  OAI211_X1 U21917 ( .C1(n19283), .C2(n18958), .A(n18950), .B(n18949), .ZN(
        P2_U3061) );
  AOI22_X1 U21918 ( .A1(n18954), .A2(n19417), .B1(n19416), .B2(n18953), .ZN(
        n18952) );
  AOI22_X1 U21919 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18955), .B1(
        n18983), .B2(n19418), .ZN(n18951) );
  OAI211_X1 U21920 ( .C1(n19421), .C2(n18958), .A(n18952), .B(n18951), .ZN(
        P2_U3062) );
  AOI22_X1 U21921 ( .A1(n18954), .A2(n19424), .B1(n19423), .B2(n18953), .ZN(
        n18957) );
  INV_X1 U21922 ( .A(n19330), .ZN(n19426) );
  AOI22_X1 U21923 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18955), .B1(
        n18983), .B2(n19426), .ZN(n18956) );
  OAI211_X1 U21924 ( .C1(n19432), .C2(n18958), .A(n18957), .B(n18956), .ZN(
        P2_U3063) );
  NOR2_X1 U21925 ( .A1(n19560), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19192) );
  NAND2_X1 U21926 ( .A1(n19192), .A2(n18988), .ZN(n18961) );
  AND2_X1 U21927 ( .A1(n18962), .A2(n18961), .ZN(n18960) );
  NAND2_X1 U21928 ( .A1(n19021), .A2(n18988), .ZN(n18964) );
  OAI22_X1 U21929 ( .A1(n18960), .A2(n19586), .B1(n19533), .B2(n18964), .ZN(
        n18982) );
  INV_X1 U21930 ( .A(n18961), .ZN(n18981) );
  AOI22_X1 U21931 ( .A1(n18982), .A2(n19371), .B1(n19370), .B2(n18981), .ZN(
        n18968) );
  AOI21_X1 U21932 ( .B1(n18962), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n18966) );
  OAI21_X1 U21933 ( .B1(n18983), .B2(n19007), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n18963) );
  NAND2_X1 U21934 ( .A1(n18964), .A2(n18963), .ZN(n18965) );
  OAI211_X1 U21935 ( .C1(n18981), .C2(n18966), .A(n18965), .B(n19377), .ZN(
        n18984) );
  AOI22_X1 U21936 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18984), .B1(
        n18983), .B2(n19303), .ZN(n18967) );
  OAI211_X1 U21937 ( .C1(n19306), .C2(n19018), .A(n18968), .B(n18967), .ZN(
        P2_U3064) );
  AOI22_X1 U21938 ( .A1(n18982), .A2(n19385), .B1(n19384), .B2(n18981), .ZN(
        n18970) );
  AOI22_X1 U21939 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18984), .B1(
        n18983), .B2(n19236), .ZN(n18969) );
  OAI211_X1 U21940 ( .C1(n19239), .C2(n19018), .A(n18970), .B(n18969), .ZN(
        P2_U3065) );
  AOI22_X1 U21941 ( .A1(n18982), .A2(n19391), .B1(n19390), .B2(n18981), .ZN(
        n18972) );
  AOI22_X1 U21942 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18984), .B1(
        n18983), .B2(n19240), .ZN(n18971) );
  OAI211_X1 U21943 ( .C1(n19243), .C2(n19018), .A(n18972), .B(n18971), .ZN(
        P2_U3066) );
  AOI22_X1 U21944 ( .A1(n18982), .A2(n19397), .B1(n19396), .B2(n18981), .ZN(
        n18974) );
  AOI22_X1 U21945 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18984), .B1(
        n18983), .B2(n19398), .ZN(n18973) );
  OAI211_X1 U21946 ( .C1(n19401), .C2(n19018), .A(n18974), .B(n18973), .ZN(
        P2_U3067) );
  AOI22_X1 U21947 ( .A1(n18982), .A2(n19403), .B1(n19402), .B2(n18981), .ZN(
        n18976) );
  AOI22_X1 U21948 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18984), .B1(
        n18983), .B2(n19316), .ZN(n18975) );
  OAI211_X1 U21949 ( .C1(n19319), .C2(n19018), .A(n18976), .B(n18975), .ZN(
        P2_U3068) );
  AOI22_X1 U21950 ( .A1(n18982), .A2(n19409), .B1(n19408), .B2(n18981), .ZN(
        n18978) );
  AOI22_X1 U21951 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18984), .B1(
        n18983), .B2(n19410), .ZN(n18977) );
  OAI211_X1 U21952 ( .C1(n19415), .C2(n19018), .A(n18978), .B(n18977), .ZN(
        P2_U3069) );
  AOI22_X1 U21953 ( .A1(n18982), .A2(n19417), .B1(n19416), .B2(n18981), .ZN(
        n18980) );
  AOI22_X1 U21954 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18984), .B1(
        n18983), .B2(n19357), .ZN(n18979) );
  OAI211_X1 U21955 ( .C1(n19360), .C2(n19018), .A(n18980), .B(n18979), .ZN(
        P2_U3070) );
  AOI22_X1 U21956 ( .A1(n18982), .A2(n19424), .B1(n19423), .B2(n18981), .ZN(
        n18986) );
  AOI22_X1 U21957 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18984), .B1(
        n18983), .B2(n19325), .ZN(n18985) );
  OAI211_X1 U21958 ( .C1(n19330), .C2(n19018), .A(n18986), .B(n18985), .ZN(
        P2_U3071) );
  NOR2_X1 U21959 ( .A1(n19227), .A2(n18987), .ZN(n19013) );
  AOI22_X1 U21960 ( .A1(n19303), .A2(n19007), .B1(n19370), .B2(n19013), .ZN(
        n18998) );
  OAI21_X1 U21961 ( .B1(n19049), .B2(n19191), .A(n19333), .ZN(n18996) );
  NAND2_X1 U21962 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18988), .ZN(
        n18995) );
  INV_X1 U21963 ( .A(n18995), .ZN(n18991) );
  INV_X1 U21964 ( .A(n19013), .ZN(n18989) );
  OAI211_X1 U21965 ( .C1(n18992), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n18989), 
        .B(n19533), .ZN(n18990) );
  OAI211_X1 U21966 ( .C1(n18996), .C2(n18991), .A(n19377), .B(n18990), .ZN(
        n19015) );
  INV_X1 U21967 ( .A(n18992), .ZN(n18993) );
  OAI21_X1 U21968 ( .B1(n18993), .B2(n19013), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n18994) );
  OAI21_X1 U21969 ( .B1(n18996), .B2(n18995), .A(n18994), .ZN(n19014) );
  AOI22_X1 U21970 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19015), .B1(
        n19371), .B2(n19014), .ZN(n18997) );
  OAI211_X1 U21971 ( .C1(n19306), .C2(n19010), .A(n18998), .B(n18997), .ZN(
        P2_U3072) );
  AOI22_X1 U21972 ( .A1(n19386), .A2(n19045), .B1(n19013), .B2(n19384), .ZN(
        n19000) );
  AOI22_X1 U21973 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19015), .B1(
        n19385), .B2(n19014), .ZN(n18999) );
  OAI211_X1 U21974 ( .C1(n19389), .C2(n19018), .A(n19000), .B(n18999), .ZN(
        P2_U3073) );
  AOI22_X1 U21975 ( .A1(n19392), .A2(n19045), .B1(n19013), .B2(n19390), .ZN(
        n19002) );
  AOI22_X1 U21976 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19015), .B1(
        n19391), .B2(n19014), .ZN(n19001) );
  OAI211_X1 U21977 ( .C1(n19395), .C2(n19018), .A(n19002), .B(n19001), .ZN(
        P2_U3074) );
  AOI22_X1 U21978 ( .A1(n19398), .A2(n19007), .B1(n19013), .B2(n19396), .ZN(
        n19004) );
  AOI22_X1 U21979 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19015), .B1(
        n19397), .B2(n19014), .ZN(n19003) );
  OAI211_X1 U21980 ( .C1(n19401), .C2(n19010), .A(n19004), .B(n19003), .ZN(
        P2_U3075) );
  AOI22_X1 U21981 ( .A1(n19404), .A2(n19045), .B1(n19013), .B2(n19402), .ZN(
        n19006) );
  AOI22_X1 U21982 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19015), .B1(
        n19403), .B2(n19014), .ZN(n19005) );
  OAI211_X1 U21983 ( .C1(n19407), .C2(n19018), .A(n19006), .B(n19005), .ZN(
        P2_U3076) );
  AOI22_X1 U21984 ( .A1(n19410), .A2(n19007), .B1(n19013), .B2(n19408), .ZN(
        n19009) );
  AOI22_X1 U21985 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19015), .B1(
        n19409), .B2(n19014), .ZN(n19008) );
  OAI211_X1 U21986 ( .C1(n19415), .C2(n19010), .A(n19009), .B(n19008), .ZN(
        P2_U3077) );
  AOI22_X1 U21987 ( .A1(n19418), .A2(n19045), .B1(n19013), .B2(n19416), .ZN(
        n19012) );
  AOI22_X1 U21988 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19015), .B1(
        n19417), .B2(n19014), .ZN(n19011) );
  OAI211_X1 U21989 ( .C1(n19421), .C2(n19018), .A(n19012), .B(n19011), .ZN(
        P2_U3078) );
  AOI22_X1 U21990 ( .A1(n19426), .A2(n19045), .B1(n19013), .B2(n19423), .ZN(
        n19017) );
  AOI22_X1 U21991 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19015), .B1(
        n19424), .B2(n19014), .ZN(n19016) );
  OAI211_X1 U21992 ( .C1(n19432), .C2(n19018), .A(n19017), .B(n19016), .ZN(
        P2_U3079) );
  OR2_X1 U21993 ( .A1(n19021), .A2(n19020), .ZN(n19261) );
  INV_X1 U21994 ( .A(n19261), .ZN(n19268) );
  NAND2_X1 U21995 ( .A1(n19268), .A2(n12827), .ZN(n19026) );
  NOR2_X1 U21996 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19056), .ZN(
        n19043) );
  OAI21_X1 U21997 ( .B1(n19023), .B2(n19043), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19022) );
  OAI21_X1 U21998 ( .B1(n19026), .B2(n19533), .A(n19022), .ZN(n19044) );
  AOI22_X1 U21999 ( .A1(n19044), .A2(n19371), .B1(n19370), .B2(n19043), .ZN(
        n19030) );
  INV_X1 U22000 ( .A(n19023), .ZN(n19024) );
  AOI21_X1 U22001 ( .B1(n19024), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19028) );
  OAI21_X1 U22002 ( .B1(n19045), .B2(n19068), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19025) );
  AOI21_X1 U22003 ( .B1(n19026), .B2(n19025), .A(n19104), .ZN(n19027) );
  AOI22_X1 U22004 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19046), .B1(
        n19045), .B2(n19303), .ZN(n19029) );
  OAI211_X1 U22005 ( .C1(n19306), .C2(n19078), .A(n19030), .B(n19029), .ZN(
        P2_U3080) );
  AOI22_X1 U22006 ( .A1(n19044), .A2(n19385), .B1(n19384), .B2(n19043), .ZN(
        n19032) );
  AOI22_X1 U22007 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19046), .B1(
        n19045), .B2(n19236), .ZN(n19031) );
  OAI211_X1 U22008 ( .C1(n19239), .C2(n19078), .A(n19032), .B(n19031), .ZN(
        P2_U3081) );
  AOI22_X1 U22009 ( .A1(n19044), .A2(n19391), .B1(n19390), .B2(n19043), .ZN(
        n19034) );
  AOI22_X1 U22010 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19046), .B1(
        n19045), .B2(n19240), .ZN(n19033) );
  OAI211_X1 U22011 ( .C1(n19243), .C2(n19078), .A(n19034), .B(n19033), .ZN(
        P2_U3082) );
  AOI22_X1 U22012 ( .A1(n19044), .A2(n19397), .B1(n19396), .B2(n19043), .ZN(
        n19036) );
  AOI22_X1 U22013 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19046), .B1(
        n19045), .B2(n19398), .ZN(n19035) );
  OAI211_X1 U22014 ( .C1(n19401), .C2(n19078), .A(n19036), .B(n19035), .ZN(
        P2_U3083) );
  AOI22_X1 U22015 ( .A1(n19044), .A2(n19403), .B1(n19402), .B2(n19043), .ZN(
        n19038) );
  AOI22_X1 U22016 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19046), .B1(
        n19045), .B2(n19316), .ZN(n19037) );
  OAI211_X1 U22017 ( .C1(n19319), .C2(n19078), .A(n19038), .B(n19037), .ZN(
        P2_U3084) );
  AOI22_X1 U22018 ( .A1(n19044), .A2(n19409), .B1(n19408), .B2(n19043), .ZN(
        n19040) );
  AOI22_X1 U22019 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19046), .B1(
        n19045), .B2(n19410), .ZN(n19039) );
  OAI211_X1 U22020 ( .C1(n19415), .C2(n19078), .A(n19040), .B(n19039), .ZN(
        P2_U3085) );
  AOI22_X1 U22021 ( .A1(n19044), .A2(n19417), .B1(n19416), .B2(n19043), .ZN(
        n19042) );
  AOI22_X1 U22022 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19046), .B1(
        n19045), .B2(n19357), .ZN(n19041) );
  OAI211_X1 U22023 ( .C1(n19360), .C2(n19078), .A(n19042), .B(n19041), .ZN(
        P2_U3086) );
  AOI22_X1 U22024 ( .A1(n19044), .A2(n19424), .B1(n19423), .B2(n19043), .ZN(
        n19048) );
  AOI22_X1 U22025 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19046), .B1(
        n19045), .B2(n19325), .ZN(n19047) );
  OAI211_X1 U22026 ( .C1(n19330), .C2(n19078), .A(n19048), .B(n19047), .ZN(
        P2_U3087) );
  AOI22_X1 U22027 ( .A1(n19380), .A2(n19095), .B1(n19370), .B2(n19073), .ZN(
        n19059) );
  OAI21_X1 U22028 ( .B1(n19049), .B2(n19297), .A(n19333), .ZN(n19057) );
  INV_X1 U22029 ( .A(n19056), .ZN(n19052) );
  INV_X1 U22030 ( .A(n19073), .ZN(n19050) );
  OAI211_X1 U22031 ( .C1(n19053), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19050), 
        .B(n19533), .ZN(n19051) );
  OAI211_X1 U22032 ( .C1(n19057), .C2(n19052), .A(n19377), .B(n19051), .ZN(
        n19075) );
  INV_X1 U22033 ( .A(n19053), .ZN(n19054) );
  OAI21_X1 U22034 ( .B1(n19054), .B2(n19073), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19055) );
  OAI21_X1 U22035 ( .B1(n19057), .B2(n19056), .A(n19055), .ZN(n19074) );
  AOI22_X1 U22036 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19075), .B1(
        n19371), .B2(n19074), .ZN(n19058) );
  OAI211_X1 U22037 ( .C1(n19383), .C2(n19078), .A(n19059), .B(n19058), .ZN(
        P2_U3088) );
  AOI22_X1 U22038 ( .A1(n19386), .A2(n19095), .B1(n19073), .B2(n19384), .ZN(
        n19061) );
  AOI22_X1 U22039 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19075), .B1(
        n19385), .B2(n19074), .ZN(n19060) );
  OAI211_X1 U22040 ( .C1(n19389), .C2(n19078), .A(n19061), .B(n19060), .ZN(
        P2_U3089) );
  AOI22_X1 U22041 ( .A1(n19240), .A2(n19068), .B1(n19390), .B2(n19073), .ZN(
        n19063) );
  AOI22_X1 U22042 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19075), .B1(
        n19391), .B2(n19074), .ZN(n19062) );
  OAI211_X1 U22043 ( .C1(n19243), .C2(n19092), .A(n19063), .B(n19062), .ZN(
        P2_U3090) );
  AOI22_X1 U22044 ( .A1(n19398), .A2(n19068), .B1(n19073), .B2(n19396), .ZN(
        n19065) );
  AOI22_X1 U22045 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19075), .B1(
        n19397), .B2(n19074), .ZN(n19064) );
  OAI211_X1 U22046 ( .C1(n19401), .C2(n19092), .A(n19065), .B(n19064), .ZN(
        P2_U3091) );
  AOI22_X1 U22047 ( .A1(n19404), .A2(n19095), .B1(n19073), .B2(n19402), .ZN(
        n19067) );
  AOI22_X1 U22048 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19075), .B1(
        n19403), .B2(n19074), .ZN(n19066) );
  OAI211_X1 U22049 ( .C1(n19407), .C2(n19078), .A(n19067), .B(n19066), .ZN(
        P2_U3092) );
  AOI22_X1 U22050 ( .A1(n19410), .A2(n19068), .B1(n19073), .B2(n19408), .ZN(
        n19070) );
  AOI22_X1 U22051 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19075), .B1(
        n19409), .B2(n19074), .ZN(n19069) );
  OAI211_X1 U22052 ( .C1(n19415), .C2(n19092), .A(n19070), .B(n19069), .ZN(
        P2_U3093) );
  AOI22_X1 U22053 ( .A1(n19418), .A2(n19095), .B1(n19073), .B2(n19416), .ZN(
        n19072) );
  AOI22_X1 U22054 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19075), .B1(
        n19417), .B2(n19074), .ZN(n19071) );
  OAI211_X1 U22055 ( .C1(n19421), .C2(n19078), .A(n19072), .B(n19071), .ZN(
        P2_U3094) );
  AOI22_X1 U22056 ( .A1(n19426), .A2(n19095), .B1(n19073), .B2(n19423), .ZN(
        n19077) );
  AOI22_X1 U22057 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19075), .B1(
        n19424), .B2(n19074), .ZN(n19076) );
  OAI211_X1 U22058 ( .C1(n19432), .C2(n19078), .A(n19077), .B(n19076), .ZN(
        P2_U3095) );
  AOI22_X1 U22059 ( .A1(n19094), .A2(n19385), .B1(n19093), .B2(n19384), .ZN(
        n19080) );
  AOI22_X1 U22060 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19096), .B1(
        n19089), .B2(n19386), .ZN(n19079) );
  OAI211_X1 U22061 ( .C1(n19389), .C2(n19092), .A(n19080), .B(n19079), .ZN(
        P2_U3097) );
  AOI22_X1 U22062 ( .A1(n19094), .A2(n19391), .B1(n19093), .B2(n19390), .ZN(
        n19082) );
  AOI22_X1 U22063 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19096), .B1(
        n19089), .B2(n19392), .ZN(n19081) );
  OAI211_X1 U22064 ( .C1(n19395), .C2(n19092), .A(n19082), .B(n19081), .ZN(
        P2_U3098) );
  AOI22_X1 U22065 ( .A1(n19094), .A2(n19397), .B1(n19093), .B2(n19396), .ZN(
        n19084) );
  AOI22_X1 U22066 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19096), .B1(
        n19095), .B2(n19398), .ZN(n19083) );
  OAI211_X1 U22067 ( .C1(n19401), .C2(n19127), .A(n19084), .B(n19083), .ZN(
        P2_U3099) );
  AOI22_X1 U22068 ( .A1(n19094), .A2(n19403), .B1(n19093), .B2(n19402), .ZN(
        n19086) );
  AOI22_X1 U22069 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19096), .B1(
        n19089), .B2(n19404), .ZN(n19085) );
  OAI211_X1 U22070 ( .C1(n19407), .C2(n19092), .A(n19086), .B(n19085), .ZN(
        P2_U3100) );
  AOI22_X1 U22071 ( .A1(n19094), .A2(n19409), .B1(n19093), .B2(n19408), .ZN(
        n19088) );
  AOI22_X1 U22072 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19096), .B1(
        n19095), .B2(n19410), .ZN(n19087) );
  OAI211_X1 U22073 ( .C1(n19415), .C2(n19127), .A(n19088), .B(n19087), .ZN(
        P2_U3101) );
  AOI22_X1 U22074 ( .A1(n19094), .A2(n19417), .B1(n19093), .B2(n19416), .ZN(
        n19091) );
  AOI22_X1 U22075 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19096), .B1(
        n19089), .B2(n19418), .ZN(n19090) );
  OAI211_X1 U22076 ( .C1(n19421), .C2(n19092), .A(n19091), .B(n19090), .ZN(
        P2_U3102) );
  AOI22_X1 U22077 ( .A1(n19094), .A2(n19424), .B1(n19093), .B2(n19423), .ZN(
        n19098) );
  AOI22_X1 U22078 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19096), .B1(
        n19095), .B2(n19325), .ZN(n19097) );
  OAI211_X1 U22079 ( .C1(n19330), .C2(n19127), .A(n19098), .B(n19097), .ZN(
        P2_U3103) );
  INV_X1 U22080 ( .A(n19099), .ZN(n19100) );
  NOR3_X1 U22081 ( .A1(n19100), .A2(n19135), .A3(n19586), .ZN(n19105) );
  AOI211_X2 U22082 ( .C1(n19106), .C2(n19586), .A(n19101), .B(n19105), .ZN(
        n19123) );
  AOI22_X1 U22083 ( .A1(n19123), .A2(n19371), .B1(n19135), .B2(n19370), .ZN(
        n19110) );
  INV_X1 U22084 ( .A(n19373), .ZN(n19102) );
  NAND2_X1 U22085 ( .A1(n19103), .A2(n19102), .ZN(n19532) );
  AOI211_X1 U22086 ( .C1(n19532), .C2(n19106), .A(n19105), .B(n19104), .ZN(
        n19107) );
  OAI21_X1 U22087 ( .B1(n19135), .B2(n19535), .A(n19107), .ZN(n19124) );
  AOI22_X1 U22088 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19124), .B1(
        n19154), .B2(n19380), .ZN(n19109) );
  OAI211_X1 U22089 ( .C1(n19383), .C2(n19127), .A(n19110), .B(n19109), .ZN(
        P2_U3104) );
  AOI22_X1 U22090 ( .A1(n19123), .A2(n19385), .B1(n19135), .B2(n19384), .ZN(
        n19112) );
  AOI22_X1 U22091 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19124), .B1(
        n19154), .B2(n19386), .ZN(n19111) );
  OAI211_X1 U22092 ( .C1(n19389), .C2(n19127), .A(n19112), .B(n19111), .ZN(
        P2_U3105) );
  AOI22_X1 U22093 ( .A1(n19123), .A2(n19391), .B1(n19135), .B2(n19390), .ZN(
        n19114) );
  AOI22_X1 U22094 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19124), .B1(
        n19154), .B2(n19392), .ZN(n19113) );
  OAI211_X1 U22095 ( .C1(n19395), .C2(n19127), .A(n19114), .B(n19113), .ZN(
        P2_U3106) );
  AOI22_X1 U22096 ( .A1(n19123), .A2(n19397), .B1(n19135), .B2(n19396), .ZN(
        n19116) );
  AOI22_X1 U22097 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19124), .B1(
        n19154), .B2(n19311), .ZN(n19115) );
  OAI211_X1 U22098 ( .C1(n19315), .C2(n19127), .A(n19116), .B(n19115), .ZN(
        P2_U3107) );
  AOI22_X1 U22099 ( .A1(n19123), .A2(n19403), .B1(n19135), .B2(n19402), .ZN(
        n19118) );
  AOI22_X1 U22100 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19124), .B1(
        n19154), .B2(n19404), .ZN(n19117) );
  OAI211_X1 U22101 ( .C1(n19407), .C2(n19127), .A(n19118), .B(n19117), .ZN(
        P2_U3108) );
  AOI22_X1 U22102 ( .A1(n19123), .A2(n19409), .B1(n19135), .B2(n19408), .ZN(
        n19120) );
  AOI22_X1 U22103 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19124), .B1(
        n19154), .B2(n19280), .ZN(n19119) );
  OAI211_X1 U22104 ( .C1(n19283), .C2(n19127), .A(n19120), .B(n19119), .ZN(
        P2_U3109) );
  AOI22_X1 U22105 ( .A1(n19123), .A2(n19417), .B1(n19135), .B2(n19416), .ZN(
        n19122) );
  AOI22_X1 U22106 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19124), .B1(
        n19154), .B2(n19418), .ZN(n19121) );
  OAI211_X1 U22107 ( .C1(n19421), .C2(n19127), .A(n19122), .B(n19121), .ZN(
        P2_U3110) );
  AOI22_X1 U22108 ( .A1(n19123), .A2(n19424), .B1(n19135), .B2(n19423), .ZN(
        n19126) );
  AOI22_X1 U22109 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19124), .B1(
        n19154), .B2(n19426), .ZN(n19125) );
  OAI211_X1 U22110 ( .C1(n19432), .C2(n19127), .A(n19126), .B(n19125), .ZN(
        P2_U3111) );
  NAND2_X1 U22111 ( .A1(n19550), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19226) );
  OR2_X1 U22112 ( .A1(n19226), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19168) );
  NOR2_X1 U22113 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19168), .ZN(
        n19153) );
  AOI22_X1 U22114 ( .A1(n19303), .A2(n19154), .B1(n19370), .B2(n19153), .ZN(
        n19140) );
  NAND2_X1 U22115 ( .A1(n19182), .A2(n19129), .ZN(n19130) );
  AOI21_X1 U22116 ( .B1(n19130), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19533), 
        .ZN(n19134) );
  OAI21_X1 U22117 ( .B1(n19136), .B2(n19586), .A(n19535), .ZN(n19131) );
  AOI21_X1 U22118 ( .B1(n19134), .B2(n19132), .A(n19131), .ZN(n19133) );
  OAI21_X1 U22119 ( .B1(n19153), .B2(n19133), .A(n19377), .ZN(n19156) );
  OAI21_X1 U22120 ( .B1(n19135), .B2(n19153), .A(n19134), .ZN(n19138) );
  OAI21_X1 U22121 ( .B1(n19136), .B2(n19153), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19137) );
  NAND2_X1 U22122 ( .A1(n19138), .A2(n19137), .ZN(n19155) );
  AOI22_X1 U22123 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19156), .B1(
        n19371), .B2(n19155), .ZN(n19139) );
  OAI211_X1 U22124 ( .C1(n19306), .C2(n19182), .A(n19140), .B(n19139), .ZN(
        P2_U3112) );
  AOI22_X1 U22125 ( .A1(n19236), .A2(n19154), .B1(n19384), .B2(n19153), .ZN(
        n19142) );
  AOI22_X1 U22126 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19156), .B1(
        n19155), .B2(n19385), .ZN(n19141) );
  OAI211_X1 U22127 ( .C1(n19239), .C2(n19182), .A(n19142), .B(n19141), .ZN(
        P2_U3113) );
  AOI22_X1 U22128 ( .A1(n19240), .A2(n19154), .B1(n19390), .B2(n19153), .ZN(
        n19144) );
  AOI22_X1 U22129 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19156), .B1(
        n19155), .B2(n19391), .ZN(n19143) );
  OAI211_X1 U22130 ( .C1(n19243), .C2(n19182), .A(n19144), .B(n19143), .ZN(
        P2_U3114) );
  AOI22_X1 U22131 ( .A1(n19398), .A2(n19154), .B1(n19396), .B2(n19153), .ZN(
        n19146) );
  AOI22_X1 U22132 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19156), .B1(
        n19155), .B2(n19397), .ZN(n19145) );
  OAI211_X1 U22133 ( .C1(n19401), .C2(n19182), .A(n19146), .B(n19145), .ZN(
        P2_U3115) );
  AOI22_X1 U22134 ( .A1(n19316), .A2(n19154), .B1(n19402), .B2(n19153), .ZN(
        n19148) );
  AOI22_X1 U22135 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19156), .B1(
        n19155), .B2(n19403), .ZN(n19147) );
  OAI211_X1 U22136 ( .C1(n19319), .C2(n19182), .A(n19148), .B(n19147), .ZN(
        P2_U3116) );
  AOI22_X1 U22137 ( .A1(n19410), .A2(n19154), .B1(n19408), .B2(n19153), .ZN(
        n19150) );
  AOI22_X1 U22138 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19156), .B1(
        n19155), .B2(n19409), .ZN(n19149) );
  OAI211_X1 U22139 ( .C1(n19415), .C2(n19182), .A(n19150), .B(n19149), .ZN(
        P2_U3117) );
  AOI22_X1 U22140 ( .A1(n19357), .A2(n19154), .B1(n9773), .B2(n19153), .ZN(
        n19152) );
  AOI22_X1 U22141 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19156), .B1(
        n19155), .B2(n19417), .ZN(n19151) );
  OAI211_X1 U22142 ( .C1(n19360), .C2(n19182), .A(n19152), .B(n19151), .ZN(
        P2_U3118) );
  AOI22_X1 U22143 ( .A1(n19325), .A2(n19154), .B1(n19423), .B2(n19153), .ZN(
        n19158) );
  AOI22_X1 U22144 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19156), .B1(
        n19155), .B2(n19424), .ZN(n19157) );
  OAI211_X1 U22145 ( .C1(n19330), .C2(n19182), .A(n19158), .B(n19157), .ZN(
        P2_U3119) );
  INV_X1 U22146 ( .A(n19182), .ZN(n19185) );
  NOR2_X1 U22147 ( .A1(n19160), .A2(n19226), .ZN(n19196) );
  AOI22_X1 U22148 ( .A1(n19303), .A2(n19185), .B1(n19370), .B2(n19196), .ZN(
        n19171) );
  AOI21_X1 U22149 ( .B1(n19165), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19163) );
  NOR2_X1 U22150 ( .A1(n19540), .A2(n19263), .ZN(n19372) );
  AOI21_X1 U22151 ( .B1(n19372), .B2(n19161), .A(n19533), .ZN(n19164) );
  NAND2_X1 U22152 ( .A1(n19164), .A2(n19168), .ZN(n19162) );
  OAI211_X1 U22153 ( .C1(n19196), .C2(n19163), .A(n19162), .B(n19377), .ZN(
        n19187) );
  INV_X1 U22154 ( .A(n19164), .ZN(n19169) );
  INV_X1 U22155 ( .A(n19165), .ZN(n19166) );
  OAI21_X1 U22156 ( .B1(n19166), .B2(n19196), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19167) );
  OAI21_X1 U22157 ( .B1(n19169), .B2(n19168), .A(n19167), .ZN(n19186) );
  AOI22_X1 U22158 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19187), .B1(
        n19371), .B2(n19186), .ZN(n19170) );
  OAI211_X1 U22159 ( .C1(n19306), .C2(n19190), .A(n19171), .B(n19170), .ZN(
        P2_U3120) );
  AOI22_X1 U22160 ( .A1(n19236), .A2(n19185), .B1(n19384), .B2(n19196), .ZN(
        n19173) );
  AOI22_X1 U22161 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19187), .B1(
        n19385), .B2(n19186), .ZN(n19172) );
  OAI211_X1 U22162 ( .C1(n19239), .C2(n19190), .A(n19173), .B(n19172), .ZN(
        P2_U3121) );
  AOI22_X1 U22163 ( .A1(n19392), .A2(n19217), .B1(n19390), .B2(n19196), .ZN(
        n19175) );
  AOI22_X1 U22164 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19187), .B1(
        n19391), .B2(n19186), .ZN(n19174) );
  OAI211_X1 U22165 ( .C1(n19395), .C2(n19182), .A(n19175), .B(n19174), .ZN(
        P2_U3122) );
  AOI22_X1 U22166 ( .A1(n19311), .A2(n19217), .B1(n19396), .B2(n19196), .ZN(
        n19177) );
  AOI22_X1 U22167 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19187), .B1(
        n19397), .B2(n19186), .ZN(n19176) );
  OAI211_X1 U22168 ( .C1(n19315), .C2(n19182), .A(n19177), .B(n19176), .ZN(
        P2_U3123) );
  AOI22_X1 U22169 ( .A1(n19316), .A2(n19185), .B1(n19402), .B2(n19196), .ZN(
        n19179) );
  AOI22_X1 U22170 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19187), .B1(
        n19403), .B2(n19186), .ZN(n19178) );
  OAI211_X1 U22171 ( .C1(n19319), .C2(n19190), .A(n19179), .B(n19178), .ZN(
        P2_U3124) );
  AOI22_X1 U22172 ( .A1(n19280), .A2(n19217), .B1(n19408), .B2(n19196), .ZN(
        n19181) );
  AOI22_X1 U22173 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19187), .B1(
        n19409), .B2(n19186), .ZN(n19180) );
  OAI211_X1 U22174 ( .C1(n19283), .C2(n19182), .A(n19181), .B(n19180), .ZN(
        P2_U3125) );
  AOI22_X1 U22175 ( .A1(n19357), .A2(n19185), .B1(n9773), .B2(n19196), .ZN(
        n19184) );
  AOI22_X1 U22176 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19187), .B1(
        n19417), .B2(n19186), .ZN(n19183) );
  OAI211_X1 U22177 ( .C1(n19360), .C2(n19190), .A(n19184), .B(n19183), .ZN(
        P2_U3126) );
  AOI22_X1 U22178 ( .A1(n19325), .A2(n19185), .B1(n19423), .B2(n19196), .ZN(
        n19189) );
  AOI22_X1 U22179 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19187), .B1(
        n19424), .B2(n19186), .ZN(n19188) );
  OAI211_X1 U22180 ( .C1(n19330), .C2(n19190), .A(n19189), .B(n19188), .ZN(
        P2_U3127) );
  INV_X1 U22181 ( .A(n19226), .ZN(n19223) );
  AND2_X1 U22182 ( .A1(n19192), .A2(n19223), .ZN(n19215) );
  OAI21_X1 U22183 ( .B1(n19195), .B2(n19215), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19193) );
  OAI21_X1 U22184 ( .B1(n19226), .B2(n19194), .A(n19193), .ZN(n19216) );
  AOI22_X1 U22185 ( .A1(n19216), .A2(n19371), .B1(n19370), .B2(n19215), .ZN(
        n19202) );
  INV_X1 U22186 ( .A(n19195), .ZN(n19198) );
  AOI221_X1 U22187 ( .B1(n19254), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19217), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19196), .ZN(n19197) );
  MUX2_X1 U22188 ( .A(n19198), .B(n19197), .S(n19586), .Z(n19199) );
  NOR2_X1 U22189 ( .A1(n19199), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19200) );
  OAI21_X1 U22190 ( .B1(n19200), .B2(n19215), .A(n19377), .ZN(n19218) );
  AOI22_X1 U22191 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19218), .B1(
        n19217), .B2(n19303), .ZN(n19201) );
  OAI211_X1 U22192 ( .C1(n19306), .C2(n19221), .A(n19202), .B(n19201), .ZN(
        P2_U3128) );
  AOI22_X1 U22193 ( .A1(n19216), .A2(n19385), .B1(n19384), .B2(n19215), .ZN(
        n19204) );
  AOI22_X1 U22194 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19218), .B1(
        n19217), .B2(n19236), .ZN(n19203) );
  OAI211_X1 U22195 ( .C1(n19239), .C2(n19221), .A(n19204), .B(n19203), .ZN(
        P2_U3129) );
  AOI22_X1 U22196 ( .A1(n19216), .A2(n19391), .B1(n19390), .B2(n19215), .ZN(
        n19206) );
  AOI22_X1 U22197 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19218), .B1(
        n19217), .B2(n19240), .ZN(n19205) );
  OAI211_X1 U22198 ( .C1(n19243), .C2(n19221), .A(n19206), .B(n19205), .ZN(
        P2_U3130) );
  AOI22_X1 U22199 ( .A1(n19216), .A2(n19397), .B1(n19396), .B2(n19215), .ZN(
        n19208) );
  AOI22_X1 U22200 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19218), .B1(
        n19217), .B2(n19398), .ZN(n19207) );
  OAI211_X1 U22201 ( .C1(n19401), .C2(n19221), .A(n19208), .B(n19207), .ZN(
        P2_U3131) );
  AOI22_X1 U22202 ( .A1(n19216), .A2(n19403), .B1(n19402), .B2(n19215), .ZN(
        n19210) );
  AOI22_X1 U22203 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19218), .B1(
        n19217), .B2(n19316), .ZN(n19209) );
  OAI211_X1 U22204 ( .C1(n19319), .C2(n19221), .A(n19210), .B(n19209), .ZN(
        P2_U3132) );
  AOI22_X1 U22205 ( .A1(n19216), .A2(n19409), .B1(n19408), .B2(n19215), .ZN(
        n19212) );
  AOI22_X1 U22206 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19218), .B1(
        n19217), .B2(n19410), .ZN(n19211) );
  OAI211_X1 U22207 ( .C1(n19415), .C2(n19221), .A(n19212), .B(n19211), .ZN(
        P2_U3133) );
  AOI22_X1 U22208 ( .A1(n19216), .A2(n19417), .B1(n19416), .B2(n19215), .ZN(
        n19214) );
  AOI22_X1 U22209 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19218), .B1(
        n19217), .B2(n19357), .ZN(n19213) );
  OAI211_X1 U22210 ( .C1(n19360), .C2(n19221), .A(n19214), .B(n19213), .ZN(
        P2_U3134) );
  AOI22_X1 U22211 ( .A1(n19216), .A2(n19424), .B1(n19423), .B2(n19215), .ZN(
        n19220) );
  AOI22_X1 U22212 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19218), .B1(
        n19217), .B2(n19325), .ZN(n19219) );
  OAI211_X1 U22213 ( .C1(n19330), .C2(n19221), .A(n19220), .B(n19219), .ZN(
        P2_U3135) );
  INV_X1 U22214 ( .A(n19292), .ZN(n19222) );
  NAND2_X1 U22215 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19223), .ZN(
        n19231) );
  INV_X1 U22216 ( .A(n19231), .ZN(n19224) );
  NAND2_X1 U22217 ( .A1(n19224), .A2(n19535), .ZN(n19229) );
  INV_X1 U22218 ( .A(n19225), .ZN(n19228) );
  NOR2_X1 U22219 ( .A1(n19227), .A2(n19226), .ZN(n19252) );
  NOR3_X1 U22220 ( .A1(n19228), .A2(n19252), .A3(n19586), .ZN(n19230) );
  AOI21_X1 U22221 ( .B1(n19586), .B2(n19229), .A(n19230), .ZN(n19253) );
  AOI22_X1 U22222 ( .A1(n19253), .A2(n19371), .B1(n19370), .B2(n19252), .ZN(
        n19235) );
  NAND2_X1 U22223 ( .A1(n19372), .A2(n19536), .ZN(n19232) );
  AOI21_X1 U22224 ( .B1(n19232), .B2(n19231), .A(n19230), .ZN(n19233) );
  OAI211_X1 U22225 ( .C1(n19252), .C2(n19535), .A(n19233), .B(n19377), .ZN(
        n19255) );
  AOI22_X1 U22226 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19255), .B1(
        n19254), .B2(n19303), .ZN(n19234) );
  OAI211_X1 U22227 ( .C1(n19306), .C2(n19291), .A(n19235), .B(n19234), .ZN(
        P2_U3136) );
  AOI22_X1 U22228 ( .A1(n19253), .A2(n19385), .B1(n19384), .B2(n19252), .ZN(
        n19238) );
  AOI22_X1 U22229 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19255), .B1(
        n19254), .B2(n19236), .ZN(n19237) );
  OAI211_X1 U22230 ( .C1(n19239), .C2(n19291), .A(n19238), .B(n19237), .ZN(
        P2_U3137) );
  AOI22_X1 U22231 ( .A1(n19253), .A2(n19391), .B1(n19390), .B2(n19252), .ZN(
        n19242) );
  AOI22_X1 U22232 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19255), .B1(
        n19254), .B2(n19240), .ZN(n19241) );
  OAI211_X1 U22233 ( .C1(n19243), .C2(n19291), .A(n19242), .B(n19241), .ZN(
        P2_U3138) );
  AOI22_X1 U22234 ( .A1(n19253), .A2(n19397), .B1(n19396), .B2(n19252), .ZN(
        n19245) );
  AOI22_X1 U22235 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19255), .B1(
        n19254), .B2(n19398), .ZN(n19244) );
  OAI211_X1 U22236 ( .C1(n19401), .C2(n19291), .A(n19245), .B(n19244), .ZN(
        P2_U3139) );
  AOI22_X1 U22237 ( .A1(n19253), .A2(n19403), .B1(n19402), .B2(n19252), .ZN(
        n19247) );
  AOI22_X1 U22238 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19255), .B1(
        n19254), .B2(n19316), .ZN(n19246) );
  OAI211_X1 U22239 ( .C1(n19319), .C2(n19291), .A(n19247), .B(n19246), .ZN(
        P2_U3140) );
  AOI22_X1 U22240 ( .A1(n19253), .A2(n19409), .B1(n19408), .B2(n19252), .ZN(
        n19249) );
  AOI22_X1 U22241 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19255), .B1(
        n19254), .B2(n19410), .ZN(n19248) );
  OAI211_X1 U22242 ( .C1(n19415), .C2(n19291), .A(n19249), .B(n19248), .ZN(
        P2_U3141) );
  AOI22_X1 U22243 ( .A1(n19253), .A2(n19417), .B1(n9773), .B2(n19252), .ZN(
        n19251) );
  AOI22_X1 U22244 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19255), .B1(
        n19254), .B2(n19357), .ZN(n19250) );
  OAI211_X1 U22245 ( .C1(n19360), .C2(n19291), .A(n19251), .B(n19250), .ZN(
        P2_U3142) );
  AOI22_X1 U22246 ( .A1(n19253), .A2(n19424), .B1(n19423), .B2(n19252), .ZN(
        n19257) );
  AOI22_X1 U22247 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19255), .B1(
        n19254), .B2(n19325), .ZN(n19256) );
  OAI211_X1 U22248 ( .C1(n19330), .C2(n19291), .A(n19257), .B(n19256), .ZN(
        P2_U3143) );
  INV_X1 U22249 ( .A(n19258), .ZN(n19262) );
  NAND3_X1 U22250 ( .A1(n19560), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19300) );
  NOR2_X1 U22251 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19300), .ZN(
        n19286) );
  OAI21_X1 U22252 ( .B1(n19259), .B2(n19286), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19260) );
  OAI21_X1 U22253 ( .B1(n19262), .B2(n19261), .A(n19260), .ZN(n19287) );
  AOI22_X1 U22254 ( .A1(n19287), .A2(n19371), .B1(n19370), .B2(n19286), .ZN(
        n19271) );
  NOR2_X2 U22255 ( .A1(n19331), .A2(n19297), .ZN(n19326) );
  INV_X1 U22256 ( .A(n19326), .ZN(n19314) );
  AOI21_X1 U22257 ( .B1(n19291), .B2(n19314), .A(n19263), .ZN(n19269) );
  INV_X1 U22258 ( .A(n19286), .ZN(n19264) );
  OAI211_X1 U22259 ( .C1(n19265), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19264), 
        .B(n19533), .ZN(n19266) );
  AND2_X1 U22260 ( .A1(n19266), .A2(n19377), .ZN(n19267) );
  OAI211_X1 U22261 ( .C1(n19269), .C2(n19268), .A(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n19267), .ZN(n19288) );
  AOI22_X1 U22262 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19288), .B1(
        n19326), .B2(n19380), .ZN(n19270) );
  OAI211_X1 U22263 ( .C1(n19383), .C2(n19291), .A(n19271), .B(n19270), .ZN(
        P2_U3144) );
  AOI22_X1 U22264 ( .A1(n19287), .A2(n19385), .B1(n19384), .B2(n19286), .ZN(
        n19273) );
  AOI22_X1 U22265 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19288), .B1(
        n19326), .B2(n19386), .ZN(n19272) );
  OAI211_X1 U22266 ( .C1(n19389), .C2(n19291), .A(n19273), .B(n19272), .ZN(
        P2_U3145) );
  AOI22_X1 U22267 ( .A1(n19287), .A2(n19391), .B1(n19390), .B2(n19286), .ZN(
        n19275) );
  AOI22_X1 U22268 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19288), .B1(
        n19326), .B2(n19392), .ZN(n19274) );
  OAI211_X1 U22269 ( .C1(n19395), .C2(n19291), .A(n19275), .B(n19274), .ZN(
        P2_U3146) );
  AOI22_X1 U22270 ( .A1(n19287), .A2(n19397), .B1(n19396), .B2(n19286), .ZN(
        n19277) );
  AOI22_X1 U22271 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19288), .B1(
        n19326), .B2(n19311), .ZN(n19276) );
  OAI211_X1 U22272 ( .C1(n19315), .C2(n19291), .A(n19277), .B(n19276), .ZN(
        P2_U3147) );
  AOI22_X1 U22273 ( .A1(n19287), .A2(n19403), .B1(n19402), .B2(n19286), .ZN(
        n19279) );
  AOI22_X1 U22274 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19288), .B1(
        n19326), .B2(n19404), .ZN(n19278) );
  OAI211_X1 U22275 ( .C1(n19407), .C2(n19291), .A(n19279), .B(n19278), .ZN(
        P2_U3148) );
  AOI22_X1 U22276 ( .A1(n19287), .A2(n19409), .B1(n19408), .B2(n19286), .ZN(
        n19282) );
  AOI22_X1 U22277 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19288), .B1(
        n19326), .B2(n19280), .ZN(n19281) );
  OAI211_X1 U22278 ( .C1(n19283), .C2(n19291), .A(n19282), .B(n19281), .ZN(
        P2_U3149) );
  AOI22_X1 U22279 ( .A1(n19287), .A2(n19417), .B1(n9773), .B2(n19286), .ZN(
        n19285) );
  AOI22_X1 U22280 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19288), .B1(
        n19326), .B2(n19418), .ZN(n19284) );
  OAI211_X1 U22281 ( .C1(n19421), .C2(n19291), .A(n19285), .B(n19284), .ZN(
        P2_U3150) );
  AOI22_X1 U22282 ( .A1(n19287), .A2(n19424), .B1(n19423), .B2(n19286), .ZN(
        n19290) );
  AOI22_X1 U22283 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19288), .B1(
        n19326), .B2(n19426), .ZN(n19289) );
  OAI211_X1 U22284 ( .C1(n19432), .C2(n19291), .A(n19290), .B(n19289), .ZN(
        P2_U3151) );
  INV_X1 U22285 ( .A(n19293), .ZN(n19294) );
  NOR2_X1 U22286 ( .A1(n19571), .A2(n19300), .ZN(n19335) );
  NOR3_X1 U22287 ( .A1(n19294), .A2(n19335), .A3(n19586), .ZN(n19299) );
  INV_X1 U22288 ( .A(n19300), .ZN(n19295) );
  AOI21_X1 U22289 ( .B1(n19535), .B2(n19295), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19296) );
  NOR2_X1 U22290 ( .A1(n19299), .A2(n19296), .ZN(n19324) );
  AOI22_X1 U22291 ( .A1(n19324), .A2(n19371), .B1(n19370), .B2(n19335), .ZN(
        n19305) );
  INV_X1 U22292 ( .A(n19297), .ZN(n19298) );
  NAND2_X1 U22293 ( .A1(n19372), .A2(n19298), .ZN(n19301) );
  AOI21_X1 U22294 ( .B1(n19301), .B2(n19300), .A(n19299), .ZN(n19302) );
  OAI211_X1 U22295 ( .C1(n19335), .C2(n19535), .A(n19302), .B(n19377), .ZN(
        n19327) );
  AOI22_X1 U22296 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19327), .B1(
        n19326), .B2(n19303), .ZN(n19304) );
  OAI211_X1 U22297 ( .C1(n19306), .C2(n19366), .A(n19305), .B(n19304), .ZN(
        P2_U3152) );
  AOI22_X1 U22298 ( .A1(n19324), .A2(n19385), .B1(n19384), .B2(n19335), .ZN(
        n19308) );
  AOI22_X1 U22299 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19327), .B1(
        n19356), .B2(n19386), .ZN(n19307) );
  OAI211_X1 U22300 ( .C1(n19389), .C2(n19314), .A(n19308), .B(n19307), .ZN(
        P2_U3153) );
  AOI22_X1 U22301 ( .A1(n19324), .A2(n19391), .B1(n19390), .B2(n19335), .ZN(
        n19310) );
  AOI22_X1 U22302 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19327), .B1(
        n19356), .B2(n19392), .ZN(n19309) );
  OAI211_X1 U22303 ( .C1(n19395), .C2(n19314), .A(n19310), .B(n19309), .ZN(
        P2_U3154) );
  AOI22_X1 U22304 ( .A1(n19324), .A2(n19397), .B1(n19396), .B2(n19335), .ZN(
        n19313) );
  AOI22_X1 U22305 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19327), .B1(
        n19356), .B2(n19311), .ZN(n19312) );
  OAI211_X1 U22306 ( .C1(n19315), .C2(n19314), .A(n19313), .B(n19312), .ZN(
        P2_U3155) );
  AOI22_X1 U22307 ( .A1(n19324), .A2(n19403), .B1(n19402), .B2(n19335), .ZN(
        n19318) );
  AOI22_X1 U22308 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19327), .B1(
        n19326), .B2(n19316), .ZN(n19317) );
  OAI211_X1 U22309 ( .C1(n19319), .C2(n19366), .A(n19318), .B(n19317), .ZN(
        P2_U3156) );
  AOI22_X1 U22310 ( .A1(n19324), .A2(n19409), .B1(n19408), .B2(n19335), .ZN(
        n19321) );
  AOI22_X1 U22311 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19327), .B1(
        n19326), .B2(n19410), .ZN(n19320) );
  OAI211_X1 U22312 ( .C1(n19415), .C2(n19366), .A(n19321), .B(n19320), .ZN(
        P2_U3157) );
  AOI22_X1 U22313 ( .A1(n19324), .A2(n19417), .B1(n9773), .B2(n19335), .ZN(
        n19323) );
  AOI22_X1 U22314 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19327), .B1(
        n19326), .B2(n19357), .ZN(n19322) );
  OAI211_X1 U22315 ( .C1(n19360), .C2(n19366), .A(n19323), .B(n19322), .ZN(
        P2_U3158) );
  AOI22_X1 U22316 ( .A1(n19324), .A2(n19424), .B1(n19423), .B2(n19335), .ZN(
        n19329) );
  AOI22_X1 U22317 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19327), .B1(
        n19326), .B2(n19325), .ZN(n19328) );
  OAI211_X1 U22318 ( .C1(n19330), .C2(n19366), .A(n19329), .B(n19328), .ZN(
        P2_U3159) );
  NAND2_X1 U22319 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19332), .ZN(
        n19375) );
  NOR2_X1 U22320 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19375), .ZN(
        n19361) );
  AOI22_X1 U22321 ( .A1(n19380), .A2(n19411), .B1(n19370), .B2(n19361), .ZN(
        n19345) );
  OAI21_X1 U22322 ( .B1(n19411), .B2(n19356), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19334) );
  NAND2_X1 U22323 ( .A1(n19334), .A2(n19333), .ZN(n19343) );
  NOR2_X1 U22324 ( .A1(n19361), .A2(n19335), .ZN(n19342) );
  INV_X1 U22325 ( .A(n19342), .ZN(n19339) );
  INV_X1 U22326 ( .A(n19340), .ZN(n19337) );
  INV_X1 U22327 ( .A(n19361), .ZN(n19336) );
  OAI211_X1 U22328 ( .C1(n19337), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19336), 
        .B(n19533), .ZN(n19338) );
  OAI211_X1 U22329 ( .C1(n19343), .C2(n19339), .A(n19377), .B(n19338), .ZN(
        n19363) );
  OAI21_X1 U22330 ( .B1(n19340), .B2(n19361), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19341) );
  AOI22_X1 U22331 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19363), .B1(
        n19371), .B2(n19362), .ZN(n19344) );
  OAI211_X1 U22332 ( .C1(n19383), .C2(n19366), .A(n19345), .B(n19344), .ZN(
        P2_U3160) );
  AOI22_X1 U22333 ( .A1(n19386), .A2(n19411), .B1(n19384), .B2(n19361), .ZN(
        n19347) );
  AOI22_X1 U22334 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19363), .B1(
        n19385), .B2(n19362), .ZN(n19346) );
  OAI211_X1 U22335 ( .C1(n19389), .C2(n19366), .A(n19347), .B(n19346), .ZN(
        P2_U3161) );
  AOI22_X1 U22336 ( .A1(n19392), .A2(n19411), .B1(n19390), .B2(n19361), .ZN(
        n19349) );
  AOI22_X1 U22337 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19363), .B1(
        n19391), .B2(n19362), .ZN(n19348) );
  OAI211_X1 U22338 ( .C1(n19395), .C2(n19366), .A(n19349), .B(n19348), .ZN(
        P2_U3162) );
  AOI22_X1 U22339 ( .A1(n19398), .A2(n19356), .B1(n19396), .B2(n19361), .ZN(
        n19351) );
  AOI22_X1 U22340 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19363), .B1(
        n19397), .B2(n19362), .ZN(n19350) );
  OAI211_X1 U22341 ( .C1(n19401), .C2(n19431), .A(n19351), .B(n19350), .ZN(
        P2_U3163) );
  AOI22_X1 U22342 ( .A1(n19404), .A2(n19411), .B1(n19402), .B2(n19361), .ZN(
        n19353) );
  AOI22_X1 U22343 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19363), .B1(
        n19403), .B2(n19362), .ZN(n19352) );
  OAI211_X1 U22344 ( .C1(n19407), .C2(n19366), .A(n19353), .B(n19352), .ZN(
        P2_U3164) );
  AOI22_X1 U22345 ( .A1(n19410), .A2(n19356), .B1(n19408), .B2(n19361), .ZN(
        n19355) );
  AOI22_X1 U22346 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19363), .B1(
        n19409), .B2(n19362), .ZN(n19354) );
  OAI211_X1 U22347 ( .C1(n19415), .C2(n19431), .A(n19355), .B(n19354), .ZN(
        P2_U3165) );
  AOI22_X1 U22348 ( .A1(n19357), .A2(n19356), .B1(n9773), .B2(n19361), .ZN(
        n19359) );
  AOI22_X1 U22349 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19363), .B1(
        n19417), .B2(n19362), .ZN(n19358) );
  OAI211_X1 U22350 ( .C1(n19360), .C2(n19431), .A(n19359), .B(n19358), .ZN(
        P2_U3166) );
  AOI22_X1 U22351 ( .A1(n19426), .A2(n19411), .B1(n19423), .B2(n19361), .ZN(
        n19365) );
  AOI22_X1 U22352 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19363), .B1(
        n19424), .B2(n19362), .ZN(n19364) );
  OAI211_X1 U22353 ( .C1(n19432), .C2(n19366), .A(n19365), .B(n19364), .ZN(
        P2_U3167) );
  INV_X1 U22354 ( .A(n19422), .ZN(n19367) );
  NAND3_X1 U22355 ( .A1(n19368), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19367), 
        .ZN(n19376) );
  OAI21_X1 U22356 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19375), .A(n19586), 
        .ZN(n19369) );
  AND2_X1 U22357 ( .A1(n19376), .A2(n19369), .ZN(n19425) );
  AOI22_X1 U22358 ( .A1(n19425), .A2(n19371), .B1(n19370), .B2(n19422), .ZN(
        n19382) );
  INV_X1 U22359 ( .A(n19372), .ZN(n19374) );
  NOR3_X1 U22360 ( .A1(n19374), .A2(P2_STATE2_REG_3__SCAN_IN), .A3(n19373), 
        .ZN(n19379) );
  AOI21_X1 U22361 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19571), .A(n19375), 
        .ZN(n19378) );
  OAI211_X1 U22362 ( .C1(n19379), .C2(n19378), .A(n19377), .B(n19376), .ZN(
        n19428) );
  AOI22_X1 U22363 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19428), .B1(
        n19427), .B2(n19380), .ZN(n19381) );
  OAI211_X1 U22364 ( .C1(n19383), .C2(n19431), .A(n19382), .B(n19381), .ZN(
        P2_U3168) );
  AOI22_X1 U22365 ( .A1(n19425), .A2(n19385), .B1(n19384), .B2(n19422), .ZN(
        n19388) );
  AOI22_X1 U22366 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19428), .B1(
        n19427), .B2(n19386), .ZN(n19387) );
  OAI211_X1 U22367 ( .C1(n19389), .C2(n19431), .A(n19388), .B(n19387), .ZN(
        P2_U3169) );
  AOI22_X1 U22368 ( .A1(n19425), .A2(n19391), .B1(n19390), .B2(n19422), .ZN(
        n19394) );
  AOI22_X1 U22369 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19428), .B1(
        n19427), .B2(n19392), .ZN(n19393) );
  OAI211_X1 U22370 ( .C1(n19395), .C2(n19431), .A(n19394), .B(n19393), .ZN(
        P2_U3170) );
  AOI22_X1 U22371 ( .A1(n19425), .A2(n19397), .B1(n19396), .B2(n19422), .ZN(
        n19400) );
  AOI22_X1 U22372 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19428), .B1(
        n19411), .B2(n19398), .ZN(n19399) );
  OAI211_X1 U22373 ( .C1(n19401), .C2(n19414), .A(n19400), .B(n19399), .ZN(
        P2_U3171) );
  AOI22_X1 U22374 ( .A1(n19425), .A2(n19403), .B1(n19402), .B2(n19422), .ZN(
        n19406) );
  AOI22_X1 U22375 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19428), .B1(
        n19427), .B2(n19404), .ZN(n19405) );
  OAI211_X1 U22376 ( .C1(n19407), .C2(n19431), .A(n19406), .B(n19405), .ZN(
        P2_U3172) );
  AOI22_X1 U22377 ( .A1(n19425), .A2(n19409), .B1(n19408), .B2(n19422), .ZN(
        n19413) );
  AOI22_X1 U22378 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19428), .B1(
        n19411), .B2(n19410), .ZN(n19412) );
  OAI211_X1 U22379 ( .C1(n19415), .C2(n19414), .A(n19413), .B(n19412), .ZN(
        P2_U3173) );
  AOI22_X1 U22380 ( .A1(n19425), .A2(n19417), .B1(n9773), .B2(n19422), .ZN(
        n19420) );
  AOI22_X1 U22381 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19428), .B1(
        n19427), .B2(n19418), .ZN(n19419) );
  OAI211_X1 U22382 ( .C1(n19421), .C2(n19431), .A(n19420), .B(n19419), .ZN(
        P2_U3174) );
  AOI22_X1 U22383 ( .A1(n19425), .A2(n19424), .B1(n19423), .B2(n19422), .ZN(
        n19430) );
  AOI22_X1 U22384 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19428), .B1(
        n19427), .B2(n19426), .ZN(n19429) );
  OAI211_X1 U22385 ( .C1(n19432), .C2(n19431), .A(n19430), .B(n19429), .ZN(
        P2_U3175) );
  OAI211_X1 U22386 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19593), .A(n19434), 
        .B(n19433), .ZN(n19439) );
  OAI21_X1 U22387 ( .B1(n19436), .B2(n19435), .A(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n19438) );
  OAI211_X1 U22388 ( .C1(n19440), .C2(n19439), .A(n19438), .B(n19437), .ZN(
        P2_U3177) );
  AND2_X1 U22389 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19441), .ZN(
        P2_U3179) );
  INV_X1 U22390 ( .A(P2_DATAWIDTH_REG_30__SCAN_IN), .ZN(n20653) );
  NOR2_X1 U22391 ( .A1(n20653), .A2(n19518), .ZN(P2_U3180) );
  AND2_X1 U22392 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19441), .ZN(
        P2_U3181) );
  AND2_X1 U22393 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19441), .ZN(
        P2_U3182) );
  AND2_X1 U22394 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19441), .ZN(
        P2_U3183) );
  AND2_X1 U22395 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19441), .ZN(
        P2_U3184) );
  AND2_X1 U22396 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19441), .ZN(
        P2_U3185) );
  AND2_X1 U22397 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19441), .ZN(
        P2_U3186) );
  AND2_X1 U22398 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19441), .ZN(
        P2_U3187) );
  AND2_X1 U22399 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19441), .ZN(
        P2_U3188) );
  AND2_X1 U22400 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19441), .ZN(
        P2_U3189) );
  AND2_X1 U22401 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19441), .ZN(
        P2_U3190) );
  AND2_X1 U22402 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19441), .ZN(
        P2_U3191) );
  AND2_X1 U22403 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19441), .ZN(
        P2_U3192) );
  AND2_X1 U22404 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19441), .ZN(
        P2_U3193) );
  AND2_X1 U22405 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19441), .ZN(
        P2_U3194) );
  AND2_X1 U22406 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19441), .ZN(
        P2_U3195) );
  AND2_X1 U22407 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19441), .ZN(
        P2_U3196) );
  AND2_X1 U22408 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19441), .ZN(
        P2_U3197) );
  AND2_X1 U22409 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19441), .ZN(
        P2_U3198) );
  AND2_X1 U22410 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19441), .ZN(
        P2_U3199) );
  AND2_X1 U22411 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19441), .ZN(
        P2_U3200) );
  AND2_X1 U22412 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19441), .ZN(P2_U3201) );
  AND2_X1 U22413 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19441), .ZN(P2_U3202) );
  AND2_X1 U22414 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19441), .ZN(P2_U3203) );
  AND2_X1 U22415 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19441), .ZN(P2_U3204) );
  AND2_X1 U22416 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19441), .ZN(P2_U3205) );
  AND2_X1 U22417 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19441), .ZN(P2_U3206) );
  AND2_X1 U22418 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19441), .ZN(P2_U3207) );
  AND2_X1 U22419 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19441), .ZN(P2_U3208) );
  NOR2_X1 U22420 ( .A1(n20458), .A2(n19447), .ZN(n19460) );
  INV_X1 U22421 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19446) );
  NOR2_X1 U22422 ( .A1(n19442), .A2(n19446), .ZN(n19443) );
  NAND2_X1 U22423 ( .A1(n19587), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19455) );
  AOI21_X1 U22424 ( .B1(n19443), .B2(n19455), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19445) );
  AOI211_X1 U22425 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n19451), .A(
        n19454), .B(n19509), .ZN(n19444) );
  OR3_X1 U22426 ( .A1(n19460), .A2(n19445), .A3(n19444), .ZN(P2_U3209) );
  AOI21_X1 U22427 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n19451), .A(n20627), 
        .ZN(n19452) );
  NOR2_X1 U22428 ( .A1(n19446), .A2(n19452), .ZN(n19448) );
  AOI21_X1 U22429 ( .B1(n19448), .B2(n19447), .A(n19582), .ZN(n19449) );
  OAI211_X1 U22430 ( .C1(n19451), .C2(n19450), .A(n19449), .B(n19455), .ZN(
        P2_U3210) );
  AOI21_X1 U22431 ( .B1(n19453), .B2(n19587), .A(n19452), .ZN(n19459) );
  INV_X1 U22432 ( .A(n19454), .ZN(n19456) );
  OAI22_X1 U22433 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19456), .B1(NA), 
        .B2(n19455), .ZN(n19457) );
  OAI211_X1 U22434 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19457), .ZN(n19458) );
  OAI21_X1 U22435 ( .B1(n19460), .B2(n19459), .A(n19458), .ZN(P2_U3211) );
  OAI222_X1 U22436 ( .A1(n19508), .A2(n19462), .B1(n19461), .B2(n19509), .C1(
        n19463), .C2(n19511), .ZN(P2_U3212) );
  OAI222_X1 U22437 ( .A1(n19511), .A2(n12102), .B1(n19464), .B2(n19509), .C1(
        n19463), .C2(n19508), .ZN(P2_U3213) );
  OAI222_X1 U22438 ( .A1(n19511), .A2(n12030), .B1(n19465), .B2(n19509), .C1(
        n12102), .C2(n19508), .ZN(P2_U3214) );
  INV_X1 U22439 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n19466) );
  OAI222_X1 U22440 ( .A1(n19511), .A2(n19466), .B1(n20626), .B2(n19509), .C1(
        n12030), .C2(n19508), .ZN(P2_U3215) );
  OAI222_X1 U22441 ( .A1(n19511), .A2(n19468), .B1(n19467), .B2(n19509), .C1(
        n19466), .C2(n19508), .ZN(P2_U3216) );
  OAI222_X1 U22442 ( .A1(n19511), .A2(n19470), .B1(n19469), .B2(n19509), .C1(
        n19468), .C2(n19508), .ZN(P2_U3217) );
  OAI222_X1 U22443 ( .A1(n19511), .A2(n12016), .B1(n19471), .B2(n19509), .C1(
        n19470), .C2(n19508), .ZN(P2_U3218) );
  OAI222_X1 U22444 ( .A1(n19511), .A2(n12156), .B1(n19472), .B2(n19509), .C1(
        n12016), .C2(n19508), .ZN(P2_U3219) );
  OAI222_X1 U22445 ( .A1(n19511), .A2(n12159), .B1(n19473), .B2(n19509), .C1(
        n12156), .C2(n19508), .ZN(P2_U3220) );
  OAI222_X1 U22446 ( .A1(n19511), .A2(n12161), .B1(n19474), .B2(n19509), .C1(
        n12159), .C2(n19508), .ZN(P2_U3221) );
  OAI222_X1 U22447 ( .A1(n19511), .A2(n12012), .B1(n19475), .B2(n19509), .C1(
        n12161), .C2(n19508), .ZN(P2_U3222) );
  OAI222_X1 U22448 ( .A1(n19511), .A2(n19477), .B1(n19476), .B2(n19509), .C1(
        n12012), .C2(n19508), .ZN(P2_U3223) );
  OAI222_X1 U22449 ( .A1(n19511), .A2(n12172), .B1(n19478), .B2(n19509), .C1(
        n19477), .C2(n19508), .ZN(P2_U3224) );
  OAI222_X1 U22450 ( .A1(n19511), .A2(n19480), .B1(n19479), .B2(n19509), .C1(
        n12172), .C2(n19508), .ZN(P2_U3225) );
  OAI222_X1 U22451 ( .A1(n19511), .A2(n12178), .B1(n19481), .B2(n19509), .C1(
        n19480), .C2(n19508), .ZN(P2_U3226) );
  OAI222_X1 U22452 ( .A1(n19511), .A2(n19483), .B1(n19482), .B2(n19509), .C1(
        n12178), .C2(n19508), .ZN(P2_U3227) );
  OAI222_X1 U22453 ( .A1(n19511), .A2(n19485), .B1(n19484), .B2(n19509), .C1(
        n19483), .C2(n19508), .ZN(P2_U3228) );
  OAI222_X1 U22454 ( .A1(n19511), .A2(n19487), .B1(n19486), .B2(n19509), .C1(
        n19485), .C2(n19508), .ZN(P2_U3229) );
  OAI222_X1 U22455 ( .A1(n19511), .A2(n14754), .B1(n19488), .B2(n19509), .C1(
        n19487), .C2(n19508), .ZN(P2_U3230) );
  OAI222_X1 U22456 ( .A1(n19511), .A2(n19490), .B1(n19489), .B2(n19509), .C1(
        n14754), .C2(n19508), .ZN(P2_U3231) );
  OAI222_X1 U22457 ( .A1(n19511), .A2(n19492), .B1(n19491), .B2(n19509), .C1(
        n19490), .C2(n19508), .ZN(P2_U3232) );
  OAI222_X1 U22458 ( .A1(n19511), .A2(n19494), .B1(n19493), .B2(n19509), .C1(
        n19492), .C2(n19508), .ZN(P2_U3233) );
  OAI222_X1 U22459 ( .A1(n19511), .A2(n19496), .B1(n19495), .B2(n19509), .C1(
        n19494), .C2(n19508), .ZN(P2_U3234) );
  INV_X1 U22460 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19498) );
  OAI222_X1 U22461 ( .A1(n19511), .A2(n19498), .B1(n19497), .B2(n19509), .C1(
        n19496), .C2(n19508), .ZN(P2_U3235) );
  INV_X1 U22462 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19500) );
  OAI222_X1 U22463 ( .A1(n19511), .A2(n19500), .B1(n19499), .B2(n19509), .C1(
        n19498), .C2(n19508), .ZN(P2_U3236) );
  OAI222_X1 U22464 ( .A1(n19511), .A2(n19503), .B1(n19501), .B2(n19509), .C1(
        n19500), .C2(n19508), .ZN(P2_U3237) );
  INV_X1 U22465 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19504) );
  OAI222_X1 U22466 ( .A1(n19508), .A2(n19503), .B1(n19502), .B2(n19509), .C1(
        n19504), .C2(n19511), .ZN(P2_U3238) );
  INV_X1 U22467 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19506) );
  OAI222_X1 U22468 ( .A1(n19511), .A2(n19506), .B1(n19505), .B2(n19509), .C1(
        n19504), .C2(n19508), .ZN(P2_U3239) );
  OAI222_X1 U22469 ( .A1(n19511), .A2(n13872), .B1(n19507), .B2(n19509), .C1(
        n19506), .C2(n19508), .ZN(P2_U3240) );
  OAI222_X1 U22470 ( .A1(n19511), .A2(n14828), .B1(n19510), .B2(n19509), .C1(
        n13872), .C2(n19508), .ZN(P2_U3241) );
  OAI22_X1 U22471 ( .A1(n19597), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n19509), .ZN(n19512) );
  INV_X1 U22472 ( .A(n19512), .ZN(P2_U3585) );
  MUX2_X1 U22473 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n19597), .Z(P2_U3586) );
  OAI22_X1 U22474 ( .A1(n19597), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n19509), .ZN(n19513) );
  INV_X1 U22475 ( .A(n19513), .ZN(P2_U3587) );
  OAI22_X1 U22476 ( .A1(n19597), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n19509), .ZN(n19514) );
  INV_X1 U22477 ( .A(n19514), .ZN(P2_U3588) );
  OAI21_X1 U22478 ( .B1(n19518), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19516), 
        .ZN(n19515) );
  INV_X1 U22479 ( .A(n19515), .ZN(P2_U3591) );
  OAI21_X1 U22480 ( .B1(n19518), .B2(n19517), .A(n19516), .ZN(P2_U3592) );
  INV_X1 U22481 ( .A(n19519), .ZN(n19520) );
  OAI22_X1 U22482 ( .A1(n19540), .A2(n19525), .B1(n19537), .B2(n19520), .ZN(
        n19522) );
  OAI22_X1 U22483 ( .A1(n19530), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n19522), .B2(n19521), .ZN(n19523) );
  INV_X1 U22484 ( .A(n19523), .ZN(P2_U3596) );
  OAI22_X1 U22485 ( .A1(n19546), .A2(n19525), .B1(n19537), .B2(n19524), .ZN(
        n19526) );
  INV_X1 U22486 ( .A(n19526), .ZN(n19527) );
  OAI21_X1 U22487 ( .B1(n19529), .B2(n19528), .A(n19527), .ZN(n19531) );
  MUX2_X1 U22488 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n19531), .S(
        n19530), .Z(P2_U3599) );
  OAI22_X1 U22489 ( .A1(n19535), .A2(n19534), .B1(n19533), .B2(n19532), .ZN(
        n19542) );
  NAND2_X1 U22490 ( .A1(n19536), .A2(n19552), .ZN(n19544) );
  NAND3_X1 U22491 ( .A1(n19538), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19537), 
        .ZN(n19539) );
  NAND2_X1 U22492 ( .A1(n19539), .A2(n19561), .ZN(n19545) );
  AOI21_X1 U22493 ( .B1(n19544), .B2(n19545), .A(n19540), .ZN(n19541) );
  OAI21_X1 U22494 ( .B1(n19542), .B2(n19541), .A(n19570), .ZN(n19543) );
  OAI21_X1 U22495 ( .B1(n19570), .B2(n12827), .A(n19543), .ZN(P2_U3602) );
  INV_X1 U22496 ( .A(n19570), .ZN(n19569) );
  OAI21_X1 U22497 ( .B1(n19546), .B2(n19545), .A(n19544), .ZN(n19547) );
  AOI21_X1 U22498 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19548), .A(n19547), 
        .ZN(n19549) );
  AOI22_X1 U22499 ( .A1(n19569), .A2(n19550), .B1(n19549), .B2(n19570), .ZN(
        P2_U3603) );
  NAND2_X1 U22500 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATEBS16_REG_SCAN_IN), .ZN(n19551) );
  NAND2_X1 U22501 ( .A1(n19561), .A2(n19551), .ZN(n19556) );
  NAND2_X1 U22502 ( .A1(n19557), .A2(n19552), .ZN(n19555) );
  NAND2_X1 U22503 ( .A1(n19553), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19554) );
  OAI211_X1 U22504 ( .C1(n19557), .C2(n19556), .A(n19555), .B(n19554), .ZN(
        n19558) );
  INV_X1 U22505 ( .A(n19558), .ZN(n19559) );
  AOI22_X1 U22506 ( .A1(n19569), .A2(n19560), .B1(n19559), .B2(n19570), .ZN(
        P2_U3604) );
  INV_X1 U22507 ( .A(n19561), .ZN(n19565) );
  INV_X1 U22508 ( .A(n19562), .ZN(n19564) );
  OAI22_X1 U22509 ( .A1(n19566), .A2(n19565), .B1(n19564), .B2(n19563), .ZN(
        n19567) );
  AOI21_X1 U22510 ( .B1(n19571), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19567), 
        .ZN(n19568) );
  OAI22_X1 U22511 ( .A1(n19571), .A2(n19570), .B1(n19569), .B2(n19568), .ZN(
        P2_U3605) );
  INV_X1 U22512 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20630) );
  AOI22_X1 U22513 ( .A1(n19509), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20630), 
        .B2(n19597), .ZN(P2_U3608) );
  INV_X1 U22514 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n19580) );
  INV_X1 U22515 ( .A(n19572), .ZN(n19576) );
  OAI22_X1 U22516 ( .A1(n19576), .A2(n19575), .B1(n19574), .B2(n19573), .ZN(
        n19578) );
  OAI21_X1 U22517 ( .B1(n19578), .B2(n19577), .A(n19581), .ZN(n19579) );
  OAI21_X1 U22518 ( .B1(n19581), .B2(n19580), .A(n19579), .ZN(P2_U3609) );
  OAI21_X1 U22519 ( .B1(n12005), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19582), 
        .ZN(n19583) );
  NAND3_X1 U22520 ( .A1(n19584), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n19583), 
        .ZN(n19589) );
  OAI21_X1 U22521 ( .B1(n19587), .B2(n19586), .A(n19585), .ZN(n19588) );
  NAND2_X1 U22522 ( .A1(n19589), .A2(n19588), .ZN(n19596) );
  OAI21_X1 U22523 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19591), .A(n19590), 
        .ZN(n19592) );
  AOI21_X1 U22524 ( .B1(n19594), .B2(n19593), .A(n19592), .ZN(n19595) );
  MUX2_X1 U22525 ( .A(n19596), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n19595), 
        .Z(P2_U3610) );
  MUX2_X1 U22526 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .B(P2_M_IO_N_REG_SCAN_IN), 
        .S(n19597), .Z(P2_U3611) );
  OAI21_X1 U22527 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n19598), .A(
        P1_STATE_REG_0__SCAN_IN), .ZN(n20459) );
  NAND2_X2 U22528 ( .A1(n20451), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20503) );
  OAI21_X1 U22529 ( .B1(n20459), .B2(P1_ADS_N_REG_SCAN_IN), .A(n20503), .ZN(
        n19599) );
  INV_X1 U22530 ( .A(n19599), .ZN(P1_U2802) );
  INV_X1 U22531 ( .A(n19600), .ZN(n19605) );
  INV_X1 U22532 ( .A(n19601), .ZN(n19603) );
  OAI21_X1 U22533 ( .B1(n19603), .B2(n19602), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19604) );
  OAI21_X1 U22534 ( .B1(n19605), .B2(n20446), .A(n19604), .ZN(P1_U2803) );
  NOR2_X1 U22535 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19607) );
  OAI21_X1 U22536 ( .B1(n19607), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20503), .ZN(
        n19606) );
  OAI21_X1 U22537 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20503), .A(n19606), 
        .ZN(P1_U2804) );
  NAND2_X1 U22538 ( .A1(n20459), .A2(n20503), .ZN(n20514) );
  INV_X1 U22539 ( .A(n20514), .ZN(n20450) );
  OAI21_X1 U22540 ( .B1(BS16), .B2(n19607), .A(n20450), .ZN(n20512) );
  OAI21_X1 U22541 ( .B1(n20450), .B2(n20347), .A(n20512), .ZN(P1_U2805) );
  OAI21_X1 U22542 ( .B1(n19610), .B2(n19609), .A(n19608), .ZN(P1_U2806) );
  NOR4_X1 U22543 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_26__SCAN_IN), .A3(P1_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_28__SCAN_IN), .ZN(n19614) );
  NOR4_X1 U22544 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_18__SCAN_IN), .A3(P1_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_17__SCAN_IN), .ZN(n19613) );
  NOR4_X1 U22545 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_24__SCAN_IN), .ZN(n19612) );
  NOR4_X1 U22546 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_19__SCAN_IN), .A3(P1_DATAWIDTH_REG_20__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_21__SCAN_IN), .ZN(n19611) );
  NAND4_X1 U22547 ( .A1(n19614), .A2(n19613), .A3(n19612), .A4(n19611), .ZN(
        n19619) );
  NOR4_X1 U22548 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n20556) );
  AOI211_X1 U22549 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n19617) );
  NOR4_X1 U22550 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_10__SCAN_IN), .A3(P1_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n19616) );
  NOR4_X1 U22551 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_6__SCAN_IN), .A3(P1_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19615) );
  NAND4_X1 U22552 ( .A1(n20556), .A2(n19617), .A3(n19616), .A4(n19615), .ZN(
        n19618) );
  NOR2_X1 U22553 ( .A1(n19619), .A2(n19618), .ZN(n20538) );
  INV_X1 U22554 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19621) );
  NOR3_X1 U22555 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19622) );
  OAI21_X1 U22556 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19622), .A(n20538), .ZN(
        n19620) );
  OAI21_X1 U22557 ( .B1(n20538), .B2(n19621), .A(n19620), .ZN(P1_U2807) );
  INV_X1 U22558 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19624) );
  NOR2_X1 U22559 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20532) );
  OAI21_X1 U22560 ( .B1(n19622), .B2(n20532), .A(n20538), .ZN(n19623) );
  OAI21_X1 U22561 ( .B1(n20538), .B2(n19624), .A(n19623), .ZN(P1_U2808) );
  OR2_X1 U22562 ( .A1(n19625), .A2(n19665), .ZN(n19635) );
  AOI22_X1 U22563 ( .A1(P1_EBX_REG_9__SCAN_IN), .A2(n19687), .B1(n19686), .B2(
        n19626), .ZN(n19627) );
  OAI21_X1 U22564 ( .B1(n19629), .B2(n19628), .A(n19627), .ZN(n19630) );
  AOI211_X1 U22565 ( .C1(n19675), .C2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n19678), .B(n19630), .ZN(n19634) );
  AOI22_X1 U22566 ( .A1(n19632), .A2(n19659), .B1(n19644), .B2(n19631), .ZN(
        n19633) );
  OAI211_X1 U22567 ( .C1(P1_REIP_REG_9__SCAN_IN), .C2(n19635), .A(n19634), .B(
        n19633), .ZN(P1_U2831) );
  NAND2_X1 U22568 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n19637) );
  OAI21_X1 U22569 ( .B1(n19637), .B2(n19667), .A(n19636), .ZN(n19657) );
  NAND2_X1 U22570 ( .A1(n19638), .A2(n19659), .ZN(n19648) );
  OAI22_X1 U22571 ( .A1(n19640), .A2(n19662), .B1(n19681), .B2(n19639), .ZN(
        n19641) );
  AOI211_X1 U22572 ( .C1(n19675), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n19678), .B(n19641), .ZN(n19647) );
  NAND4_X1 U22573 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .A3(n19651), .A4(n19650), .ZN(n19646) );
  INV_X1 U22574 ( .A(n19642), .ZN(n19643) );
  NAND2_X1 U22575 ( .A1(n19644), .A2(n19643), .ZN(n19645) );
  AND4_X1 U22576 ( .A1(n19648), .A2(n19647), .A3(n19646), .A4(n19645), .ZN(
        n19649) );
  OAI21_X1 U22577 ( .B1(n19657), .B2(n19650), .A(n19649), .ZN(P1_U2833) );
  INV_X1 U22578 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20596) );
  NAND3_X1 U22579 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n19651), .A3(n20596), 
        .ZN(n19652) );
  OAI211_X1 U22580 ( .C1(n19691), .C2(n19654), .A(n19653), .B(n19652), .ZN(
        n19655) );
  AOI21_X1 U22581 ( .B1(n19686), .B2(n19704), .A(n19655), .ZN(n19661) );
  OAI22_X1 U22582 ( .A1(n19657), .A2(n20596), .B1(n19656), .B2(n19690), .ZN(
        n19658) );
  AOI21_X1 U22583 ( .B1(n19659), .B2(n19707), .A(n19658), .ZN(n19660) );
  OAI211_X1 U22584 ( .C1(n19709), .C2(n19662), .A(n19661), .B(n19660), .ZN(
        P1_U2834) );
  AOI22_X1 U22585 ( .A1(P1_EBX_REG_5__SCAN_IN), .A2(n19687), .B1(n19686), .B2(
        n19663), .ZN(n19664) );
  OAI21_X1 U22586 ( .B1(P1_REIP_REG_5__SCAN_IN), .B2(n19665), .A(n19664), .ZN(
        n19666) );
  AOI211_X1 U22587 ( .C1(n19675), .C2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n19678), .B(n19666), .ZN(n19672) );
  INV_X1 U22588 ( .A(n19667), .ZN(n19668) );
  NOR2_X1 U22589 ( .A1(n19669), .A2(n19668), .ZN(n19674) );
  AOI22_X1 U22590 ( .A1(n19670), .A2(n19699), .B1(n19674), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n19671) );
  OAI211_X1 U22591 ( .C1(n19673), .C2(n19690), .A(n19672), .B(n19671), .ZN(
        P1_U2835) );
  AOI22_X1 U22592 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19675), .B1(
        P1_REIP_REG_4__SCAN_IN), .B2(n19674), .ZN(n19676) );
  INV_X1 U22593 ( .A(n19676), .ZN(n19677) );
  AOI211_X1 U22594 ( .C1(n19687), .C2(P1_EBX_REG_4__SCAN_IN), .A(n19678), .B(
        n19677), .ZN(n19685) );
  OAI22_X1 U22595 ( .A1(n19681), .A2(n19799), .B1(n19680), .B2(n19679), .ZN(
        n19683) );
  NAND2_X1 U22596 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n19688) );
  NOR3_X1 U22597 ( .A1(n19696), .A2(P1_REIP_REG_4__SCAN_IN), .A3(n19688), .ZN(
        n19682) );
  AOI211_X1 U22598 ( .C1(n19786), .C2(n19699), .A(n19683), .B(n19682), .ZN(
        n19684) );
  OAI211_X1 U22599 ( .C1(n19792), .C2(n19690), .A(n19685), .B(n19684), .ZN(
        P1_U2836) );
  AOI22_X1 U22600 ( .A1(P1_EBX_REG_3__SCAN_IN), .A2(n19687), .B1(n19686), .B2(
        n19806), .ZN(n19702) );
  OAI21_X1 U22601 ( .B1(P1_REIP_REG_3__SCAN_IN), .B2(P1_REIP_REG_2__SCAN_IN), 
        .A(n19688), .ZN(n19697) );
  OAI22_X1 U22602 ( .A1(n19692), .A2(n19691), .B1(n19690), .B2(n19689), .ZN(
        n19693) );
  AOI21_X1 U22603 ( .B1(n19694), .B2(n20517), .A(n19693), .ZN(n19695) );
  OAI21_X1 U22604 ( .B1(n19697), .B2(n19696), .A(n19695), .ZN(n19698) );
  AOI21_X1 U22605 ( .B1(n19700), .B2(n19699), .A(n19698), .ZN(n19701) );
  OAI211_X1 U22606 ( .C1(n19703), .C2(n12998), .A(n19702), .B(n19701), .ZN(
        P1_U2837) );
  AOI22_X1 U22607 ( .A1(n19707), .A2(n19706), .B1(n19705), .B2(n19704), .ZN(
        n19708) );
  OAI21_X1 U22608 ( .B1(n19710), .B2(n19709), .A(n19708), .ZN(P1_U2866) );
  INV_X1 U22609 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n19749) );
  INV_X1 U22610 ( .A(n19846), .ZN(n19711) );
  OAI222_X1 U22611 ( .A1(n19715), .A2(n19714), .B1(n19749), .B2(n19713), .C1(
        n19712), .C2(n19711), .ZN(P1_U2904) );
  AOI22_X1 U22612 ( .A1(P1_LWORD_REG_15__SCAN_IN), .A2(n19746), .B1(n19745), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n19717) );
  OAI21_X1 U22613 ( .B1(n12646), .B2(n19748), .A(n19717), .ZN(P1_U2921) );
  INV_X1 U22614 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n19719) );
  AOI22_X1 U22615 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n19746), .B1(n19745), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n19718) );
  OAI21_X1 U22616 ( .B1(n19719), .B2(n19748), .A(n19718), .ZN(P1_U2922) );
  INV_X1 U22617 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n19721) );
  AOI22_X1 U22618 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n19746), .B1(n19745), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n19720) );
  OAI21_X1 U22619 ( .B1(n19721), .B2(n19748), .A(n19720), .ZN(P1_U2923) );
  INV_X1 U22620 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n19723) );
  AOI22_X1 U22621 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n19746), .B1(n19745), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n19722) );
  OAI21_X1 U22622 ( .B1(n19723), .B2(n19748), .A(n19722), .ZN(P1_U2924) );
  INV_X1 U22623 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n19725) );
  AOI22_X1 U22624 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n19746), .B1(n19745), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n19724) );
  OAI21_X1 U22625 ( .B1(n19725), .B2(n19748), .A(n19724), .ZN(P1_U2925) );
  INV_X1 U22626 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n19727) );
  AOI22_X1 U22627 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n19746), .B1(n19745), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n19726) );
  OAI21_X1 U22628 ( .B1(n19727), .B2(n19748), .A(n19726), .ZN(P1_U2926) );
  INV_X1 U22629 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n19729) );
  AOI22_X1 U22630 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n19736), .B1(n19745), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n19728) );
  OAI21_X1 U22631 ( .B1(n19729), .B2(n19748), .A(n19728), .ZN(P1_U2927) );
  INV_X1 U22632 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n19731) );
  AOI22_X1 U22633 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n19736), .B1(n19745), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n19730) );
  OAI21_X1 U22634 ( .B1(n19731), .B2(n19748), .A(n19730), .ZN(P1_U2928) );
  AOI22_X1 U22635 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n19736), .B1(n19745), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n19732) );
  OAI21_X1 U22636 ( .B1(n10647), .B2(n19748), .A(n19732), .ZN(P1_U2929) );
  AOI22_X1 U22637 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n19736), .B1(n19745), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n19733) );
  OAI21_X1 U22638 ( .B1(n19734), .B2(n19748), .A(n19733), .ZN(P1_U2930) );
  AOI22_X1 U22639 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n19736), .B1(n19745), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n19735) );
  OAI21_X1 U22640 ( .B1(n10616), .B2(n19748), .A(n19735), .ZN(P1_U2931) );
  AOI22_X1 U22641 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n19736), .B1(n19745), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n19737) );
  OAI21_X1 U22642 ( .B1(n19738), .B2(n19748), .A(n19737), .ZN(P1_U2932) );
  AOI22_X1 U22643 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n19746), .B1(n19745), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n19739) );
  OAI21_X1 U22644 ( .B1(n19740), .B2(n19748), .A(n19739), .ZN(P1_U2933) );
  AOI22_X1 U22645 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n19746), .B1(n19745), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n19741) );
  OAI21_X1 U22646 ( .B1(n19742), .B2(n19748), .A(n19741), .ZN(P1_U2934) );
  AOI22_X1 U22647 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n19746), .B1(n19745), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n19743) );
  OAI21_X1 U22648 ( .B1(n19744), .B2(n19748), .A(n19743), .ZN(P1_U2935) );
  AOI22_X1 U22649 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n19746), .B1(n19745), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n19747) );
  OAI21_X1 U22650 ( .B1(n19749), .B2(n19748), .A(n19747), .ZN(P1_U2936) );
  AOI22_X1 U22651 ( .A1(n19774), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n19773), .ZN(n19751) );
  NAND2_X1 U22652 ( .A1(n19763), .A2(n19750), .ZN(n19765) );
  NAND2_X1 U22653 ( .A1(n19751), .A2(n19765), .ZN(P1_U2945) );
  AOI22_X1 U22654 ( .A1(n19774), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n19773), .ZN(n19753) );
  NAND2_X1 U22655 ( .A1(n19763), .A2(n19752), .ZN(n19767) );
  NAND2_X1 U22656 ( .A1(n19753), .A2(n19767), .ZN(P1_U2946) );
  AOI22_X1 U22657 ( .A1(n19774), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n19773), .ZN(n19755) );
  NAND2_X1 U22658 ( .A1(n19763), .A2(n19754), .ZN(n19769) );
  NAND2_X1 U22659 ( .A1(n19755), .A2(n19769), .ZN(P1_U2947) );
  AOI22_X1 U22660 ( .A1(n19774), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n19773), .ZN(n19757) );
  NAND2_X1 U22661 ( .A1(n19763), .A2(n19756), .ZN(n19771) );
  NAND2_X1 U22662 ( .A1(n19757), .A2(n19771), .ZN(P1_U2948) );
  AOI22_X1 U22663 ( .A1(n19774), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n19773), .ZN(n19759) );
  NAND2_X1 U22664 ( .A1(n19763), .A2(n19758), .ZN(n19775) );
  NAND2_X1 U22665 ( .A1(n19759), .A2(n19775), .ZN(P1_U2949) );
  AOI22_X1 U22666 ( .A1(n19774), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n19773), .ZN(n19761) );
  NAND2_X1 U22667 ( .A1(n19763), .A2(n19760), .ZN(n19777) );
  NAND2_X1 U22668 ( .A1(n19761), .A2(n19777), .ZN(P1_U2950) );
  AOI22_X1 U22669 ( .A1(n19774), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n19773), .ZN(n19764) );
  NAND2_X1 U22670 ( .A1(n19763), .A2(n19762), .ZN(n19779) );
  NAND2_X1 U22671 ( .A1(n19764), .A2(n19779), .ZN(P1_U2951) );
  AOI22_X1 U22672 ( .A1(n19774), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n19773), .ZN(n19766) );
  NAND2_X1 U22673 ( .A1(n19766), .A2(n19765), .ZN(P1_U2960) );
  AOI22_X1 U22674 ( .A1(n19774), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n19773), .ZN(n19768) );
  NAND2_X1 U22675 ( .A1(n19768), .A2(n19767), .ZN(P1_U2961) );
  AOI22_X1 U22676 ( .A1(n19774), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n19773), .ZN(n19770) );
  NAND2_X1 U22677 ( .A1(n19770), .A2(n19769), .ZN(P1_U2962) );
  AOI22_X1 U22678 ( .A1(n19774), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n19773), .ZN(n19772) );
  NAND2_X1 U22679 ( .A1(n19772), .A2(n19771), .ZN(P1_U2963) );
  AOI22_X1 U22680 ( .A1(n19774), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n19773), .ZN(n19776) );
  NAND2_X1 U22681 ( .A1(n19776), .A2(n19775), .ZN(P1_U2964) );
  AOI22_X1 U22682 ( .A1(n19774), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n19773), .ZN(n19778) );
  NAND2_X1 U22683 ( .A1(n19778), .A2(n19777), .ZN(P1_U2965) );
  AOI22_X1 U22684 ( .A1(n19774), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n19773), .ZN(n19780) );
  NAND2_X1 U22685 ( .A1(n19780), .A2(n19779), .ZN(P1_U2966) );
  AOI22_X1 U22686 ( .A1(n19782), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n19781), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n19791) );
  OAI21_X1 U22687 ( .B1(n19785), .B2(n19784), .A(n19783), .ZN(n19797) );
  INV_X1 U22688 ( .A(n19797), .ZN(n19789) );
  AOI22_X1 U22689 ( .A1(n19789), .A2(n19788), .B1(n19787), .B2(n19786), .ZN(
        n19790) );
  OAI211_X1 U22690 ( .C1(n19793), .C2(n19792), .A(n19791), .B(n19790), .ZN(
        P1_U2995) );
  OAI22_X1 U22691 ( .A1(n19795), .A2(n19794), .B1(n19824), .B2(n19826), .ZN(
        n19796) );
  NOR2_X1 U22692 ( .A1(n19817), .A2(n19796), .ZN(n19815) );
  INV_X1 U22693 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20471) );
  OAI222_X1 U22694 ( .A1(n19799), .A2(n19823), .B1(n19798), .B2(n20471), .C1(
        n19820), .C2(n19797), .ZN(n19800) );
  INV_X1 U22695 ( .A(n19800), .ZN(n19803) );
  OAI211_X1 U22696 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n19809), .B(n19801), .ZN(n19802) );
  OAI211_X1 U22697 ( .C1(n19815), .C2(n19804), .A(n19803), .B(n19802), .ZN(
        P1_U3027) );
  AOI21_X1 U22698 ( .B1(n19807), .B2(n19806), .A(n19805), .ZN(n19813) );
  INV_X1 U22699 ( .A(n19808), .ZN(n19811) );
  AOI22_X1 U22700 ( .A1(n19811), .A2(n19810), .B1(n19809), .B2(n19814), .ZN(
        n19812) );
  OAI211_X1 U22701 ( .C1(n19815), .C2(n19814), .A(n19813), .B(n19812), .ZN(
        P1_U3028) );
  NAND2_X1 U22702 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n19816), .ZN(
        n19832) );
  AOI21_X1 U22703 ( .B1(n19819), .B2(n19818), .A(n19817), .ZN(n19830) );
  NOR2_X1 U22704 ( .A1(n19821), .A2(n19820), .ZN(n19829) );
  OAI22_X1 U22705 ( .A1(n19823), .A2(n19822), .B1(n13058), .B2(n19798), .ZN(
        n19828) );
  NAND2_X1 U22706 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19825) );
  AOI221_X1 U22707 ( .B1(n19831), .B2(n19826), .C1(n19825), .C2(n19826), .A(
        n19824), .ZN(n19827) );
  OAI221_X1 U22708 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n19832), .C1(
        n19831), .C2(n19830), .A(n9743), .ZN(P1_U3029) );
  NOR2_X1 U22709 ( .A1(n19833), .A2(n20526), .ZN(P1_U3032) );
  NOR2_X2 U22710 ( .A1(n19835), .A2(n19834), .ZN(n19883) );
  NOR2_X2 U22711 ( .A1(n19836), .A2(n19835), .ZN(n19884) );
  AOI22_X1 U22712 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19883), .B1(DATAI_24_), 
        .B2(n19884), .ZN(n20227) );
  NAND2_X1 U22713 ( .A1(n19839), .A2(n19885), .ZN(n20263) );
  NOR3_X1 U22714 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19900) );
  NAND2_X1 U22715 ( .A1(n20315), .A2(n19900), .ZN(n19887) );
  OAI22_X1 U22716 ( .A1(n20443), .A2(n20227), .B1(n20263), .B2(n19887), .ZN(
        n19840) );
  INV_X1 U22717 ( .A(n19840), .ZN(n19852) );
  INV_X1 U22718 ( .A(n20443), .ZN(n20423) );
  OAI21_X1 U22719 ( .B1(n19918), .B2(n20423), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n19841) );
  NAND2_X1 U22720 ( .A1(n19841), .A2(n20316), .ZN(n19850) );
  OR2_X1 U22721 ( .A1(n19842), .A2(n20517), .ZN(n19962) );
  NOR2_X1 U22722 ( .A1(n19962), .A2(n20349), .ZN(n19847) );
  INV_X1 U22723 ( .A(n19848), .ZN(n19843) );
  NOR2_X1 U22724 ( .A1(n19843), .A2(n20448), .ZN(n20261) );
  NOR2_X1 U22725 ( .A1(n19897), .A2(n20261), .ZN(n20180) );
  INV_X1 U22726 ( .A(n19844), .ZN(n20121) );
  NAND2_X1 U22727 ( .A1(n20121), .A2(n20178), .ZN(n19997) );
  AOI22_X1 U22728 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n19997), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n19887), .ZN(n19845) );
  OAI211_X1 U22729 ( .C1(n19850), .C2(n19847), .A(n20180), .B(n19845), .ZN(
        n19891) );
  NAND2_X1 U22730 ( .A1(n19846), .A2(n20000), .ZN(n20274) );
  INV_X1 U22731 ( .A(n19847), .ZN(n19849) );
  OR2_X1 U22732 ( .A1(n19848), .A2(n20448), .ZN(n20172) );
  AOI22_X1 U22733 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19891), .B1(
        n20386), .B2(n19890), .ZN(n19851) );
  OAI211_X1 U22734 ( .C1(n20395), .C2(n19915), .A(n19852), .B(n19851), .ZN(
        P1_U3033) );
  AOI22_X1 U22735 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19883), .B1(DATAI_25_), 
        .B2(n19884), .ZN(n20231) );
  NAND2_X1 U22736 ( .A1(n19853), .A2(n19885), .ZN(n20275) );
  OAI22_X1 U22737 ( .A1(n20443), .A2(n20231), .B1(n20275), .B2(n19887), .ZN(
        n19854) );
  INV_X1 U22738 ( .A(n19854), .ZN(n19857) );
  NAND2_X1 U22739 ( .A1(n19855), .A2(n20000), .ZN(n20279) );
  AOI22_X1 U22740 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19891), .B1(
        n20397), .B2(n19890), .ZN(n19856) );
  OAI211_X1 U22741 ( .C1(n20401), .C2(n19915), .A(n19857), .B(n19856), .ZN(
        P1_U3034) );
  AOI22_X1 U22742 ( .A1(DATAI_18_), .A2(n19884), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n19883), .ZN(n20363) );
  AOI22_X1 U22743 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19883), .B1(DATAI_26_), 
        .B2(n19884), .ZN(n20407) );
  NAND2_X1 U22744 ( .A1(n19858), .A2(n19885), .ZN(n20280) );
  OAI22_X1 U22745 ( .A1(n20443), .A2(n20407), .B1(n20280), .B2(n19887), .ZN(
        n19859) );
  INV_X1 U22746 ( .A(n19859), .ZN(n19862) );
  NAND2_X1 U22747 ( .A1(n19860), .A2(n20000), .ZN(n20284) );
  AOI22_X1 U22748 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19891), .B1(
        n20403), .B2(n19890), .ZN(n19861) );
  OAI211_X1 U22749 ( .C1(n20363), .C2(n19915), .A(n19862), .B(n19861), .ZN(
        P1_U3035) );
  AOI22_X1 U22750 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19883), .B1(DATAI_27_), 
        .B2(n19884), .ZN(n20237) );
  NAND2_X1 U22751 ( .A1(n19863), .A2(n19885), .ZN(n20285) );
  OAI22_X1 U22752 ( .A1(n20443), .A2(n20237), .B1(n20285), .B2(n19887), .ZN(
        n19864) );
  INV_X1 U22753 ( .A(n19864), .ZN(n19867) );
  NAND2_X1 U22754 ( .A1(n19865), .A2(n20000), .ZN(n20289) );
  AOI22_X1 U22755 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19891), .B1(
        n20409), .B2(n19890), .ZN(n19866) );
  OAI211_X1 U22756 ( .C1(n20413), .C2(n19915), .A(n19867), .B(n19866), .ZN(
        P1_U3036) );
  AOI22_X1 U22757 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19883), .B1(DATAI_28_), 
        .B2(n19884), .ZN(n20419) );
  NAND2_X1 U22758 ( .A1(n10396), .A2(n19885), .ZN(n20290) );
  OAI22_X1 U22759 ( .A1(n20443), .A2(n20419), .B1(n20290), .B2(n19887), .ZN(
        n19869) );
  INV_X1 U22760 ( .A(n19869), .ZN(n19872) );
  NAND2_X1 U22761 ( .A1(n19870), .A2(n20000), .ZN(n20294) );
  AOI22_X1 U22762 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19891), .B1(
        n20415), .B2(n19890), .ZN(n19871) );
  OAI211_X1 U22763 ( .C1(n20369), .C2(n19915), .A(n19872), .B(n19871), .ZN(
        P1_U3037) );
  AOI22_X1 U22764 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19883), .B1(DATAI_21_), 
        .B2(n19884), .ZN(n20373) );
  AOI22_X1 U22765 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19883), .B1(DATAI_29_), 
        .B2(n19884), .ZN(n20427) );
  NAND2_X1 U22766 ( .A1(n19873), .A2(n19885), .ZN(n20295) );
  OAI22_X1 U22767 ( .A1(n20443), .A2(n20427), .B1(n20295), .B2(n19887), .ZN(
        n19874) );
  INV_X1 U22768 ( .A(n19874), .ZN(n19877) );
  NAND2_X1 U22769 ( .A1(n19875), .A2(n20000), .ZN(n20299) );
  AOI22_X1 U22770 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19891), .B1(
        n20421), .B2(n19890), .ZN(n19876) );
  OAI211_X1 U22771 ( .C1(n20373), .C2(n19915), .A(n19877), .B(n19876), .ZN(
        P1_U3038) );
  AOI22_X1 U22772 ( .A1(DATAI_22_), .A2(n19884), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n19883), .ZN(n20433) );
  AOI22_X1 U22773 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19883), .B1(DATAI_30_), 
        .B2(n19884), .ZN(n20245) );
  NAND2_X1 U22774 ( .A1(n19878), .A2(n19885), .ZN(n20300) );
  OAI22_X1 U22775 ( .A1(n20443), .A2(n20245), .B1(n20300), .B2(n19887), .ZN(
        n19879) );
  INV_X1 U22776 ( .A(n19879), .ZN(n19882) );
  NAND2_X1 U22777 ( .A1(n19880), .A2(n20000), .ZN(n20304) );
  AOI22_X1 U22778 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19891), .B1(
        n20429), .B2(n19890), .ZN(n19881) );
  OAI211_X1 U22779 ( .C1(n20433), .C2(n19915), .A(n19882), .B(n19881), .ZN(
        P1_U3039) );
  AOI22_X1 U22780 ( .A1(DATAI_31_), .A2(n19884), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n19883), .ZN(n20253) );
  NAND2_X1 U22781 ( .A1(n19886), .A2(n19885), .ZN(n20306) );
  OAI22_X1 U22782 ( .A1(n20443), .A2(n20253), .B1(n20306), .B2(n19887), .ZN(
        n19888) );
  INV_X1 U22783 ( .A(n19888), .ZN(n19893) );
  NAND2_X1 U22784 ( .A1(n19889), .A2(n20000), .ZN(n20312) );
  AOI22_X1 U22785 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19891), .B1(
        n20436), .B2(n19890), .ZN(n19892) );
  OAI211_X1 U22786 ( .C1(n20444), .C2(n19915), .A(n19893), .B(n19892), .ZN(
        P1_U3040) );
  INV_X1 U22787 ( .A(n20314), .ZN(n19894) );
  INV_X1 U22788 ( .A(n19962), .ZN(n19895) );
  INV_X1 U22789 ( .A(n20317), .ZN(n20146) );
  INV_X1 U22790 ( .A(n19900), .ZN(n19896) );
  NOR2_X1 U22791 ( .A1(n20315), .A2(n19896), .ZN(n19916) );
  AOI21_X1 U22792 ( .B1(n19895), .B2(n20146), .A(n19916), .ZN(n19898) );
  OAI22_X1 U22793 ( .A1(n19898), .A2(n20516), .B1(n19896), .B2(n20448), .ZN(
        n19917) );
  AOI22_X1 U22794 ( .A1(n19917), .A2(n20386), .B1(n20385), .B2(n19916), .ZN(
        n19902) );
  AOI21_X1 U22795 ( .B1(n20315), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n19897), 
        .ZN(n20390) );
  INV_X1 U22796 ( .A(n19958), .ZN(n19964) );
  OR2_X1 U22797 ( .A1(n9631), .A2(n20347), .ZN(n20320) );
  OAI211_X1 U22798 ( .C1(n19964), .C2(n20320), .A(n20316), .B(n19898), .ZN(
        n19899) );
  OAI211_X1 U22799 ( .C1(n20316), .C2(n19900), .A(n20390), .B(n19899), .ZN(
        n19919) );
  INV_X1 U22800 ( .A(n20227), .ZN(n20392) );
  AOI22_X1 U22801 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19919), .B1(
        n19918), .B2(n20392), .ZN(n19901) );
  OAI211_X1 U22802 ( .C1(n20395), .C2(n19957), .A(n19902), .B(n19901), .ZN(
        P1_U3041) );
  AOI22_X1 U22803 ( .A1(n19917), .A2(n20397), .B1(n20396), .B2(n19916), .ZN(
        n19904) );
  INV_X1 U22804 ( .A(n19957), .ZN(n19925) );
  INV_X1 U22805 ( .A(n20401), .ZN(n20228) );
  AOI22_X1 U22806 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19919), .B1(
        n19925), .B2(n20228), .ZN(n19903) );
  OAI211_X1 U22807 ( .C1(n20231), .C2(n19915), .A(n19904), .B(n19903), .ZN(
        P1_U3042) );
  AOI22_X1 U22808 ( .A1(n19917), .A2(n20403), .B1(n20402), .B2(n19916), .ZN(
        n19906) );
  INV_X1 U22809 ( .A(n20407), .ZN(n20360) );
  AOI22_X1 U22810 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19919), .B1(
        n19918), .B2(n20360), .ZN(n19905) );
  OAI211_X1 U22811 ( .C1(n20363), .C2(n19957), .A(n19906), .B(n19905), .ZN(
        P1_U3043) );
  AOI22_X1 U22812 ( .A1(n19917), .A2(n20409), .B1(n20408), .B2(n19916), .ZN(
        n19908) );
  INV_X1 U22813 ( .A(n20237), .ZN(n20410) );
  AOI22_X1 U22814 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19919), .B1(
        n19918), .B2(n20410), .ZN(n19907) );
  OAI211_X1 U22815 ( .C1(n20413), .C2(n19957), .A(n19908), .B(n19907), .ZN(
        P1_U3044) );
  AOI22_X1 U22816 ( .A1(n19917), .A2(n20415), .B1(n20414), .B2(n19916), .ZN(
        n19910) );
  INV_X1 U22817 ( .A(n20419), .ZN(n20366) );
  AOI22_X1 U22818 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19919), .B1(
        n19918), .B2(n20366), .ZN(n19909) );
  OAI211_X1 U22819 ( .C1(n20369), .C2(n19957), .A(n19910), .B(n19909), .ZN(
        P1_U3045) );
  AOI22_X1 U22820 ( .A1(n19917), .A2(n20421), .B1(n20420), .B2(n19916), .ZN(
        n19912) );
  INV_X1 U22821 ( .A(n20427), .ZN(n20370) );
  AOI22_X1 U22822 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19919), .B1(
        n19918), .B2(n20370), .ZN(n19911) );
  OAI211_X1 U22823 ( .C1(n20373), .C2(n19957), .A(n19912), .B(n19911), .ZN(
        P1_U3046) );
  AOI22_X1 U22824 ( .A1(n19917), .A2(n20429), .B1(n20428), .B2(n19916), .ZN(
        n19914) );
  INV_X1 U22825 ( .A(n20433), .ZN(n20242) );
  AOI22_X1 U22826 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19919), .B1(
        n19925), .B2(n20242), .ZN(n19913) );
  OAI211_X1 U22827 ( .C1(n20245), .C2(n19915), .A(n19914), .B(n19913), .ZN(
        P1_U3047) );
  AOI22_X1 U22828 ( .A1(n19917), .A2(n20436), .B1(n20434), .B2(n19916), .ZN(
        n19921) );
  INV_X1 U22829 ( .A(n20253), .ZN(n20438) );
  AOI22_X1 U22830 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19919), .B1(
        n19918), .B2(n20438), .ZN(n19920) );
  OAI211_X1 U22831 ( .C1(n20444), .C2(n19957), .A(n19921), .B(n19920), .ZN(
        P1_U3048) );
  NOR3_X1 U22832 ( .A1(n19923), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19965) );
  NAND2_X1 U22833 ( .A1(n20315), .A2(n19965), .ZN(n19951) );
  OAI22_X1 U22834 ( .A1(n19957), .A2(n20227), .B1(n20263), .B2(n19951), .ZN(
        n19924) );
  INV_X1 U22835 ( .A(n19924), .ZN(n19932) );
  OAI21_X1 U22836 ( .B1(n19984), .B2(n19925), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n19926) );
  NAND2_X1 U22837 ( .A1(n19926), .A2(n20316), .ZN(n19930) );
  NOR2_X1 U22838 ( .A1(n19962), .A2(n12952), .ZN(n19928) );
  OR2_X1 U22839 ( .A1(n20178), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20055) );
  AND2_X1 U22840 ( .A1(n20055), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20051) );
  AOI21_X1 U22841 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n19951), .A(n20051), 
        .ZN(n19927) );
  OAI211_X1 U22842 ( .C1(n19930), .C2(n19928), .A(n20180), .B(n19927), .ZN(
        n19954) );
  INV_X1 U22843 ( .A(n19928), .ZN(n19929) );
  AOI22_X1 U22844 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19954), .B1(
        n20386), .B2(n19953), .ZN(n19931) );
  OAI211_X1 U22845 ( .C1(n20395), .C2(n19988), .A(n19932), .B(n19931), .ZN(
        P1_U3049) );
  OAI22_X1 U22846 ( .A1(n19988), .A2(n20401), .B1(n20275), .B2(n19951), .ZN(
        n19933) );
  INV_X1 U22847 ( .A(n19933), .ZN(n19935) );
  AOI22_X1 U22848 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19954), .B1(
        n20397), .B2(n19953), .ZN(n19934) );
  OAI211_X1 U22849 ( .C1(n20231), .C2(n19957), .A(n19935), .B(n19934), .ZN(
        P1_U3050) );
  OAI22_X1 U22850 ( .A1(n19988), .A2(n20363), .B1(n20280), .B2(n19951), .ZN(
        n19936) );
  INV_X1 U22851 ( .A(n19936), .ZN(n19938) );
  AOI22_X1 U22852 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19954), .B1(
        n20403), .B2(n19953), .ZN(n19937) );
  OAI211_X1 U22853 ( .C1(n20407), .C2(n19957), .A(n19938), .B(n19937), .ZN(
        P1_U3051) );
  OAI22_X1 U22854 ( .A1(n19988), .A2(n20413), .B1(n20285), .B2(n19951), .ZN(
        n19939) );
  INV_X1 U22855 ( .A(n19939), .ZN(n19941) );
  AOI22_X1 U22856 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19954), .B1(
        n20409), .B2(n19953), .ZN(n19940) );
  OAI211_X1 U22857 ( .C1(n20237), .C2(n19957), .A(n19941), .B(n19940), .ZN(
        P1_U3052) );
  OAI22_X1 U22858 ( .A1(n19957), .A2(n20419), .B1(n20290), .B2(n19951), .ZN(
        n19942) );
  INV_X1 U22859 ( .A(n19942), .ZN(n19944) );
  AOI22_X1 U22860 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19954), .B1(
        n20415), .B2(n19953), .ZN(n19943) );
  OAI211_X1 U22861 ( .C1(n20369), .C2(n19988), .A(n19944), .B(n19943), .ZN(
        P1_U3053) );
  OAI22_X1 U22862 ( .A1(n19988), .A2(n20373), .B1(n20295), .B2(n19951), .ZN(
        n19945) );
  INV_X1 U22863 ( .A(n19945), .ZN(n19947) );
  AOI22_X1 U22864 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19954), .B1(
        n20421), .B2(n19953), .ZN(n19946) );
  OAI211_X1 U22865 ( .C1(n20427), .C2(n19957), .A(n19947), .B(n19946), .ZN(
        P1_U3054) );
  OAI22_X1 U22866 ( .A1(n19957), .A2(n20245), .B1(n20300), .B2(n19951), .ZN(
        n19948) );
  INV_X1 U22867 ( .A(n19948), .ZN(n19950) );
  AOI22_X1 U22868 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19954), .B1(
        n20429), .B2(n19953), .ZN(n19949) );
  OAI211_X1 U22869 ( .C1(n20433), .C2(n19988), .A(n19950), .B(n19949), .ZN(
        P1_U3055) );
  OAI22_X1 U22870 ( .A1(n19988), .A2(n20444), .B1(n20306), .B2(n19951), .ZN(
        n19952) );
  INV_X1 U22871 ( .A(n19952), .ZN(n19956) );
  AOI22_X1 U22872 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19954), .B1(
        n20436), .B2(n19953), .ZN(n19955) );
  OAI211_X1 U22873 ( .C1(n20253), .C2(n19957), .A(n19956), .B(n19955), .ZN(
        P1_U3056) );
  OR2_X1 U22874 ( .A1(n19958), .A2(n20516), .ZN(n19959) );
  INV_X1 U22875 ( .A(n20216), .ZN(n20089) );
  INV_X1 U22876 ( .A(n19969), .ZN(n19963) );
  NAND2_X1 U22877 ( .A1(n19961), .A2(n19960), .ZN(n20383) );
  OR2_X1 U22878 ( .A1(n20211), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19987) );
  OAI21_X1 U22879 ( .B1(n19962), .B2(n20383), .A(n19987), .ZN(n19968) );
  INV_X1 U22880 ( .A(n20395), .ZN(n20224) );
  INV_X1 U22881 ( .A(n19987), .ZN(n19983) );
  AOI22_X1 U22882 ( .A1(n20018), .A2(n20224), .B1(n20385), .B2(n19983), .ZN(
        n19971) );
  INV_X1 U22883 ( .A(n19965), .ZN(n19966) );
  INV_X1 U22884 ( .A(n20390), .ZN(n20217) );
  AOI21_X1 U22885 ( .B1(n20516), .B2(n19966), .A(n20217), .ZN(n19967) );
  AOI22_X1 U22886 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19990), .B1(
        n19984), .B2(n20392), .ZN(n19970) );
  OAI211_X1 U22887 ( .C1(n19993), .C2(n20274), .A(n19971), .B(n19970), .ZN(
        P1_U3057) );
  AOI22_X1 U22888 ( .A1(n20018), .A2(n20228), .B1(n20396), .B2(n19983), .ZN(
        n19973) );
  INV_X1 U22889 ( .A(n20231), .ZN(n20398) );
  AOI22_X1 U22890 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19990), .B1(
        n19984), .B2(n20398), .ZN(n19972) );
  OAI211_X1 U22891 ( .C1(n19993), .C2(n20279), .A(n19973), .B(n19972), .ZN(
        P1_U3058) );
  INV_X1 U22892 ( .A(n20363), .ZN(n20404) );
  AOI22_X1 U22893 ( .A1(n20018), .A2(n20404), .B1(n20402), .B2(n19983), .ZN(
        n19975) );
  AOI22_X1 U22894 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19990), .B1(
        n19984), .B2(n20360), .ZN(n19974) );
  OAI211_X1 U22895 ( .C1(n19993), .C2(n20284), .A(n19975), .B(n19974), .ZN(
        P1_U3059) );
  INV_X1 U22896 ( .A(n20413), .ZN(n20234) );
  AOI22_X1 U22897 ( .A1(n20018), .A2(n20234), .B1(n20408), .B2(n19983), .ZN(
        n19977) );
  AOI22_X1 U22898 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19990), .B1(
        n19984), .B2(n20410), .ZN(n19976) );
  OAI211_X1 U22899 ( .C1(n19993), .C2(n20289), .A(n19977), .B(n19976), .ZN(
        P1_U3060) );
  INV_X1 U22900 ( .A(n20369), .ZN(n20416) );
  AOI22_X1 U22901 ( .A1(n20018), .A2(n20416), .B1(n20414), .B2(n19983), .ZN(
        n19979) );
  AOI22_X1 U22902 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19990), .B1(
        n19984), .B2(n20366), .ZN(n19978) );
  OAI211_X1 U22903 ( .C1(n19993), .C2(n20294), .A(n19979), .B(n19978), .ZN(
        P1_U3061) );
  OAI22_X1 U22904 ( .A1(n19988), .A2(n20427), .B1(n20295), .B2(n19987), .ZN(
        n19980) );
  INV_X1 U22905 ( .A(n19980), .ZN(n19982) );
  INV_X1 U22906 ( .A(n20373), .ZN(n20422) );
  AOI22_X1 U22907 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19990), .B1(
        n20018), .B2(n20422), .ZN(n19981) );
  OAI211_X1 U22908 ( .C1(n19993), .C2(n20299), .A(n19982), .B(n19981), .ZN(
        P1_U3062) );
  AOI22_X1 U22909 ( .A1(n20018), .A2(n20242), .B1(n20428), .B2(n19983), .ZN(
        n19986) );
  INV_X1 U22910 ( .A(n20245), .ZN(n20430) );
  AOI22_X1 U22911 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19990), .B1(
        n19984), .B2(n20430), .ZN(n19985) );
  OAI211_X1 U22912 ( .C1(n19993), .C2(n20304), .A(n19986), .B(n19985), .ZN(
        P1_U3063) );
  OAI22_X1 U22913 ( .A1(n19988), .A2(n20253), .B1(n20306), .B2(n19987), .ZN(
        n19989) );
  INV_X1 U22914 ( .A(n19989), .ZN(n19992) );
  INV_X1 U22915 ( .A(n20444), .ZN(n20248) );
  AOI22_X1 U22916 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19990), .B1(
        n20018), .B2(n20248), .ZN(n19991) );
  OAI211_X1 U22917 ( .C1(n19993), .C2(n20312), .A(n19992), .B(n19991), .ZN(
        P1_U3064) );
  INV_X1 U22918 ( .A(n20261), .ZN(n20345) );
  NOR2_X1 U22919 ( .A1(n20259), .A2(n19995), .ZN(n20087) );
  NAND3_X1 U22920 ( .A1(n20087), .A2(n20316), .A3(n12952), .ZN(n19996) );
  OAI21_X1 U22921 ( .B1(n20345), .B2(n19997), .A(n19996), .ZN(n20017) );
  NOR3_X1 U22922 ( .A1(n20262), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20025) );
  INV_X1 U22923 ( .A(n20025), .ZN(n20022) );
  NOR2_X1 U22924 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20022), .ZN(
        n20016) );
  AOI22_X1 U22925 ( .A1(n20017), .A2(n20386), .B1(n20385), .B2(n20016), .ZN(
        n20003) );
  INV_X1 U22926 ( .A(n20047), .ZN(n20034) );
  OAI21_X1 U22927 ( .B1(n20018), .B2(n20034), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n19999) );
  NAND2_X1 U22928 ( .A1(n20087), .A2(n12952), .ZN(n19998) );
  AOI21_X1 U22929 ( .B1(n19999), .B2(n19998), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20001) );
  AOI22_X1 U22930 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20019), .B1(
        n20018), .B2(n20392), .ZN(n20002) );
  OAI211_X1 U22931 ( .C1(n20395), .C2(n20047), .A(n20003), .B(n20002), .ZN(
        P1_U3065) );
  AOI22_X1 U22932 ( .A1(n20017), .A2(n20397), .B1(n20396), .B2(n20016), .ZN(
        n20005) );
  AOI22_X1 U22933 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20019), .B1(
        n20018), .B2(n20398), .ZN(n20004) );
  OAI211_X1 U22934 ( .C1(n20401), .C2(n20047), .A(n20005), .B(n20004), .ZN(
        P1_U3066) );
  AOI22_X1 U22935 ( .A1(n20017), .A2(n20403), .B1(n20402), .B2(n20016), .ZN(
        n20007) );
  AOI22_X1 U22936 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20019), .B1(
        n20018), .B2(n20360), .ZN(n20006) );
  OAI211_X1 U22937 ( .C1(n20363), .C2(n20047), .A(n20007), .B(n20006), .ZN(
        P1_U3067) );
  AOI22_X1 U22938 ( .A1(n20017), .A2(n20409), .B1(n20408), .B2(n20016), .ZN(
        n20009) );
  AOI22_X1 U22939 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20019), .B1(
        n20018), .B2(n20410), .ZN(n20008) );
  OAI211_X1 U22940 ( .C1(n20413), .C2(n20047), .A(n20009), .B(n20008), .ZN(
        P1_U3068) );
  AOI22_X1 U22941 ( .A1(n20017), .A2(n20415), .B1(n20414), .B2(n20016), .ZN(
        n20011) );
  AOI22_X1 U22942 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20019), .B1(
        n20018), .B2(n20366), .ZN(n20010) );
  OAI211_X1 U22943 ( .C1(n20369), .C2(n20047), .A(n20011), .B(n20010), .ZN(
        P1_U3069) );
  AOI22_X1 U22944 ( .A1(n20017), .A2(n20421), .B1(n20420), .B2(n20016), .ZN(
        n20013) );
  AOI22_X1 U22945 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20019), .B1(
        n20018), .B2(n20370), .ZN(n20012) );
  OAI211_X1 U22946 ( .C1(n20373), .C2(n20047), .A(n20013), .B(n20012), .ZN(
        P1_U3070) );
  AOI22_X1 U22947 ( .A1(n20017), .A2(n20429), .B1(n20428), .B2(n20016), .ZN(
        n20015) );
  AOI22_X1 U22948 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20019), .B1(
        n20018), .B2(n20430), .ZN(n20014) );
  OAI211_X1 U22949 ( .C1(n20433), .C2(n20047), .A(n20015), .B(n20014), .ZN(
        P1_U3071) );
  AOI22_X1 U22950 ( .A1(n20017), .A2(n20436), .B1(n20434), .B2(n20016), .ZN(
        n20021) );
  AOI22_X1 U22951 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20019), .B1(
        n20018), .B2(n20438), .ZN(n20020) );
  OAI211_X1 U22952 ( .C1(n20444), .C2(n20047), .A(n20021), .B(n20020), .ZN(
        P1_U3072) );
  NOR2_X1 U22953 ( .A1(n20315), .A2(n20022), .ZN(n20041) );
  AOI21_X1 U22954 ( .B1(n20087), .B2(n20146), .A(n20041), .ZN(n20023) );
  OAI22_X1 U22955 ( .A1(n20023), .A2(n20516), .B1(n20022), .B2(n20448), .ZN(
        n20042) );
  AOI22_X1 U22956 ( .A1(n20042), .A2(n20386), .B1(n20385), .B2(n20041), .ZN(
        n20027) );
  OAI211_X1 U22957 ( .C1(n20521), .C2(n20320), .A(n20316), .B(n20023), .ZN(
        n20024) );
  OAI211_X1 U22958 ( .C1(n20316), .C2(n20025), .A(n20390), .B(n20024), .ZN(
        n20044) );
  AOI22_X1 U22959 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20044), .B1(
        n20034), .B2(n20392), .ZN(n20026) );
  OAI211_X1 U22960 ( .C1(n20395), .C2(n20084), .A(n20027), .B(n20026), .ZN(
        P1_U3073) );
  AOI22_X1 U22961 ( .A1(n20042), .A2(n20397), .B1(n20396), .B2(n20041), .ZN(
        n20029) );
  AOI22_X1 U22962 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20044), .B1(
        n20034), .B2(n20398), .ZN(n20028) );
  OAI211_X1 U22963 ( .C1(n20401), .C2(n20084), .A(n20029), .B(n20028), .ZN(
        P1_U3074) );
  AOI22_X1 U22964 ( .A1(n20042), .A2(n20403), .B1(n20402), .B2(n20041), .ZN(
        n20031) );
  INV_X1 U22965 ( .A(n20084), .ZN(n20043) );
  AOI22_X1 U22966 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20044), .B1(
        n20043), .B2(n20404), .ZN(n20030) );
  OAI211_X1 U22967 ( .C1(n20407), .C2(n20047), .A(n20031), .B(n20030), .ZN(
        P1_U3075) );
  AOI22_X1 U22968 ( .A1(n20042), .A2(n20409), .B1(n20408), .B2(n20041), .ZN(
        n20033) );
  AOI22_X1 U22969 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20044), .B1(
        n20043), .B2(n20234), .ZN(n20032) );
  OAI211_X1 U22970 ( .C1(n20237), .C2(n20047), .A(n20033), .B(n20032), .ZN(
        P1_U3076) );
  AOI22_X1 U22971 ( .A1(n20042), .A2(n20415), .B1(n20414), .B2(n20041), .ZN(
        n20036) );
  AOI22_X1 U22972 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20044), .B1(
        n20034), .B2(n20366), .ZN(n20035) );
  OAI211_X1 U22973 ( .C1(n20369), .C2(n20084), .A(n20036), .B(n20035), .ZN(
        P1_U3077) );
  AOI22_X1 U22974 ( .A1(n20042), .A2(n20421), .B1(n20420), .B2(n20041), .ZN(
        n20038) );
  AOI22_X1 U22975 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20044), .B1(
        n20043), .B2(n20422), .ZN(n20037) );
  OAI211_X1 U22976 ( .C1(n20427), .C2(n20047), .A(n20038), .B(n20037), .ZN(
        P1_U3078) );
  AOI22_X1 U22977 ( .A1(n20042), .A2(n20429), .B1(n20428), .B2(n20041), .ZN(
        n20040) );
  AOI22_X1 U22978 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20044), .B1(
        n20043), .B2(n20242), .ZN(n20039) );
  OAI211_X1 U22979 ( .C1(n20245), .C2(n20047), .A(n20040), .B(n20039), .ZN(
        P1_U3079) );
  AOI22_X1 U22980 ( .A1(n20042), .A2(n20436), .B1(n20434), .B2(n20041), .ZN(
        n20046) );
  AOI22_X1 U22981 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20044), .B1(
        n20043), .B2(n20248), .ZN(n20045) );
  OAI211_X1 U22982 ( .C1(n20253), .C2(n20047), .A(n20046), .B(n20045), .ZN(
        P1_U3080) );
  INV_X1 U22983 ( .A(n20048), .ZN(n20343) );
  NOR2_X1 U22984 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20088), .ZN(
        n20053) );
  INV_X1 U22985 ( .A(n20053), .ZN(n20078) );
  OAI22_X1 U22986 ( .A1(n20084), .A2(n20227), .B1(n20263), .B2(n20078), .ZN(
        n20049) );
  INV_X1 U22987 ( .A(n20049), .ZN(n20059) );
  NAND2_X1 U22988 ( .A1(n20109), .A2(n20084), .ZN(n20050) );
  AOI21_X1 U22989 ( .B1(n20050), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20516), 
        .ZN(n20054) );
  NAND2_X1 U22990 ( .A1(n20087), .A2(n20349), .ZN(n20056) );
  AOI21_X1 U22991 ( .B1(n20054), .B2(n20056), .A(n20051), .ZN(n20052) );
  OAI211_X1 U22992 ( .C1(n20053), .C2(n20270), .A(n20353), .B(n20052), .ZN(
        n20081) );
  INV_X1 U22993 ( .A(n20054), .ZN(n20057) );
  OAI22_X1 U22994 ( .A1(n20057), .A2(n20056), .B1(n20055), .B2(n20345), .ZN(
        n20080) );
  AOI22_X1 U22995 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20081), .B1(
        n20386), .B2(n20080), .ZN(n20058) );
  OAI211_X1 U22996 ( .C1(n20395), .C2(n20109), .A(n20059), .B(n20058), .ZN(
        P1_U3081) );
  OAI22_X1 U22997 ( .A1(n20109), .A2(n20401), .B1(n20275), .B2(n20078), .ZN(
        n20060) );
  INV_X1 U22998 ( .A(n20060), .ZN(n20062) );
  AOI22_X1 U22999 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20081), .B1(
        n20397), .B2(n20080), .ZN(n20061) );
  OAI211_X1 U23000 ( .C1(n20231), .C2(n20084), .A(n20062), .B(n20061), .ZN(
        P1_U3082) );
  OAI22_X1 U23001 ( .A1(n20084), .A2(n20407), .B1(n20280), .B2(n20078), .ZN(
        n20063) );
  INV_X1 U23002 ( .A(n20063), .ZN(n20065) );
  AOI22_X1 U23003 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20081), .B1(
        n20403), .B2(n20080), .ZN(n20064) );
  OAI211_X1 U23004 ( .C1(n20363), .C2(n20109), .A(n20065), .B(n20064), .ZN(
        P1_U3083) );
  OAI22_X1 U23005 ( .A1(n20084), .A2(n20237), .B1(n20285), .B2(n20078), .ZN(
        n20066) );
  INV_X1 U23006 ( .A(n20066), .ZN(n20068) );
  AOI22_X1 U23007 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20081), .B1(
        n20409), .B2(n20080), .ZN(n20067) );
  OAI211_X1 U23008 ( .C1(n20413), .C2(n20109), .A(n20068), .B(n20067), .ZN(
        P1_U3084) );
  OAI22_X1 U23009 ( .A1(n20109), .A2(n20369), .B1(n20290), .B2(n20078), .ZN(
        n20069) );
  INV_X1 U23010 ( .A(n20069), .ZN(n20071) );
  AOI22_X1 U23011 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20081), .B1(
        n20415), .B2(n20080), .ZN(n20070) );
  OAI211_X1 U23012 ( .C1(n20419), .C2(n20084), .A(n20071), .B(n20070), .ZN(
        P1_U3085) );
  OAI22_X1 U23013 ( .A1(n20109), .A2(n20373), .B1(n20295), .B2(n20078), .ZN(
        n20072) );
  INV_X1 U23014 ( .A(n20072), .ZN(n20074) );
  AOI22_X1 U23015 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20081), .B1(
        n20421), .B2(n20080), .ZN(n20073) );
  OAI211_X1 U23016 ( .C1(n20427), .C2(n20084), .A(n20074), .B(n20073), .ZN(
        P1_U3086) );
  OAI22_X1 U23017 ( .A1(n20109), .A2(n20433), .B1(n20300), .B2(n20078), .ZN(
        n20075) );
  INV_X1 U23018 ( .A(n20075), .ZN(n20077) );
  AOI22_X1 U23019 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20081), .B1(
        n20429), .B2(n20080), .ZN(n20076) );
  OAI211_X1 U23020 ( .C1(n20245), .C2(n20084), .A(n20077), .B(n20076), .ZN(
        P1_U3087) );
  OAI22_X1 U23021 ( .A1(n20109), .A2(n20444), .B1(n20306), .B2(n20078), .ZN(
        n20079) );
  INV_X1 U23022 ( .A(n20079), .ZN(n20083) );
  AOI22_X1 U23023 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20081), .B1(
        n20436), .B2(n20080), .ZN(n20082) );
  OAI211_X1 U23024 ( .C1(n20253), .C2(n20084), .A(n20083), .B(n20082), .ZN(
        P1_U3088) );
  INV_X1 U23025 ( .A(n20383), .ZN(n20086) );
  INV_X1 U23026 ( .A(n20085), .ZN(n20110) );
  AOI21_X1 U23027 ( .B1(n20087), .B2(n20086), .A(n20110), .ZN(n20091) );
  OAI22_X1 U23028 ( .A1(n20091), .A2(n20516), .B1(n20088), .B2(n20448), .ZN(
        n20111) );
  AOI22_X1 U23029 ( .A1(n20111), .A2(n20386), .B1(n20110), .B2(n20385), .ZN(
        n20096) );
  INV_X1 U23030 ( .A(n20521), .ZN(n20090) );
  OAI21_X1 U23031 ( .B1(n20090), .B2(n20516), .A(n20089), .ZN(n20092) );
  NAND2_X1 U23032 ( .A1(n20092), .A2(n20091), .ZN(n20093) );
  OAI211_X1 U23033 ( .C1(n20094), .C2(n20316), .A(n20390), .B(n20093), .ZN(
        n20113) );
  INV_X1 U23034 ( .A(n20109), .ZN(n20112) );
  AOI22_X1 U23035 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20113), .B1(
        n20112), .B2(n20392), .ZN(n20095) );
  OAI211_X1 U23036 ( .C1(n20395), .C2(n20116), .A(n20096), .B(n20095), .ZN(
        P1_U3089) );
  AOI22_X1 U23037 ( .A1(n20111), .A2(n20397), .B1(n20110), .B2(n20396), .ZN(
        n20098) );
  AOI22_X1 U23038 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20113), .B1(
        n20142), .B2(n20228), .ZN(n20097) );
  OAI211_X1 U23039 ( .C1(n20231), .C2(n20109), .A(n20098), .B(n20097), .ZN(
        P1_U3090) );
  AOI22_X1 U23040 ( .A1(n20111), .A2(n20403), .B1(n20110), .B2(n20402), .ZN(
        n20100) );
  AOI22_X1 U23041 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20113), .B1(
        n20142), .B2(n20404), .ZN(n20099) );
  OAI211_X1 U23042 ( .C1(n20407), .C2(n20109), .A(n20100), .B(n20099), .ZN(
        P1_U3091) );
  AOI22_X1 U23043 ( .A1(n20111), .A2(n20409), .B1(n20110), .B2(n20408), .ZN(
        n20102) );
  AOI22_X1 U23044 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20113), .B1(
        n20112), .B2(n20410), .ZN(n20101) );
  OAI211_X1 U23045 ( .C1(n20413), .C2(n20116), .A(n20102), .B(n20101), .ZN(
        P1_U3092) );
  AOI22_X1 U23046 ( .A1(n20111), .A2(n20415), .B1(n20110), .B2(n20414), .ZN(
        n20104) );
  AOI22_X1 U23047 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20113), .B1(
        n20112), .B2(n20366), .ZN(n20103) );
  OAI211_X1 U23048 ( .C1(n20369), .C2(n20116), .A(n20104), .B(n20103), .ZN(
        P1_U3093) );
  AOI22_X1 U23049 ( .A1(n20111), .A2(n20421), .B1(n20110), .B2(n20420), .ZN(
        n20106) );
  AOI22_X1 U23050 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20113), .B1(
        n20112), .B2(n20370), .ZN(n20105) );
  OAI211_X1 U23051 ( .C1(n20373), .C2(n20116), .A(n20106), .B(n20105), .ZN(
        P1_U3094) );
  AOI22_X1 U23052 ( .A1(n20111), .A2(n20429), .B1(n20110), .B2(n20428), .ZN(
        n20108) );
  AOI22_X1 U23053 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20113), .B1(
        n20142), .B2(n20242), .ZN(n20107) );
  OAI211_X1 U23054 ( .C1(n20245), .C2(n20109), .A(n20108), .B(n20107), .ZN(
        P1_U3095) );
  AOI22_X1 U23055 ( .A1(n20111), .A2(n20436), .B1(n20110), .B2(n20434), .ZN(
        n20115) );
  AOI22_X1 U23056 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20113), .B1(
        n20112), .B2(n20438), .ZN(n20114) );
  OAI211_X1 U23057 ( .C1(n20444), .C2(n20116), .A(n20115), .B(n20114), .ZN(
        P1_U3096) );
  INV_X1 U23058 ( .A(n20223), .ZN(n20119) );
  AND2_X1 U23059 ( .A1(n20517), .A2(n20259), .ZN(n20210) );
  NOR3_X1 U23060 ( .A1(n20528), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20150) );
  INV_X1 U23061 ( .A(n20150), .ZN(n20147) );
  NOR2_X1 U23062 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20147), .ZN(
        n20140) );
  AOI21_X1 U23063 ( .B1(n20210), .B2(n12952), .A(n20140), .ZN(n20123) );
  INV_X1 U23064 ( .A(n20178), .ZN(n20120) );
  NOR2_X1 U23065 ( .A1(n20121), .A2(n20120), .ZN(n20260) );
  INV_X1 U23066 ( .A(n20260), .ZN(n20266) );
  OAI22_X1 U23067 ( .A1(n20123), .A2(n20516), .B1(n20172), .B2(n20266), .ZN(
        n20141) );
  AOI22_X1 U23068 ( .A1(n20141), .A2(n20386), .B1(n20385), .B2(n20140), .ZN(
        n20127) );
  INV_X1 U23069 ( .A(n20170), .ZN(n20122) );
  OAI21_X1 U23070 ( .B1(n20122), .B2(n20142), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20124) );
  NAND2_X1 U23071 ( .A1(n20124), .A2(n20123), .ZN(n20125) );
  AOI22_X1 U23072 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20143), .B1(
        n20142), .B2(n20392), .ZN(n20126) );
  OAI211_X1 U23073 ( .C1(n20395), .C2(n20170), .A(n20127), .B(n20126), .ZN(
        P1_U3097) );
  AOI22_X1 U23074 ( .A1(n20141), .A2(n20397), .B1(n20396), .B2(n20140), .ZN(
        n20129) );
  AOI22_X1 U23075 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20143), .B1(
        n20142), .B2(n20398), .ZN(n20128) );
  OAI211_X1 U23076 ( .C1(n20401), .C2(n20170), .A(n20129), .B(n20128), .ZN(
        P1_U3098) );
  AOI22_X1 U23077 ( .A1(n20141), .A2(n20403), .B1(n20402), .B2(n20140), .ZN(
        n20131) );
  AOI22_X1 U23078 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20143), .B1(
        n20142), .B2(n20360), .ZN(n20130) );
  OAI211_X1 U23079 ( .C1(n20363), .C2(n20170), .A(n20131), .B(n20130), .ZN(
        P1_U3099) );
  AOI22_X1 U23080 ( .A1(n20141), .A2(n20409), .B1(n20408), .B2(n20140), .ZN(
        n20133) );
  AOI22_X1 U23081 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20143), .B1(
        n20142), .B2(n20410), .ZN(n20132) );
  OAI211_X1 U23082 ( .C1(n20413), .C2(n20170), .A(n20133), .B(n20132), .ZN(
        P1_U3100) );
  AOI22_X1 U23083 ( .A1(n20141), .A2(n20415), .B1(n20414), .B2(n20140), .ZN(
        n20135) );
  AOI22_X1 U23084 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20143), .B1(
        n20142), .B2(n20366), .ZN(n20134) );
  OAI211_X1 U23085 ( .C1(n20369), .C2(n20170), .A(n20135), .B(n20134), .ZN(
        P1_U3101) );
  AOI22_X1 U23086 ( .A1(n20141), .A2(n20421), .B1(n20420), .B2(n20140), .ZN(
        n20137) );
  AOI22_X1 U23087 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20143), .B1(
        n20142), .B2(n20370), .ZN(n20136) );
  OAI211_X1 U23088 ( .C1(n20373), .C2(n20170), .A(n20137), .B(n20136), .ZN(
        P1_U3102) );
  AOI22_X1 U23089 ( .A1(n20141), .A2(n20429), .B1(n20428), .B2(n20140), .ZN(
        n20139) );
  AOI22_X1 U23090 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20143), .B1(
        n20142), .B2(n20430), .ZN(n20138) );
  OAI211_X1 U23091 ( .C1(n20433), .C2(n20170), .A(n20139), .B(n20138), .ZN(
        P1_U3103) );
  AOI22_X1 U23092 ( .A1(n20141), .A2(n20436), .B1(n20434), .B2(n20140), .ZN(
        n20145) );
  AOI22_X1 U23093 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20143), .B1(
        n20142), .B2(n20438), .ZN(n20144) );
  OAI211_X1 U23094 ( .C1(n20444), .C2(n20170), .A(n20145), .B(n20144), .ZN(
        P1_U3104) );
  NOR2_X1 U23095 ( .A1(n20315), .A2(n20147), .ZN(n20165) );
  AOI21_X1 U23096 ( .B1(n20210), .B2(n20146), .A(n20165), .ZN(n20148) );
  OAI22_X1 U23097 ( .A1(n20148), .A2(n20516), .B1(n20147), .B2(n20448), .ZN(
        n20166) );
  AOI22_X1 U23098 ( .A1(n20166), .A2(n20386), .B1(n20385), .B2(n20165), .ZN(
        n20152) );
  OAI211_X1 U23099 ( .C1(n20223), .C2(n20320), .A(n20316), .B(n20148), .ZN(
        n20149) );
  OAI211_X1 U23100 ( .C1(n20316), .C2(n20150), .A(n20390), .B(n20149), .ZN(
        n20167) );
  AOI22_X1 U23101 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20167), .B1(
        n20205), .B2(n20224), .ZN(n20151) );
  OAI211_X1 U23102 ( .C1(n20227), .C2(n20170), .A(n20152), .B(n20151), .ZN(
        P1_U3105) );
  AOI22_X1 U23103 ( .A1(n20166), .A2(n20397), .B1(n20396), .B2(n20165), .ZN(
        n20154) );
  AOI22_X1 U23104 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20167), .B1(
        n20205), .B2(n20228), .ZN(n20153) );
  OAI211_X1 U23105 ( .C1(n20231), .C2(n20170), .A(n20154), .B(n20153), .ZN(
        P1_U3106) );
  AOI22_X1 U23106 ( .A1(n20166), .A2(n20403), .B1(n20402), .B2(n20165), .ZN(
        n20156) );
  AOI22_X1 U23107 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20167), .B1(
        n20205), .B2(n20404), .ZN(n20155) );
  OAI211_X1 U23108 ( .C1(n20407), .C2(n20170), .A(n20156), .B(n20155), .ZN(
        P1_U3107) );
  AOI22_X1 U23109 ( .A1(n20166), .A2(n20409), .B1(n20408), .B2(n20165), .ZN(
        n20158) );
  AOI22_X1 U23110 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20167), .B1(
        n20205), .B2(n20234), .ZN(n20157) );
  OAI211_X1 U23111 ( .C1(n20237), .C2(n20170), .A(n20158), .B(n20157), .ZN(
        P1_U3108) );
  AOI22_X1 U23112 ( .A1(n20166), .A2(n20415), .B1(n20414), .B2(n20165), .ZN(
        n20160) );
  AOI22_X1 U23113 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20167), .B1(
        n20205), .B2(n20416), .ZN(n20159) );
  OAI211_X1 U23114 ( .C1(n20419), .C2(n20170), .A(n20160), .B(n20159), .ZN(
        P1_U3109) );
  AOI22_X1 U23115 ( .A1(n20166), .A2(n20421), .B1(n20420), .B2(n20165), .ZN(
        n20162) );
  AOI22_X1 U23116 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20167), .B1(
        n20205), .B2(n20422), .ZN(n20161) );
  OAI211_X1 U23117 ( .C1(n20427), .C2(n20170), .A(n20162), .B(n20161), .ZN(
        P1_U3110) );
  AOI22_X1 U23118 ( .A1(n20166), .A2(n20429), .B1(n20428), .B2(n20165), .ZN(
        n20164) );
  AOI22_X1 U23119 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20167), .B1(
        n20205), .B2(n20242), .ZN(n20163) );
  OAI211_X1 U23120 ( .C1(n20245), .C2(n20170), .A(n20164), .B(n20163), .ZN(
        P1_U3111) );
  AOI22_X1 U23121 ( .A1(n20166), .A2(n20436), .B1(n20434), .B2(n20165), .ZN(
        n20169) );
  AOI22_X1 U23122 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20167), .B1(
        n20205), .B2(n20248), .ZN(n20168) );
  OAI211_X1 U23123 ( .C1(n20253), .C2(n20170), .A(n20169), .B(n20168), .ZN(
        P1_U3112) );
  NAND3_X1 U23124 ( .A1(n20252), .A2(n20198), .A3(n20316), .ZN(n20171) );
  NAND2_X1 U23125 ( .A1(n20171), .A2(n20256), .ZN(n20177) );
  AND2_X1 U23126 ( .A1(n20210), .A2(n20349), .ZN(n20175) );
  NOR2_X1 U23127 ( .A1(n20178), .A2(n20528), .ZN(n20344) );
  INV_X1 U23128 ( .A(n20172), .ZN(n20173) );
  NAND3_X1 U23129 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n20262), .ZN(n20218) );
  OR2_X1 U23130 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20218), .ZN(
        n20203) );
  OAI22_X1 U23131 ( .A1(n20252), .A2(n20395), .B1(n20203), .B2(n20263), .ZN(
        n20174) );
  INV_X1 U23132 ( .A(n20174), .ZN(n20182) );
  INV_X1 U23133 ( .A(n20175), .ZN(n20176) );
  AOI22_X1 U23134 ( .A1(n20177), .A2(n20176), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20203), .ZN(n20179) );
  OAI21_X1 U23135 ( .B1(n20528), .B2(n20178), .A(P1_STATE2_REG_2__SCAN_IN), 
        .ZN(n20352) );
  NAND3_X1 U23136 ( .A1(n20180), .A2(n20179), .A3(n20352), .ZN(n20206) );
  AOI22_X1 U23137 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20206), .B1(
        n20205), .B2(n20392), .ZN(n20181) );
  OAI211_X1 U23138 ( .C1(n20209), .C2(n20274), .A(n20182), .B(n20181), .ZN(
        P1_U3113) );
  OAI22_X1 U23139 ( .A1(n20252), .A2(n20401), .B1(n20203), .B2(n20275), .ZN(
        n20183) );
  INV_X1 U23140 ( .A(n20183), .ZN(n20185) );
  AOI22_X1 U23141 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20206), .B1(
        n20205), .B2(n20398), .ZN(n20184) );
  OAI211_X1 U23142 ( .C1(n20209), .C2(n20279), .A(n20185), .B(n20184), .ZN(
        P1_U3114) );
  OAI22_X1 U23143 ( .A1(n20252), .A2(n20363), .B1(n20203), .B2(n20280), .ZN(
        n20186) );
  INV_X1 U23144 ( .A(n20186), .ZN(n20188) );
  AOI22_X1 U23145 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20206), .B1(
        n20205), .B2(n20360), .ZN(n20187) );
  OAI211_X1 U23146 ( .C1(n20209), .C2(n20284), .A(n20188), .B(n20187), .ZN(
        P1_U3115) );
  OAI22_X1 U23147 ( .A1(n20198), .A2(n20237), .B1(n20285), .B2(n20203), .ZN(
        n20189) );
  INV_X1 U23148 ( .A(n20189), .ZN(n20191) );
  INV_X1 U23149 ( .A(n20252), .ZN(n20200) );
  AOI22_X1 U23150 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20206), .B1(
        n20200), .B2(n20234), .ZN(n20190) );
  OAI211_X1 U23151 ( .C1(n20209), .C2(n20289), .A(n20191), .B(n20190), .ZN(
        P1_U3116) );
  OAI22_X1 U23152 ( .A1(n20252), .A2(n20369), .B1(n20203), .B2(n20290), .ZN(
        n20192) );
  INV_X1 U23153 ( .A(n20192), .ZN(n20194) );
  AOI22_X1 U23154 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20206), .B1(
        n20205), .B2(n20366), .ZN(n20193) );
  OAI211_X1 U23155 ( .C1(n20209), .C2(n20294), .A(n20194), .B(n20193), .ZN(
        P1_U3117) );
  OAI22_X1 U23156 ( .A1(n20198), .A2(n20427), .B1(n20203), .B2(n20295), .ZN(
        n20195) );
  INV_X1 U23157 ( .A(n20195), .ZN(n20197) );
  AOI22_X1 U23158 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20206), .B1(
        n20200), .B2(n20422), .ZN(n20196) );
  OAI211_X1 U23159 ( .C1(n20209), .C2(n20299), .A(n20197), .B(n20196), .ZN(
        P1_U3118) );
  OAI22_X1 U23160 ( .A1(n20198), .A2(n20245), .B1(n20203), .B2(n20300), .ZN(
        n20199) );
  INV_X1 U23161 ( .A(n20199), .ZN(n20202) );
  AOI22_X1 U23162 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20206), .B1(
        n20200), .B2(n20242), .ZN(n20201) );
  OAI211_X1 U23163 ( .C1(n20209), .C2(n20304), .A(n20202), .B(n20201), .ZN(
        P1_U3119) );
  OAI22_X1 U23164 ( .A1(n20252), .A2(n20444), .B1(n20203), .B2(n20306), .ZN(
        n20204) );
  INV_X1 U23165 ( .A(n20204), .ZN(n20208) );
  AOI22_X1 U23166 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20206), .B1(
        n20205), .B2(n20438), .ZN(n20207) );
  OAI211_X1 U23167 ( .C1(n20209), .C2(n20312), .A(n20208), .B(n20207), .ZN(
        P1_U3120) );
  INV_X1 U23168 ( .A(n20210), .ZN(n20213) );
  INV_X1 U23169 ( .A(n20211), .ZN(n20212) );
  NAND2_X1 U23170 ( .A1(n20212), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20215) );
  OAI21_X1 U23171 ( .B1(n20213), .B2(n20383), .A(n20215), .ZN(n20220) );
  INV_X1 U23172 ( .A(n20220), .ZN(n20214) );
  OAI22_X1 U23173 ( .A1(n20214), .A2(n20516), .B1(n20218), .B2(n20448), .ZN(
        n20247) );
  INV_X1 U23174 ( .A(n20215), .ZN(n20246) );
  AOI22_X1 U23175 ( .A1(n20247), .A2(n20386), .B1(n20246), .B2(n20385), .ZN(
        n20226) );
  AOI21_X1 U23176 ( .B1(n20223), .B2(n20316), .A(n20216), .ZN(n20221) );
  AOI21_X1 U23177 ( .B1(n20218), .B2(n20516), .A(n20217), .ZN(n20219) );
  OAI21_X1 U23178 ( .B1(n20221), .B2(n20220), .A(n20219), .ZN(n20249) );
  AOI22_X1 U23179 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20249), .B1(
        n20308), .B2(n20224), .ZN(n20225) );
  OAI211_X1 U23180 ( .C1(n20227), .C2(n20252), .A(n20226), .B(n20225), .ZN(
        P1_U3121) );
  AOI22_X1 U23181 ( .A1(n20247), .A2(n20397), .B1(n20246), .B2(n20396), .ZN(
        n20230) );
  AOI22_X1 U23182 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20249), .B1(
        n20308), .B2(n20228), .ZN(n20229) );
  OAI211_X1 U23183 ( .C1(n20231), .C2(n20252), .A(n20230), .B(n20229), .ZN(
        P1_U3122) );
  AOI22_X1 U23184 ( .A1(n20247), .A2(n20403), .B1(n20246), .B2(n20402), .ZN(
        n20233) );
  AOI22_X1 U23185 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20249), .B1(
        n20308), .B2(n20404), .ZN(n20232) );
  OAI211_X1 U23186 ( .C1(n20407), .C2(n20252), .A(n20233), .B(n20232), .ZN(
        P1_U3123) );
  AOI22_X1 U23187 ( .A1(n20247), .A2(n20409), .B1(n20246), .B2(n20408), .ZN(
        n20236) );
  AOI22_X1 U23188 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20249), .B1(
        n20308), .B2(n20234), .ZN(n20235) );
  OAI211_X1 U23189 ( .C1(n20237), .C2(n20252), .A(n20236), .B(n20235), .ZN(
        P1_U3124) );
  AOI22_X1 U23190 ( .A1(n20247), .A2(n20415), .B1(n20246), .B2(n20414), .ZN(
        n20239) );
  AOI22_X1 U23191 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20249), .B1(
        n20308), .B2(n20416), .ZN(n20238) );
  OAI211_X1 U23192 ( .C1(n20419), .C2(n20252), .A(n20239), .B(n20238), .ZN(
        P1_U3125) );
  AOI22_X1 U23193 ( .A1(n20247), .A2(n20421), .B1(n20246), .B2(n20420), .ZN(
        n20241) );
  AOI22_X1 U23194 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20249), .B1(
        n20308), .B2(n20422), .ZN(n20240) );
  OAI211_X1 U23195 ( .C1(n20427), .C2(n20252), .A(n20241), .B(n20240), .ZN(
        P1_U3126) );
  AOI22_X1 U23196 ( .A1(n20247), .A2(n20429), .B1(n20246), .B2(n20428), .ZN(
        n20244) );
  AOI22_X1 U23197 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20249), .B1(
        n20308), .B2(n20242), .ZN(n20243) );
  OAI211_X1 U23198 ( .C1(n20245), .C2(n20252), .A(n20244), .B(n20243), .ZN(
        P1_U3127) );
  AOI22_X1 U23199 ( .A1(n20247), .A2(n20436), .B1(n20246), .B2(n20434), .ZN(
        n20251) );
  AOI22_X1 U23200 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20249), .B1(
        n20308), .B2(n20248), .ZN(n20250) );
  OAI211_X1 U23201 ( .C1(n20253), .C2(n20252), .A(n20251), .B(n20250), .ZN(
        P1_U3128) );
  NAND3_X1 U23202 ( .A1(n20255), .A2(n20316), .A3(n20322), .ZN(n20257) );
  NAND2_X1 U23203 ( .A1(n20257), .A2(n20256), .ZN(n20268) );
  NOR2_X1 U23204 ( .A1(n20259), .A2(n20258), .ZN(n20350) );
  AND2_X1 U23205 ( .A1(n20350), .A2(n12952), .ZN(n20265) );
  NOR3_X1 U23206 ( .A1(n20262), .A2(n20528), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20321) );
  INV_X1 U23207 ( .A(n20321), .ZN(n20318) );
  NOR2_X1 U23208 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20318), .ZN(
        n20271) );
  INV_X1 U23209 ( .A(n20271), .ZN(n20305) );
  OAI22_X1 U23210 ( .A1(n20322), .A2(n20395), .B1(n20263), .B2(n20305), .ZN(
        n20264) );
  INV_X1 U23211 ( .A(n20264), .ZN(n20273) );
  INV_X1 U23212 ( .A(n20265), .ZN(n20267) );
  AOI22_X1 U23213 ( .A1(n20268), .A2(n20267), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20266), .ZN(n20269) );
  OAI211_X1 U23214 ( .C1(n20271), .C2(n20270), .A(n20353), .B(n20269), .ZN(
        n20309) );
  AOI22_X1 U23215 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20309), .B1(
        n20308), .B2(n20392), .ZN(n20272) );
  OAI211_X1 U23216 ( .C1(n20313), .C2(n20274), .A(n20273), .B(n20272), .ZN(
        P1_U3129) );
  OAI22_X1 U23217 ( .A1(n20322), .A2(n20401), .B1(n20275), .B2(n20305), .ZN(
        n20276) );
  INV_X1 U23218 ( .A(n20276), .ZN(n20278) );
  AOI22_X1 U23219 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20309), .B1(
        n20308), .B2(n20398), .ZN(n20277) );
  OAI211_X1 U23220 ( .C1(n20313), .C2(n20279), .A(n20278), .B(n20277), .ZN(
        P1_U3130) );
  OAI22_X1 U23221 ( .A1(n20322), .A2(n20363), .B1(n20280), .B2(n20305), .ZN(
        n20281) );
  INV_X1 U23222 ( .A(n20281), .ZN(n20283) );
  AOI22_X1 U23223 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20309), .B1(
        n20308), .B2(n20360), .ZN(n20282) );
  OAI211_X1 U23224 ( .C1(n20313), .C2(n20284), .A(n20283), .B(n20282), .ZN(
        P1_U3131) );
  OAI22_X1 U23225 ( .A1(n20322), .A2(n20413), .B1(n20285), .B2(n20305), .ZN(
        n20286) );
  INV_X1 U23226 ( .A(n20286), .ZN(n20288) );
  AOI22_X1 U23227 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20309), .B1(
        n20308), .B2(n20410), .ZN(n20287) );
  OAI211_X1 U23228 ( .C1(n20313), .C2(n20289), .A(n20288), .B(n20287), .ZN(
        P1_U3132) );
  OAI22_X1 U23229 ( .A1(n20322), .A2(n20369), .B1(n20290), .B2(n20305), .ZN(
        n20291) );
  INV_X1 U23230 ( .A(n20291), .ZN(n20293) );
  AOI22_X1 U23231 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20309), .B1(
        n20308), .B2(n20366), .ZN(n20292) );
  OAI211_X1 U23232 ( .C1(n20313), .C2(n20294), .A(n20293), .B(n20292), .ZN(
        P1_U3133) );
  OAI22_X1 U23233 ( .A1(n20322), .A2(n20373), .B1(n20295), .B2(n20305), .ZN(
        n20296) );
  INV_X1 U23234 ( .A(n20296), .ZN(n20298) );
  AOI22_X1 U23235 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20309), .B1(
        n20308), .B2(n20370), .ZN(n20297) );
  OAI211_X1 U23236 ( .C1(n20313), .C2(n20299), .A(n20298), .B(n20297), .ZN(
        P1_U3134) );
  OAI22_X1 U23237 ( .A1(n20322), .A2(n20433), .B1(n20300), .B2(n20305), .ZN(
        n20301) );
  INV_X1 U23238 ( .A(n20301), .ZN(n20303) );
  AOI22_X1 U23239 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20309), .B1(
        n20308), .B2(n20430), .ZN(n20302) );
  OAI211_X1 U23240 ( .C1(n20313), .C2(n20304), .A(n20303), .B(n20302), .ZN(
        P1_U3135) );
  OAI22_X1 U23241 ( .A1(n20322), .A2(n20444), .B1(n20306), .B2(n20305), .ZN(
        n20307) );
  INV_X1 U23242 ( .A(n20307), .ZN(n20311) );
  AOI22_X1 U23243 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20309), .B1(
        n20308), .B2(n20438), .ZN(n20310) );
  OAI211_X1 U23244 ( .C1(n20313), .C2(n20312), .A(n20311), .B(n20310), .ZN(
        P1_U3136) );
  NOR2_X1 U23245 ( .A1(n20315), .A2(n20318), .ZN(n20337) );
  INV_X1 U23246 ( .A(n20337), .ZN(n20319) );
  NAND2_X1 U23247 ( .A1(n20350), .A2(n20316), .ZN(n20382) );
  OAI222_X1 U23248 ( .A1(n20319), .A2(n20516), .B1(n20448), .B2(n20318), .C1(
        n20317), .C2(n20382), .ZN(n20338) );
  AOI22_X1 U23249 ( .A1(n20338), .A2(n20386), .B1(n20385), .B2(n20337), .ZN(
        n20324) );
  NOR3_X1 U23250 ( .A1(n20389), .A2(n20320), .A3(n20516), .ZN(n20522) );
  OAI21_X1 U23251 ( .B1(n20321), .B2(n20522), .A(n20390), .ZN(n20340) );
  INV_X1 U23252 ( .A(n20322), .ZN(n20339) );
  AOI22_X1 U23253 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20340), .B1(
        n20339), .B2(n20392), .ZN(n20323) );
  OAI211_X1 U23254 ( .C1(n20395), .C2(n20355), .A(n20324), .B(n20323), .ZN(
        P1_U3137) );
  AOI22_X1 U23255 ( .A1(n20338), .A2(n20397), .B1(n20396), .B2(n20337), .ZN(
        n20326) );
  AOI22_X1 U23256 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20340), .B1(
        n20339), .B2(n20398), .ZN(n20325) );
  OAI211_X1 U23257 ( .C1(n20401), .C2(n20355), .A(n20326), .B(n20325), .ZN(
        P1_U3138) );
  AOI22_X1 U23258 ( .A1(n20338), .A2(n20403), .B1(n20402), .B2(n20337), .ZN(
        n20328) );
  AOI22_X1 U23259 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20340), .B1(
        n20339), .B2(n20360), .ZN(n20327) );
  OAI211_X1 U23260 ( .C1(n20363), .C2(n20355), .A(n20328), .B(n20327), .ZN(
        P1_U3139) );
  AOI22_X1 U23261 ( .A1(n20338), .A2(n20409), .B1(n20408), .B2(n20337), .ZN(
        n20330) );
  AOI22_X1 U23262 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20340), .B1(
        n20339), .B2(n20410), .ZN(n20329) );
  OAI211_X1 U23263 ( .C1(n20413), .C2(n20355), .A(n20330), .B(n20329), .ZN(
        P1_U3140) );
  AOI22_X1 U23264 ( .A1(n20338), .A2(n20415), .B1(n20414), .B2(n20337), .ZN(
        n20332) );
  AOI22_X1 U23265 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20340), .B1(
        n20339), .B2(n20366), .ZN(n20331) );
  OAI211_X1 U23266 ( .C1(n20369), .C2(n20355), .A(n20332), .B(n20331), .ZN(
        P1_U3141) );
  AOI22_X1 U23267 ( .A1(n20338), .A2(n20421), .B1(n20420), .B2(n20337), .ZN(
        n20334) );
  AOI22_X1 U23268 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20340), .B1(
        n20339), .B2(n20370), .ZN(n20333) );
  OAI211_X1 U23269 ( .C1(n20373), .C2(n20355), .A(n20334), .B(n20333), .ZN(
        P1_U3142) );
  AOI22_X1 U23270 ( .A1(n20338), .A2(n20429), .B1(n20428), .B2(n20337), .ZN(
        n20336) );
  AOI22_X1 U23271 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20340), .B1(
        n20339), .B2(n20430), .ZN(n20335) );
  OAI211_X1 U23272 ( .C1(n20433), .C2(n20355), .A(n20336), .B(n20335), .ZN(
        P1_U3143) );
  AOI22_X1 U23273 ( .A1(n20338), .A2(n20436), .B1(n20434), .B2(n20337), .ZN(
        n20342) );
  AOI22_X1 U23274 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20340), .B1(
        n20339), .B2(n20438), .ZN(n20341) );
  OAI211_X1 U23275 ( .C1(n20444), .C2(n20355), .A(n20342), .B(n20341), .ZN(
        P1_U3144) );
  INV_X1 U23276 ( .A(n20344), .ZN(n20346) );
  OAI22_X1 U23277 ( .A1(n20382), .A2(n12952), .B1(n20346), .B2(n20345), .ZN(
        n20377) );
  NOR2_X1 U23278 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20388), .ZN(
        n20376) );
  AOI22_X1 U23279 ( .A1(n20377), .A2(n20386), .B1(n20385), .B2(n20376), .ZN(
        n20357) );
  AOI21_X1 U23280 ( .B1(n20426), .B2(n20355), .A(n20347), .ZN(n20348) );
  AOI21_X1 U23281 ( .B1(n20350), .B2(n20349), .A(n20348), .ZN(n20351) );
  NOR2_X1 U23282 ( .A1(n20351), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20354) );
  AOI22_X1 U23283 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20379), .B1(
        n20378), .B2(n20392), .ZN(n20356) );
  OAI211_X1 U23284 ( .C1(n20395), .C2(n20426), .A(n20357), .B(n20356), .ZN(
        P1_U3145) );
  AOI22_X1 U23285 ( .A1(n20377), .A2(n20397), .B1(n20396), .B2(n20376), .ZN(
        n20359) );
  AOI22_X1 U23286 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20379), .B1(
        n20378), .B2(n20398), .ZN(n20358) );
  OAI211_X1 U23287 ( .C1(n20401), .C2(n20426), .A(n20359), .B(n20358), .ZN(
        P1_U3146) );
  AOI22_X1 U23288 ( .A1(n20377), .A2(n20403), .B1(n20402), .B2(n20376), .ZN(
        n20362) );
  AOI22_X1 U23289 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20379), .B1(
        n20378), .B2(n20360), .ZN(n20361) );
  OAI211_X1 U23290 ( .C1(n20363), .C2(n20426), .A(n20362), .B(n20361), .ZN(
        P1_U3147) );
  AOI22_X1 U23291 ( .A1(n20377), .A2(n20409), .B1(n20408), .B2(n20376), .ZN(
        n20365) );
  AOI22_X1 U23292 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20379), .B1(
        n20378), .B2(n20410), .ZN(n20364) );
  OAI211_X1 U23293 ( .C1(n20413), .C2(n20426), .A(n20365), .B(n20364), .ZN(
        P1_U3148) );
  AOI22_X1 U23294 ( .A1(n20377), .A2(n20415), .B1(n20414), .B2(n20376), .ZN(
        n20368) );
  AOI22_X1 U23295 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20379), .B1(
        n20378), .B2(n20366), .ZN(n20367) );
  OAI211_X1 U23296 ( .C1(n20369), .C2(n20426), .A(n20368), .B(n20367), .ZN(
        P1_U3149) );
  AOI22_X1 U23297 ( .A1(n20377), .A2(n20421), .B1(n20420), .B2(n20376), .ZN(
        n20372) );
  AOI22_X1 U23298 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20379), .B1(
        n20378), .B2(n20370), .ZN(n20371) );
  OAI211_X1 U23299 ( .C1(n20373), .C2(n20426), .A(n20372), .B(n20371), .ZN(
        P1_U3150) );
  AOI22_X1 U23300 ( .A1(n20377), .A2(n20429), .B1(n20428), .B2(n20376), .ZN(
        n20375) );
  AOI22_X1 U23301 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20379), .B1(
        n20378), .B2(n20430), .ZN(n20374) );
  OAI211_X1 U23302 ( .C1(n20433), .C2(n20426), .A(n20375), .B(n20374), .ZN(
        P1_U3151) );
  AOI22_X1 U23303 ( .A1(n20377), .A2(n20436), .B1(n20434), .B2(n20376), .ZN(
        n20381) );
  AOI22_X1 U23304 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20379), .B1(
        n20378), .B2(n20438), .ZN(n20380) );
  OAI211_X1 U23305 ( .C1(n20444), .C2(n20426), .A(n20381), .B(n20380), .ZN(
        P1_U3152) );
  OAI222_X1 U23306 ( .A1(n20516), .A2(n20384), .B1(n20448), .B2(n20388), .C1(
        n20383), .C2(n20382), .ZN(n20437) );
  INV_X1 U23307 ( .A(n20384), .ZN(n20435) );
  AOI22_X1 U23308 ( .A1(n20437), .A2(n20386), .B1(n20435), .B2(n20385), .ZN(
        n20394) );
  INV_X1 U23309 ( .A(n20387), .ZN(n20520) );
  OAI21_X1 U23310 ( .B1(n20389), .B2(n20520), .A(n20388), .ZN(n20391) );
  NAND2_X1 U23311 ( .A1(n20391), .A2(n20390), .ZN(n20440) );
  INV_X1 U23312 ( .A(n20426), .ZN(n20439) );
  AOI22_X1 U23313 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20440), .B1(
        n20439), .B2(n20392), .ZN(n20393) );
  OAI211_X1 U23314 ( .C1(n20395), .C2(n20443), .A(n20394), .B(n20393), .ZN(
        P1_U3153) );
  AOI22_X1 U23315 ( .A1(n20437), .A2(n20397), .B1(n20435), .B2(n20396), .ZN(
        n20400) );
  AOI22_X1 U23316 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20440), .B1(
        n20439), .B2(n20398), .ZN(n20399) );
  OAI211_X1 U23317 ( .C1(n20401), .C2(n20443), .A(n20400), .B(n20399), .ZN(
        P1_U3154) );
  AOI22_X1 U23318 ( .A1(n20437), .A2(n20403), .B1(n20435), .B2(n20402), .ZN(
        n20406) );
  AOI22_X1 U23319 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20440), .B1(
        n20423), .B2(n20404), .ZN(n20405) );
  OAI211_X1 U23320 ( .C1(n20407), .C2(n20426), .A(n20406), .B(n20405), .ZN(
        P1_U3155) );
  AOI22_X1 U23321 ( .A1(n20437), .A2(n20409), .B1(n20435), .B2(n20408), .ZN(
        n20412) );
  AOI22_X1 U23322 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20440), .B1(
        n20439), .B2(n20410), .ZN(n20411) );
  OAI211_X1 U23323 ( .C1(n20413), .C2(n20443), .A(n20412), .B(n20411), .ZN(
        P1_U3156) );
  AOI22_X1 U23324 ( .A1(n20437), .A2(n20415), .B1(n20435), .B2(n20414), .ZN(
        n20418) );
  AOI22_X1 U23325 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20440), .B1(
        n20423), .B2(n20416), .ZN(n20417) );
  OAI211_X1 U23326 ( .C1(n20419), .C2(n20426), .A(n20418), .B(n20417), .ZN(
        P1_U3157) );
  AOI22_X1 U23327 ( .A1(n20437), .A2(n20421), .B1(n20435), .B2(n20420), .ZN(
        n20425) );
  AOI22_X1 U23328 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20440), .B1(
        n20423), .B2(n20422), .ZN(n20424) );
  OAI211_X1 U23329 ( .C1(n20427), .C2(n20426), .A(n20425), .B(n20424), .ZN(
        P1_U3158) );
  AOI22_X1 U23330 ( .A1(n20437), .A2(n20429), .B1(n20435), .B2(n20428), .ZN(
        n20432) );
  AOI22_X1 U23331 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20440), .B1(
        n20439), .B2(n20430), .ZN(n20431) );
  OAI211_X1 U23332 ( .C1(n20433), .C2(n20443), .A(n20432), .B(n20431), .ZN(
        P1_U3159) );
  AOI22_X1 U23333 ( .A1(n20437), .A2(n20436), .B1(n20435), .B2(n20434), .ZN(
        n20442) );
  AOI22_X1 U23334 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20440), .B1(
        n20439), .B2(n20438), .ZN(n20441) );
  OAI211_X1 U23335 ( .C1(n20444), .C2(n20443), .A(n20442), .B(n20441), .ZN(
        P1_U3160) );
  NOR2_X1 U23336 ( .A1(n20446), .A2(n20445), .ZN(n20449) );
  OAI21_X1 U23337 ( .B1(n20449), .B2(n20448), .A(n20447), .ZN(P1_U3163) );
  AND2_X1 U23338 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20514), .ZN(
        P1_U3164) );
  INV_X1 U23339 ( .A(P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n20607) );
  NOR2_X1 U23340 ( .A1(n20450), .A2(n20607), .ZN(P1_U3165) );
  AND2_X1 U23341 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20514), .ZN(
        P1_U3166) );
  AND2_X1 U23342 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20514), .ZN(
        P1_U3167) );
  AND2_X1 U23343 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20514), .ZN(
        P1_U3168) );
  AND2_X1 U23344 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20514), .ZN(
        P1_U3169) );
  AND2_X1 U23345 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20514), .ZN(
        P1_U3170) );
  AND2_X1 U23346 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20514), .ZN(
        P1_U3171) );
  AND2_X1 U23347 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20514), .ZN(
        P1_U3172) );
  AND2_X1 U23348 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20514), .ZN(
        P1_U3173) );
  AND2_X1 U23349 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20514), .ZN(
        P1_U3174) );
  AND2_X1 U23350 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20514), .ZN(
        P1_U3175) );
  AND2_X1 U23351 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20514), .ZN(
        P1_U3176) );
  AND2_X1 U23352 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20514), .ZN(
        P1_U3177) );
  AND2_X1 U23353 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20514), .ZN(
        P1_U3178) );
  AND2_X1 U23354 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20514), .ZN(
        P1_U3179) );
  AND2_X1 U23355 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20514), .ZN(
        P1_U3180) );
  AND2_X1 U23356 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20514), .ZN(
        P1_U3181) );
  INV_X1 U23357 ( .A(P1_DATAWIDTH_REG_13__SCAN_IN), .ZN(n20671) );
  NOR2_X1 U23358 ( .A1(n20450), .A2(n20671), .ZN(P1_U3182) );
  INV_X1 U23359 ( .A(P1_DATAWIDTH_REG_12__SCAN_IN), .ZN(n20639) );
  NOR2_X1 U23360 ( .A1(n20450), .A2(n20639), .ZN(P1_U3183) );
  AND2_X1 U23361 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20514), .ZN(
        P1_U3184) );
  AND2_X1 U23362 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20514), .ZN(
        P1_U3185) );
  AND2_X1 U23363 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20514), .ZN(P1_U3186) );
  AND2_X1 U23364 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20514), .ZN(P1_U3187) );
  AND2_X1 U23365 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20514), .ZN(P1_U3188) );
  AND2_X1 U23366 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20514), .ZN(P1_U3189) );
  AND2_X1 U23367 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20514), .ZN(P1_U3190) );
  INV_X1 U23368 ( .A(P1_DATAWIDTH_REG_4__SCAN_IN), .ZN(n20665) );
  NOR2_X1 U23369 ( .A1(n20450), .A2(n20665), .ZN(P1_U3191) );
  AND2_X1 U23370 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20514), .ZN(P1_U3192) );
  AND2_X1 U23371 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20514), .ZN(P1_U3193) );
  AOI21_X1 U23372 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20457), .A(n20451), 
        .ZN(n20466) );
  OAI211_X1 U23373 ( .C1(P1_STATE_REG_0__SCAN_IN), .C2(n20458), .A(
        P1_REQUESTPENDING_REG_SCAN_IN), .B(n20452), .ZN(n20453) );
  NOR2_X1 U23374 ( .A1(n20454), .A2(n20453), .ZN(n20455) );
  OAI22_X1 U23375 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20466), .B1(n20540), 
        .B2(n20455), .ZN(P1_U3194) );
  OAI21_X1 U23376 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n20456), .A(n20458), 
        .ZN(n20464) );
  NAND3_X1 U23377 ( .A1(n20458), .A2(n20457), .A3(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20460) );
  NAND2_X1 U23378 ( .A1(n20460), .A2(n20459), .ZN(n20461) );
  OAI211_X1 U23379 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20462), .A(HOLD), .B(
        n20461), .ZN(n20463) );
  OAI221_X1 U23380 ( .B1(n20466), .B2(n20465), .C1(n20466), .C2(n20464), .A(
        n20463), .ZN(P1_U3196) );
  OR2_X1 U23381 ( .A1(n20503), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20506) );
  INV_X1 U23382 ( .A(n20506), .ZN(n20499) );
  NAND2_X1 U23383 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20540), .ZN(n20501) );
  INV_X1 U23384 ( .A(n20501), .ZN(n20504) );
  AOI222_X1 U23385 ( .A1(n20499), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n20503), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n20504), .ZN(n20467) );
  INV_X1 U23386 ( .A(n20467), .ZN(P1_U3197) );
  AOI222_X1 U23387 ( .A1(n20504), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n20503), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n20499), .ZN(n20468) );
  INV_X1 U23388 ( .A(n20468), .ZN(P1_U3198) );
  OAI222_X1 U23389 ( .A1(n20501), .A2(n12998), .B1(n20469), .B2(n20540), .C1(
        n20471), .C2(n20506), .ZN(P1_U3199) );
  AOI22_X1 U23390 ( .A1(P1_ADDRESS_REG_3__SCAN_IN), .A2(n20503), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n20499), .ZN(n20470) );
  OAI21_X1 U23391 ( .B1(n20471), .B2(n20501), .A(n20470), .ZN(P1_U3200) );
  AOI22_X1 U23392 ( .A1(P1_ADDRESS_REG_4__SCAN_IN), .A2(n20503), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n20504), .ZN(n20472) );
  OAI21_X1 U23393 ( .B1(n20596), .B2(n20506), .A(n20472), .ZN(P1_U3201) );
  AOI222_X1 U23394 ( .A1(n20504), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20503), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n20499), .ZN(n20473) );
  INV_X1 U23395 ( .A(n20473), .ZN(P1_U3202) );
  AOI222_X1 U23396 ( .A1(n20504), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n20503), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20499), .ZN(n20474) );
  INV_X1 U23397 ( .A(n20474), .ZN(P1_U3203) );
  AOI222_X1 U23398 ( .A1(n20504), .A2(P1_REIP_REG_8__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n20503), .C1(P1_REIP_REG_9__SCAN_IN), 
        .C2(n20499), .ZN(n20475) );
  INV_X1 U23399 ( .A(n20475), .ZN(P1_U3204) );
  AOI222_X1 U23400 ( .A1(n20504), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20503), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20499), .ZN(n20476) );
  INV_X1 U23401 ( .A(n20476), .ZN(P1_U3205) );
  AOI222_X1 U23402 ( .A1(n20499), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20503), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20504), .ZN(n20477) );
  INV_X1 U23403 ( .A(n20477), .ZN(P1_U3206) );
  AOI222_X1 U23404 ( .A1(n20504), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20503), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20499), .ZN(n20478) );
  INV_X1 U23405 ( .A(n20478), .ZN(P1_U3207) );
  AOI222_X1 U23406 ( .A1(n20504), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20503), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n20499), .ZN(n20479) );
  INV_X1 U23407 ( .A(n20479), .ZN(P1_U3208) );
  AOI222_X1 U23408 ( .A1(n20504), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n20503), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20499), .ZN(n20480) );
  INV_X1 U23409 ( .A(n20480), .ZN(P1_U3209) );
  AOI222_X1 U23410 ( .A1(n20499), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n20503), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20504), .ZN(n20481) );
  INV_X1 U23411 ( .A(n20481), .ZN(P1_U3210) );
  AOI222_X1 U23412 ( .A1(n20504), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20503), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n20499), .ZN(n20482) );
  INV_X1 U23413 ( .A(n20482), .ZN(P1_U3211) );
  AOI222_X1 U23414 ( .A1(n20504), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n20503), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n20499), .ZN(n20483) );
  INV_X1 U23415 ( .A(n20483), .ZN(P1_U3212) );
  AOI222_X1 U23416 ( .A1(n20504), .A2(P1_REIP_REG_17__SCAN_IN), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n20503), .C1(P1_REIP_REG_18__SCAN_IN), 
        .C2(n20499), .ZN(n20484) );
  INV_X1 U23417 ( .A(n20484), .ZN(P1_U3213) );
  AOI222_X1 U23418 ( .A1(n20504), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n20503), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20499), .ZN(n20485) );
  INV_X1 U23419 ( .A(n20485), .ZN(P1_U3214) );
  AOI22_X1 U23420 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n20503), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n20499), .ZN(n20486) );
  OAI21_X1 U23421 ( .B1(n14355), .B2(n20501), .A(n20486), .ZN(P1_U3215) );
  AOI22_X1 U23422 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(n20503), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n20504), .ZN(n20487) );
  OAI21_X1 U23423 ( .B1(n20488), .B2(n20506), .A(n20487), .ZN(P1_U3216) );
  AOI222_X1 U23424 ( .A1(n20499), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20503), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n20504), .ZN(n20489) );
  INV_X1 U23425 ( .A(n20489), .ZN(P1_U3217) );
  AOI222_X1 U23426 ( .A1(n20504), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n20503), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n20499), .ZN(n20490) );
  INV_X1 U23427 ( .A(n20490), .ZN(P1_U3218) );
  AOI222_X1 U23428 ( .A1(n20504), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n20503), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n20499), .ZN(n20491) );
  INV_X1 U23429 ( .A(n20491), .ZN(P1_U3219) );
  AOI222_X1 U23430 ( .A1(n20504), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20503), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20499), .ZN(n20492) );
  INV_X1 U23431 ( .A(n20492), .ZN(P1_U3220) );
  AOI22_X1 U23432 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n20499), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20503), .ZN(n20493) );
  OAI21_X1 U23433 ( .B1(n20494), .B2(n20501), .A(n20493), .ZN(P1_U3221) );
  AOI22_X1 U23434 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n20504), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20503), .ZN(n20495) );
  OAI21_X1 U23435 ( .B1(n20496), .B2(n20506), .A(n20495), .ZN(P1_U3222) );
  AOI222_X1 U23436 ( .A1(n20504), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20503), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20499), .ZN(n20497) );
  INV_X1 U23437 ( .A(n20497), .ZN(P1_U3223) );
  AOI222_X1 U23438 ( .A1(n20504), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20503), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20499), .ZN(n20498) );
  INV_X1 U23439 ( .A(n20498), .ZN(P1_U3224) );
  AOI22_X1 U23440 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20499), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20503), .ZN(n20500) );
  OAI21_X1 U23441 ( .B1(n20502), .B2(n20501), .A(n20500), .ZN(P1_U3225) );
  AOI22_X1 U23442 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20504), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20503), .ZN(n20505) );
  OAI21_X1 U23443 ( .B1(n20507), .B2(n20506), .A(n20505), .ZN(P1_U3226) );
  OAI22_X1 U23444 ( .A1(n20503), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20540), .ZN(n20508) );
  INV_X1 U23445 ( .A(n20508), .ZN(P1_U3458) );
  OAI22_X1 U23446 ( .A1(n20503), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20540), .ZN(n20509) );
  INV_X1 U23447 ( .A(n20509), .ZN(P1_U3459) );
  OAI22_X1 U23448 ( .A1(n20503), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20540), .ZN(n20510) );
  INV_X1 U23449 ( .A(n20510), .ZN(P1_U3460) );
  OAI22_X1 U23450 ( .A1(n20503), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20540), .ZN(n20511) );
  INV_X1 U23451 ( .A(n20511), .ZN(P1_U3461) );
  INV_X1 U23452 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20531) );
  INV_X1 U23453 ( .A(n20512), .ZN(n20513) );
  AOI21_X1 U23454 ( .B1(n20531), .B2(n20514), .A(n20513), .ZN(P1_U3464) );
  AOI21_X1 U23455 ( .B1(n20514), .B2(P1_DATAWIDTH_REG_1__SCAN_IN), .A(n20513), 
        .ZN(n20515) );
  INV_X1 U23456 ( .A(n20515), .ZN(P1_U3465) );
  INV_X1 U23457 ( .A(n20517), .ZN(n20519) );
  OAI22_X1 U23458 ( .A1(n20521), .A2(n20520), .B1(n20519), .B2(n20518), .ZN(
        n20523) );
  AOI211_X1 U23459 ( .C1(n20525), .C2(n20524), .A(n20523), .B(n20522), .ZN(
        n20527) );
  AOI22_X1 U23460 ( .A1(n20529), .A2(n20528), .B1(n20527), .B2(n20526), .ZN(
        P1_U3475) );
  NOR3_X1 U23461 ( .A1(n20531), .A2(P1_REIP_REG_0__SCAN_IN), .A3(
        P1_REIP_REG_1__SCAN_IN), .ZN(n20530) );
  AOI221_X1 U23462 ( .B1(n20532), .B2(n20531), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(P1_REIP_REG_0__SCAN_IN), .A(n20530), .ZN(n20534) );
  INV_X1 U23463 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20533) );
  INV_X1 U23464 ( .A(n20538), .ZN(n20535) );
  AOI22_X1 U23465 ( .A1(n20538), .A2(n20534), .B1(n20533), .B2(n20535), .ZN(
        P1_U3481) );
  NOR2_X1 U23466 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n20537) );
  INV_X1 U23467 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20536) );
  AOI22_X1 U23468 ( .A1(n20538), .A2(n20537), .B1(n20536), .B2(n20535), .ZN(
        P1_U3482) );
  AOI22_X1 U23469 ( .A1(n20540), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20539), 
        .B2(n20503), .ZN(P1_U3483) );
  OAI21_X1 U23470 ( .B1(n20541), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n20543) );
  OAI22_X1 U23471 ( .A1(n20544), .A2(n20543), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n20542), .ZN(n20545) );
  INV_X1 U23472 ( .A(n20545), .ZN(n20552) );
  AND3_X1 U23473 ( .A1(n20547), .A2(P1_STATE2_REG_2__SCAN_IN), .A3(n20546), 
        .ZN(n20549) );
  NOR3_X1 U23474 ( .A1(n20550), .A2(n20549), .A3(n20548), .ZN(n20551) );
  MUX2_X1 U23475 ( .A(n20552), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n20551), 
        .Z(P1_U3485) );
  MUX2_X1 U23476 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(P1_M_IO_N_REG_SCAN_IN), 
        .S(n20503), .Z(P1_U3486) );
  NOR4_X1 U23477 ( .A1(P2_ADDRESS_REG_3__SCAN_IN), .A2(
        P2_LWORD_REG_14__SCAN_IN), .A3(P2_LWORD_REG_12__SCAN_IN), .A4(
        P3_ADDRESS_REG_16__SCAN_IN), .ZN(n20555) );
  NOR4_X1 U23478 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_REIP_REG_16__SCAN_IN), .A3(BUF1_REG_14__SCAN_IN), .A4(
        P2_LWORD_REG_0__SCAN_IN), .ZN(n20554) );
  NOR4_X1 U23479 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(
        P3_STATE_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20553) );
  NAND4_X1 U23480 ( .A1(n20556), .A2(n20555), .A3(n20554), .A4(n20553), .ZN(
        n20572) );
  NOR4_X1 U23481 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(P3_EAX_REG_8__SCAN_IN), .A4(
        P3_EAX_REG_6__SCAN_IN), .ZN(n20560) );
  NOR4_X1 U23482 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_5__3__SCAN_IN), .A3(P3_INSTQUEUE_REG_5__5__SCAN_IN), 
        .A4(P3_EBX_REG_17__SCAN_IN), .ZN(n20559) );
  NOR4_X1 U23483 ( .A1(BUF1_REG_7__SCAN_IN), .A2(P3_EBX_REG_24__SCAN_IN), .A3(
        P1_DATAO_REG_8__SCAN_IN), .A4(P2_DATAO_REG_17__SCAN_IN), .ZN(n20558)
         );
  NOR4_X1 U23484 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_12__7__SCAN_IN), .A3(BUF1_REG_29__SCAN_IN), .A4(
        BUF2_REG_18__SCAN_IN), .ZN(n20557) );
  NAND4_X1 U23485 ( .A1(n20560), .A2(n20559), .A3(n20558), .A4(n20557), .ZN(
        n20571) );
  NOR4_X1 U23486 ( .A1(n13301), .A2(n20620), .A3(n20623), .A4(n20637), .ZN(
        n20564) );
  INV_X1 U23487 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20602) );
  NOR4_X1 U23488 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n20602), .A4(n20600), .ZN(
        n20563) );
  NOR4_X1 U23489 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A4(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n20561) );
  AND4_X1 U23490 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20561), .A3(
        P1_INSTQUEUE_REG_10__4__SCAN_IN), .A4(P1_REIP_REG_6__SCAN_IN), .ZN(
        n20562) );
  INV_X1 U23491 ( .A(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n20608) );
  NAND4_X1 U23492 ( .A1(n20564), .A2(n20563), .A3(n20562), .A4(
        P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n20570) );
  NAND4_X1 U23493 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(
        P2_STATE_REG_2__SCAN_IN), .A3(P3_LWORD_REG_10__SCAN_IN), .A4(
        P2_W_R_N_REG_SCAN_IN), .ZN(n20568) );
  NAND4_X1 U23494 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_9__2__SCAN_IN), .A3(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A4(P1_LWORD_REG_14__SCAN_IN), .ZN(n20567) );
  NAND4_X1 U23495 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(DATAI_26_), .A3(
        BUF1_REG_8__SCAN_IN), .A4(P2_DATAO_REG_7__SCAN_IN), .ZN(n20566) );
  NAND4_X1 U23496 ( .A1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A3(P1_DATAO_REG_24__SCAN_IN), 
        .A4(P1_DATAO_REG_18__SCAN_IN), .ZN(n20565) );
  OR4_X1 U23497 ( .A1(n20568), .A2(n20567), .A3(n20566), .A4(n20565), .ZN(
        n20569) );
  NOR4_X1 U23498 ( .A1(n20572), .A2(n20571), .A3(n20570), .A4(n20569), .ZN(
        n20711) );
  INV_X1 U23499 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n20575) );
  AOI22_X1 U23500 ( .A1(n20575), .A2(keyinput16), .B1(keyinput32), .B2(n20574), 
        .ZN(n20573) );
  OAI221_X1 U23501 ( .B1(n20575), .B2(keyinput16), .C1(n20574), .C2(keyinput32), .A(n20573), .ZN(n20588) );
  AOI22_X1 U23502 ( .A1(n20578), .A2(keyinput57), .B1(n20577), .B2(keyinput44), 
        .ZN(n20576) );
  OAI221_X1 U23503 ( .B1(n20578), .B2(keyinput57), .C1(n20577), .C2(keyinput44), .A(n20576), .ZN(n20587) );
  INV_X1 U23504 ( .A(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n20581) );
  AOI22_X1 U23505 ( .A1(n20581), .A2(keyinput37), .B1(keyinput6), .B2(n20580), 
        .ZN(n20579) );
  OAI221_X1 U23506 ( .B1(n20581), .B2(keyinput37), .C1(n20580), .C2(keyinput6), 
        .A(n20579), .ZN(n20586) );
  INV_X1 U23507 ( .A(DATAI_26_), .ZN(n20583) );
  AOI22_X1 U23508 ( .A1(n20584), .A2(keyinput3), .B1(n20583), .B2(keyinput36), 
        .ZN(n20582) );
  OAI221_X1 U23509 ( .B1(n20584), .B2(keyinput3), .C1(n20583), .C2(keyinput36), 
        .A(n20582), .ZN(n20585) );
  NOR4_X1 U23510 ( .A1(n20588), .A2(n20587), .A3(n20586), .A4(n20585), .ZN(
        n20704) );
  INV_X1 U23511 ( .A(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n20590) );
  AOI22_X1 U23512 ( .A1(n20591), .A2(keyinput0), .B1(n20590), .B2(keyinput9), 
        .ZN(n20589) );
  OAI221_X1 U23513 ( .B1(n20591), .B2(keyinput0), .C1(n20590), .C2(keyinput9), 
        .A(n20589), .ZN(n20686) );
  INV_X1 U23514 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20594) );
  AOI22_X1 U23515 ( .A1(n20594), .A2(keyinput41), .B1(keyinput25), .B2(n20593), 
        .ZN(n20592) );
  OAI221_X1 U23516 ( .B1(n20594), .B2(keyinput41), .C1(n20593), .C2(keyinput25), .A(n20592), .ZN(n20685) );
  INV_X1 U23517 ( .A(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n20597) );
  OAI22_X1 U23518 ( .A1(n20597), .A2(keyinput50), .B1(n20596), .B2(keyinput59), 
        .ZN(n20595) );
  AOI221_X1 U23519 ( .B1(n20597), .B2(keyinput50), .C1(keyinput59), .C2(n20596), .A(n20595), .ZN(n20618) );
  INV_X1 U23520 ( .A(P2_LWORD_REG_14__SCAN_IN), .ZN(n20599) );
  OAI22_X1 U23521 ( .A1(n20600), .A2(keyinput34), .B1(n20599), .B2(keyinput52), 
        .ZN(n20598) );
  AOI221_X1 U23522 ( .B1(n20600), .B2(keyinput34), .C1(keyinput52), .C2(n20599), .A(n20598), .ZN(n20617) );
  AOI22_X1 U23523 ( .A1(n20602), .A2(keyinput40), .B1(n11754), .B2(keyinput13), 
        .ZN(n20601) );
  OAI221_X1 U23524 ( .B1(n20602), .B2(keyinput40), .C1(n11754), .C2(keyinput13), .A(n20601), .ZN(n20615) );
  INV_X1 U23525 ( .A(P2_LWORD_REG_12__SCAN_IN), .ZN(n20605) );
  AOI22_X1 U23526 ( .A1(n20605), .A2(keyinput4), .B1(n20604), .B2(keyinput19), 
        .ZN(n20603) );
  OAI221_X1 U23527 ( .B1(n20605), .B2(keyinput4), .C1(n20604), .C2(keyinput19), 
        .A(n20603), .ZN(n20614) );
  AOI22_X1 U23528 ( .A1(n20608), .A2(keyinput48), .B1(keyinput15), .B2(n20607), 
        .ZN(n20606) );
  OAI221_X1 U23529 ( .B1(n20608), .B2(keyinput48), .C1(n20607), .C2(keyinput15), .A(n20606), .ZN(n20613) );
  AOI22_X1 U23530 ( .A1(n20611), .A2(keyinput7), .B1(keyinput39), .B2(n20610), 
        .ZN(n20609) );
  OAI221_X1 U23531 ( .B1(n20611), .B2(keyinput7), .C1(n20610), .C2(keyinput39), 
        .A(n20609), .ZN(n20612) );
  NOR4_X1 U23532 ( .A1(n20615), .A2(n20614), .A3(n20613), .A4(n20612), .ZN(
        n20616) );
  NAND3_X1 U23533 ( .A1(n20618), .A2(n20617), .A3(n20616), .ZN(n20684) );
  INV_X1 U23534 ( .A(P3_LWORD_REG_10__SCAN_IN), .ZN(n20621) );
  AOI22_X1 U23535 ( .A1(n20621), .A2(keyinput20), .B1(n20620), .B2(keyinput12), 
        .ZN(n20619) );
  OAI221_X1 U23536 ( .B1(n20621), .B2(keyinput20), .C1(n20620), .C2(keyinput12), .A(n20619), .ZN(n20634) );
  AOI22_X1 U23537 ( .A1(n20624), .A2(keyinput54), .B1(n20623), .B2(keyinput38), 
        .ZN(n20622) );
  OAI221_X1 U23538 ( .B1(n20624), .B2(keyinput54), .C1(n20623), .C2(keyinput38), .A(n20622), .ZN(n20633) );
  AOI22_X1 U23539 ( .A1(n20627), .A2(keyinput35), .B1(keyinput28), .B2(n20626), 
        .ZN(n20625) );
  OAI221_X1 U23540 ( .B1(n20627), .B2(keyinput35), .C1(n20626), .C2(keyinput28), .A(n20625), .ZN(n20632) );
  AOI22_X1 U23541 ( .A1(n20630), .A2(keyinput11), .B1(n20629), .B2(keyinput61), 
        .ZN(n20628) );
  OAI221_X1 U23542 ( .B1(n20630), .B2(keyinput11), .C1(n20629), .C2(keyinput61), .A(n20628), .ZN(n20631) );
  NOR4_X1 U23543 ( .A1(n20634), .A2(n20633), .A3(n20632), .A4(n20631), .ZN(
        n20682) );
  AOI22_X1 U23544 ( .A1(n20637), .A2(keyinput22), .B1(keyinput58), .B2(n20636), 
        .ZN(n20635) );
  OAI221_X1 U23545 ( .B1(n20637), .B2(keyinput22), .C1(n20636), .C2(keyinput58), .A(n20635), .ZN(n20648) );
  AOI22_X1 U23546 ( .A1(n20640), .A2(keyinput1), .B1(keyinput21), .B2(n20639), 
        .ZN(n20638) );
  OAI221_X1 U23547 ( .B1(n20640), .B2(keyinput1), .C1(n20639), .C2(keyinput21), 
        .A(n20638), .ZN(n20647) );
  AOI22_X1 U23548 ( .A1(n20642), .A2(keyinput33), .B1(n13301), .B2(keyinput23), 
        .ZN(n20641) );
  OAI221_X1 U23549 ( .B1(n20642), .B2(keyinput33), .C1(n13301), .C2(keyinput23), .A(n20641), .ZN(n20646) );
  XNOR2_X1 U23550 ( .A(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B(keyinput26), .ZN(
        n20644) );
  XNOR2_X1 U23551 ( .A(keyinput17), .B(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n20643) );
  NAND2_X1 U23552 ( .A1(n20644), .A2(n20643), .ZN(n20645) );
  NOR4_X1 U23553 ( .A1(n20648), .A2(n20647), .A3(n20646), .A4(n20645), .ZN(
        n20681) );
  AOI22_X1 U23554 ( .A1(n10109), .A2(keyinput29), .B1(n20650), .B2(keyinput56), 
        .ZN(n20649) );
  OAI221_X1 U23555 ( .B1(n10109), .B2(keyinput29), .C1(n20650), .C2(keyinput56), .A(n20649), .ZN(n20663) );
  INV_X1 U23556 ( .A(P1_LWORD_REG_14__SCAN_IN), .ZN(n20652) );
  AOI22_X1 U23557 ( .A1(n20653), .A2(keyinput14), .B1(n20652), .B2(keyinput43), 
        .ZN(n20651) );
  OAI221_X1 U23558 ( .B1(n20653), .B2(keyinput14), .C1(n20652), .C2(keyinput43), .A(n20651), .ZN(n20662) );
  INV_X1 U23559 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n20656) );
  AOI22_X1 U23560 ( .A1(n20656), .A2(keyinput18), .B1(keyinput51), .B2(n20655), 
        .ZN(n20654) );
  OAI221_X1 U23561 ( .B1(n20656), .B2(keyinput18), .C1(n20655), .C2(keyinput51), .A(n20654), .ZN(n20661) );
  AOI22_X1 U23562 ( .A1(n20659), .A2(keyinput53), .B1(n20658), .B2(keyinput47), 
        .ZN(n20657) );
  OAI221_X1 U23563 ( .B1(n20659), .B2(keyinput53), .C1(n20658), .C2(keyinput47), .A(n20657), .ZN(n20660) );
  NOR4_X1 U23564 ( .A1(n20663), .A2(n20662), .A3(n20661), .A4(n20660), .ZN(
        n20680) );
  AOI22_X1 U23565 ( .A1(n20666), .A2(keyinput60), .B1(keyinput10), .B2(n20665), 
        .ZN(n20664) );
  OAI221_X1 U23566 ( .B1(n20666), .B2(keyinput60), .C1(n20665), .C2(keyinput10), .A(n20664), .ZN(n20678) );
  AOI22_X1 U23567 ( .A1(n20668), .A2(keyinput2), .B1(n12178), .B2(keyinput42), 
        .ZN(n20667) );
  OAI221_X1 U23568 ( .B1(n20668), .B2(keyinput2), .C1(n12178), .C2(keyinput42), 
        .A(n20667), .ZN(n20677) );
  INV_X1 U23569 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n20670) );
  AOI22_X1 U23570 ( .A1(n20671), .A2(keyinput30), .B1(n20670), .B2(keyinput62), 
        .ZN(n20669) );
  OAI221_X1 U23571 ( .B1(n20671), .B2(keyinput30), .C1(n20670), .C2(keyinput62), .A(n20669), .ZN(n20676) );
  XOR2_X1 U23572 ( .A(n20672), .B(keyinput55), .Z(n20674) );
  XNOR2_X1 U23573 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B(keyinput46), .ZN(
        n20673) );
  NAND2_X1 U23574 ( .A1(n20674), .A2(n20673), .ZN(n20675) );
  NOR4_X1 U23575 ( .A1(n20678), .A2(n20677), .A3(n20676), .A4(n20675), .ZN(
        n20679) );
  NAND4_X1 U23576 ( .A1(n20682), .A2(n20681), .A3(n20680), .A4(n20679), .ZN(
        n20683) );
  NOR4_X1 U23577 ( .A1(n20686), .A2(n20685), .A3(n20684), .A4(n20683), .ZN(
        n20703) );
  INV_X1 U23578 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n20689) );
  INV_X1 U23579 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n20688) );
  AOI22_X1 U23580 ( .A1(n20689), .A2(keyinput49), .B1(n20688), .B2(keyinput63), 
        .ZN(n20687) );
  OAI221_X1 U23581 ( .B1(n20689), .B2(keyinput49), .C1(n20688), .C2(keyinput63), .A(n20687), .ZN(n20693) );
  XOR2_X1 U23582 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B(keyinput24), .Z(
        n20692) );
  XNOR2_X1 U23583 ( .A(n20690), .B(keyinput27), .ZN(n20691) );
  OR3_X1 U23584 ( .A1(n20693), .A2(n20692), .A3(n20691), .ZN(n20701) );
  AOI22_X1 U23585 ( .A1(n12402), .A2(keyinput5), .B1(keyinput31), .B2(n20695), 
        .ZN(n20694) );
  OAI221_X1 U23586 ( .B1(n12402), .B2(keyinput5), .C1(n20695), .C2(keyinput31), 
        .A(n20694), .ZN(n20700) );
  INV_X1 U23587 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n20698) );
  AOI22_X1 U23588 ( .A1(n20698), .A2(keyinput45), .B1(n20697), .B2(keyinput8), 
        .ZN(n20696) );
  OAI221_X1 U23589 ( .B1(n20698), .B2(keyinput45), .C1(n20697), .C2(keyinput8), 
        .A(n20696), .ZN(n20699) );
  NOR3_X1 U23590 ( .A1(n20701), .A2(n20700), .A3(n20699), .ZN(n20702) );
  NAND3_X1 U23591 ( .A1(n20704), .A2(n20703), .A3(n20702), .ZN(n20709) );
  OAI222_X1 U23592 ( .A1(n18380), .A2(n20707), .B1(n18328), .B2(n20706), .C1(
        n20705), .C2(n18318), .ZN(n20708) );
  XOR2_X1 U23593 ( .A(n20709), .B(n20708), .Z(n20710) );
  XNOR2_X1 U23594 ( .A(n20711), .B(n20710), .ZN(P3_U3044) );
  AND2_X1 U13220 ( .A1(n12918), .A2(n14428), .ZN(n10464) );
  OR2_X1 U13234 ( .A1(n10313), .A2(n10312), .ZN(n19863) );
  BUF_X1 U16760 ( .A(n13606), .Z(n16739) );
  NAND2_X1 U13321 ( .A1(n12478), .A2(n13056), .ZN(n11247) );
  CLKBUF_X2 U11136 ( .A(n15128), .Z(n9613) );
  BUF_X1 U11048 ( .A(n14368), .Z(n9603) );
  CLKBUF_X1 U11333 ( .A(n13606), .Z(n15248) );
  XNOR2_X1 U11128 ( .A(n13860), .B(n13472), .ZN(n13856) );
  CLKBUF_X1 U12345 ( .A(n13187), .Z(n13263) );
  CLKBUF_X1 U12382 ( .A(n16072), .Z(n16079) );
  CLKBUF_X1 U12536 ( .A(n17030), .Z(n17038) );
endmodule

